/** @file vj_weights.vh
 *  @brief Viola-Jones weights data structure
 */

// assume we use haarcascade_frontalface_default.xml
`define NUM_STAGE 25
`define NUM_FEATURE 2913
`define WINDOW_SIZE 24
`define LAPTOP_WIDTH 160
`define LAPTOP_HEIGHT 120
`define PYRAMID_LEVELS 9

`define PYRAMID_WIDTHS {32'd37,32'd44,32'd53,32'd64,32'd77,32'd92,32'd111,32'd133,32'd160}
`define PYRAMID_HEIGHTS {32'd27,32'd33,32'd40,32'd48,32'd57,32'd69,32'd83,32'd99,32'd120}

`define PYRAMID_X_MAPPINGS {{8'd687,8'd683,8'd678,8'd674,8'd670,8'd665,8'd661,8'd657,8'd652,8'd648,8'd644,8'd640,8'd635,8'd631,8'd627,8'd622,8'd618,8'd614,8'd609,8'd605,8'd601,8'd596,8'd592,8'd588,8'd583,8'd579,8'd575,8'd570,8'd566,8'd562,8'd557,8'd553,8'd549,8'd544,8'd540,8'd536,8'd531,8'd527,8'd523,8'd518,8'd514,8'd510,8'd505,8'd501,8'd497,8'd492,8'd488,8'd484,8'd480,8'd475,8'd471,8'd467,8'd462,8'd458,8'd454,8'd449,8'd445,8'd441,8'd436,8'd432,8'd428,8'd423,8'd419,8'd415,8'd410,8'd406,8'd402,8'd397,8'd393,8'd389,8'd384,8'd380,8'd376,8'd371,8'd367,8'd363,8'd358,8'd354,8'd350,8'd345,8'd341,8'd337,8'd332,8'd328,8'd324,8'd320,8'd315,8'd311,8'd307,8'd302,8'd298,8'd294,8'd289,8'd285,8'd281,8'd276,8'd272,8'd268,8'd263,8'd259,8'd255,8'd250,8'd246,8'd242,8'd237,8'd233,8'd229,8'd224,8'd220,8'd216,8'd211,8'd207,8'd203,8'd198,8'd194,8'd190,8'd185,8'd181,8'd177,8'd172,8'd168,8'd164,8'd160,8'd155,8'd151,8'd147,8'd142,8'd138,8'd134,8'd129,8'd125,8'd121,8'd116,8'd112,8'd108,8'd103,8'd99,8'd95,8'd90,8'd86,8'd82,8'd77,8'd73,8'd69,8'd64,8'd60,8'd56,8'd51,8'd47,8'd43,8'd38,8'd34,8'd30,8'd25,8'd21,8'd17,8'd12,8'd8,8'd4,8'd0},{8'd578,8'd574,8'd570,8'd567,8'd563,8'd560,8'd556,8'd552,8'd549,8'd545,8'd541,8'd538,8'd534,8'd530,8'd527,8'd523,8'd520,8'd516,8'd512,8'd509,8'd505,8'd501,8'd498,8'd494,8'd490,8'd487,8'd483,8'd480,8'd476,8'd472,8'd469,8'd465,8'd461,8'd458,8'd454,8'd450,8'd447,8'd443,8'd440,8'd436,8'd432,8'd429,8'd425,8'd421,8'd418,8'd414,8'd410,8'd407,8'd403,8'd400,8'd396,8'd392,8'd389,8'd385,8'd381,8'd378,8'd374,8'd370,8'd367,8'd363,8'd360,8'd356,8'd352,8'd349,8'd345,8'd341,8'd338,8'd334,8'd330,8'd327,8'd323,8'd320,8'd316,8'd312,8'd309,8'd305,8'd301,8'd298,8'd294,8'd290,8'd287,8'd283,8'd280,8'd276,8'd272,8'd269,8'd265,8'd261,8'd258,8'd254,8'd250,8'd247,8'd243,8'd240,8'd236,8'd232,8'd229,8'd225,8'd221,8'd218,8'd214,8'd210,8'd207,8'd203,8'd200,8'd196,8'd192,8'd189,8'd185,8'd181,8'd178,8'd174,8'd170,8'd167,8'd163,8'd160,8'd156,8'd152,8'd149,8'd145,8'd141,8'd138,8'd134,8'd130,8'd127,8'd123,8'd120,8'd116,8'd112,8'd109,8'd105,8'd101,8'd98,8'd94,8'd90,8'd87,8'd83,8'd80,8'd76,8'd72,8'd69,8'd65,8'd61,8'd58,8'd54,8'd50,8'd47,8'd43,8'd40,8'd36,8'd32,8'd29,8'd25,8'd21,8'd18,8'd14,8'd10,8'd7,8'd3,8'd0},{8'd480,8'd476,8'd473,8'd470,8'd467,8'd464,8'd461,8'd458,8'd455,8'd452,8'd449,8'd446,8'd443,8'd440,8'd437,8'd434,8'd431,8'd428,8'd425,8'd422,8'd419,8'd416,8'd413,8'd410,8'd407,8'd404,8'd401,8'd398,8'd395,8'd392,8'd389,8'd386,8'd383,8'd380,8'd377,8'd374,8'd371,8'd368,8'd365,8'd362,8'd359,8'd356,8'd353,8'd350,8'd347,8'd344,8'd341,8'd338,8'd335,8'd332,8'd329,8'd326,8'd323,8'd320,8'd316,8'd313,8'd310,8'd307,8'd304,8'd301,8'd298,8'd295,8'd292,8'd289,8'd286,8'd283,8'd280,8'd277,8'd274,8'd271,8'd268,8'd265,8'd262,8'd259,8'd256,8'd253,8'd250,8'd247,8'd244,8'd241,8'd238,8'd235,8'd232,8'd229,8'd226,8'd223,8'd220,8'd217,8'd214,8'd211,8'd208,8'd205,8'd202,8'd199,8'd196,8'd193,8'd190,8'd187,8'd184,8'd181,8'd178,8'd175,8'd172,8'd169,8'd166,8'd163,8'd160,8'd156,8'd153,8'd150,8'd147,8'd144,8'd141,8'd138,8'd135,8'd132,8'd129,8'd126,8'd123,8'd120,8'd117,8'd114,8'd111,8'd108,8'd105,8'd102,8'd99,8'd96,8'd93,8'd90,8'd87,8'd84,8'd81,8'd78,8'd75,8'd72,8'd69,8'd66,8'd63,8'd60,8'd57,8'd54,8'd51,8'd48,8'd45,8'd42,8'd39,8'd36,8'd33,8'd30,8'd27,8'd24,8'd21,8'd18,8'd15,8'd12,8'd9,8'd6,8'd3,8'd0},{8'd397,8'd395,8'd392,8'd390,8'd387,8'd385,8'd382,8'd380,8'd377,8'd375,8'd372,8'd370,8'd367,8'd365,8'd362,8'd360,8'd357,8'd355,8'd352,8'd350,8'd347,8'd345,8'd342,8'd340,8'd337,8'd335,8'd332,8'd330,8'd327,8'd325,8'd322,8'd320,8'd317,8'd315,8'd312,8'd310,8'd307,8'd305,8'd302,8'd300,8'd297,8'd295,8'd292,8'd290,8'd287,8'd285,8'd282,8'd280,8'd277,8'd275,8'd272,8'd270,8'd267,8'd265,8'd262,8'd260,8'd257,8'd255,8'd252,8'd250,8'd247,8'd245,8'd242,8'd240,8'd237,8'd235,8'd232,8'd230,8'd227,8'd225,8'd222,8'd220,8'd217,8'd215,8'd212,8'd210,8'd207,8'd205,8'd202,8'd200,8'd197,8'd195,8'd192,8'd190,8'd187,8'd185,8'd182,8'd180,8'd177,8'd175,8'd172,8'd170,8'd167,8'd165,8'd162,8'd160,8'd157,8'd155,8'd152,8'd150,8'd147,8'd145,8'd142,8'd140,8'd137,8'd135,8'd132,8'd130,8'd127,8'd125,8'd122,8'd120,8'd117,8'd115,8'd112,8'd110,8'd107,8'd105,8'd102,8'd100,8'd97,8'd95,8'd92,8'd90,8'd87,8'd85,8'd82,8'd80,8'd77,8'd75,8'd72,8'd70,8'd67,8'd65,8'd62,8'd60,8'd57,8'd55,8'd52,8'd50,8'd47,8'd45,8'd42,8'd40,8'd37,8'd35,8'd32,8'd30,8'd27,8'd25,8'd22,8'd20,8'd17,8'd15,8'd12,8'd10,8'd7,8'd5,8'd2,8'd0},{8'd330,8'd328,8'd326,8'd324,8'd322,8'd320,8'd317,8'd315,8'd313,8'd311,8'd309,8'd307,8'd305,8'd303,8'd301,8'd299,8'd297,8'd295,8'd292,8'd290,8'd288,8'd286,8'd284,8'd282,8'd280,8'd278,8'd276,8'd274,8'd272,8'd270,8'd268,8'd265,8'd263,8'd261,8'd259,8'd257,8'd255,8'd253,8'd251,8'd249,8'd247,8'd245,8'd243,8'd241,8'd238,8'd236,8'd234,8'd232,8'd230,8'd228,8'd226,8'd224,8'd222,8'd220,8'd218,8'd216,8'd214,8'd211,8'd209,8'd207,8'd205,8'd203,8'd201,8'd199,8'd197,8'd195,8'd193,8'd191,8'd189,8'd187,8'd184,8'd182,8'd180,8'd178,8'd176,8'd174,8'd172,8'd170,8'd168,8'd166,8'd164,8'd162,8'd160,8'd157,8'd155,8'd153,8'd151,8'd149,8'd147,8'd145,8'd143,8'd141,8'd139,8'd137,8'd135,8'd132,8'd130,8'd128,8'd126,8'd124,8'd122,8'd120,8'd118,8'd116,8'd114,8'd112,8'd110,8'd108,8'd105,8'd103,8'd101,8'd99,8'd97,8'd95,8'd93,8'd91,8'd89,8'd87,8'd85,8'd83,8'd81,8'd78,8'd76,8'd74,8'd72,8'd70,8'd68,8'd66,8'd64,8'd62,8'd60,8'd58,8'd56,8'd54,8'd51,8'd49,8'd47,8'd45,8'd43,8'd41,8'd39,8'd37,8'd35,8'd33,8'd31,8'd29,8'd27,8'd24,8'd22,8'd20,8'd18,8'd16,8'd14,8'd12,8'd10,8'd8,8'd6,8'd4,8'd2,8'd0},{8'd276,8'd274,8'd273,8'd271,8'd269,8'd267,8'd266,8'd264,8'd262,8'd260,8'd259,8'd257,8'd255,8'd253,8'd252,8'd250,8'd248,8'd246,8'd245,8'd243,8'd241,8'd240,8'd238,8'd236,8'd234,8'd233,8'd231,8'd229,8'd227,8'd226,8'd224,8'd222,8'd220,8'd219,8'd217,8'd215,8'd213,8'd212,8'd210,8'd208,8'd206,8'd205,8'd203,8'd201,8'd200,8'd198,8'd196,8'd194,8'd193,8'd191,8'd189,8'd187,8'd186,8'd184,8'd182,8'd180,8'd179,8'd177,8'd175,8'd173,8'd172,8'd170,8'd168,8'd166,8'd165,8'd163,8'd161,8'd160,8'd158,8'd156,8'd154,8'd153,8'd151,8'd149,8'd147,8'd146,8'd144,8'd142,8'd140,8'd139,8'd137,8'd135,8'd133,8'd132,8'd130,8'd128,8'd126,8'd125,8'd123,8'd121,8'd120,8'd118,8'd116,8'd114,8'd113,8'd111,8'd109,8'd107,8'd106,8'd104,8'd102,8'd100,8'd99,8'd97,8'd95,8'd93,8'd92,8'd90,8'd88,8'd86,8'd85,8'd83,8'd81,8'd80,8'd78,8'd76,8'd74,8'd73,8'd71,8'd69,8'd67,8'd66,8'd64,8'd62,8'd60,8'd59,8'd57,8'd55,8'd53,8'd52,8'd50,8'd48,8'd46,8'd45,8'd43,8'd41,8'd40,8'd38,8'd36,8'd34,8'd33,8'd31,8'd29,8'd27,8'd26,8'd24,8'd22,8'd20,8'd19,8'd17,8'd15,8'd13,8'd12,8'd10,8'd8,8'd6,8'd5,8'd3,8'd1,8'd0},{8'd229,8'd227,8'd226,8'd224,8'd223,8'd221,8'd220,8'd219,8'd217,8'd216,8'd214,8'd213,8'd211,8'd210,8'd209,8'd207,8'd206,8'd204,8'd203,8'd201,8'd200,8'd198,8'd197,8'd196,8'd194,8'd193,8'd191,8'd190,8'd188,8'd187,8'd185,8'd184,8'd183,8'd181,8'd180,8'd178,8'd177,8'd175,8'd174,8'd172,8'd171,8'd170,8'd168,8'd167,8'd165,8'd164,8'd162,8'd161,8'd160,8'd158,8'd157,8'd155,8'd154,8'd152,8'd151,8'd149,8'd148,8'd147,8'd145,8'd144,8'd142,8'd141,8'd139,8'd138,8'd136,8'd135,8'd134,8'd132,8'd131,8'd129,8'd128,8'd126,8'd125,8'd123,8'd122,8'd121,8'd119,8'd118,8'd116,8'd115,8'd113,8'd112,8'd110,8'd109,8'd108,8'd106,8'd105,8'd103,8'd102,8'd100,8'd99,8'd98,8'd96,8'd95,8'd93,8'd92,8'd90,8'd89,8'd87,8'd86,8'd85,8'd83,8'd82,8'd80,8'd79,8'd77,8'd76,8'd74,8'd73,8'd72,8'd70,8'd69,8'd67,8'd66,8'd64,8'd63,8'd61,8'd60,8'd59,8'd57,8'd56,8'd54,8'd53,8'd51,8'd50,8'd49,8'd47,8'd46,8'd44,8'd43,8'd41,8'd40,8'd38,8'd37,8'd36,8'd34,8'd33,8'd31,8'd30,8'd28,8'd27,8'd25,8'd24,8'd23,8'd21,8'd20,8'd18,8'd17,8'd15,8'd14,8'd12,8'd11,8'd10,8'd8,8'd7,8'd5,8'd4,8'd2,8'd1,8'd0},{8'd191,8'd190,8'd188,8'd187,8'd186,8'd185,8'd184,8'd182,8'd181,8'd180,8'd179,8'd178,8'd176,8'd175,8'd174,8'd173,8'd172,8'd170,8'd169,8'd168,8'd167,8'd166,8'd164,8'd163,8'd162,8'd161,8'd160,8'd158,8'd157,8'd156,8'd155,8'd153,8'd152,8'd151,8'd150,8'd149,8'd147,8'd146,8'd145,8'd144,8'd143,8'd141,8'd140,8'd139,8'd138,8'd137,8'd135,8'd134,8'd133,8'd132,8'd131,8'd129,8'd128,8'd127,8'd126,8'd125,8'd123,8'd122,8'd121,8'd120,8'd119,8'd117,8'd116,8'd115,8'd114,8'd113,8'd111,8'd110,8'd109,8'd108,8'd107,8'd105,8'd104,8'd103,8'd102,8'd101,8'd99,8'd98,8'd97,8'd96,8'd95,8'd93,8'd92,8'd91,8'd90,8'd89,8'd87,8'd86,8'd85,8'd84,8'd83,8'd81,8'd80,8'd79,8'd78,8'd76,8'd75,8'd74,8'd73,8'd72,8'd70,8'd69,8'd68,8'd67,8'd66,8'd64,8'd63,8'd62,8'd61,8'd60,8'd58,8'd57,8'd56,8'd55,8'd54,8'd52,8'd51,8'd50,8'd49,8'd48,8'd46,8'd45,8'd44,8'd43,8'd42,8'd40,8'd39,8'd38,8'd37,8'd36,8'd34,8'd33,8'd32,8'd31,8'd30,8'd28,8'd27,8'd26,8'd25,8'd24,8'd22,8'd21,8'd20,8'd19,8'd18,8'd16,8'd15,8'd14,8'd13,8'd12,8'd10,8'd9,8'd8,8'd7,8'd6,8'd4,8'd3,8'd2,8'd1,8'd0}}
`define PYRAMID_Y_MAPPINGS {{8'd528,8'd524,8'd520,8'd515,8'd511,8'd506,8'd502,8'd497,8'd493,8'd488,8'd484,8'd480,8'd475,8'd471,8'd466,8'd462,8'd457,8'd453,8'd448,8'd444,8'd440,8'd435,8'd431,8'd426,8'd422,8'd417,8'd413,8'd408,8'd404,8'd400,8'd395,8'd391,8'd386,8'd382,8'd377,8'd373,8'd368,8'd364,8'd360,8'd355,8'd351,8'd346,8'd342,8'd337,8'd333,8'd328,8'd324,8'd320,8'd315,8'd311,8'd306,8'd302,8'd297,8'd293,8'd288,8'd284,8'd280,8'd275,8'd271,8'd266,8'd262,8'd257,8'd253,8'd248,8'd244,8'd240,8'd235,8'd231,8'd226,8'd222,8'd217,8'd213,8'd208,8'd204,8'd200,8'd195,8'd191,8'd186,8'd182,8'd177,8'd173,8'd168,8'd164,8'd160,8'd155,8'd151,8'd146,8'd142,8'd137,8'd133,8'd128,8'd124,8'd120,8'd115,8'd111,8'd106,8'd102,8'd97,8'd93,8'd88,8'd84,8'd80,8'd75,8'd71,8'd66,8'd62,8'd57,8'd53,8'd48,8'd44,8'd40,8'd35,8'd31,8'd26,8'd22,8'd17,8'd13,8'd8,8'd4,8'd0},{8'd432,8'd429,8'd425,8'd421,8'd418,8'd414,8'd410,8'd407,8'd403,8'd400,8'd396,8'd392,8'd389,8'd385,8'd381,8'd378,8'd374,8'd370,8'd367,8'd363,8'd360,8'd356,8'd352,8'd349,8'd345,8'd341,8'd338,8'd334,8'd330,8'd327,8'd323,8'd320,8'd316,8'd312,8'd309,8'd305,8'd301,8'd298,8'd294,8'd290,8'd287,8'd283,8'd280,8'd276,8'd272,8'd269,8'd265,8'd261,8'd258,8'd254,8'd250,8'd247,8'd243,8'd240,8'd236,8'd232,8'd229,8'd225,8'd221,8'd218,8'd214,8'd210,8'd207,8'd203,8'd200,8'd196,8'd192,8'd189,8'd185,8'd181,8'd178,8'd174,8'd170,8'd167,8'd163,8'd160,8'd156,8'd152,8'd149,8'd145,8'd141,8'd138,8'd134,8'd130,8'd127,8'd123,8'd120,8'd116,8'd112,8'd109,8'd105,8'd101,8'd98,8'd94,8'd90,8'd87,8'd83,8'd80,8'd76,8'd72,8'd69,8'd65,8'd61,8'd58,8'd54,8'd50,8'd47,8'd43,8'd40,8'd36,8'd32,8'd29,8'd25,8'd21,8'd18,8'd14,8'd10,8'd7,8'd3,8'd0},{8'd357,8'd354,8'd351,8'd348,8'd345,8'd342,8'd339,8'd336,8'd333,8'd330,8'd327,8'd324,8'd321,8'd318,8'd315,8'd312,8'd309,8'd306,8'd303,8'd300,8'd297,8'd294,8'd291,8'd288,8'd285,8'd282,8'd279,8'd276,8'd273,8'd270,8'd267,8'd264,8'd261,8'd258,8'd255,8'd252,8'd249,8'd246,8'd243,8'd240,8'd237,8'd234,8'd231,8'd228,8'd225,8'd222,8'd219,8'd216,8'd213,8'd210,8'd207,8'd204,8'd201,8'd198,8'd195,8'd192,8'd189,8'd186,8'd183,8'd180,8'd177,8'd174,8'd171,8'd168,8'd165,8'd162,8'd159,8'd156,8'd153,8'd150,8'd147,8'd144,8'd141,8'd138,8'd135,8'd132,8'd129,8'd126,8'd123,8'd120,8'd117,8'd114,8'd111,8'd108,8'd105,8'd102,8'd99,8'd96,8'd93,8'd90,8'd87,8'd84,8'd81,8'd78,8'd75,8'd72,8'd69,8'd66,8'd63,8'd60,8'd57,8'd54,8'd51,8'd48,8'd45,8'd42,8'd39,8'd36,8'd33,8'd30,8'd27,8'd24,8'd21,8'd18,8'd15,8'd12,8'd9,8'd6,8'd3,8'd0},{8'd297,8'd295,8'd292,8'd290,8'd287,8'd285,8'd282,8'd280,8'd277,8'd275,8'd272,8'd270,8'd267,8'd265,8'd262,8'd260,8'd257,8'd255,8'd252,8'd250,8'd247,8'd245,8'd242,8'd240,8'd237,8'd235,8'd232,8'd230,8'd227,8'd225,8'd222,8'd220,8'd217,8'd215,8'd212,8'd210,8'd207,8'd205,8'd202,8'd200,8'd197,8'd195,8'd192,8'd190,8'd187,8'd185,8'd182,8'd180,8'd177,8'd175,8'd172,8'd170,8'd167,8'd165,8'd162,8'd160,8'd157,8'd155,8'd152,8'd150,8'd147,8'd145,8'd142,8'd140,8'd137,8'd135,8'd132,8'd130,8'd127,8'd125,8'd122,8'd120,8'd117,8'd115,8'd112,8'd110,8'd107,8'd105,8'd102,8'd100,8'd97,8'd95,8'd92,8'd90,8'd87,8'd85,8'd82,8'd80,8'd77,8'd75,8'd72,8'd70,8'd67,8'd65,8'd62,8'd60,8'd57,8'd55,8'd52,8'd50,8'd47,8'd45,8'd42,8'd40,8'd37,8'd35,8'd32,8'd30,8'd27,8'd25,8'd22,8'd20,8'd17,8'd15,8'd12,8'd10,8'd7,8'd5,8'd2,8'd0},{8'd250,8'd248,8'd246,8'd244,8'd242,8'd240,8'd237,8'd235,8'd233,8'd231,8'd229,8'd227,8'd225,8'd223,8'd221,8'd218,8'd216,8'd214,8'd212,8'd210,8'd208,8'd206,8'd204,8'd202,8'd200,8'd197,8'd195,8'd193,8'd191,8'd189,8'd187,8'd185,8'd183,8'd181,8'd178,8'd176,8'd174,8'd172,8'd170,8'd168,8'd166,8'd164,8'd162,8'd160,8'd157,8'd155,8'd153,8'd151,8'd149,8'd147,8'd145,8'd143,8'd141,8'd138,8'd136,8'd134,8'd132,8'd130,8'd128,8'd126,8'd124,8'd122,8'd120,8'd117,8'd115,8'd113,8'd111,8'd109,8'd107,8'd105,8'd103,8'd101,8'd98,8'd96,8'd94,8'd92,8'd90,8'd88,8'd86,8'd84,8'd82,8'd80,8'd77,8'd75,8'd73,8'd71,8'd69,8'd67,8'd65,8'd63,8'd61,8'd58,8'd56,8'd54,8'd52,8'd50,8'd48,8'd46,8'd44,8'd42,8'd40,8'd37,8'd35,8'd33,8'd31,8'd29,8'd27,8'd25,8'd23,8'd21,8'd18,8'd16,8'd14,8'd12,8'd10,8'd8,8'd6,8'd4,8'd2,8'd0},{8'd206,8'd205,8'd203,8'd201,8'd200,8'd198,8'd196,8'd194,8'd193,8'd191,8'd189,8'd187,8'd186,8'd184,8'd182,8'd180,8'd179,8'd177,8'd175,8'd173,8'd172,8'd170,8'd168,8'd166,8'd165,8'd163,8'd161,8'd160,8'd158,8'd156,8'd154,8'd153,8'd151,8'd149,8'd147,8'd146,8'd144,8'd142,8'd140,8'd139,8'd137,8'd135,8'd133,8'd132,8'd130,8'd128,8'd126,8'd125,8'd123,8'd121,8'd120,8'd118,8'd116,8'd114,8'd113,8'd111,8'd109,8'd107,8'd106,8'd104,8'd102,8'd100,8'd99,8'd97,8'd95,8'd93,8'd92,8'd90,8'd88,8'd86,8'd85,8'd83,8'd81,8'd80,8'd78,8'd76,8'd74,8'd73,8'd71,8'd69,8'd67,8'd66,8'd64,8'd62,8'd60,8'd59,8'd57,8'd55,8'd53,8'd52,8'd50,8'd48,8'd46,8'd45,8'd43,8'd41,8'd40,8'd38,8'd36,8'd34,8'd33,8'd31,8'd29,8'd27,8'd26,8'd24,8'd22,8'd20,8'd19,8'd17,8'd15,8'd13,8'd12,8'd10,8'd8,8'd6,8'd5,8'd3,8'd1,8'd0},{8'd172,8'd170,8'd169,8'd167,8'd166,8'd164,8'd163,8'd161,8'd160,8'd159,8'd157,8'd156,8'd154,8'd153,8'd151,8'd150,8'd148,8'd147,8'd146,8'd144,8'd143,8'd141,8'd140,8'd138,8'd137,8'd135,8'd134,8'd133,8'd131,8'd130,8'd128,8'd127,8'd125,8'd124,8'd122,8'd121,8'd120,8'd118,8'd117,8'd115,8'd114,8'd112,8'd111,8'd109,8'd108,8'd106,8'd105,8'd104,8'd102,8'd101,8'd99,8'd98,8'd96,8'd95,8'd93,8'd92,8'd91,8'd89,8'd88,8'd86,8'd85,8'd83,8'd82,8'd80,8'd79,8'd78,8'd76,8'd75,8'd73,8'd72,8'd70,8'd69,8'd67,8'd66,8'd65,8'd63,8'd62,8'd60,8'd59,8'd57,8'd56,8'd54,8'd53,8'd52,8'd50,8'd49,8'd47,8'd46,8'd44,8'd43,8'd41,8'd40,8'd39,8'd37,8'd36,8'd34,8'd33,8'd31,8'd30,8'd28,8'd27,8'd26,8'd24,8'd23,8'd21,8'd20,8'd18,8'd17,8'd15,8'd14,8'd13,8'd11,8'd10,8'd8,8'd7,8'd5,8'd4,8'd2,8'd1,8'd0},{8'd144,8'd143,8'd141,8'd140,8'd139,8'd138,8'd136,8'd135,8'd134,8'd133,8'd132,8'd130,8'd129,8'd128,8'd127,8'd126,8'd124,8'd123,8'd122,8'd121,8'd120,8'd118,8'd117,8'd116,8'd115,8'd113,8'd112,8'd111,8'd110,8'd109,8'd107,8'd106,8'd105,8'd104,8'd103,8'd101,8'd100,8'd99,8'd98,8'd96,8'd95,8'd94,8'd93,8'd92,8'd90,8'd89,8'd88,8'd87,8'd86,8'd84,8'd83,8'd82,8'd81,8'd80,8'd78,8'd77,8'd76,8'd75,8'd73,8'd72,8'd71,8'd70,8'd69,8'd67,8'd66,8'd65,8'd64,8'd63,8'd61,8'd60,8'd59,8'd58,8'd56,8'd55,8'd54,8'd53,8'd52,8'd50,8'd49,8'd48,8'd47,8'd46,8'd44,8'd43,8'd42,8'd41,8'd40,8'd38,8'd37,8'd36,8'd35,8'd33,8'd32,8'd31,8'd30,8'd29,8'd27,8'd26,8'd25,8'd24,8'd23,8'd21,8'd20,8'd19,8'd18,8'd16,8'd15,8'd14,8'd13,8'd12,8'd10,8'd9,8'd8,8'd7,8'd6,8'd4,8'd3,8'd2,8'd1,8'd0}}

`define STAGE_NUM_FEATURE {32'd2913,32'd2713,32'd2502,32'd2303,32'd2122,32'd1925,32'd1729,32'd1560,32'd1405,32'd1246,32'd1109,32'd973,32'd838,32'd711,32'd596,32'd497,32'd406,32'd323,32'd251,32'd189,32'd136,32'd84,32'd52,32'd25,32'd9,32'd0}
// thresholds are negative values
`define STAGE_THRESHOLD {32'd4294966913,32'd4294966865,32'd4294966879,32'd4294966871,32'd4294966877,32'd4294966885,32'd4294966881,32'd4294966862,32'd4294966836,32'd4294966846,32'd4294966857,32'd4294966822,32'd4294966840,32'd4294966820,32'd4294966801,32'd4294966829,32'd4294966804,32'd4294966799,32'd4294966781,32'd4294966767,32'd4294966735,32'd4294966726,32'd4294966700,32'd4294966658,32'd4294966651}

`define RECTANGLE1_X1 {5'd9,5'd0,5'd16,5'd3,5'd12,5'd0,5'd15,5'd0,5'd3,5'd0,5'd15,5'd1,5'd15,5'd0,5'd18,5'd6,5'd0,5'd0,5'd11,5'd3,5'd13,5'd3,5'd13,5'd10,5'd14,5'd2,5'd6,5'd5,5'd15,5'd1,5'd13,5'd0,5'd16,5'd5,5'd3,5'd3,5'd15,5'd2,5'd11,5'd9,5'd5,5'd5,5'd9,5'd6,5'd12,5'd9,5'd6,5'd4,5'd5,5'd3,5'd9,5'd8,5'd14,5'd7,5'd10,5'd2,5'd6,5'd9,5'd5,5'd8,5'd8,5'd1,5'd9,5'd0,5'd5,5'd1,5'd0,5'd1,5'd10,5'd1,5'd8,5'd4,5'd4,5'd5,5'd8,5'd6,5'd0,5'd1,5'd9,5'd8,5'd10,5'd9,5'd10,5'd0,5'd7,5'd1,5'd6,5'd1,5'd9,5'd10,5'd11,5'd0,5'd12,5'd5,5'd6,5'd3,5'd15,5'd6,5'd12,5'd4,5'd0,5'd0,5'd6,5'd0,5'd2,5'd0,5'd6,5'd9,5'd12,5'd0,5'd12,5'd0,5'd6,5'd6,5'd10,5'd5,5'd12,5'd3,5'd13,5'd6,5'd16,5'd4,5'd4,5'd3,5'd4,5'd5,5'd3,5'd0,5'd5,5'd0,5'd14,5'd0,5'd15,5'd0,5'd14,5'd2,5'd12,5'd7,5'd12,5'd0,5'd3,5'd1,5'd19,5'd4,5'd19,5'd0,5'd6,5'd0,5'd0,5'd0,5'd18,5'd1,5'd11,5'd7,5'd6,5'd5,5'd9,5'd4,5'd6,5'd0,5'd11,5'd5,5'd9,5'd0,5'd17,5'd5,5'd3,5'd6,5'd10,5'd0,5'd18,5'd5,5'd6,5'd2,5'd5,5'd9,5'd9,5'd9,5'd2,5'd0,5'd5,5'd0,5'd0,5'd8,5'd6,5'd3,5'd16,5'd8,5'd9,5'd4,5'd5,5'd3,5'd11,5'd4,5'd9,5'd3,5'd12,5'd1,5'd6,5'd6,5'd9,5'd14,5'd6,5'd8,5'd0,5'd5,5'd3,5'd12,5'd9,5'd11,5'd0,5'd12,5'd3,5'd15,5'd0,5'd18,5'd0,5'd15,5'd4,5'd10,5'd2,5'd15,5'd2,5'd3,5'd7,5'd2,5'd2,5'd10,5'd5,5'd16,5'd0,5'd12,5'd10,5'd4,5'd7,5'd14,5'd9,5'd8,5'd4,5'd12,5'd0,5'd7,5'd4,5'd8,5'd8,5'd8,5'd9,5'd7,5'd6,5'd7,5'd4,5'd8,5'd0,5'd18,5'd1,5'd20,5'd0,5'd4,5'd3,5'd0,5'd0,5'd16,5'd1,5'd6,5'd3,5'd9,5'd3,5'd7,5'd7,5'd7,5'd1,5'd9,5'd0,5'd17,5'd0,5'd6,5'd8,5'd16,5'd8,5'd12,5'd9,5'd6,5'd0,5'd15,5'd3,5'd10,5'd4,5'd8,5'd3,5'd7,5'd4,5'd3,5'd2,5'd19,5'd0,5'd11,5'd0,5'd8,5'd1,5'd17,5'd2,5'd4,5'd0,5'd18,5'd3,5'd15,5'd1,5'd16,5'd4,5'd16,5'd2,5'd3,5'd0,5'd4,5'd6,5'd8,5'd3,5'd13,5'd1,5'd9,5'd7,5'd7,5'd3,5'd10,5'd7,5'd2,5'd1,5'd6,5'd5,5'd11,5'd1,5'd15,5'd9,5'd8,5'd6,5'd2,5'd5,5'd10,5'd8,5'd12,5'd3,5'd9,5'd0,5'd0,5'd0,5'd4,5'd8,5'd5,5'd7,5'd11,5'd7,5'd13,5'd7,5'd12,5'd3,5'd13,5'd3,5'd6,5'd8,5'd5,5'd6,5'd9,5'd8,5'd5,5'd5,5'd3,5'd1,5'd14,5'd2,5'd14,5'd0,5'd14,5'd7,5'd12,5'd0,5'd13,5'd0,5'd18,5'd1,5'd5,5'd10,5'd7,5'd5,5'd4,5'd8,5'd15,5'd6,5'd14,5'd0,5'd6,5'd0,5'd14,5'd0,5'd14,5'd0,5'd3,5'd5,5'd13,5'd0,5'd7,5'd4,5'd4,5'd6,5'd4,5'd0,5'd18,5'd8,5'd2,5'd0,5'd6,5'd5,5'd3,5'd5,5'd5,5'd9,5'd3,5'd6,5'd0,5'd4,5'd7,5'd10,5'd0,5'd13,5'd3,5'd12,5'd0,5'd15,5'd8,5'd15,5'd0,5'd16,5'd2,5'd9,5'd6,5'd2,5'd2,5'd16,5'd6,5'd15,5'd6,5'd15,5'd10,5'd15,5'd1,5'd15,5'd3,5'd10,5'd7,5'd6,5'd1,5'd8,5'd6,5'd6,5'd0,5'd15,5'd2,5'd4,5'd0,5'd7,5'd8,5'd12,5'd6,5'd12,5'd2,5'd1,5'd9,5'd9,5'd9,5'd14,5'd5,5'd4,5'd4,5'd12,5'd9,5'd5,5'd6,5'd12,5'd4,5'd15,5'd5,5'd11,5'd6,5'd11,5'd5,5'd15,5'd7,5'd0,5'd2,5'd17,5'd2,5'd5,5'd3,5'd14,5'd2,5'd3,5'd3,5'd13,5'd8,5'd10,5'd2,5'd2,5'd6,5'd10,5'd2,5'd13,5'd3,5'd3,5'd3,5'd0,5'd0,5'd1,5'd7,5'd13,5'd2,5'd4,5'd3,5'd10,5'd10,5'd6,5'd7,5'd12,5'd6,5'd15,5'd9,5'd6,5'd4,5'd7,5'd5,5'd16,5'd1,5'd7,5'd8,5'd6,5'd0,5'd7,5'd1,5'd13,5'd0,5'd7,5'd0,5'd10,5'd4,5'd7,5'd0,5'd20,5'd0,5'd19,5'd3,5'd9,5'd5,5'd3,5'd5,5'd13,5'd7,5'd15,5'd2,5'd7,5'd7,5'd20,5'd3,5'd14,5'd7,5'd11,5'd3,5'd15,5'd1,5'd19,5'd0,5'd6,5'd2,5'd13,5'd0,5'd14,5'd4,5'd14,5'd6,5'd10,5'd5,5'd14,5'd6,5'd9,5'd2,5'd12,5'd3,5'd13,5'd0,5'd7,5'd6,5'd0,5'd0,5'd4,5'd7,5'd13,5'd10,5'd13,5'd0,5'd8,5'd1,5'd7,5'd0,5'd9,5'd10,5'd5,5'd0,5'd18,5'd0,5'd19,5'd6,5'd0,5'd4,5'd4,5'd19,5'd0,5'd10,5'd3,5'd11,5'd0,5'd14,5'd8,5'd10,5'd2,5'd16,5'd6,5'd12,5'd8,5'd10,5'd7,5'd3,5'd0,5'd0,5'd3,5'd10,5'd6,5'd1,5'd0,5'd13,5'd7,5'd11,5'd7,5'd6,5'd5,5'd14,5'd5,5'd12,5'd2,5'd8,5'd6,5'd0,5'd9,5'd3,5'd0,5'd0,5'd5,5'd10,5'd0,5'd4,5'd7,5'd14,5'd2,5'd8,5'd3,5'd4,5'd4,5'd3,5'd2,5'd16,5'd3,5'd13,5'd7,5'd10,5'd4,5'd0,5'd0,5'd16,5'd3,5'd10,5'd2,5'd7,5'd5,5'd4,5'd4,5'd14,5'd3,5'd10,5'd7,5'd11,5'd5,5'd13,5'd2,5'd13,5'd0,5'd6,5'd0,5'd6,5'd1,5'd15,5'd2,5'd9,5'd0,5'd5,5'd10,5'd9,5'd7,5'd9,5'd7,5'd9,5'd7,5'd9,5'd1,5'd15,5'd0,5'd9,5'd7,5'd19,5'd3,5'd19,5'd1,5'd5,5'd0,5'd3,5'd0,5'd6,5'd2,5'd3,5'd2,5'd4,5'd0,5'd11,5'd0,5'd5,5'd5,5'd16,5'd0,5'd0,5'd7,5'd5,5'd2,5'd7,5'd7,5'd9,5'd5,5'd6,5'd4,5'd11,5'd1,5'd10,5'd2,5'd14,5'd9,5'd8,5'd5,5'd2,5'd9,5'd6,5'd8,5'd1,5'd5,5'd5,5'd0,5'd19,5'd2,5'd6,5'd9,5'd3,5'd0,5'd6,5'd4,5'd10,5'd7,5'd9,5'd5,5'd10,5'd2,5'd9,5'd0,5'd18,5'd5,5'd18,5'd1,5'd7,5'd9,5'd11,5'd0,5'd18,5'd2,5'd6,5'd0,5'd9,5'd3,5'd0,5'd4,5'd1,5'd4,5'd0,5'd14,5'd0,5'd14,5'd6,5'd12,5'd8,5'd12,5'd0,5'd13,5'd7,5'd11,5'd2,5'd7,5'd8,5'd7,5'd10,5'd13,5'd8,5'd1,5'd0,5'd14,5'd4,5'd6,5'd0,5'd10,5'd6,5'd5,5'd9,5'd11,5'd10,5'd10,5'd2,5'd3,5'd0,5'd6,5'd0,5'd16,5'd5,5'd17,5'd7,5'd3,5'd0,5'd11,5'd1,5'd11,5'd1,5'd11,5'd6,5'd11,5'd0,5'd20,5'd4,5'd3,5'd0,5'd6,5'd4,5'd6,5'd0,5'd4,5'd3,5'd15,5'd1,5'd6,5'd1,5'd1,5'd7,5'd0,5'd3,5'd15,5'd4,5'd14,5'd1,5'd15,5'd0,5'd7,5'd9,5'd4,5'd7,5'd13,5'd3,5'd14,5'd1,5'd13,5'd2,5'd16,5'd9,5'd9,5'd3,5'd9,5'd1,5'd1,5'd0,5'd9,5'd1,5'd7,5'd0,5'd9,5'd7,5'd7,5'd6,5'd11,5'd1,5'd7,5'd0,5'd4,5'd7,5'd11,5'd8,5'd7,5'd8,5'd10,5'd4,5'd9,5'd0,5'd5,5'd3,5'd8,5'd6,5'd14,5'd7,5'd10,5'd6,5'd10,5'd1,5'd14,5'd1,5'd4,5'd0,5'd0,5'd8,5'd6,5'd1,5'd13,5'd1,5'd9,5'd3,5'd15,5'd0,5'd14,5'd1,5'd5,5'd3,5'd15,5'd3,5'd8,5'd3,5'd15,5'd4,5'd6,5'd4,5'd2,5'd1,5'd3,5'd0,5'd19,5'd1,5'd9,5'd6,5'd7,5'd1,5'd17,5'd9,5'd4,5'd9,5'd11,5'd7,5'd11,5'd5,5'd15,5'd3,5'd14,5'd2,5'd6,5'd8,5'd7,5'd1,5'd12,5'd0,5'd11,5'd0,5'd18,5'd5,5'd13,5'd0,5'd1,5'd1,5'd11,5'd2,5'd13,5'd6,5'd10,5'd6,5'd6,5'd0,5'd9,5'd1,5'd13,5'd4,5'd12,5'd4,5'd11,5'd1,5'd0,5'd1,5'd3,5'd0,5'd11,5'd1,5'd11,5'd5,5'd6,5'd1,5'd5,5'd1,5'd12,5'd0,5'd20,5'd0,5'd10,5'd0,5'd8,5'd7,5'd11,5'd5,5'd7,5'd4,5'd9,5'd6,5'd15,5'd3,5'd11,5'd1,5'd6,5'd0,5'd12,5'd4,5'd2,5'd0,5'd14,5'd0,5'd6,5'd3,5'd16,5'd0,5'd8,5'd9,5'd10,5'd5,5'd0,5'd0,5'd12,5'd3,5'd6,5'd6,5'd10,5'd5,5'd8,5'd0,5'd5,5'd0,5'd12,5'd5,5'd16,5'd0,5'd18,5'd0,5'd15,5'd2,5'd16,5'd0,5'd12,5'd3,5'd15,5'd4,5'd17,5'd8,5'd13,5'd4,5'd14,5'd4,5'd6,5'd7,5'd11,5'd2,5'd14,5'd0,5'd11,5'd7,5'd0,5'd4,5'd9,5'd3,5'd14,5'd2,5'd5,5'd0,5'd8,5'd2,5'd10,5'd9,5'd7,5'd1,5'd1,5'd0,5'd14,5'd0,5'd3,5'd3,5'd5,5'd6,5'd7,5'd6,5'd12,5'd7,5'd8,5'd5,5'd15,5'd7,5'd10,5'd5,5'd13,5'd3,5'd13,5'd10,5'd7,5'd4,5'd10,5'd1,5'd15,5'd1,5'd11,5'd2,5'd14,5'd7,5'd10,5'd9,5'd6,5'd6,5'd12,5'd3,5'd6,5'd0,5'd15,5'd0,5'd4,5'd0,5'd6,5'd0,5'd6,5'd3,5'd5,5'd6,5'd9,5'd10,5'd6,5'd4,5'd16,5'd4,5'd3,5'd9,5'd4,5'd5,5'd14,5'd10,5'd14,5'd7,5'd7,5'd4,5'd14,5'd3,5'd9,5'd0,5'd14,5'd1,5'd17,5'd4,5'd14,5'd7,5'd14,5'd9,5'd9,5'd4,5'd2,5'd0,5'd3,5'd8,5'd5,5'd1,5'd6,5'd3,5'd8,5'd3,5'd7,5'd3,5'd7,5'd9,5'd7,5'd10,5'd1,5'd2,5'd2,5'd0,5'd1,5'd10,5'd6,5'd0,5'd0,5'd13,5'd0,5'd8,5'd4,5'd16,5'd0,5'd14,5'd5,5'd14,5'd5,5'd10,5'd9,5'd6,5'd9,5'd9,5'd0,5'd4,5'd5,5'd7,5'd6,5'd5,5'd8,5'd10,5'd5,5'd2,5'd3,5'd1,5'd0,5'd12,5'd9,5'd9,5'd0,5'd2,5'd0,5'd6,5'd5,5'd11,5'd6,5'd6,5'd7,5'd1,5'd5,5'd11,5'd5,5'd6,5'd4,5'd11,5'd9,5'd5,5'd6,5'd3,5'd1,5'd12,5'd1,5'd15,5'd0,5'd13,5'd5,5'd17,5'd3,5'd2,5'd1,5'd7,5'd5,5'd16,5'd3,5'd11,5'd5,5'd13,5'd0,5'd18,5'd3,5'd18,5'd6,5'd12,5'd7,5'd9,5'd9,5'd3,5'd4,5'd3,5'd8,5'd14,5'd3,5'd4,5'd8,5'd13,5'd7,5'd1,5'd8,5'd4,5'd2,5'd14,5'd4,5'd11,5'd8,5'd10,5'd4,5'd8,5'd5,5'd0,5'd0,5'd13,5'd0,5'd16,5'd3,5'd9,5'd0,5'd15,5'd0,5'd17,5'd4,5'd15,5'd2,5'd9,5'd0,5'd15,5'd2,5'd9,5'd1,5'd13,5'd6,5'd12,5'd1,5'd9,5'd0,5'd9,5'd11,5'd8,5'd8,5'd12,5'd8,5'd9,5'd2,5'd13,5'd5,5'd13,5'd3,5'd3,5'd0,5'd0,5'd8,5'd20,5'd4,5'd13,5'd2,5'd9,5'd0,5'd9,5'd0,5'd2,5'd7,5'd1,5'd13,5'd6,5'd10,5'd8,5'd12,5'd3,5'd12,5'd3,5'd12,5'd1,5'd16,5'd0,5'd17,5'd9,5'd7,5'd10,5'd4,5'd2,5'd0,5'd0,5'd8,5'd2,5'd11,5'd0,5'd8,5'd6,5'd4,5'd3,5'd9,5'd8,5'd10,5'd5,5'd6,5'd4,5'd9,5'd7,5'd10,5'd0,5'd12,5'd2,5'd1,5'd1,5'd6,5'd4,5'd18,5'd1,5'd6,5'd0,5'd10,5'd4,5'd0,5'd4,5'd10,5'd5,5'd11,5'd1,5'd15,5'd7,5'd15,5'd4,5'd3,5'd2,5'd10,5'd3,5'd17,5'd4,5'd7,5'd8,5'd10,5'd9,5'd7,5'd6,5'd10,5'd0,5'd14,5'd8,5'd6,5'd6,5'd15,5'd1,5'd10,5'd0,5'd12,5'd0,5'd14,5'd1,5'd3,5'd7,5'd14,5'd1,5'd17,5'd8,5'd9,5'd6,5'd14,5'd6,5'd10,5'd6,5'd13,5'd1,5'd2,5'd9,5'd11,5'd6,5'd10,5'd10,5'd0,5'd2,5'd2,5'd0,5'd1,5'd0,5'd3,5'd3,5'd0,5'd0,5'd15,5'd4,5'd14,5'd6,5'd5,5'd0,5'd18,5'd1,5'd3,5'd1,5'd14,5'd3,5'd14,5'd8,5'd14,5'd2,5'd10,5'd10,5'd7,5'd7,5'd15,5'd11,5'd5,5'd2,5'd18,5'd0,5'd18,5'd5,5'd6,5'd7,5'd9,5'd6,5'd2,5'd4,5'd14,5'd6,5'd7,5'd0,5'd0,5'd2,5'd2,5'd8,5'd6,5'd14,5'd6,5'd8,5'd8,5'd5,5'd9,5'd7,5'd8,5'd10,5'd5,5'd9,5'd2,5'd3,5'd0,5'd18,5'd1,5'd17,5'd0,5'd19,5'd3,5'd0,5'd4,5'd10,5'd7,5'd10,5'd6,5'd9,5'd1,5'd15,5'd1,5'd9,5'd3,5'd11,5'd2,5'd3,5'd5,5'd9,5'd5,5'd13,5'd2,5'd8,5'd0,5'd12,5'd6,5'd7,5'd7,5'd4,5'd2,5'd18,5'd3,5'd4,5'd9,5'd4,5'd2,5'd7,5'd6,5'd3,5'd0,5'd18,5'd0,5'd22,5'd7,5'd15,5'd0,5'd11,5'd1,5'd18,5'd3,5'd16,5'd4,5'd14,5'd1,5'd8,5'd0,5'd15,5'd5,5'd4,5'd0,5'd9,5'd8,5'd14,5'd3,5'd16,5'd2,5'd12,5'd4,5'd13,5'd1,5'd14,5'd0,5'd6,5'd0,5'd3,5'd0,5'd8,5'd0,5'd16,5'd1,5'd6,5'd9,5'd11,5'd7,5'd9,5'd5,5'd10,5'd8,5'd9,5'd5,5'd9,5'd3,5'd9,5'd0,5'd5,5'd0,5'd15,5'd0,5'd15,5'd3,5'd15,5'd7,5'd10,5'd0,5'd0,5'd0,5'd17,5'd0,5'd18,5'd1,5'd2,5'd0,5'd11,5'd0,5'd18,5'd0,5'd6,5'd6,5'd10,5'd0,5'd3,5'd6,5'd11,5'd5,5'd13,5'd1,5'd7,5'd2,5'd4,5'd5,5'd11,5'd6,5'd3,5'd9,5'd0,5'd4,5'd10,5'd10,5'd0,5'd0,5'd0,5'd16,5'd3,5'd6,5'd5,5'd5,5'd7,5'd10,5'd0,5'd7,5'd3,5'd8,5'd10,5'd7,5'd1,5'd10,5'd0,5'd15,5'd0,5'd15,5'd4,5'd15,5'd3,5'd15,5'd2,5'd10,5'd4,5'd8,5'd7,5'd2,5'd1,5'd9,5'd0,5'd18,5'd0,5'd8,5'd2,5'd8,5'd10,5'd4,5'd5,5'd9,5'd3,5'd0,5'd6,5'd12,5'd0,5'd18,5'd0,5'd6,5'd5,5'd13,5'd6,5'd6,5'd5,5'd2,5'd2,5'd3,5'd0,5'd18,5'd5,5'd5,5'd5,5'd13,5'd0,5'd2,5'd0,5'd3,5'd3,5'd17,5'd7,5'd15,5'd9,5'd9,5'd3,5'd16,5'd3,5'd12,5'd0,5'd2,5'd1,5'd18,5'd4,5'd14,5'd4,5'd14,5'd1,5'd5,5'd1,5'd5,5'd2,5'd13,5'd0,5'd15,5'd7,5'd16,5'd3,5'd10,5'd9,5'd15,5'd1,5'd11,5'd6,5'd12,5'd5,5'd14,5'd7,5'd10,5'd10,5'd11,5'd5,5'd16,5'd7,5'd8,5'd0,5'd20,5'd1,5'd0,5'd4,5'd14,5'd6,5'd14,5'd4,5'd14,5'd1,5'd19,5'd2,5'd3,5'd8,5'd15,5'd9,5'd6,5'd3,5'd2,5'd0,5'd7,5'd2,5'd4,5'd5,5'd2,5'd9,5'd1,5'd5,5'd0,5'd0,5'd0,5'd2,5'd12,5'd6,5'd7,5'd5,5'd10,5'd3,5'd12,5'd3,5'd10,5'd10,5'd7,5'd3,5'd8,5'd1,5'd9,5'd9,5'd12,5'd4,5'd8,5'd0,5'd12,5'd3,5'd8,5'd1,5'd9,5'd5,5'd14,5'd6,5'd5,5'd0,5'd12,5'd1,5'd12,5'd2,5'd12,5'd0,5'd1,5'd7,5'd10,5'd10,5'd5,5'd5,5'd11,5'd8,5'd5,5'd0,5'd10,5'd0,5'd4,5'd3,5'd3,5'd2,5'd3,5'd9,5'd11,5'd6,5'd11,5'd6,5'd10,5'd6,5'd15,5'd1,5'd15,5'd3,5'd15,5'd8,5'd12,5'd9,5'd7,5'd4,5'd16,5'd0,5'd9,5'd1,5'd15,5'd0,5'd7,5'd1,5'd17,5'd2,5'd2,5'd1,5'd8,5'd0,5'd13,5'd5,5'd12,5'd5,5'd11,5'd1,5'd10,5'd6,5'd6,5'd3,5'd5,5'd5,5'd13,5'd0,5'd15,5'd0,5'd20,5'd0,5'd6,5'd0,5'd6,5'd8,5'd20,5'd0,5'd6,5'd0,5'd4,5'd5,5'd8,5'd0,5'd16,5'd0,5'd16,5'd3,5'd9,5'd1,5'd1,5'd7,5'd2,5'd17,5'd6,5'd9,5'd1,5'd8,5'd6,5'd10,5'd9,5'd6,5'd1,5'd18,5'd2,5'd5,5'd7,5'd10,5'd8,5'd8,5'd9,5'd16,5'd0,5'd4,5'd5,5'd9,5'd9,5'd1,5'd5,5'd13,5'd0,5'd6,5'd0,5'd9,5'd8,5'd5,5'd3,5'd8,5'd1,5'd3,5'd7,5'd13,5'd2,5'd4,5'd7,5'd11,5'd9,5'd10,5'd4,5'd18,5'd9,5'd10,5'd5,5'd7,5'd2,5'd3,5'd0,5'd0,5'd7,5'd6,5'd4,5'd5,5'd3,5'd8,5'd1,5'd10,5'd6,5'd8,5'd3,5'd1,5'd5,5'd2,5'd0,5'd5,5'd1,5'd19,5'd2,5'd13,5'd7,5'd3,5'd5,5'd5,5'd5,5'd12,5'd0,5'd12,5'd0,5'd6,5'd4,5'd11,5'd5,5'd13,5'd0,5'd13,5'd0,5'd6,5'd9,5'd18,5'd7,5'd9,5'd6,5'd13,5'd2,5'd3,5'd2,5'd18,5'd0,5'd10,5'd6,5'd8,5'd9,5'd5,5'd2,5'd11,5'd2,5'd6,5'd8,5'd4,5'd5,5'd1,5'd0,5'd14,5'd0,5'd0,5'd0,5'd20,5'd0,5'd6,5'd0,5'd8,5'd3,5'd8,5'd2,5'd9,5'd7,5'd2,5'd4,5'd5,5'd11,5'd5,5'd11,5'd7,5'd11,5'd2,5'd8,5'd1,5'd6,5'd1,5'd9,5'd9,5'd11,5'd1,5'd3,5'd0,5'd11,5'd3,5'd7,5'd2,5'd12,5'd8,5'd13,5'd2,5'd5,5'd9,5'd4,5'd10,5'd3,5'd8,5'd10,5'd9,5'd11,5'd0,5'd6,5'd5,5'd13,5'd6,5'd15,5'd1,5'd13,5'd6,5'd12,5'd8,5'd10,5'd8,5'd6,5'd0,5'd15,5'd1,5'd0,5'd2,5'd0,5'd5,5'd13,5'd0,5'd15,5'd0,5'd13,5'd0,5'd12,5'd7,5'd3,5'd1,5'd13,5'd2,5'd3,5'd1,5'd15,5'd4,5'd12,5'd0,5'd13,5'd1,5'd1,5'd0,5'd9,5'd7,5'd12,5'd0,5'd16,5'd0,5'd19,5'd1,5'd0,5'd5,5'd13,5'd8,5'd9,5'd0,5'd4,5'd9,5'd10,5'd8,5'd12,5'd0,5'd3,5'd10,5'd3,5'd3,5'd11,5'd1,5'd10,5'd2,5'd16,5'd0,5'd15,5'd1,5'd20,5'd0,5'd10,5'd2,5'd15,5'd7,5'd17,5'd8,5'd17,5'd1,5'd8,5'd5,5'd15,5'd0,5'd12,5'd1,5'd6,5'd2,5'd4,5'd10,5'd5,5'd16,5'd3,5'd7,5'd2,5'd4,5'd8,5'd10,5'd0,5'd7,5'd0,5'd18,5'd0,5'd19,5'd0,5'd1,5'd2,5'd20,5'd3,5'd18,5'd2,5'd9,5'd3,5'd7,5'd1,5'd5,5'd6,5'd2,5'd2,5'd14,5'd0,5'd2,5'd8,5'd12,5'd3,5'd9,5'd1,5'd8,5'd5,5'd11,5'd9,5'd12,5'd4,5'd14,5'd5,5'd13,5'd1,5'd8,5'd7,5'd7,5'd0,5'd12,5'd7,5'd13,5'd1,5'd5,5'd0,5'd14,5'd6,5'd14,5'd2,5'd12,5'd7,5'd11,5'd10,5'd11,5'd1,5'd14,5'd6,5'd6,5'd3,5'd1,5'd1,5'd5,5'd1,5'd3,5'd0,5'd5,5'd0,5'd3,5'd5,5'd8,5'd7,5'd8,5'd6,5'd14,5'd8,5'd10,5'd2,5'd13,5'd0,5'd11,5'd4,5'd14,5'd6,5'd7,5'd5,5'd13,5'd4,5'd13,5'd0,5'd13,5'd0,5'd9,5'd3,5'd18,5'd0,5'd11,5'd5,5'd6,5'd3,5'd0,5'd7,5'd2,5'd12,5'd0,5'd0,5'd3,5'd3,5'd0,5'd10,5'd6,5'd11,5'd0,5'd15,5'd6,5'd12,5'd9,5'd12,5'd0,5'd15,5'd0,5'd10,5'd10,5'd5,5'd6,5'd8,5'd3,5'd15,5'd0,5'd15,5'd6,5'd4,5'd1,5'd19,5'd1,5'd17,5'd3,5'd15,5'd2,5'd8,5'd3,5'd6,5'd0,5'd5,5'd7,5'd13,5'd0,5'd10,5'd0,5'd16,5'd3,5'd16,5'd6,5'd11,5'd10,5'd0,5'd3,5'd3,5'd6,5'd14,5'd6,5'd12,5'd7,5'd11,5'd0,5'd15,5'd10,5'd21,5'd7,5'd8,5'd6,5'd21,5'd5,5'd18,5'd0,5'd14,5'd2,5'd4,5'd0,5'd18,5'd9,5'd3,5'd2,5'd17,5'd0,5'd15,5'd1,5'd14,5'd9,5'd14,5'd0,5'd5,5'd8,5'd10,5'd0,5'd3,5'd3,5'd1,5'd0,5'd6,5'd6,5'd8,5'd10,5'd5,5'd2,5'd4,5'd16,5'd10,5'd12,5'd7,5'd6,5'd3,5'd12,5'd8,5'd9,5'd11,5'd12,5'd0,5'd15,5'd2,5'd12,5'd5,5'd0,5'd4,5'd16,5'd5,5'd13,5'd1,5'd9,5'd7,5'd13,5'd0,5'd6,5'd3,5'd5,5'd0,5'd0,5'd0,5'd14,5'd0,5'd14,5'd6,5'd2,5'd3,5'd0,5'd5,5'd1,5'd4,5'd6,5'd1,5'd0,5'd0,5'd5,5'd5,5'd10,5'd1,5'd6,5'd6,5'd12,5'd9,5'd3,5'd6,5'd14,5'd1,5'd17,5'd0,5'd9,5'd0,5'd18,5'd7,5'd18,5'd6,5'd18,5'd2,5'd14,5'd7,5'd13,5'd7,5'd9,5'd1,5'd9,5'd6,5'd8,5'd0,5'd20,5'd3,5'd3,5'd0,5'd9,5'd5,5'd14,5'd0,5'd8,5'd6,5'd3,5'd9,5'd9,5'd10,5'd0,5'd16,5'd4,5'd5,5'd1,5'd14,5'd0,5'd16,5'd0,5'd6,5'd9,5'd8,5'd0,5'd6,5'd1,5'd6,5'd0,5'd15,5'd2,5'd10,5'd4,5'd12,5'd7,5'd16,5'd1,5'd17,5'd6,5'd14,5'd2,5'd4,5'd0,5'd15,5'd3,5'd15,5'd3,5'd15,5'd0,5'd10,5'd1,5'd4,5'd1,5'd14,5'd1,5'd18,5'd7,5'd13,5'd4,5'd15,5'd8,5'd8,5'd2,5'd15,5'd3,5'd15,5'd8,5'd10,5'd6,5'd5,5'd0,5'd18,5'd3,5'd18,5'd0,5'd18,5'd7,5'd16,5'd8,5'd3,5'd2,5'd3,5'd7,5'd11,5'd4,5'd5,5'd6,5'd6,5'd0,5'd10,5'd3,5'd10,5'd1,5'd12,5'd1,5'd12,5'd6,5'd3,5'd9,5'd12,5'd9,5'd5,5'd2,5'd14,5'd7,5'd9,5'd5,5'd15,5'd6,5'd12,5'd7,5'd11,5'd8,5'd8,5'd0,5'd18,5'd0,5'd9,5'd4,5'd0,5'd2,5'd14,5'd5,5'd7,5'd10,5'd9,5'd0,5'd3,5'd0,5'd8,5'd0,5'd15,5'd7,5'd15,5'd0,5'd15,5'd0,5'd7,5'd8,5'd7,5'd7,5'd6,5'd6,5'd12,5'd7,5'd13,5'd1,5'd14,5'd6,5'd12,5'd3,5'd15,5'd0,5'd10,5'd1,5'd7,5'd3,5'd17,5'd9,5'd15,5'd3,5'd14,5'd1,5'd17,5'd5,5'd9,5'd2,5'd0,5'd4,5'd1,5'd0,5'd10,5'd1,5'd5,5'd9,5'd13,5'd4,5'd3,5'd0,5'd3,5'd7,5'd7,5'd0,5'd7,5'd4,5'd9,5'd0,5'd3,5'd2,5'd13,5'd8,5'd11,5'd7,5'd13,5'd0,5'd11,5'd1,5'd18,5'd3,5'd18,5'd6,5'd11,5'd7,5'd9,5'd0,5'd2,5'd2,5'd1,5'd0,5'd6,5'd0,5'd5,5'd0,5'd5,5'd2,5'd20,5'd9,5'd5,5'd1,5'd10,5'd7,5'd6,5'd0,5'd0,5'd9,5'd3,5'd13,5'd6,5'd17,5'd8,5'd14,5'd8,5'd14,5'd2,5'd2,5'd0,5'd7,5'd6,5'd12,5'd5,5'd1,5'd0,5'd7,5'd6,5'd8,5'd5,5'd10,5'd1,5'd10,5'd4,5'd10,5'd7,5'd14,5'd1,5'd0,5'd7,5'd8,5'd0,5'd15,5'd5,5'd14,5'd2,5'd9,5'd2,5'd16,5'd0,5'd18,5'd0,5'd18,5'd7,5'd4,5'd0,5'd9,5'd7,5'd6,5'd0,5'd19,5'd0,5'd12,5'd0,5'd8,5'd1,5'd3,5'd6,5'd6,5'd0,5'd3,5'd6,5'd4,5'd4,5'd9,5'd5,5'd3,5'd2,5'd2,5'd3,5'd10,5'd0,5'd8,5'd6,5'd12,5'd0,5'd11,5'd5,5'd12,5'd0,5'd2,5'd0,5'd20,5'd2,5'd6,5'd1,5'd6,5'd0,5'd7,5'd6,5'd10,5'd1,5'd9,5'd9,5'd11,5'd4,5'd11,5'd0,5'd11,5'd4,5'd0,5'd6,5'd3,5'd8,5'd10,5'd7,5'd9,5'd9,5'd6,5'd5,5'd11,5'd1,5'd14,5'd3,5'd5,5'd1,5'd3,5'd0,5'd4,5'd1,5'd15,5'd8,5'd6,5'd3,5'd14,5'd1,5'd0,5'd1,5'd19,5'd2,5'd4,5'd0,5'd6,5'd6,5'd0,5'd17,5'd1,5'd5,5'd8,5'd12,5'd0,5'd12,5'd0,5'd18,5'd0,5'd20,5'd0,5'd2,5'd8,5'd2,5'd5,5'd0,5'd1,5'd18,5'd5,5'd3,5'd6,5'd9,5'd9,5'd5,5'd0,5'd5,5'd7,5'd9,5'd0,5'd18,5'd2,5'd10,5'd7,5'd13,5'd5,5'd5,5'd9,5'd0,5'd1,5'd6,5'd6,5'd4,5'd11,5'd5,5'd6,5'd3,5'd8,5'd3,5'd6,5'd6}
`define RECTANGLE1_Y1 {5'd1,5'd13,5'd2,5'd17,5'd17,5'd17,5'd17,5'd13,5'd15,5'd18,5'd17,5'd6,5'd17,5'd12,5'd12,5'd20,5'd16,5'd18,5'd14,5'd8,5'd8,5'd10,5'd11,5'd1,5'd12,5'd11,5'd11,5'd8,5'd8,5'd13,5'd13,5'd8,5'd8,5'd0,5'd20,5'd1,5'd1,5'd0,5'd9,5'd9,5'd8,5'd9,5'd1,5'd0,5'd0,5'd0,5'd9,5'd0,5'd2,5'd1,5'd2,5'd5,5'd5,5'd5,5'd6,5'd6,5'd8,5'd3,5'd4,5'd6,5'd14,5'd20,5'd17,5'd16,5'd17,5'd14,5'd4,5'd5,5'd5,5'd7,5'd5,5'd4,5'd4,5'd2,5'd9,5'd14,5'd3,5'd0,5'd1,5'd0,5'd6,5'd5,5'd0,5'd0,5'd7,5'd8,5'd9,5'd10,5'd12,5'd2,5'd2,5'd11,5'd11,5'd8,5'd12,5'd10,5'd10,5'd14,5'd8,5'd10,5'd12,5'd3,5'd3,5'd0,5'd5,5'd5,5'd14,5'd6,5'd6,5'd14,5'd6,5'd8,5'd8,5'd4,5'd5,5'd11,5'd6,5'd14,5'd14,5'd4,5'd4,5'd3,5'd12,5'd0,5'd0,5'd3,5'd5,5'd18,5'd18,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd16,5'd16,5'd18,5'd18,5'd19,5'd21,5'd6,5'd6,5'd6,5'd0,5'd0,5'd7,5'd5,5'd6,5'd8,5'd8,5'd11,5'd5,5'd9,5'd1,5'd6,5'd7,5'd6,5'd16,5'd16,5'd6,5'd11,5'd11,5'd0,5'd0,5'd2,5'd2,5'd5,5'd5,5'd3,5'd3,5'd0,5'd0,5'd6,5'd11,5'd12,5'd15,5'd13,5'd1,5'd6,5'd10,5'd20,5'd16,5'd6,5'd6,5'd9,5'd9,5'd6,5'd6,5'd2,5'd3,5'd9,5'd3,5'd13,5'd18,5'd12,5'd12,5'd1,5'd5,5'd4,5'd1,5'd1,5'd2,5'd14,5'd13,5'd5,5'd4,5'd1,5'd0,5'd6,5'd2,5'd2,5'd0,5'd0,5'd0,5'd0,5'd8,5'd8,5'd4,5'd9,5'd2,5'd6,5'd7,5'd2,5'd6,5'd8,5'd18,5'd15,5'd0,5'd0,5'd0,5'd1,5'd2,5'd7,5'd0,5'd0,5'd1,5'd11,5'd7,5'd17,5'd2,5'd6,5'd3,5'd2,5'd14,5'd2,5'd8,5'd6,5'd3,5'd6,5'd6,5'd18,5'd8,5'd8,5'd3,5'd2,5'd1,5'd2,5'd2,5'd9,5'd7,5'd7,5'd10,5'd10,5'd2,5'd8,5'd8,5'd8,5'd7,5'd6,5'd6,5'd6,5'd13,5'd0,5'd18,5'd6,5'd1,5'd6,5'd15,5'd1,5'd10,5'd7,5'd10,5'd10,5'd8,5'd14,5'd14,5'd15,5'd13,5'd13,5'd4,5'd10,5'd1,5'd1,5'd4,5'd12,5'd6,5'd8,5'd6,5'd0,5'd1,5'd7,5'd5,5'd5,5'd9,5'd12,5'd4,5'd0,5'd0,5'd0,5'd4,5'd17,5'd17,5'd6,5'd7,5'd7,5'd16,5'd4,5'd0,5'd19,5'd12,5'd8,5'd9,5'd5,5'd6,5'd8,5'd12,5'd1,5'd0,5'd0,5'd14,5'd14,5'd6,5'd7,5'd11,5'd0,5'd0,5'd6,5'd0,5'd1,5'd3,5'd0,5'd15,5'd1,5'd3,5'd17,5'd9,5'd7,5'd15,5'd9,5'd0,5'd0,5'd7,5'd1,5'd3,5'd0,5'd1,5'd11,5'd2,5'd6,5'd1,5'd1,5'd2,5'd0,5'd13,5'd15,5'd13,5'd13,5'd4,5'd4,5'd9,5'd0,5'd3,5'd9,5'd2,5'd3,5'd1,5'd1,5'd20,5'd20,5'd6,5'd7,5'd8,5'd20,5'd13,5'd8,5'd2,5'd13,5'd18,5'd16,5'd16,5'd13,5'd16,5'd16,5'd2,5'd10,5'd11,5'd11,5'd1,5'd9,5'd12,5'd7,5'd0,5'd6,5'd0,5'd1,5'd17,5'd12,5'd1,5'd6,5'd0,5'd0,5'd1,5'd9,5'd1,5'd4,5'd9,5'd21,5'd1,5'd0,5'd0,5'd1,5'd15,5'd10,5'd10,5'd15,5'd15,5'd6,5'd17,5'd7,5'd7,5'd11,5'd0,5'd5,5'd1,5'd4,5'd7,5'd5,5'd17,5'd1,5'd17,5'd3,5'd17,5'd12,5'd17,5'd14,5'd12,5'd7,5'd6,5'd9,5'd7,5'd6,5'd0,5'd15,5'd15,5'd13,5'd13,5'd1,5'd2,5'd7,5'd7,5'd5,5'd6,5'd7,5'd4,5'd4,5'd5,5'd10,5'd8,5'd4,5'd6,5'd5,5'd6,5'd1,5'd9,5'd6,5'd6,5'd7,5'd7,5'd8,5'd4,5'd1,5'd13,5'd1,5'd1,5'd16,5'd17,5'd12,5'd8,5'd15,5'd4,5'd21,5'd17,5'd4,5'd9,5'd11,5'd8,5'd8,5'd8,5'd11,5'd2,5'd0,5'd2,5'd0,5'd0,5'd1,5'd6,5'd2,5'd0,5'd0,5'd4,5'd0,5'd0,5'd15,5'd14,5'd18,5'd8,5'd6,5'd0,5'd2,5'd7,5'd0,5'd0,5'd2,5'd5,5'd9,5'd6,5'd4,5'd4,5'd1,5'd1,5'd10,5'd19,5'd10,5'd1,5'd11,5'd0,5'd13,5'd2,5'd1,5'd11,5'd19,5'd7,5'd4,5'd4,5'd8,5'd8,5'd16,5'd5,5'd6,5'd5,5'd12,5'd12,5'd0,5'd0,5'd1,5'd0,5'd6,5'd4,5'd6,5'd6,5'd9,5'd6,5'd20,5'd0,5'd2,5'd2,5'd16,5'd16,5'd18,5'd18,5'd20,5'd15,5'd9,5'd9,5'd6,5'd8,5'd14,5'd6,5'd6,5'd6,5'd15,5'd14,5'd18,5'd15,5'd3,5'd8,5'd4,5'd18,5'd0,5'd13,5'd11,5'd9,5'd5,5'd9,5'd10,5'd2,5'd7,5'd3,5'd21,5'd6,5'd7,5'd15,5'd0,5'd0,5'd6,5'd3,5'd8,5'd1,5'd7,5'd12,5'd2,5'd15,5'd1,5'd2,5'd17,5'd20,5'd20,5'd15,5'd15,5'd12,5'd12,5'd10,5'd10,5'd6,5'd16,5'd12,5'd3,5'd11,5'd6,5'd8,5'd0,5'd6,5'd12,5'd12,5'd14,5'd0,5'd2,5'd7,5'd9,5'd8,5'd2,5'd0,5'd0,5'd7,5'd8,5'd18,5'd5,5'd11,5'd0,5'd5,5'd8,5'd0,5'd13,5'd13,5'd10,5'd14,5'd14,5'd16,5'd18,5'd10,5'd9,5'd12,5'd6,5'd1,5'd1,5'd0,5'd10,5'd0,5'd8,5'd7,5'd7,5'd0,5'd0,5'd4,5'd0,5'd2,5'd2,5'd6,5'd5,5'd0,5'd0,5'd4,5'd0,5'd5,5'd5,5'd1,5'd1,5'd15,5'd15,5'd16,5'd18,5'd18,5'd4,5'd10,5'd16,5'd17,5'd10,5'd1,5'd5,5'd5,5'd8,5'd6,5'd8,5'd8,5'd8,5'd8,5'd8,5'd5,5'd16,5'd6,5'd13,5'd15,5'd4,5'd7,5'd4,5'd21,5'd21,5'd14,5'd14,5'd9,5'd7,5'd3,5'd0,5'd16,5'd16,5'd0,5'd4,5'd1,5'd6,5'd1,5'd0,5'd2,5'd10,5'd1,5'd1,5'd5,5'd6,5'd8,5'd16,5'd4,5'd5,5'd6,5'd3,5'd3,5'd18,5'd14,5'd14,5'd12,5'd6,5'd4,5'd0,5'd6,5'd17,5'd15,5'd2,5'd2,5'd0,5'd1,5'd4,5'd3,5'd2,5'd6,5'd20,5'd7,5'd7,5'd1,5'd6,5'd0,5'd0,5'd6,5'd6,5'd2,5'd12,5'd2,5'd2,5'd1,5'd1,5'd3,5'd7,5'd6,5'd14,5'd12,5'd12,5'd12,5'd22,5'd17,5'd6,5'd6,5'd1,5'd0,5'd6,5'd6,5'd12,5'd12,5'd6,5'd5,5'd8,5'd8,5'd1,5'd8,5'd19,5'd4,5'd16,5'd16,5'd14,5'd1,5'd1,5'd8,5'd6,5'd2,5'd9,5'd10,5'd11,5'd12,5'd3,5'd5,5'd0,5'd16,5'd4,5'd9,5'd1,5'd1,5'd6,5'd5,5'd11,5'd7,5'd14,5'd0,5'd1,5'd1,5'd0,5'd1,5'd14,5'd7,5'd1,5'd1,5'd0,5'd1,5'd16,5'd1,5'd21,5'd1,5'd14,5'd14,5'd6,5'd2,5'd10,5'd10,5'd12,5'd18,5'd10,5'd14,5'd15,5'd15,5'd17,5'd18,5'd17,5'd0,5'd1,5'd2,5'd0,5'd0,5'd5,5'd5,5'd0,5'd0,5'd3,5'd7,5'd10,5'd7,5'd1,5'd1,5'd12,5'd7,5'd8,5'd1,5'd0,5'd0,5'd6,5'd14,5'd19,5'd1,5'd6,5'd5,5'd5,5'd12,5'd13,5'd3,5'd6,5'd1,5'd8,5'd5,5'd0,5'd16,5'd10,5'd3,5'd16,5'd22,5'd7,5'd2,5'd2,5'd3,5'd3,5'd14,5'd1,5'd1,5'd0,5'd4,5'd6,5'd7,5'd4,5'd4,5'd5,5'd5,5'd8,5'd10,5'd10,5'd0,5'd15,5'd9,5'd1,5'd0,5'd14,5'd19,5'd19,5'd19,5'd18,5'd5,5'd13,5'd13,5'd15,5'd15,5'd13,5'd9,5'd7,5'd7,5'd15,5'd18,5'd18,5'd6,5'd4,5'd0,5'd1,5'd1,5'd5,5'd5,5'd0,5'd4,5'd1,5'd14,5'd18,5'd13,5'd17,5'd1,5'd13,5'd1,5'd5,5'd5,5'd0,5'd0,5'd6,5'd6,5'd5,5'd15,5'd19,5'd6,5'd2,5'd6,5'd13,5'd14,5'd1,5'd7,5'd2,5'd2,5'd0,5'd0,5'd17,5'd10,5'd20,5'd2,5'd10,5'd0,5'd12,5'd10,5'd5,5'd4,5'd1,5'd10,5'd15,5'd10,5'd12,5'd12,5'd12,5'd12,5'd12,5'd9,5'd10,5'd10,5'd8,5'd14,5'd15,5'd12,5'd6,5'd10,5'd12,5'd7,5'd8,5'd6,5'd9,5'd2,5'd13,5'd13,5'd2,5'd1,5'd0,5'd0,5'd0,5'd7,5'd4,5'd5,5'd3,5'd3,5'd0,5'd9,5'd6,5'd13,5'd15,5'd8,5'd3,5'd3,5'd12,5'd3,5'd0,5'd18,5'd16,5'd16,5'd4,5'd2,5'd3,5'd0,5'd1,5'd14,5'd15,5'd0,5'd2,5'd9,5'd0,5'd2,5'd4,5'd10,5'd15,5'd7,5'd9,5'd9,5'd10,5'd0,5'd1,5'd1,5'd6,5'd6,5'd0,5'd0,5'd2,5'd2,5'd0,5'd0,5'd12,5'd0,5'd3,5'd9,5'd10,5'd10,5'd13,5'd6,5'd6,5'd14,5'd7,5'd12,5'd12,5'd0,5'd8,5'd5,5'd8,5'd2,5'd6,5'd2,5'd6,5'd5,5'd5,5'd3,5'd18,5'd18,5'd15,5'd8,5'd16,5'd19,5'd16,5'd16,5'd0,5'd8,5'd1,5'd6,5'd3,5'd7,5'd2,5'd2,5'd2,5'd1,5'd4,5'd1,5'd3,5'd6,5'd15,5'd15,5'd21,5'd15,5'd14,5'd17,5'd0,5'd1,5'd2,5'd1,5'd4,5'd1,5'd0,5'd9,5'd8,5'd7,5'd0,5'd16,5'd0,5'd0,5'd17,5'd15,5'd14,5'd14,5'd3,5'd3,5'd15,5'd18,5'd0,5'd0,5'd6,5'd6,5'd7,5'd15,5'd5,5'd6,5'd0,5'd16,5'd13,5'd0,5'd6,5'd4,5'd20,5'd13,5'd6,5'd13,5'd2,5'd6,5'd10,5'd7,5'd10,5'd5,5'd0,5'd13,5'd1,5'd1,5'd0,5'd0,5'd16,5'd0,5'd0,5'd6,5'd6,5'd0,5'd0,5'd21,5'd8,5'd8,5'd0,5'd0,5'd0,5'd0,5'd12,5'd7,5'd14,5'd1,5'd8,5'd7,5'd14,5'd18,5'd11,5'd15,5'd2,5'd1,5'd16,5'd16,5'd9,5'd11,5'd11,5'd17,5'd18,5'd15,5'd0,5'd2,5'd11,5'd9,5'd9,5'd6,5'd0,5'd4,5'd17,5'd10,5'd15,5'd8,5'd1,5'd2,5'd4,5'd0,5'd18,5'd14,5'd14,5'd0,5'd5,5'd0,5'd1,5'd0,5'd0,5'd1,5'd0,5'd4,5'd7,5'd5,5'd4,5'd2,5'd2,5'd7,5'd11,5'd9,5'd10,5'd15,5'd18,5'd1,5'd0,5'd1,5'd2,5'd3,5'd10,5'd3,5'd21,5'd13,5'd1,5'd0,5'd13,5'd12,5'd0,5'd2,5'd0,5'd10,5'd5,5'd21,5'd21,5'd6,5'd4,5'd9,5'd9,5'd7,5'd11,5'd2,5'd2,5'd5,5'd2,5'd1,5'd1,5'd0,5'd7,5'd1,5'd21,5'd13,5'd2,5'd0,5'd0,5'd10,5'd22,5'd1,5'd3,5'd0,5'd9,5'd7,5'd4,5'd4,5'd6,5'd5,5'd5,5'd4,5'd2,5'd3,5'd9,5'd2,5'd14,5'd13,5'd18,5'd14,5'd13,5'd15,5'd18,5'd17,5'd17,5'd3,5'd2,5'd0,5'd17,5'd17,5'd13,5'd8,5'd17,5'd16,5'd7,5'd5,5'd6,5'd0,5'd0,5'd8,5'd14,5'd2,5'd2,5'd1,5'd3,5'd3,5'd3,5'd6,5'd2,5'd2,5'd5,5'd6,5'd6,5'd17,5'd6,5'd4,5'd1,5'd6,5'd4,5'd5,5'd2,5'd8,5'd18,5'd3,5'd6,5'd8,5'd0,5'd5,5'd5,5'd5,5'd4,5'd5,5'd1,5'd1,5'd4,5'd2,5'd2,5'd2,5'd0,5'd1,5'd0,5'd0,5'd15,5'd3,5'd2,5'd5,5'd9,5'd11,5'd0,5'd16,5'd11,5'd6,5'd7,5'd1,5'd2,5'd2,5'd6,5'd11,5'd15,5'd15,5'd4,5'd15,5'd13,5'd8,5'd13,5'd15,5'd8,5'd8,5'd8,5'd10,5'd10,5'd21,5'd3,5'd5,5'd2,5'd0,5'd2,5'd2,5'd2,5'd13,5'd13,5'd13,5'd8,5'd8,5'd4,5'd4,5'd2,5'd4,5'd10,5'd6,5'd5,5'd1,5'd3,5'd3,5'd8,5'd4,5'd9,5'd9,5'd6,5'd6,5'd16,5'd12,5'd16,5'd16,5'd10,5'd0,5'd1,5'd0,5'd18,5'd9,5'd6,5'd6,5'd3,5'd3,5'd20,5'd17,5'd4,5'd0,5'd0,5'd0,5'd3,5'd10,5'd15,5'd3,5'd0,5'd1,5'd7,5'd2,5'd18,5'd1,5'd7,5'd0,5'd6,5'd7,5'd2,5'd5,5'd18,5'd10,5'd16,5'd16,5'd16,5'd17,5'd1,5'd20,5'd21,5'd1,5'd15,5'd15,5'd16,5'd11,5'd4,5'd4,5'd7,5'd7,5'd12,5'd12,5'd12,5'd15,5'd7,5'd15,5'd9,5'd0,5'd6,5'd11,5'd4,5'd4,5'd0,5'd18,5'd4,5'd4,5'd0,5'd4,5'd11,5'd5,5'd10,5'd17,5'd7,5'd0,5'd11,5'd0,5'd7,5'd8,5'd2,5'd4,5'd20,5'd12,5'd0,5'd12,5'd12,5'd11,5'd1,5'd4,5'd18,5'd6,5'd8,5'd11,5'd11,5'd3,5'd3,5'd3,5'd3,5'd2,5'd2,5'd3,5'd3,5'd8,5'd8,5'd7,5'd6,5'd6,5'd4,5'd8,5'd15,5'd7,5'd11,5'd9,5'd10,5'd15,5'd12,5'd16,5'd0,5'd5,5'd2,5'd16,5'd15,5'd10,5'd10,5'd9,5'd0,5'd2,5'd12,5'd7,5'd13,5'd7,5'd14,5'd12,5'd4,5'd6,5'd6,5'd12,5'd21,5'd18,5'd9,5'd10,5'd6,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd2,5'd15,5'd7,5'd4,5'd5,5'd5,5'd8,5'd8,5'd1,5'd2,5'd0,5'd0,5'd2,5'd17,5'd16,5'd1,5'd0,5'd13,5'd12,5'd14,5'd12,5'd10,5'd7,5'd6,5'd7,5'd6,5'd11,5'd16,5'd16,5'd6,5'd6,5'd18,5'd9,5'd14,5'd9,5'd12,5'd5,5'd10,5'd8,5'd8,5'd7,5'd6,5'd5,5'd8,5'd0,5'd8,5'd7,5'd8,5'd14,5'd15,5'd15,5'd14,5'd17,5'd17,5'd0,5'd0,5'd0,5'd6,5'd2,5'd6,5'd7,5'd3,5'd0,5'd7,5'd10,5'd2,5'd0,5'd0,5'd2,5'd2,5'd0,5'd0,5'd5,5'd2,5'd10,5'd0,5'd7,5'd0,5'd0,5'd0,5'd4,5'd15,5'd10,5'd3,5'd6,5'd6,5'd5,5'd21,5'd6,5'd1,5'd4,5'd2,5'd14,5'd13,5'd3,5'd2,5'd2,5'd9,5'd2,5'd10,5'd7,5'd16,5'd1,5'd0,5'd7,5'd22,5'd4,5'd12,5'd6,5'd0,5'd0,5'd15,5'd15,5'd12,5'd12,5'd0,5'd12,5'd4,5'd4,5'd0,5'd6,5'd5,5'd5,5'd8,5'd8,5'd20,5'd18,5'd18,5'd5,5'd10,5'd4,5'd9,5'd15,5'd0,5'd14,5'd8,5'd7,5'd13,5'd2,5'd0,5'd0,5'd0,5'd0,5'd2,5'd4,5'd11,5'd11,5'd5,5'd7,5'd12,5'd1,5'd13,5'd4,5'd2,5'd2,5'd16,5'd6,5'd5,5'd17,5'd3,5'd7,5'd3,5'd18,5'd18,5'd3,5'd0,5'd0,5'd8,5'd11,5'd7,5'd3,5'd10,5'd2,5'd12,5'd0,5'd2,5'd2,5'd2,5'd2,5'd15,5'd2,5'd1,5'd0,5'd16,5'd16,5'd16,5'd16,5'd13,5'd13,5'd13,5'd3,5'd4,5'd1,5'd0,5'd13,5'd10,5'd13,5'd6,5'd8,5'd5,5'd14,5'd5,5'd6,5'd5,5'd5,5'd21,5'd12,5'd0,5'd16,5'd4,5'd0,5'd2,5'd2,5'd5,5'd5,5'd5,5'd5,5'd14,5'd14,5'd7,5'd0,5'd15,5'd22,5'd0,5'd8,5'd1,5'd4,5'd0,5'd10,5'd9,5'd1,5'd3,5'd2,5'd2,5'd9,5'd6,5'd1,5'd0,5'd4,5'd6,5'd0,5'd16,5'd16,5'd4,5'd5,5'd7,5'd1,5'd17,5'd17,5'd8,5'd15,5'd7,5'd8,5'd4,5'd7,5'd9,5'd9,5'd12,5'd17,5'd13,5'd5,5'd15,5'd10,5'd10,5'd8,5'd10,5'd9,5'd20,5'd13,5'd14,5'd0,5'd0,5'd17,5'd17,5'd17,5'd18,5'd17,5'd5,5'd5,5'd9,5'd7,5'd2,5'd0,5'd12,5'd12,5'd15,5'd5,5'd2,5'd15,5'd1,5'd1,5'd5,5'd13,5'd7,5'd7,5'd3,5'd3,5'd7,5'd1,5'd0,5'd5,5'd3,5'd0,5'd3,5'd1,5'd15,5'd15,5'd1,5'd1,5'd6,5'd6,5'd3,5'd14,5'd15,5'd11,5'd1,5'd14,5'd12,5'd6,5'd10,5'd10,5'd2,5'd2,5'd0,5'd1,5'd13,5'd12,5'd5,5'd0,5'd0,5'd12,5'd5,5'd3,5'd0,5'd6,5'd20,5'd11,5'd11,5'd11,5'd0,5'd0,5'd3,5'd3,5'd14,5'd17,5'd8,5'd11,5'd6,5'd3,5'd0,5'd0,5'd12,5'd1,5'd7,5'd12,5'd8,5'd8,5'd19,5'd8,5'd18,5'd6,5'd1,5'd3,5'd4,5'd9,5'd9,5'd0,5'd9,5'd5,5'd9,5'd4,5'd4,5'd12,5'd9,5'd11,5'd8,5'd11,5'd6,5'd10,5'd4,5'd0,5'd10,5'd12,5'd10,5'd7,5'd6,5'd5,5'd5,5'd0,5'd16,5'd8,5'd13,5'd16,5'd4,5'd7,5'd14,5'd6,5'd10,5'd9,5'd18,5'd11,5'd1,5'd0,5'd0,5'd11,5'd8,5'd14,5'd14,5'd9,5'd5,5'd7,5'd8,5'd0,5'd7,5'd2,5'd6,5'd5,5'd18,5'd17,5'd1,5'd6,5'd3,5'd3,5'd6,5'd6,5'd3,5'd12,5'd4,5'd7,5'd7,5'd4,5'd9,5'd3,5'd16,5'd3,5'd16,5'd1,5'd1,5'd0,5'd3,5'd0,5'd18,5'd4,5'd10,5'd7,5'd16,5'd6,5'd16,5'd11,5'd11,5'd6,5'd6,5'd0,5'd2,5'd10,5'd0,5'd12,5'd11,5'd14,5'd8,5'd8,5'd7,5'd4,5'd6,5'd0,5'd21,5'd12,5'd8,5'd0,5'd7,5'd6,5'd2,5'd1,5'd16,5'd12,5'd8,5'd13,5'd12,5'd14,5'd2,5'd13,5'd5,5'd15,5'd13,5'd16,5'd1,5'd2,5'd2,5'd3,5'd7,5'd17,5'd0,5'd0,5'd17,5'd2,5'd0,5'd6,5'd0,5'd7,5'd10,5'd9,5'd11,5'd10,5'd2,5'd1,5'd19,5'd1,5'd5,5'd16,5'd13,5'd6,5'd12,5'd17,5'd15,5'd20,5'd21,5'd12,5'd10,5'd11,5'd10,5'd10,5'd4,5'd0,5'd5,5'd0,5'd4,5'd3,5'd0,5'd10,5'd3,5'd0,5'd0,5'd2,5'd0,5'd11,5'd8,5'd8,5'd9,5'd5,5'd7,5'd6,5'd5,5'd8,5'd8,5'd6,5'd8,5'd17,5'd15,5'd15,5'd16,5'd0,5'd4,5'd3,5'd11,5'd11,5'd16,5'd16,5'd16,5'd10,5'd6,5'd17,5'd0,5'd4,5'd2,5'd11,5'd0,5'd10,5'd12,5'd14,5'd6,5'd10,5'd13,5'd17,5'd15,5'd2,5'd5,5'd13,5'd6,5'd5,5'd6,5'd6,5'd5,5'd5,5'd11,5'd0,5'd9,5'd10,5'd13,5'd9,5'd16,5'd16,5'd4,5'd5,5'd5,5'd5,5'd0,5'd9,5'd0,5'd6,5'd8,5'd8,5'd5,5'd2,5'd8,5'd8,5'd13,5'd15,5'd3,5'd0,5'd1,5'd10,5'd22,5'd5,5'd0,5'd0,5'd2,5'd3,5'd2,5'd18,5'd7,5'd6,5'd12,5'd7,5'd1,5'd3,5'd0,5'd10,5'd10,5'd5,5'd5,5'd6,5'd6,5'd5,5'd11,5'd9,5'd14,5'd3,5'd0,5'd5,5'd2,5'd3,5'd0,5'd2,5'd9,5'd18,5'd2,5'd7,5'd10,5'd6,5'd4,5'd5,5'd5,5'd19,5'd6,5'd9,5'd11,5'd14,5'd14,5'd5,5'd7,5'd8,5'd5,5'd2,5'd2,5'd18,5'd18,5'd4,5'd4,5'd4,5'd4,5'd2,5'd2,5'd10,5'd10,5'd4,5'd4,5'd5,5'd6,5'd6,5'd9,5'd8,5'd4,5'd10,5'd21,5'd3,5'd5,5'd6,5'd5,5'd11,5'd10,5'd0,5'd0,5'd6,5'd3,5'd18,5'd17,5'd2,5'd8,5'd7,5'd9,5'd13,5'd17,5'd16,5'd3,5'd11,5'd2,5'd0,5'd16,5'd2,5'd8,5'd4,5'd8,5'd6,5'd3,5'd2,5'd14,5'd7,5'd18,5'd0,5'd2,5'd0,5'd0,5'd15,5'd4,5'd11,5'd11,5'd12,5'd11,5'd20,5'd11,5'd0,5'd6,5'd1,5'd0,5'd6,5'd14,5'd13,5'd5,5'd8,5'd0,5'd0,5'd16,5'd16,5'd2,5'd12,5'd14,5'd14,5'd0,5'd6,5'd7,5'd9,5'd0,5'd3,5'd6,5'd6,5'd7,5'd6,5'd0,5'd0,5'd7,5'd7,5'd2,5'd2,5'd5,5'd17,5'd0,5'd0,5'd2,5'd2,5'd9,5'd15,5'd1,5'd1,5'd5,5'd5,5'd5,5'd5,5'd13,5'd14,5'd12,5'd16,5'd9,5'd5,5'd1,5'd1,5'd7,5'd14,5'd10,5'd10,5'd4,5'd10,5'd2,5'd1,5'd5,5'd13,5'd0,5'd0,5'd1,5'd3,5'd4,5'd1,5'd6,5'd7,5'd2,5'd0,5'd6,5'd0,5'd12,5'd8,5'd0,5'd0,5'd11,5'd3,5'd0,5'd0,5'd0,5'd0,5'd3,5'd3,5'd17,5'd15,5'd17,5'd3,5'd9,5'd9,5'd18,5'd18,5'd6,5'd18,5'd17,5'd7,5'd7,5'd2,5'd5,5'd6,5'd21,5'd10,5'd0,5'd6,5'd0,5'd4,5'd3,5'd4,5'd2,5'd0,5'd14,5'd6,5'd7,5'd7,5'd7,5'd3,5'd0,5'd6,5'd5,5'd6,5'd2,5'd2,5'd2,5'd7,5'd0,5'd13,5'd5,5'd7,5'd7,5'd0,5'd0,5'd4,5'd5,5'd4,5'd0,5'd13,5'd16,5'd15,5'd15,5'd17,5'd1,5'd0,5'd0,5'd7,5'd5,5'd3,5'd10,5'd13,5'd0,5'd20,5'd2,5'd12,5'd8,5'd15,5'd0,5'd0,5'd4,5'd6,5'd6,5'd17,5'd17,5'd0,5'd0,5'd12,5'd9,5'd11,5'd11,5'd14,5'd14,5'd22,5'd4,5'd4,5'd4,5'd6,5'd4,5'd5,5'd3,5'd8,5'd15,5'd0,5'd0,5'd2,5'd12,5'd20,5'd2,5'd7,5'd7,5'd16,5'd4,5'd18,5'd1,5'd1,5'd6,5'd7,5'd7,5'd2,5'd5,5'd8,5'd1,5'd15,5'd8,5'd6,5'd7,5'd5,5'd3,5'd0,5'd13,5'd17,5'd3,5'd10,5'd14,5'd8,5'd12,5'd7,5'd15,5'd15,5'd0,5'd9,5'd1,5'd15,5'd10,5'd6,5'd0,5'd1,5'd3,5'd14,5'd1,5'd1,5'd0,5'd15,5'd13,5'd14,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd4,5'd7,5'd0,5'd6,5'd13,5'd13,5'd21,5'd9,5'd1,5'd1,5'd12,5'd12,5'd6,5'd8,5'd5,5'd12,5'd6,5'd12,5'd0,5'd0,5'd0,5'd10,5'd2,5'd2,5'd18,5'd2,5'd6,5'd6,5'd9,5'd6,5'd6,5'd12,5'd3,5'd7,5'd6,5'd6,5'd14,5'd8,5'd6,5'd4,5'd2,5'd14,5'd21,5'd14,5'd2,5'd5,5'd3,5'd16,5'd1,5'd3,5'd4,5'd4,5'd0,5'd18,5'd17,5'd5,5'd13,5'd14,5'd10,5'd2,5'd3,5'd3,5'd0,5'd0,5'd7,5'd7,5'd12,5'd12,5'd12,5'd8,5'd9,5'd11,5'd0,5'd0,5'd0,5'd9,5'd6,5'd1,5'd0,5'd10,5'd14,5'd14,5'd8,5'd8,5'd0,5'd3,5'd3,5'd2,5'd1,5'd4,5'd3,5'd7,5'd6,5'd18,5'd2,5'd2,5'd0,5'd1,5'd12,5'd6,5'd13,5'd13,5'd1,5'd7,5'd17,5'd4,5'd2,5'd6,5'd14,5'd2,5'd1,5'd6,5'd0,5'd15,5'd15,5'd8,5'd7,5'd7,5'd21,5'd0,5'd0,5'd1,5'd2,5'd5,5'd20,5'd7,5'd0,5'd0,5'd6,5'd16,5'd10,5'd6,5'd6,5'd9,5'd14,5'd6,5'd4,5'd15,5'd20,5'd18,5'd18,5'd17,5'd7,5'd6,5'd0,5'd0,5'd4,5'd0,5'd5,5'd5,5'd15,5'd1,5'd4,5'd2,5'd1,5'd7,5'd12,5'd12,5'd8,5'd2,5'd1,5'd5,5'd1,5'd6,5'd0,5'd22,5'd0,5'd0,5'd15,5'd0,5'd4,5'd5,5'd5,5'd8,5'd2,5'd17,5'd4,5'd18,5'd14,5'd14,5'd6,5'd1,5'd1,5'd0,5'd0,5'd0,5'd4,5'd13,5'd10,5'd11,5'd11,5'd11,5'd10,5'd10,5'd3,5'd3,5'd18,5'd0,5'd0,5'd1,5'd0,5'd3,5'd0,5'd0,5'd12,5'd10,5'd14,5'd7,5'd6,5'd8,5'd8,5'd6,5'd7,5'd15,5'd9,5'd10,5'd7,5'd0,5'd0,5'd1,5'd1,5'd5,5'd1,5'd7,5'd17,5'd5,5'd8,5'd2,5'd1,5'd16,5'd16,5'd12,5'd9,5'd8,5'd2,5'd1,5'd6,5'd0,5'd16,5'd13,5'd14,5'd5,5'd5,5'd6,5'd0,5'd9,5'd10,5'd19,5'd8,5'd16,5'd14,5'd0,5'd0,5'd8,5'd8,5'd10,5'd0,5'd12,5'd16,5'd4,5'd4,5'd4,5'd16,5'd1,5'd18,5'd14,5'd6,5'd7,5'd7,5'd22,5'd12,5'd6,5'd6,5'd13,5'd6,5'd20,5'd6,5'd7,5'd0,5'd0,5'd8,5'd6,5'd6,5'd0,5'd6,5'd0,5'd0,5'd5,5'd6,5'd15,5'd15,5'd14,5'd8,5'd5,5'd0,5'd1,5'd4,5'd17,5'd15,5'd7,5'd6,5'd12,5'd7,5'd7,5'd1,5'd3,5'd3,5'd17,5'd10,5'd1,5'd5,5'd4,5'd4,5'd13,5'd10,5'd5,5'd1,5'd1,5'd6,5'd1,5'd3,5'd4,5'd5,5'd2,5'd1,5'd13,5'd1,5'd12,5'd6,5'd8,5'd1,5'd1,5'd6,5'd21,5'd6,5'd5,5'd6,5'd8,5'd3,5'd7,5'd18,5'd6,5'd6,5'd0,5'd5,5'd8,5'd5,5'd11,5'd0,5'd6,5'd9,5'd2,5'd8,5'd4,5'd6,5'd0,5'd14,5'd8,5'd5,5'd5,5'd18,5'd9,5'd4,5'd4}
`define RECTANGLE1_X2 {5'd15,5'd24,5'd19,5'd12,5'd21,5'd9,5'd24,5'd18,5'd22,5'd18,5'd24,5'd23,5'd24,5'd6,5'd24,5'd18,5'd24,5'd22,5'd21,5'd11,5'd21,5'd20,5'd22,5'd13,5'd21,5'd18,5'd22,5'd9,5'd19,5'd11,5'd23,5'd8,5'd24,5'd9,5'd21,5'd9,5'd21,5'd8,5'd15,5'd15,5'd24,5'd18,5'd15,5'd12,5'd18,5'd14,5'd22,5'd16,5'd22,5'd21,5'd19,5'd10,5'd16,5'd13,5'd14,5'd20,5'd18,5'd14,5'd23,5'd16,5'd16,5'd23,5'd18,5'd18,5'd23,5'd11,5'd24,5'd14,5'd23,5'd17,5'd17,5'd18,5'd20,5'd18,5'd16,5'd15,5'd24,5'd19,5'd15,5'd14,5'd14,5'd15,5'd16,5'd18,5'd23,5'd10,5'd22,5'd7,5'd15,5'd13,5'd14,5'd9,5'd21,5'd15,5'd24,5'd9,5'd21,5'd14,5'd18,5'd20,5'd24,5'd18,5'd24,5'd21,5'd24,5'd18,5'd24,5'd12,5'd15,5'd18,5'd15,5'd18,5'd24,5'd18,5'd18,5'd17,5'd15,5'd11,5'd21,5'd8,5'd18,5'd16,5'd20,5'd19,5'd23,5'd12,5'd21,5'd18,5'd23,5'd10,5'd24,5'd9,5'd24,5'd10,5'd24,5'd12,5'd22,5'd16,5'd24,5'd9,5'd21,5'd5,5'd23,5'd16,5'd22,5'd10,5'd24,5'd10,5'd24,5'd6,5'd24,5'd23,5'd24,5'd13,5'd18,5'd17,5'd24,5'd13,5'd24,5'd18,5'd14,5'd15,5'd19,5'd7,5'd24,5'd18,5'd23,5'd14,5'd18,5'd6,5'd24,5'd8,5'd24,5'd17,5'd23,5'd15,5'd15,5'd15,5'd22,5'd6,5'd23,5'd20,5'd24,5'd11,5'd20,5'd8,5'd21,5'd14,5'd15,5'd16,5'd24,5'd21,5'd18,5'd10,5'd21,5'd15,5'd18,5'd9,5'd18,5'd18,5'd12,5'd24,5'd15,5'd17,5'd10,5'd21,5'd21,5'd15,5'd15,5'd15,5'd12,5'd24,5'd9,5'd21,5'd6,5'd24,5'd9,5'd24,5'd10,5'd24,5'd20,5'd24,5'd21,5'd22,5'd16,5'd22,5'd20,5'd15,5'd8,5'd19,5'd18,5'd15,5'd14,5'd22,5'd10,5'd17,5'd13,5'd16,5'd16,5'd23,5'd7,5'd17,5'd20,5'd17,5'd14,5'd17,5'd15,5'd19,5'd15,5'd19,5'd16,5'd19,5'd6,5'd24,5'd4,5'd23,5'd18,5'd22,5'd18,5'd24,5'd8,5'd24,5'd18,5'd23,5'd9,5'd22,5'd17,5'd21,5'd16,5'd19,5'd9,5'd19,5'd15,5'd23,5'd19,5'd20,5'd12,5'd23,5'd14,5'd15,5'd14,5'd18,5'd9,5'd24,5'd8,5'd14,5'd12,5'd17,5'd17,5'd21,5'd14,5'd21,5'd5,5'd22,5'd3,5'd23,5'd20,5'd18,5'd3,5'd23,5'd14,5'd22,5'd6,5'd24,5'd21,5'd24,5'd19,5'd24,5'd12,5'd24,5'd8,5'd21,5'd18,5'd22,5'd16,5'd18,5'd21,5'd23,5'd19,5'd24,5'd17,5'd17,5'd19,5'd18,5'd16,5'd22,5'd19,5'd18,5'd13,5'd19,5'd9,5'd23,5'd15,5'd17,5'd18,5'd23,5'd11,5'd16,5'd14,5'd15,5'd17,5'd15,5'd18,5'd24,5'd18,5'd21,5'd13,5'd23,5'd16,5'd16,5'd11,5'd17,5'd13,5'd15,5'd19,5'd19,5'd21,5'd18,5'd14,5'd19,5'd15,5'd18,5'd14,5'd23,5'd14,5'd21,5'd10,5'd23,5'd10,5'd22,5'd12,5'd20,5'd11,5'd24,5'd6,5'd17,5'd6,5'd24,5'd19,5'd23,5'd14,5'd19,5'd9,5'd22,5'd16,5'd19,5'd12,5'd23,5'd9,5'd24,5'd18,5'd23,5'd10,5'd24,5'd6,5'd22,5'd11,5'd19,5'd24,5'd17,5'd14,5'd22,5'd18,5'd21,5'd6,5'd24,5'd14,5'd24,5'd8,5'd18,5'd12,5'd11,5'd19,5'd11,5'd15,5'd12,5'd24,5'd19,5'd20,5'd17,5'd16,5'd6,5'd23,5'd12,5'd21,5'd9,5'd24,5'd16,5'd24,5'd8,5'd24,5'd10,5'd15,5'd18,5'd23,5'd22,5'd24,5'd17,5'd24,5'd17,5'd24,5'd13,5'd24,5'd11,5'd24,5'd21,5'd16,5'd16,5'd24,5'd19,5'd18,5'd12,5'd24,5'd9,5'd24,5'd20,5'd22,5'd3,5'd17,5'd12,5'd16,5'd15,5'd18,5'd20,5'd23,5'd12,5'd18,5'd15,5'd22,5'd12,5'd20,5'd8,5'd18,5'd12,5'd19,5'd12,5'd18,5'd9,5'd20,5'd17,5'd14,5'd12,5'd19,5'd9,5'd19,5'd16,5'd24,5'd22,5'd23,5'd14,5'd20,5'd21,5'd22,5'd4,5'd21,5'd12,5'd17,5'd14,5'd16,5'd21,5'd22,5'd13,5'd14,5'd11,5'd22,5'd9,5'd21,5'd19,5'd24,5'd9,5'd23,5'd11,5'd17,5'd11,5'd24,5'd13,5'd16,5'd14,5'd19,5'd16,5'd16,5'd17,5'd24,5'd14,5'd18,5'd10,5'd17,5'd8,5'd19,5'd17,5'd23,5'd14,5'd21,5'd21,5'd23,5'd15,5'd17,5'd6,5'd21,5'd24,5'd22,5'd18,5'd17,5'd4,5'd24,5'd5,5'd24,5'd13,5'd18,5'd14,5'd21,5'd11,5'd19,5'd9,5'd17,5'd20,5'd17,5'd13,5'd24,5'd10,5'd20,5'd17,5'd15,5'd19,5'd17,5'd5,5'd23,5'd18,5'd24,5'd11,5'd22,5'd18,5'd23,5'd10,5'd20,5'd10,5'd16,5'd11,5'd20,5'd13,5'd15,5'd17,5'd18,5'd15,5'd20,5'd6,5'd17,5'd14,5'd24,5'd19,5'd22,5'd17,5'd21,5'd14,5'd21,5'd24,5'd17,5'd19,5'd17,5'd18,5'd15,5'd14,5'd24,5'd6,5'd24,5'd9,5'd23,5'd18,5'd24,5'd9,5'd13,5'd22,5'd10,5'd20,5'd17,5'd20,5'd10,5'd24,5'd14,5'd16,5'd8,5'd22,5'd12,5'd18,5'd14,5'd20,5'd11,5'd21,5'd24,5'd24,5'd21,5'd14,5'd15,5'd23,5'd22,5'd22,5'd13,5'd23,5'd10,5'd18,5'd15,5'd16,5'd12,5'd19,5'd22,5'd18,5'd15,5'd24,5'd15,5'd22,5'd5,5'd24,5'd8,5'd19,5'd19,5'd20,5'd16,5'd23,5'd14,5'd24,5'd11,5'd20,5'd20,5'd21,5'd8,5'd22,5'd7,5'd21,5'd17,5'd18,5'd18,5'd24,5'd8,5'd24,5'd9,5'd14,5'd17,5'd22,5'd11,5'd22,5'd10,5'd20,5'd7,5'd16,5'd13,5'd17,5'd11,5'd19,5'd11,5'd22,5'd9,5'd24,5'd18,5'd18,5'd19,5'd24,5'd13,5'd15,5'd11,5'd19,5'd14,5'd21,5'd16,5'd21,5'd16,5'd21,5'd15,5'd17,5'd5,5'd24,5'd4,5'd20,5'd17,5'd23,5'd21,5'd23,5'd19,5'd23,5'd21,5'd24,5'd12,5'd20,5'd22,5'd21,5'd20,5'd22,5'd8,5'd17,5'd24,5'd23,5'd15,5'd24,5'd6,5'd24,5'd15,5'd20,5'd20,5'd17,5'd13,5'd24,5'd9,5'd18,5'd18,5'd14,5'd7,5'd22,5'd10,5'd22,5'd15,5'd20,5'd10,5'd22,5'd12,5'd24,5'd14,5'd23,5'd19,5'd20,5'd19,5'd23,5'd20,5'd18,5'd15,5'd21,5'd18,5'd24,5'd16,5'd16,5'd16,5'd15,5'd17,5'd14,5'd22,5'd24,5'd6,5'd24,5'd11,5'd24,5'd7,5'd17,5'd15,5'd15,5'd6,5'd24,5'd8,5'd24,5'd18,5'd15,5'd9,5'd24,5'd20,5'd20,5'd23,5'd10,5'd24,5'd24,5'd20,5'd12,5'd18,5'd16,5'd18,5'd19,5'd17,5'd13,5'd17,5'd14,5'd19,5'd16,5'd17,5'd14,5'd19,5'd14,5'd23,5'd4,5'd24,5'd19,5'd20,5'd18,5'd18,5'd12,5'd23,5'd13,5'd15,5'd14,5'd16,5'd8,5'd21,5'd9,5'd24,5'd8,5'd24,5'd19,5'd24,5'd16,5'd22,5'd6,5'd15,5'd4,5'd15,5'd11,5'd15,5'd18,5'd15,5'd4,5'd24,5'd14,5'd21,5'd18,5'd24,5'd13,5'd24,5'd6,5'd24,5'd9,5'd21,5'd10,5'd24,5'd20,5'd24,5'd17,5'd24,5'd9,5'd21,5'd10,5'd20,5'd9,5'd23,5'd4,5'd17,5'd15,5'd24,5'd11,5'd17,5'd21,5'd21,5'd9,5'd17,5'd8,5'd22,5'd13,5'd15,5'd21,5'd15,5'd20,5'd24,5'd9,5'd21,5'd23,5'd19,5'd24,5'd18,5'd17,5'd21,5'd16,5'd17,5'd9,5'd19,5'd24,5'd24,5'd16,5'd14,5'd12,5'd19,5'd16,5'd17,5'd18,5'd18,5'd24,5'd21,5'd19,5'd17,5'd10,5'd18,5'd13,5'd14,5'd16,5'd18,5'd22,5'd24,5'd20,5'd24,5'd6,5'd24,5'd12,5'd24,5'd11,5'd23,5'd13,5'd17,5'd9,5'd21,5'd10,5'd24,5'd13,5'd23,5'd9,5'd21,5'd9,5'd20,5'd21,5'd19,5'd14,5'd24,5'd20,5'd23,5'd13,5'd22,5'd8,5'd24,5'd7,5'd18,5'd16,5'd17,5'd19,5'd23,5'd15,5'd20,5'd15,5'd17,5'd13,5'd17,5'd9,5'd19,5'd21,5'd20,5'd22,5'd18,5'd11,5'd22,5'd10,5'd21,5'd4,5'd17,5'd6,5'd24,5'd11,5'd19,5'd18,5'd23,5'd22,5'd20,5'd20,5'd19,5'd11,5'd20,5'd18,5'd19,5'd21,5'd15,5'd21,5'd17,5'd12,5'd20,5'd13,5'd20,5'd21,5'd24,5'd21,5'd23,5'd18,5'd17,5'd19,5'd20,5'd19,5'd20,5'd10,5'd24,5'd21,5'd24,5'd5,5'd23,5'd14,5'd24,5'd18,5'd18,5'd13,5'd17,5'd14,5'd19,5'd20,5'd19,5'd9,5'd18,5'd18,5'd20,5'd16,5'd24,5'd16,5'd24,5'd10,5'd23,5'd6,5'd20,5'd12,5'd24,5'd8,5'd21,5'd17,5'd20,5'd13,5'd14,5'd8,5'd24,5'd18,5'd24,5'd18,5'd18,5'd12,5'd16,5'd18,5'd16,5'd20,5'd19,5'd12,5'd24,5'd17,5'd20,5'd6,5'd24,5'd9,5'd24,5'd8,5'd22,5'd12,5'd24,5'd9,5'd21,5'd20,5'd20,5'd12,5'd21,5'd10,5'd20,5'd13,5'd20,5'd17,5'd21,5'd20,5'd24,5'd6,5'd17,5'd13,5'd24,5'd19,5'd24,5'd21,5'd24,5'd11,5'd23,5'd10,5'd24,5'd14,5'd22,5'd15,5'd17,5'd10,5'd23,5'd24,5'd23,5'd24,5'd21,5'd21,5'd21,5'd18,5'd19,5'd12,5'd18,5'd15,5'd23,5'd19,5'd24,5'd13,5'd14,5'd11,5'd19,5'd21,5'd19,5'd14,5'd17,5'd18,5'd15,5'd9,5'd24,5'd13,5'd16,5'd12,5'd20,5'd17,5'd14,5'd12,5'd24,5'd14,5'd15,5'd21,5'd24,5'd9,5'd24,5'd24,5'd23,5'd9,5'd24,5'd24,5'd24,5'd21,5'd19,5'd18,5'd21,5'd14,5'd20,5'd20,5'd21,5'd10,5'd24,5'd15,5'd20,5'd19,5'd20,5'd14,5'd20,5'd11,5'd19,5'd18,5'd17,5'd12,5'd15,5'd6,5'd20,5'd7,5'd23,5'd10,5'd20,5'd16,5'd20,5'd15,5'd15,5'd19,5'd22,5'd6,5'd21,5'd13,5'd21,5'd7,5'd18,5'd20,5'd14,5'd21,5'd17,5'd22,5'd16,5'd15,5'd11,5'd14,5'd13,5'd23,5'd10,5'd24,5'd22,5'd24,5'd14,5'd24,5'd11,5'd24,5'd18,5'd17,5'd10,5'd24,5'd23,5'd23,5'd10,5'd19,5'd15,5'd16,5'd15,5'd24,5'd15,5'd15,5'd6,5'd22,5'd17,5'd19,5'd12,5'd23,5'd14,5'd16,5'd11,5'd24,5'd21,5'd23,5'd12,5'd24,5'd12,5'd15,5'd22,5'd23,5'd10,5'd24,5'd13,5'd19,5'd16,5'd18,5'd16,5'd23,5'd17,5'd23,5'd15,5'd24,5'd20,5'd15,5'd14,5'd23,5'd10,5'd22,5'd9,5'd15,5'd7,5'd23,5'd7,5'd19,5'd11,5'd23,5'd11,5'd24,5'd17,5'd23,5'd15,5'd22,5'd13,5'd21,5'd15,5'd24,5'd6,5'd24,5'd21,5'd24,5'd12,5'd18,5'd17,5'd19,5'd13,5'd21,5'd19,5'd21,5'd10,5'd16,5'd12,5'd22,5'd14,5'd17,5'd13,5'd24,5'd15,5'd21,5'd22,5'd20,5'd13,5'd20,5'd13,5'd14,5'd20,5'd17,5'd17,5'd24,5'd8,5'd19,5'd24,5'd24,5'd9,5'd21,5'd9,5'd24,5'd6,5'd23,5'd19,5'd24,5'd22,5'd16,5'd12,5'd24,5'd20,5'd23,5'd19,5'd17,5'd12,5'd18,5'd19,5'd18,5'd19,5'd18,5'd13,5'd16,5'd12,5'd16,5'd14,5'd18,5'd22,5'd21,5'd19,5'd19,5'd19,5'd21,5'd4,5'd24,5'd16,5'd24,5'd9,5'd23,5'd22,5'd21,5'd6,5'd15,5'd9,5'd23,5'd17,5'd13,5'd19,5'd18,5'd18,5'd12,5'd16,5'd21,5'd22,5'd12,5'd21,5'd20,5'd22,5'd7,5'd24,5'd15,5'd17,5'd14,5'd20,5'd22,5'd24,5'd9,5'd17,5'd20,5'd20,5'd24,5'd17,5'd18,5'd21,5'd17,5'd21,5'd14,5'd16,5'd9,5'd24,5'd13,5'd16,5'd16,5'd16,5'd12,5'd24,5'd14,5'd23,5'd19,5'd24,5'd12,5'd24,5'd13,5'd18,5'd24,5'd18,5'd12,5'd24,5'd11,5'd15,5'd13,5'd19,5'd9,5'd23,5'd16,5'd23,5'd20,5'd21,5'd18,5'd18,5'd7,5'd21,5'd10,5'd18,5'd14,5'd16,5'd13,5'd19,5'd16,5'd22,5'd10,5'd24,5'd16,5'd18,5'd18,5'd24,5'd22,5'd15,5'd12,5'd24,5'd10,5'd24,5'd23,5'd21,5'd11,5'd20,5'd7,5'd23,5'd12,5'd15,5'd18,5'd24,5'd9,5'd14,5'd18,5'd17,5'd13,5'd22,5'd15,5'd17,5'd12,5'd16,5'd14,5'd24,5'd14,5'd23,5'd9,5'd23,5'd18,5'd21,5'd9,5'd24,5'd24,5'd21,5'd10,5'd20,5'd15,5'd21,5'd6,5'd24,5'd23,5'd21,5'd10,5'd23,5'd15,5'd20,5'd14,5'd20,5'd18,5'd16,5'd14,5'd17,5'd9,5'd17,5'd13,5'd24,5'd6,5'd22,5'd6,5'd22,5'd11,5'd18,5'd17,5'd15,5'd18,5'd22,5'd9,5'd20,5'd14,5'd17,5'd24,5'd2,5'd24,5'd12,5'd20,5'd10,5'd18,5'd12,5'd17,5'd14,5'd23,5'd15,5'd17,5'd14,5'd16,5'd15,5'd19,5'd11,5'd21,5'd6,5'd24,5'd7,5'd23,5'd5,5'd24,5'd9,5'd24,5'd10,5'd18,5'd16,5'd16,5'd18,5'd18,5'd9,5'd23,5'd13,5'd15,5'd18,5'd14,5'd14,5'd23,5'd17,5'd18,5'd11,5'd19,5'd14,5'd17,5'd4,5'd18,5'd18,5'd19,5'd13,5'd22,5'd11,5'd24,5'd21,5'd22,5'd15,5'd24,5'd20,5'd19,5'd13,5'd21,5'd6,5'd24,5'd2,5'd24,5'd9,5'd17,5'd24,5'd23,5'd7,5'd24,5'd8,5'd21,5'd10,5'd20,5'd7,5'd16,5'd8,5'd23,5'd18,5'd22,5'd9,5'd15,5'd14,5'd20,5'd9,5'd22,5'd11,5'd22,5'd15,5'd20,5'd23,5'd20,5'd19,5'd24,5'd10,5'd23,5'd20,5'd20,5'd22,5'd24,5'd19,5'd18,5'd15,5'd17,5'd15,5'd17,5'd17,5'd14,5'd14,5'd17,5'd11,5'd17,5'd18,5'd17,5'd9,5'd23,5'd23,5'd24,5'd18,5'd24,5'd9,5'd21,5'd13,5'd16,5'd6,5'd24,5'd6,5'd23,5'd22,5'd24,5'd19,5'd22,5'd20,5'd17,5'd6,5'd24,5'd18,5'd24,5'd12,5'd14,5'd20,5'd21,5'd15,5'd17,5'd11,5'd19,5'd5,5'd17,5'd20,5'd24,5'd14,5'd15,5'd9,5'd21,5'd14,5'd24,5'd19,5'd14,5'd14,5'd8,5'd24,5'd8,5'd24,5'd15,5'd18,5'd17,5'd20,5'd16,5'd22,5'd12,5'd18,5'd21,5'd18,5'd14,5'd17,5'd5,5'd18,5'd9,5'd24,5'd9,5'd24,5'd19,5'd24,5'd9,5'd21,5'd8,5'd16,5'd16,5'd20,5'd13,5'd22,5'd21,5'd23,5'd16,5'd24,5'd6,5'd20,5'd17,5'd17,5'd14,5'd23,5'd17,5'd19,5'd21,5'd24,5'd12,5'd18,5'd6,5'd24,5'd6,5'd24,5'd11,5'd19,5'd15,5'd18,5'd19,5'd23,5'd11,5'd23,5'd6,5'd24,5'd19,5'd19,5'd17,5'd22,5'd24,5'd24,5'd7,5'd24,5'd12,5'd24,5'd9,5'd17,5'd15,5'd15,5'd21,5'd24,5'd21,5'd18,5'd18,5'd23,5'd23,5'd24,5'd10,5'd20,5'd19,5'd20,5'd20,5'd23,5'd19,5'd23,5'd11,5'd22,5'd9,5'd24,5'd13,5'd24,5'd19,5'd15,5'd15,5'd24,5'd21,5'd17,5'd18,5'd24,5'd19,5'd24,5'd13,5'd16,5'd14,5'd17,5'd19,5'd23,5'd13,5'd17,5'd4,5'd24,5'd7,5'd24,5'd10,5'd20,5'd10,5'd18,5'd10,5'd20,5'd9,5'd23,5'd22,5'd22,5'd12,5'd24,5'd15,5'd20,5'd9,5'd23,5'd4,5'd17,5'd21,5'd20,5'd19,5'd22,5'd15,5'd23,5'd16,5'd24,5'd9,5'd24,5'd12,5'd22,5'd15,5'd19,5'd9,5'd19,5'd12,5'd21,5'd9,5'd16,5'd14,5'd17,5'd9,5'd17,5'd15,5'd23,5'd15,5'd21,5'd10,5'd17,5'd24,5'd22,5'd12,5'd17,5'd22,5'd15,5'd18,5'd20,5'd15,5'd19,5'd24,5'd21,5'd19,5'd21,5'd21,5'd21,5'd6,5'd23,5'd15,5'd15,5'd14,5'd19,5'd13,5'd19,5'd14,5'd23,5'd24,5'd16,5'd20,5'd24,5'd9,5'd21,5'd20,5'd22,5'd15,5'd14,5'd16,5'd14,5'd9,5'd14,5'd18,5'd18,5'd7,5'd18,5'd9,5'd21,5'd12,5'd16,5'd13,5'd19,5'd20,5'd23,5'd18,5'd18,5'd23,5'd23,5'd9,5'd21,5'd7,5'd23,5'd21,5'd23,5'd7,5'd16,5'd21,5'd24,5'd17,5'd18,5'd11,5'd19,5'd16,5'd14,5'd15,5'd22,5'd21,5'd24,5'd11,5'd19,5'd9,5'd24,5'd4,5'd24,5'd9,5'd24,5'd12,5'd18,5'd14,5'd24,5'd24,5'd19,5'd24,5'd23,5'd10,5'd16,5'd8,5'd24,5'd24,5'd24,5'd15,5'd15,5'd22,5'd24,5'd17,5'd7,5'd22,5'd9,5'd15,5'd17,5'd17,5'd14,5'd18,5'd15,5'd18,5'd13,5'd22,5'd22,5'd19,5'd17,5'd18,5'd12,5'd16,5'd15,5'd24,5'd6,5'd20,5'd15,5'd19,5'd15,5'd23,5'd19,5'd22,5'd12,5'd24,5'd8,5'd18,5'd15,5'd24,5'd18,5'd17,5'd7,5'd21,5'd11,5'd17,5'd22,5'd20,5'd13,5'd17,5'd15,5'd16,5'd19,5'd24,5'd13,5'd14,5'd17,5'd18,5'd8,5'd21,5'd10,5'd24,5'd16,5'd24,5'd13,5'd19,5'd19,5'd16,5'd10,5'd16,5'd16,5'd18,5'd17,5'd23,5'd18,5'd22,5'd11,5'd23,5'd5,5'd23,5'd11,5'd24,5'd11,5'd21,5'd19,5'd24,5'd11,5'd24,5'd21,5'd24,5'd18,5'd24,5'd13,5'd20,5'd11,5'd23,5'd12,5'd19,5'd23,5'd18,5'd15,5'd22,5'd13,5'd15,5'd10,5'd20,5'd18,5'd24,5'd8,5'd24,5'd8,5'd16,5'd18,5'd16,5'd13,5'd21,5'd18,5'd17,5'd10,5'd22,5'd14,5'd24,5'd11,5'd23,5'd19,5'd23,5'd9,5'd24,5'd4,5'd24,5'd6,5'd18,5'd18,5'd17,5'd21,5'd16,5'd20,5'd15,5'd17,5'd23,5'd9,5'd11,5'd20,5'd17,5'd20,5'd15,5'd15,5'd11,5'd17,5'd21,5'd18,5'd7,5'd18,5'd13,5'd21,5'd10,5'd21,5'd24,5'd20,5'd11,5'd19,5'd12,5'd22,5'd16,5'd19,5'd20,5'd21,5'd15,5'd20,5'd13,5'd21,5'd14,5'd16,5'd15,5'd17,5'd22,5'd24,5'd17,5'd23,5'd17,5'd18,5'd22,5'd21,5'd12,5'd18,5'd13,5'd16,5'd14,5'd24,5'd9,5'd24,5'd19,5'd24,5'd20,5'd24,5'd11,5'd19,5'd9,5'd24,5'd18,5'd21,5'd23,5'd24,5'd17,5'd24,5'd9,5'd22,5'd11,5'd23,5'd10,5'd24,5'd13,5'd22,5'd8,5'd24,5'd20,5'd24,5'd12,5'd15,5'd13,5'd24,5'd8,5'd24,5'd5,5'd24,5'd19,5'd24,5'd19,5'd16,5'd16,5'd15,5'd20,5'd22,5'd13,5'd16,5'd12,5'd16,5'd4,5'd21,5'd14,5'd21,5'd15,5'd20,5'd20,5'd14,5'd8,5'd22,5'd8,5'd24,5'd7,5'd24,5'd4,5'd22,5'd20,5'd24,5'd13,5'd23,5'd16,5'd23,5'd23,5'd17,5'd12,5'd19,5'd22,5'd19,5'd9,5'd18,5'd20,5'd13,5'd24,5'd8,5'd19,5'd17,5'd21,5'd20,5'd21,5'd12,5'd14,5'd24,5'd19,5'd10,5'd24,5'd6,5'd23,5'd4,5'd23,5'd22,5'd24,5'd21,5'd24,5'd21,5'd18,5'd17,5'd19,5'd10,5'd21,5'd18,5'd22,5'd10,5'd22,5'd12,5'd22,5'd14,5'd24,5'd15,5'd21,5'd22,5'd18,5'd13,5'd19,5'd15,5'd18,5'd10,5'd20,5'd11,5'd19,5'd16,5'd23,5'd10,5'd21,5'd5,5'd21,5'd16,5'd21,5'd19,5'd23,5'd6,5'd17,5'd15,5'd17,5'd8,5'd21,5'd13,5'd17,5'd14,5'd17,5'd11,5'd24,5'd9,5'd18,5'd21,5'd24,5'd10,5'd23,5'd19,5'd21,5'd24,5'd21,5'd10,5'd22,5'd19,5'd17,5'd11,5'd16,5'd18,5'd24,5'd12,5'd20,5'd8,5'd23,5'd20,5'd15,5'd10,5'd20,5'd16,5'd18,5'd11,5'd19,5'd14,5'd19,5'd24,5'd19,5'd6,5'd23,5'd21,5'd24,5'd6,5'd15,5'd19,5'd18,5'd18,5'd24,5'd17,5'd12,5'd22,5'd3,5'd24,5'd11,5'd21,5'd6,5'd14,5'd16,5'd19,5'd9,5'd23,5'd12,5'd18,5'd15,5'd18,5'd9,5'd24,5'd14,5'd24,5'd13,5'd19,5'd9,5'd17,5'd9,5'd21,5'd9,5'd24,5'd18,5'd22,5'd5,5'd23,5'd7,5'd23,5'd21,5'd18,5'd10,5'd17,5'd9,5'd24,5'd6,5'd21,5'd11,5'd17,5'd24,5'd21,5'd8,5'd24,5'd19,5'd24,5'd12,5'd17,5'd14,5'd24,5'd21,5'd21,5'd18,5'd16,5'd18,5'd18,5'd13,5'd17,5'd24,5'd24,5'd14,5'd24,5'd15,5'd17,5'd12,5'd24,5'd17,5'd24,5'd10,5'd24,5'd12,5'd20,5'd6,5'd24,5'd15,5'd24,5'd20,5'd23,5'd9,5'd24,5'd10,5'd23,5'd15,5'd23,5'd10,5'd20,5'd16,5'd14,5'd6,5'd24,5'd21,5'd24,5'd24,5'd18,5'd17,5'd13,5'd14,5'd10,5'd23,5'd10,5'd22,5'd14,5'd19,5'd15,5'd20,5'd12,5'd18,5'd14,5'd24,5'd13,5'd22,5'd6,5'd24,5'd8,5'd18,5'd15,5'd24,5'd8,5'd22,5'd11,5'd19,5'd3,5'd18,5'd13,5'd19,5'd21,5'd24,5'd19,5'd21,5'd18,5'd24,5'd10,5'd24,5'd24,5'd20,5'd17,5'd24,5'd21,5'd24,5'd19,5'd23,5'd11,5'd18,5'd19,5'd24,5'd22,5'd20,5'd19,5'd21,5'd19,5'd24,5'd12,5'd18,5'd15,5'd21,5'd10,5'd18,5'd7,5'd23,5'd19,5'd18,5'd6,5'd24,5'd16,5'd24,5'd17,5'd24,5'd20,5'd23,5'd11,5'd17,5'd16,5'd18,5'd22,5'd18,5'd16,5'd18,5'd10,5'd24,5'd15,5'd22,5'd6,5'd15,5'd10,5'd19,5'd24,5'd14,5'd18,5'd21,5'd15,5'd15,5'd16,5'd18,5'd19,5'd20,5'd23,5'd19,5'd24,5'd24,5'd19,5'd24,5'd24,5'd15,5'd23,5'd9,5'd19,5'd12,5'd23,5'd21,5'd24,5'd20,5'd16,5'd18,5'd16,5'd16,5'd22,5'd7,5'd23,5'd16,5'd24,5'd21,5'd23,5'd9,5'd24,5'd9,5'd21,5'd9,5'd21,5'd6,5'd18,5'd19,5'd20,5'd23,5'd24,5'd19,5'd24,5'd11,5'd17,5'd14,5'd24,5'd11,5'd17,5'd8,5'd24,5'd16,5'd24,5'd14,5'd16,5'd18,5'd23,5'd6,5'd24,5'd18,5'd24,5'd6,5'd24,5'd13,5'd22,5'd14,5'd22,5'd22,5'd21,5'd10,5'd16,5'd12,5'd19,5'd18,5'd18,5'd24,5'd16,5'd21,5'd15,5'd23,5'd18,5'd21,5'd21,5'd12,5'd21,5'd12,5'd15,5'd15,5'd24,5'd20,5'd17,5'd12,5'd15,5'd11,5'd24,5'd12,5'd18,5'd13,5'd17,5'd14,5'd18,5'd6,5'd24,5'd16,5'd15,5'd17,5'd24,5'd8,5'd20,5'd8,5'd17,5'd14,5'd17,5'd24,5'd21,5'd9,5'd17,5'd9,5'd24,5'd9,5'd17,5'd6,5'd17,5'd6,5'd17,5'd16,5'd19,5'd13,5'd18,5'd12,5'd18,5'd16,5'd17,5'd14,5'd17,5'd12,5'd18,5'd9,5'd20,5'd24,5'd15,5'd7,5'd17,5'd15,5'd23,5'd15,5'd22,5'd19,5'd24,5'd21,5'd23,5'd15,5'd19,5'd20,5'd24,5'd19,5'd23,5'd24,5'd15,5'd22,5'd20,5'd11,5'd15,5'd18,5'd21,5'd18,5'd21,5'd13,5'd17,5'd15,5'd17,5'd20,5'd24,5'd15,5'd21,5'd16,5'd22,5'd14,5'd17,5'd11,5'd17,5'd24,5'd17,5'd17,5'd24,5'd21,5'd24,5'd18,5'd15,5'd16,5'd15,5'd22,5'd24,5'd9,5'd23,5'd20,5'd20,5'd6,5'd24,5'd4,5'd24,5'd20,5'd24,5'd14,5'd23,5'd10,5'd16,5'd13,5'd20,5'd12,5'd18,5'd17,5'd21,5'd22,5'd15,5'd20,5'd10,5'd16,5'd10,5'd16,5'd22,5'd24,5'd24,5'd18,5'd12,5'd18,5'd13,5'd23,5'd18,5'd19,5'd12,5'd18,5'd14,5'd19,5'd21,5'd19,5'd20,5'd19,5'd17,5'd20,5'd19,5'd24,5'd10,5'd18,5'd9,5'd24,5'd13,5'd17,5'd19,5'd15,5'd21,5'd24,5'd6,5'd24,5'd6,5'd24,5'd13,5'd21,5'd22,5'd15,5'd16,5'd18,5'd24,5'd24,5'd12,5'd24,5'd15,5'd19,5'd23,5'd22,5'd10,5'd18,5'd6,5'd21,5'd14,5'd22,5'd16,5'd19,5'd19,5'd21,5'd20,5'd22,5'd15,5'd16,5'd9,5'd17,5'd12,5'd18,5'd12,5'd23,5'd11,5'd18,5'd8,5'd22,5'd4,5'd24,5'd8,5'd24,5'd23,5'd24,5'd10,5'd17,5'd14,5'd14,5'd19,5'd15,5'd13,5'd15,5'd19,5'd15,5'd24,5'd17,5'd20,5'd24,5'd18,5'd21,5'd14,5'd16,5'd13,5'd15,5'd15,5'd18,5'd19,5'd19,5'd10,5'd23,5'd10,5'd19,5'd21,5'd21,5'd4,5'd20,5'd19,5'd24,5'd14,5'd18,5'd19,5'd17,5'd9,5'd24,5'd5,5'd23,5'd14,5'd22,5'd24,5'd18,5'd18,5'd6,5'd21,5'd19,5'd19,5'd12,5'd16,5'd19,5'd16,5'd6,5'd24,5'd22,5'd24,5'd6,5'd22,5'd12,5'd23,5'd19,5'd24,5'd7,5'd24,5'd18,5'd21,5'd9,5'd15,5'd14,5'd20,5'd24,5'd19,5'd17,5'd15,5'd24,5'd24,5'd6,5'd16,5'd13,5'd22,5'd19,5'd19,5'd15,5'd24,5'd20,5'd18,5'd18,5'd11,5'd15,5'd17,5'd18,5'd7,5'd17,5'd21,5'd18,5'd18}
`define RECTANGLE1_Y2 {5'd23,5'd21,5'd22,5'd23,5'd23,5'd23,5'd23,5'd16,5'd18,5'd20,5'd23,5'd16,5'd23,5'd24,5'd24,5'd23,5'd20,5'd24,5'd22,5'd23,5'd23,5'd19,5'd15,5'd22,5'd21,5'd23,5'd23,5'd23,5'd23,5'd21,5'd21,5'd20,5'd20,5'd20,5'd24,5'd15,5'd15,5'd14,5'd24,5'd17,5'd11,5'd13,5'd13,5'd9,5'd9,5'd18,5'd15,5'd6,5'd24,5'd13,5'd8,5'd23,5'd23,5'd11,5'd24,5'd12,5'd11,5'd13,5'd7,5'd21,5'd20,5'd24,5'd23,5'd19,5'd20,5'd23,5'd10,5'd14,5'd14,5'd13,5'd11,5'd13,5'd13,5'd11,5'd19,5'd18,5'd6,5'd9,5'd10,5'd9,5'd24,5'd11,5'd9,5'd3,5'd13,5'd14,5'd15,5'd19,5'd22,5'd20,5'd20,5'd17,5'd15,5'd14,5'd14,5'd24,5'd24,5'd21,5'd16,5'd16,5'd23,5'd20,5'd20,5'd10,5'd8,5'd8,5'd17,5'd24,5'd24,5'd17,5'd24,5'd18,5'd18,5'd14,5'd15,5'd17,5'd24,5'd24,5'd24,5'd23,5'd23,5'd18,5'd24,5'd4,5'd15,5'd12,5'd17,5'd21,5'd20,5'd20,5'd20,5'd20,5'd20,5'd12,5'd12,5'd24,5'd24,5'd22,5'd24,5'd23,5'd24,5'd24,5'd24,5'd22,5'd19,5'd6,5'd10,5'd11,5'd9,5'd14,5'd14,5'd24,5'd11,5'd21,5'd10,5'd12,5'd11,5'd16,5'd19,5'd19,5'd24,5'd17,5'd17,5'd14,5'd14,5'd6,5'd5,5'd14,5'd14,5'd13,5'd13,5'd18,5'd3,5'd12,5'd13,5'd21,5'd23,5'd24,5'd4,5'd16,5'd12,5'd23,5'd21,5'd20,5'd12,5'd24,5'd24,5'd15,5'd15,5'd8,5'd5,5'd12,5'd21,5'd19,5'd24,5'd18,5'd20,5'd6,5'd11,5'd13,5'd13,5'd9,5'd8,5'd20,5'd19,5'd13,5'd10,5'd13,5'd16,5'd15,5'd22,5'd22,5'd22,5'd22,5'd14,5'd14,5'd24,5'd24,5'd20,5'd13,5'd10,5'd10,5'd10,5'd12,5'd12,5'd11,5'd20,5'd23,5'd24,5'd24,5'd13,5'd13,5'd17,5'd11,5'd22,5'd22,5'd10,5'd21,5'd15,5'd23,5'd14,5'd18,5'd23,5'd8,5'd23,5'd8,5'd15,5'd11,5'd9,5'd11,5'd11,5'd24,5'd24,5'd24,5'd22,5'd20,5'd5,5'd10,5'd10,5'd19,5'd16,5'd16,5'd16,5'd16,5'd14,5'd12,5'd22,5'd22,5'd13,5'd11,5'd16,5'd20,5'd19,5'd24,5'd21,5'd9,5'd23,5'd12,5'd24,5'd13,5'd18,5'd16,5'd16,5'd16,5'd24,5'd24,5'd24,5'd21,5'd20,5'd20,5'd13,5'd13,5'd19,5'd19,5'd23,5'd17,5'd12,5'd14,5'd24,5'd23,5'd21,5'd11,5'd14,5'd14,5'd15,5'd18,5'd13,5'd24,5'd15,5'd24,5'd14,5'd20,5'd20,5'd13,5'd19,5'd19,5'd20,5'd12,5'd9,5'd23,5'd20,5'd12,5'd17,5'd21,5'd13,5'd14,5'd14,5'd6,5'd10,5'd10,5'd24,5'd24,5'd24,5'd15,5'd16,5'd7,5'd9,5'd16,5'd9,5'd13,5'd15,5'd9,5'd18,5'd3,5'd17,5'd23,5'd21,5'd13,5'd21,5'd21,5'd24,5'd24,5'd16,5'd13,5'd9,5'd7,5'd16,5'd17,5'd15,5'd12,5'd7,5'd7,5'd9,5'd3,5'd19,5'd18,5'd19,5'd19,5'd24,5'd24,5'd15,5'd9,5'd21,5'd15,5'd14,5'd21,5'd21,5'd21,5'd23,5'd23,5'd15,5'd10,5'd20,5'd23,5'd21,5'd20,5'd11,5'd19,5'd24,5'd19,5'd19,5'd19,5'd22,5'd22,5'd11,5'd13,5'd17,5'd17,5'd4,5'd21,5'd18,5'd11,5'd6,5'd24,5'd6,5'd8,5'd23,5'd16,5'd15,5'd11,5'd9,5'd20,5'd10,5'd15,5'd16,5'd10,5'd13,5'd24,5'd9,5'd12,5'd12,5'd13,5'd23,5'd17,5'd17,5'd24,5'd24,5'd16,5'd24,5'd12,5'd12,5'd16,5'd9,5'd19,5'd7,5'd23,5'd12,5'd11,5'd24,5'd10,5'd24,5'd22,5'd24,5'd18,5'd24,5'd17,5'd24,5'd15,5'd9,5'd15,5'd11,5'd18,5'd24,5'd21,5'd21,5'd17,5'd17,5'd21,5'd24,5'd19,5'd19,5'd12,5'd18,5'd9,5'd18,5'd22,5'd11,5'd24,5'd20,5'd24,5'd24,5'd23,5'd18,5'd15,5'd17,5'd18,5'd18,5'd15,5'd15,5'd14,5'd22,5'd10,5'd22,5'd23,5'd23,5'd20,5'd23,5'd16,5'd17,5'd21,5'd10,5'd23,5'd23,5'd24,5'd14,5'd20,5'd17,5'd17,5'd17,5'd14,5'd6,5'd10,5'd17,5'd6,5'd6,5'd11,5'd12,5'd10,5'd18,5'd6,5'd6,5'd19,5'd19,5'd21,5'd17,5'd24,5'd17,5'd24,5'd6,5'd6,5'd19,5'd10,5'd6,5'd17,5'd9,5'd15,5'd14,5'd16,5'd16,5'd21,5'd21,5'd16,5'd24,5'd19,5'd21,5'd14,5'd19,5'd22,5'd22,5'd4,5'd14,5'd23,5'd11,5'd24,5'd24,5'd23,5'd23,5'd24,5'd11,5'd12,5'd24,5'd19,5'd19,5'd24,5'd24,5'd7,5'd14,5'd15,5'd24,5'd15,5'd15,5'd23,5'd24,5'd24,5'd24,5'd24,5'd24,5'd19,5'd19,5'd24,5'd24,5'd24,5'd21,5'd21,5'd21,5'd24,5'd17,5'd23,5'd15,5'd18,5'd22,5'd23,5'd23,5'd24,5'd24,5'd12,5'd12,5'd20,5'd24,5'd2,5'd17,5'd21,5'd19,5'd14,5'd19,5'd24,5'd8,5'd10,5'd18,5'd24,5'd15,5'd22,5'd18,5'd22,5'd22,5'd12,5'd13,5'd12,5'd4,5'd19,5'd20,5'd21,5'd19,5'd5,5'd6,5'd23,5'd24,5'd24,5'd24,5'd24,5'd24,5'd24,5'd22,5'd22,5'd15,5'd24,5'd22,5'd24,5'd21,5'd12,5'd15,5'd9,5'd12,5'd18,5'd16,5'd18,5'd9,5'd18,5'd21,5'd17,5'd20,5'd20,5'd20,5'd20,5'd10,5'd14,5'd22,5'd13,5'd23,5'd18,5'd17,5'd14,5'd23,5'd19,5'd19,5'd22,5'd20,5'd18,5'd21,5'd24,5'd20,5'd24,5'd16,5'd18,5'd9,5'd9,5'd9,5'd20,5'd14,5'd23,5'd10,5'd13,5'd18,5'd18,5'd16,5'd9,5'd10,5'd10,5'd15,5'd10,5'd9,5'd9,5'd24,5'd24,5'd15,5'd15,5'd17,5'd17,5'd21,5'd21,5'd22,5'd21,5'd21,5'd17,5'd12,5'd22,5'd23,5'd20,5'd5,5'd17,5'd23,5'd13,5'd13,5'd13,5'd15,5'd13,5'd18,5'd18,5'd23,5'd22,5'd16,5'd22,5'd21,5'd22,5'd10,5'd22,5'd24,5'd24,5'd18,5'd18,5'd15,5'd10,5'd24,5'd10,5'd19,5'd19,5'd10,5'd15,5'd4,5'd9,5'd10,5'd10,5'd15,5'd13,5'd19,5'd9,5'd8,5'd12,5'd22,5'd20,5'd19,5'd18,5'd12,5'd23,5'd12,5'd24,5'd24,5'd24,5'd24,5'd11,5'd16,5'd3,5'd24,5'd20,5'd24,5'd16,5'd7,5'd4,5'd4,5'd22,5'd6,5'd17,5'd15,5'd23,5'd10,5'd10,5'd21,5'd15,5'd6,5'd9,5'd20,5'd15,5'd5,5'd18,5'd13,5'd13,5'd10,5'd14,5'd16,5'd17,5'd22,5'd24,5'd21,5'd21,5'd21,5'd24,5'd20,5'd15,5'd21,5'd6,5'd9,5'd9,5'd9,5'd18,5'd18,5'd10,5'd14,5'd16,5'd16,5'd23,5'd16,5'd22,5'd14,5'd22,5'd22,5'd20,5'd15,5'd13,5'd24,5'd24,5'd14,5'd19,5'd13,5'd21,5'd18,5'd10,5'd17,5'd8,5'd22,5'd13,5'd15,5'd21,5'd21,5'd24,5'd14,5'd20,5'd15,5'd20,5'd4,5'd7,5'd7,5'd8,5'd7,5'd20,5'd11,5'd10,5'd21,5'd19,5'd21,5'd24,5'd21,5'd24,5'd21,5'd23,5'd23,5'd16,5'd11,5'd15,5'd15,5'd19,5'd21,5'd24,5'd20,5'd24,5'd24,5'd23,5'd20,5'd20,5'd8,5'd5,5'd5,5'd16,5'd16,5'd21,5'd21,5'd12,5'd12,5'd18,5'd11,5'd17,5'd11,5'd23,5'd23,5'd16,5'd16,5'd20,5'd23,5'd9,5'd9,5'd18,5'd23,5'd22,5'd22,5'd18,5'd11,5'd11,5'd18,5'd17,5'd8,5'd9,5'd7,5'd16,5'd19,5'd24,5'd22,5'd24,5'd8,5'd20,5'd24,5'd13,5'd21,5'd15,5'd8,5'd13,5'd23,5'd5,5'd7,5'd4,5'd18,5'd12,5'd13,5'd17,5'd17,5'd15,5'd14,5'd12,5'd18,5'd24,5'd6,5'd23,5'd15,5'd10,5'd6,5'd24,5'd22,5'd23,5'd23,5'd24,5'd13,5'd22,5'd22,5'd21,5'd21,5'd19,5'd15,5'd15,5'd15,5'd24,5'd24,5'd21,5'd16,5'd18,5'd3,5'd9,5'd9,5'd11,5'd8,5'd8,5'd16,5'd13,5'd18,5'd24,5'd21,5'd20,5'd13,5'd24,5'd7,5'd11,5'd14,5'd9,5'd9,5'd24,5'd24,5'd19,5'd24,5'd23,5'd12,5'd20,5'd12,5'd17,5'd18,5'd10,5'd21,5'd22,5'd22,5'd9,5'd9,5'd20,5'd12,5'd23,5'd6,5'd16,5'd9,5'd20,5'd16,5'd10,5'd13,5'd4,5'd16,5'd17,5'd20,5'd17,5'd17,5'd19,5'd19,5'd20,5'd11,5'd16,5'd16,5'd12,5'd23,5'd19,5'd19,5'd24,5'd22,5'd18,5'd10,5'd11,5'd12,5'd21,5'd23,5'd19,5'd19,5'd4,5'd10,5'd9,5'd9,5'd13,5'd10,5'd12,5'd13,5'd21,5'd21,5'd11,5'd15,5'd12,5'd18,5'd24,5'd14,5'd15,5'd6,5'd24,5'd15,5'd5,5'd20,5'd24,5'd24,5'd8,5'd8,5'd12,5'd14,5'd19,5'd19,5'd18,5'd5,5'd14,5'd13,5'd9,5'd20,5'd13,5'd20,5'd18,5'd16,5'd15,5'd15,5'd17,5'd9,5'd14,5'd14,5'd12,5'd12,5'd17,5'd17,5'd22,5'd22,5'd14,5'd14,5'd24,5'd18,5'd17,5'd15,5'd22,5'd22,5'd20,5'd12,5'd14,5'd23,5'd16,5'd18,5'd24,5'd9,5'd20,5'd9,5'd14,5'd8,5'd9,5'd11,5'd12,5'd8,5'd11,5'd12,5'd24,5'd24,5'd24,5'd12,5'd22,5'd23,5'd24,5'd22,5'd22,5'd13,5'd10,5'd12,5'd13,5'd11,5'd14,5'd14,5'd12,5'd10,5'd12,5'd5,5'd14,5'd24,5'd24,5'd24,5'd24,5'd24,5'd24,5'd21,5'd24,5'd13,5'd12,5'd5,5'd14,5'd13,5'd9,5'd23,5'd20,5'd17,5'd23,5'd19,5'd6,5'd23,5'd20,5'd17,5'd18,5'd18,5'd5,5'd5,5'd21,5'd21,5'd21,5'd21,5'd16,5'd12,5'd11,5'd23,5'd20,5'd12,5'd16,5'd24,5'd22,5'd4,5'd15,5'd16,5'd24,5'd22,5'd15,5'd22,5'd22,5'd12,5'd22,5'd23,5'd16,5'd11,5'd9,5'd22,5'd17,5'd17,5'd9,5'd9,5'd22,5'd9,5'd9,5'd15,5'd16,5'd3,5'd6,5'd24,5'd20,5'd14,5'd13,5'd11,5'd9,5'd12,5'd24,5'd17,5'd16,5'd7,5'd20,5'd17,5'd24,5'd24,5'd14,5'd20,5'd5,5'd4,5'd22,5'd24,5'd15,5'd17,5'd17,5'd20,5'd22,5'd24,5'd12,5'd17,5'd17,5'd17,5'd17,5'd14,5'd9,5'd13,5'd19,5'd23,5'd24,5'd20,5'd4,5'd8,5'd8,5'd13,5'd21,5'd23,5'd23,5'd9,5'd11,5'd4,5'd5,5'd18,5'd18,5'd13,5'd22,5'd20,5'd13,5'd14,5'd10,5'd12,5'd12,5'd14,5'd16,5'd15,5'd14,5'd18,5'd24,5'd9,5'd3,5'd5,5'd17,5'd15,5'd13,5'd16,5'd23,5'd23,5'd13,5'd12,5'd23,5'd21,5'd9,5'd20,5'd12,5'd20,5'd19,5'd24,5'd24,5'd14,5'd10,5'd16,5'd16,5'd11,5'd17,5'd8,5'd8,5'd7,5'd8,5'd17,5'd17,5'd18,5'd11,5'd12,5'd24,5'd19,5'd12,5'd24,5'd24,5'd16,5'd24,5'd14,5'd12,5'd9,5'd11,5'd13,5'd20,5'd16,5'd15,5'd17,5'd17,5'd12,5'd12,5'd7,5'd15,5'd10,5'd20,5'd23,5'd24,5'd18,5'd23,5'd24,5'd24,5'd23,5'd23,5'd12,5'd8,5'd4,5'd23,5'd20,5'd21,5'd14,5'd23,5'd19,5'd13,5'd8,5'd21,5'd9,5'd9,5'd13,5'd20,5'd5,5'd8,5'd19,5'd13,5'd14,5'd14,5'd15,5'd8,5'd5,5'd15,5'd12,5'd15,5'd23,5'd9,5'd13,5'd7,5'd20,5'd13,5'd23,5'd6,5'd14,5'd24,5'd10,5'd15,5'd17,5'd5,5'd11,5'd8,5'd11,5'd17,5'd15,5'd10,5'd10,5'd6,5'd8,5'd6,5'd6,5'd8,5'd13,5'd10,5'd10,5'd23,5'd7,5'd17,5'd17,5'd15,5'd17,5'd6,5'd20,5'd14,5'd16,5'd10,5'd10,5'd23,5'd10,5'd12,5'd21,5'd24,5'd24,5'd20,5'd19,5'd19,5'd20,5'd19,5'd24,5'd14,5'd14,5'd17,5'd13,5'd12,5'd24,5'd13,5'd14,5'd14,5'd9,5'd8,5'd18,5'd13,5'd23,5'd22,5'd21,5'd22,5'd22,5'd24,5'd24,5'd8,5'd24,5'd22,5'd18,5'd13,5'd19,5'd24,5'd24,5'd24,5'd16,5'd23,5'd23,5'd24,5'd12,5'd24,5'd17,5'd24,5'd24,5'd22,5'd12,5'd5,5'd6,5'd20,5'd24,5'd22,5'd22,5'd8,5'd8,5'd24,5'd23,5'd14,5'd16,5'd14,5'd14,5'd12,5'd19,5'd23,5'd8,5'd18,5'd14,5'd11,5'd15,5'd24,5'd4,5'd16,5'd9,5'd15,5'd19,5'd17,5'd9,5'd24,5'd13,5'd22,5'd20,5'd19,5'd20,5'd24,5'd24,5'd24,5'd24,5'd24,5'd24,5'd20,5'd17,5'd10,5'd10,5'd13,5'd10,5'd18,5'd18,5'd18,5'd24,5'd16,5'd24,5'd17,5'd9,5'd15,5'd19,5'd22,5'd22,5'd18,5'd21,5'd21,5'd21,5'd6,5'd21,5'd19,5'd14,5'd14,5'd23,5'd15,5'd9,5'd19,5'd14,5'd17,5'd12,5'd6,5'd24,5'd23,5'd17,5'd18,5'd23,5'd23,5'd17,5'd8,5'd13,5'd21,5'd13,5'd12,5'd22,5'd23,5'd11,5'd11,5'd9,5'd9,5'd11,5'd11,5'd9,5'd9,5'd16,5'd16,5'd21,5'd18,5'd15,5'd14,5'd15,5'd24,5'd13,5'd21,5'd23,5'd24,5'd23,5'd24,5'd20,5'd24,5'd11,5'd5,5'd22,5'd21,5'd19,5'd19,5'd15,5'd6,5'd12,5'd18,5'd16,5'd19,5'd21,5'd18,5'd18,5'd13,5'd9,5'd9,5'd24,5'd24,5'd23,5'd21,5'd18,5'd20,5'd23,5'd23,5'd21,5'd21,5'd20,5'd20,5'd6,5'd23,5'd22,5'd13,5'd20,5'd20,5'd20,5'd20,5'd10,5'd9,5'd12,5'd12,5'd16,5'd20,5'd22,5'd24,5'd9,5'd19,5'd24,5'd23,5'd19,5'd18,5'd16,5'd18,5'd11,5'd15,5'd14,5'd19,5'd24,5'd18,5'd24,5'd24,5'd17,5'd24,5'd15,5'd18,5'd24,5'd24,5'd18,5'd18,5'd11,5'd24,5'd14,5'd18,5'd12,5'd18,5'd13,5'd18,5'd20,5'd18,5'd21,5'd20,5'd20,5'd23,5'd9,5'd9,5'd9,5'd15,5'd12,5'd12,5'd16,5'd12,5'd9,5'd16,5'd12,5'd4,5'd3,5'd9,5'd13,5'd13,5'd22,5'd22,5'd17,5'd14,5'd14,5'd2,5'd13,5'd9,5'd9,5'd9,5'd22,5'd21,5'd13,5'd5,5'd14,5'd15,5'd17,5'd24,5'd22,5'd7,5'd13,5'd23,5'd24,5'd23,5'd14,5'd8,5'd8,5'd18,5'd8,5'd23,5'd23,5'd20,5'd7,5'd10,5'd13,5'd24,5'd10,5'd22,5'd12,5'd16,5'd10,5'd21,5'd21,5'd18,5'd18,5'd22,5'd18,5'd16,5'd16,5'd16,5'd15,5'd13,5'd13,5'd17,5'd14,5'd24,5'd24,5'd24,5'd14,5'd19,5'd11,5'd13,5'd21,5'd20,5'd17,5'd11,5'd11,5'd17,5'd6,5'd9,5'd9,5'd13,5'd15,5'd13,5'd6,5'd17,5'd17,5'd11,5'd11,5'd20,5'd16,5'd21,5'd14,5'd11,5'd11,5'd22,5'd12,5'd13,5'd21,5'd19,5'd10,5'd12,5'd21,5'd24,5'd12,5'd18,5'd18,5'd17,5'd20,5'd10,5'd12,5'd13,5'd11,5'd15,5'd12,5'd6,5'd11,5'd13,5'd13,5'd21,5'd13,5'd3,5'd3,5'd19,5'd19,5'd22,5'd22,5'd19,5'd19,5'd23,5'd12,5'd10,5'd15,5'd9,5'd19,5'd18,5'd23,5'd18,5'd14,5'd19,5'd18,5'd14,5'd15,5'd15,5'd14,5'd24,5'd21,5'd9,5'd22,5'd24,5'd21,5'd15,5'd23,5'd11,5'd11,5'd15,5'd15,5'd23,5'd23,5'd15,5'd13,5'd18,5'd24,5'd21,5'd17,5'd10,5'd13,5'd6,5'd13,5'd24,5'd5,5'd6,5'd8,5'd16,5'd13,5'd24,5'd5,5'd4,5'd10,5'd12,5'd4,5'd24,5'd24,5'd12,5'd11,5'd17,5'd7,5'd21,5'd21,5'd24,5'd24,5'd16,5'd12,5'd24,5'd24,5'd19,5'd19,5'd18,5'd21,5'd22,5'd11,5'd18,5'd18,5'd17,5'd14,5'd13,5'd21,5'd24,5'd22,5'd20,5'd4,5'd3,5'd21,5'd20,5'd21,5'd21,5'd21,5'd11,5'd11,5'd23,5'd19,5'd17,5'd6,5'd17,5'd17,5'd21,5'd8,5'd10,5'd21,5'd5,5'd5,5'd14,5'd17,5'd10,5'd10,5'd15,5'd21,5'd12,5'd13,5'd19,5'd14,5'd7,5'd19,5'd12,5'd20,5'd24,5'd24,5'd11,5'd11,5'd15,5'd11,5'd7,5'd23,5'd18,5'd17,5'd5,5'd23,5'd18,5'd20,5'd24,5'd24,5'd5,5'd4,5'd12,5'd13,5'd16,5'd18,5'd13,5'd9,5'd9,5'd17,5'd17,5'd17,5'd6,5'd12,5'd24,5'd14,5'd19,5'd19,5'd19,5'd19,5'd12,5'd12,5'd20,5'd20,5'd14,5'd19,5'd15,5'd14,5'd3,5'd8,5'd21,5'd3,5'd15,5'd22,5'd24,5'd24,5'd23,5'd24,5'd24,5'd15,5'd4,5'd21,5'd10,5'd23,5'd23,5'd18,5'd17,5'd17,5'd15,5'd20,5'd20,5'd19,5'd13,5'd21,5'd24,5'd13,5'd20,5'd16,5'd20,5'd9,5'd22,5'd24,5'd24,5'd16,5'd12,5'd15,5'd15,5'd9,5'd22,5'd22,5'd17,5'd22,5'd7,5'd19,5'd20,5'd22,5'd12,5'd15,5'd24,5'd20,5'd8,5'd13,5'd13,5'd14,5'd17,5'd24,5'd24,5'd19,5'd14,5'd17,5'd17,5'd18,5'd17,5'd24,5'd12,5'd21,5'd21,5'd23,5'd4,5'd12,5'd5,5'd9,5'd12,5'd12,5'd13,5'd18,5'd13,5'd11,5'd11,5'd7,5'd24,5'd7,5'd19,5'd7,5'd19,5'd24,5'd24,5'd6,5'd7,5'd9,5'd22,5'd8,5'd12,5'd21,5'd22,5'd9,5'd22,5'd24,5'd24,5'd12,5'd12,5'd12,5'd6,5'd15,5'd12,5'd15,5'd16,5'd24,5'd24,5'd22,5'd16,5'd18,5'd12,5'd6,5'd24,5'd18,5'd17,5'd12,5'd16,5'd12,5'd12,5'd13,5'd24,5'd18,5'd22,5'd22,5'd18,5'd24,5'd5,5'd19,5'd17,5'd18,5'd19,5'd22,5'd5,5'd11,5'd11,5'd12,5'd12,5'd20,5'd6,5'd2,5'd23,5'd4,5'd15,5'd12,5'd6,5'd19,5'd19,5'd15,5'd16,5'd18,5'd14,5'd19,5'd23,5'd10,5'd8,5'd20,5'd22,5'd12,5'd24,5'd21,5'd21,5'd24,5'd24,5'd20,5'd20,5'd16,5'd14,5'd14,5'd9,5'd9,5'd9,5'd4,5'd14,5'd23,5'd14,5'd18,5'd17,5'd9,5'd9,5'd10,5'd22,5'd15,5'd11,5'd16,5'd21,5'd17,5'd13,5'd15,5'd16,5'd16,5'd16,5'd15,5'd18,5'd20,5'd21,5'd21,5'd19,5'd4,5'd7,5'd9,5'd17,5'd17,5'd20,5'd20,5'd19,5'd20,5'd10,5'd21,5'd14,5'd10,5'd7,5'd21,5'd18,5'd18,5'd18,5'd20,5'd15,5'd14,5'd18,5'd21,5'd18,5'd5,5'd17,5'd24,5'd15,5'd17,5'd24,5'd24,5'd17,5'd17,5'd13,5'd10,5'd23,5'd22,5'd21,5'd21,5'd19,5'd19,5'd15,5'd15,5'd23,5'd23,5'd9,5'd23,5'd12,5'd9,5'd17,5'd15,5'd8,5'd17,5'd20,5'd20,5'd22,5'd21,5'd20,5'd10,5'd12,5'd16,5'd24,5'd17,5'd9,5'd12,5'd20,5'd20,5'd6,5'd22,5'd15,5'd21,5'd16,5'd15,5'd6,5'd11,5'd9,5'd14,5'd14,5'd23,5'd23,5'd12,5'd12,5'd13,5'd17,5'd24,5'd24,5'd9,5'd12,5'd11,5'd11,5'd22,5'd23,5'd20,5'd12,5'd21,5'd20,5'd9,5'd19,5'd9,5'd10,5'd17,5'd10,5'd23,5'd12,5'd14,5'd24,5'd24,5'd24,5'd11,5'd13,5'd17,5'd11,5'd8,5'd8,5'd24,5'd24,5'd14,5'd14,5'd13,5'd11,5'd16,5'd16,5'd16,5'd16,5'd24,5'd24,5'd24,5'd12,5'd18,5'd17,5'd14,5'd14,5'd14,5'd24,5'd12,5'd24,5'd12,5'd24,5'd20,5'd16,5'd9,5'd9,5'd15,5'd15,5'd24,5'd23,5'd24,5'd11,5'd10,5'd19,5'd19,5'd20,5'd19,5'd8,5'd22,5'd20,5'd8,5'd24,5'd11,5'd12,5'd20,5'd18,5'd12,5'd7,5'd11,5'd23,5'd18,5'd24,5'd3,5'd17,5'd9,5'd9,5'd19,5'd16,5'd18,5'd17,5'd18,5'd18,5'd23,5'd17,5'd6,5'd24,5'd4,5'd6,5'd13,5'd24,5'd19,5'd11,5'd12,5'd3,5'd9,5'd24,5'd24,5'd22,5'd16,5'd24,5'd17,5'd9,5'd24,5'd19,5'd21,5'd21,5'd12,5'd21,5'd21,5'd16,5'd20,5'd6,5'd6,5'd22,5'd22,5'd14,5'd14,5'd23,5'd21,5'd17,5'd17,5'd8,5'd8,5'd13,5'd24,5'd10,5'd10,5'd16,5'd16,5'd8,5'd23,5'd23,5'd20,5'd21,5'd19,5'd18,5'd13,5'd17,5'd17,5'd16,5'd20,5'd24,5'd24,5'd19,5'd24,5'd24,5'd10,5'd14,5'd17,5'd3,5'd8,5'd9,5'd24,5'd16,5'd13,5'd16,5'd16,5'd5,5'd6,5'd15,5'd18,5'd22,5'd15,5'd9,5'd18,5'd17,5'd13,5'd5,5'd5,5'd16,5'd10,5'd12,5'd12,5'd23,5'd21,5'd20,5'd12,5'd15,5'd15,5'd24,5'd24,5'd22,5'd24,5'd23,5'd19,5'd17,5'd17,5'd17,5'd12,5'd24,5'd16,5'd5,5'd11,5'd9,5'd12,5'd13,5'd16,5'd5,5'd13,5'd23,5'd24,5'd19,5'd13,5'd10,5'd10,5'd9,5'd16,5'd11,5'd24,5'd16,5'd11,5'd17,5'd21,5'd9,5'd19,5'd19,5'd19,5'd21,5'd24,5'd24,5'd24,5'd11,5'd15,5'd24,5'd23,5'd19,5'd21,5'd21,5'd20,5'd5,5'd10,5'd10,5'd13,5'd11,5'd11,5'd12,5'd17,5'd16,5'd23,5'd8,5'd24,5'd17,5'd19,5'd24,5'd2,5'd8,5'd12,5'd18,5'd20,5'd20,5'd9,5'd9,5'd22,5'd16,5'd20,5'd20,5'd23,5'd23,5'd24,5'd8,5'd13,5'd13,5'd12,5'd13,5'd19,5'd14,5'd13,5'd21,5'd14,5'd14,5'd8,5'd18,5'd24,5'd8,5'd19,5'd19,5'd23,5'd23,5'd24,5'd10,5'd18,5'd15,5'd19,5'd19,5'd6,5'd14,5'd15,5'd22,5'd24,5'd18,5'd15,5'd11,5'd17,5'd12,5'd9,5'd16,5'd23,5'd6,5'd22,5'd18,5'd11,5'd21,5'd11,5'd21,5'd21,5'd18,5'd13,5'd24,5'd21,5'd13,5'd15,5'd8,5'd13,5'd15,5'd23,5'd13,5'd13,5'd12,5'd21,5'd16,5'd17,5'd18,5'd18,5'd24,5'd24,5'd9,5'd9,5'd24,5'd21,5'd22,5'd12,5'd17,5'd22,5'd24,5'd18,5'd20,5'd20,5'd16,5'd18,5'd20,5'd14,5'd20,5'd18,5'd12,5'd18,5'd9,5'd9,5'd6,5'd12,5'd11,5'd11,5'd24,5'd11,5'd24,5'd24,5'd21,5'd20,5'd15,5'd18,5'd5,5'd15,5'd22,5'd20,5'd24,5'd20,5'd11,5'd13,5'd6,5'd24,5'd24,5'd24,5'd18,5'd17,5'd19,5'd22,5'd15,5'd12,5'd22,5'd22,5'd9,5'd21,5'd20,5'd21,5'd21,5'd24,5'd17,5'd6,5'd18,5'd18,5'd9,5'd9,5'd16,5'd11,5'd21,5'd21,5'd16,5'd17,5'd13,5'd13,5'd12,5'd10,5'd19,5'd21,5'd16,5'd13,5'd19,5'd14,5'd20,5'd20,5'd12,5'd12,5'd23,5'd24,5'd12,5'd22,5'd10,5'd16,5'd24,5'd10,5'd15,5'd24,5'd11,5'd11,5'd6,5'd10,5'd18,5'd22,5'd19,5'd19,5'd13,5'd19,5'd22,5'd16,5'd16,5'd12,5'd24,5'd16,5'd14,5'd21,5'd9,5'd21,5'd19,5'd24,5'd11,5'd11,5'd24,5'd19,5'd9,5'd9,5'd8,5'd23,5'd24,5'd17,5'd18,5'd18,5'd12,5'd20,5'd13,5'd9,5'd15,5'd23,5'd24,5'd12,5'd8,5'd24,5'd24,5'd22,5'd24,5'd23,5'd16,5'd15,5'd13,5'd13,5'd18,5'd9,5'd11,5'd14,5'd18,5'd16,5'd16,5'd12,5'd7,5'd18,5'd16,5'd16,5'd17,5'd5,5'd3,5'd17,5'd10,5'd24,5'd9,5'd24,5'd3,5'd9,5'd23,5'd9,5'd20,5'd21,5'd11,5'd14,5'd6,5'd20,5'd22,5'd21,5'd18,5'd20,5'd24,5'd23,5'd23,5'd24,5'd24,5'd17,5'd16,5'd17,5'd16,5'd17,5'd17,5'd19,5'd13,5'd13,5'd9,5'd12,5'd24,5'd6,5'd6,5'd5,5'd6,5'd7,5'd6,5'd16,5'd18,5'd24,5'd22,5'd21,5'd24,5'd19,5'd19,5'd16,5'd21,5'd21,5'd21,5'd16,5'd23,5'd22,5'd22,5'd8,5'd9,5'd15,5'd10,5'd22,5'd23,5'd11,5'd12,5'd6,5'd13,5'd22,5'd22,5'd22,5'd13,5'd21,5'd4,5'd15,5'd24,5'd6,5'd22,5'd21,5'd17,5'd17,5'd17,5'd16,5'd24,5'd21,5'd12,5'd22,5'd18,5'd22,5'd20,5'd9,5'd9,5'd14,5'd14,5'd16,5'd9,5'd21,5'd22,5'd14,5'd14,5'd19,5'd19,5'd4,5'd20,5'd18,5'd12,5'd17,5'd17,5'd24,5'd24,5'd15,5'd15,5'd17,5'd15,5'd23,5'd12,5'd19,5'd6,5'd9,5'd12,5'd15,5'd15,5'd9,5'd15,5'd9,5'd5,5'd19,5'd16,5'd21,5'd21,5'd23,5'd20,5'd19,5'd2,5'd21,5'd16,5'd20,5'd21,5'd19,5'd12,5'd18,5'd21,5'd19,5'd24,5'd16,5'd16,5'd23,5'd16,5'd6,5'd11,5'd13,5'd13,5'd24,5'd12,5'd19,5'd10,5'd10,5'd9,5'd10,5'd14,5'd13,5'd24,5'd15,5'd14,5'd23,5'd11,5'd24,5'd18,5'd23,5'd16,5'd16,5'd12,5'd24,5'd18,5'd15,5'd20,5'd14,5'd6,5'd19,5'd24,5'd15,5'd19,5'd11,5'd14,5'd18,5'd15,5'd17,5'd9,5'd16,5'd24,5'd5,5'd20,5'd11,5'd12,5'd6,5'd24,5'd14,5'd21,5'd24,5'd24,5'd18,5'd11,5'd13}
`define RECTANGLE1_WEIGHTS {32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168}
`define RECTANGLE2_X1 {5'd12,5'd0,5'd17,5'd3,5'd12,5'd0,5'd15,5'd0,5'd3,5'd0,5'd15,5'd1,5'd15,5'd0,5'd21,5'd12,5'd0,5'd0,5'd16,5'd3,5'd13,5'd3,5'd13,5'd10,5'd14,5'd2,5'd6,5'd5,5'd15,5'd1,5'd18,5'd0,5'd20,5'd5,5'd12,5'd3,5'd18,5'd2,5'd11,5'd9,5'd5,5'd5,5'd11,5'd8,5'd14,5'd9,5'd14,5'd4,5'd5,5'd12,5'd9,5'd8,5'd14,5'd10,5'd12,5'd2,5'd6,5'd9,5'd5,5'd8,5'd8,5'd1,5'd9,5'd0,5'd5,5'd1,5'd12,5'd1,5'd10,5'd1,5'd8,5'd4,5'd4,5'd5,5'd12,5'd6,5'd0,5'd1,5'd9,5'd10,5'd12,5'd12,5'd12,5'd0,5'd7,5'd1,5'd14,5'd1,5'd11,5'd11,5'd12,5'd0,5'd12,5'd5,5'd6,5'd3,5'd18,5'd10,5'd12,5'd4,5'd8,5'd6,5'd12,5'd7,5'd2,5'd0,5'd6,5'd9,5'd12,5'd0,5'd12,5'd0,5'd15,5'd6,5'd14,5'd5,5'd12,5'd3,5'd17,5'd7,5'd16,5'd10,5'd4,5'd3,5'd4,5'd5,5'd12,5'd0,5'd5,5'd0,5'd14,5'd0,5'd15,5'd0,5'd19,5'd2,5'd17,5'd7,5'd18,5'd0,5'd3,5'd1,5'd21,5'd4,5'd20,5'd0,5'd6,5'd0,5'd0,5'd0,5'd18,5'd12,5'd11,5'd7,5'd6,5'd5,5'd9,5'd4,5'd6,5'd0,5'd11,5'd10,5'd9,5'd0,5'd17,5'd5,5'd3,5'd10,5'd10,5'd2,5'd20,5'd6,5'd6,5'd2,5'd5,5'd9,5'd9,5'd11,5'd2,5'd2,5'd5,5'd10,5'd8,5'd8,5'd13,5'd3,5'd16,5'd10,5'd11,5'd4,5'd5,5'd9,5'd11,5'd4,5'd15,5'd3,5'd12,5'd5,5'd10,5'd6,5'd9,5'd19,5'd9,5'd8,5'd0,5'd13,5'd3,5'd12,5'd12,5'd11,5'd4,5'd16,5'd5,5'd17,5'd2,5'd20,5'd3,5'd18,5'd7,5'd10,5'd8,5'd15,5'd2,5'd3,5'd7,5'd2,5'd2,5'd10,5'd6,5'd17,5'd9,5'd12,5'd10,5'd13,5'd8,5'd15,5'd11,5'd12,5'd4,5'd12,5'd0,5'd12,5'd4,5'd11,5'd8,5'd11,5'd12,5'd7,5'd9,5'd11,5'd8,5'd8,5'd2,5'd20,5'd2,5'd21,5'd0,5'd10,5'd8,5'd12,5'd0,5'd16,5'd1,5'd6,5'd3,5'd9,5'd3,5'd14,5'd10,5'd7,5'd1,5'd14,5'd5,5'd17,5'd0,5'd6,5'd10,5'd16,5'd10,5'd12,5'd9,5'd6,5'd0,5'd15,5'd3,5'd10,5'd4,5'd11,5'd10,5'd7,5'd9,5'd9,5'd3,5'd20,5'd1,5'd15,5'd0,5'd8,5'd1,5'd17,5'd2,5'd13,5'd0,5'd18,5'd3,5'd15,5'd7,5'd16,5'd8,5'd16,5'd4,5'd3,5'd0,5'd10,5'd6,5'd13,5'd9,5'd18,5'd7,5'd14,5'd7,5'd7,5'd3,5'd14,5'd10,5'd12,5'd10,5'd6,5'd5,5'd15,5'd1,5'd19,5'd9,5'd11,5'd10,5'd9,5'd7,5'd12,5'd10,5'd12,5'd3,5'd11,5'd0,5'd0,5'd0,5'd4,5'd8,5'd5,5'd7,5'd11,5'd9,5'd13,5'd9,5'd12,5'd3,5'd13,5'd9,5'd12,5'd10,5'd12,5'd9,5'd12,5'd11,5'd5,5'd5,5'd9,5'd1,5'd14,5'd2,5'd18,5'd0,5'd16,5'd7,5'd18,5'd0,5'd15,5'd0,5'd21,5'd7,5'd11,5'd12,5'd7,5'd7,5'd10,5'd8,5'd15,5'd8,5'd14,5'd0,5'd6,5'd0,5'd14,5'd0,5'd14,5'd0,5'd3,5'd8,5'd13,5'd8,5'd12,5'd4,5'd13,5'd6,5'd4,5'd3,5'd18,5'd8,5'd2,5'd4,5'd10,5'd5,5'd3,5'd5,5'd8,5'd9,5'd3,5'd15,5'd0,5'd4,5'd7,5'd13,5'd0,5'd18,5'd6,5'd15,5'd3,5'd18,5'd8,5'd18,5'd4,5'd16,5'd6,5'd11,5'd6,5'd9,5'd12,5'd16,5'd6,5'd18,5'd6,5'd18,5'd11,5'd18,5'd1,5'd18,5'd3,5'd12,5'd10,5'd6,5'd1,5'd8,5'd6,5'd15,5'd0,5'd15,5'd2,5'd13,5'd1,5'd7,5'd8,5'd12,5'd9,5'd12,5'd2,5'd12,5'd10,5'd12,5'd9,5'd14,5'd5,5'd4,5'd4,5'd12,5'd9,5'd12,5'd6,5'd15,5'd4,5'd15,5'd5,5'd11,5'd8,5'd11,5'd5,5'd17,5'd7,5'd0,5'd2,5'd17,5'd2,5'd10,5'd3,5'd14,5'd2,5'd9,5'd6,5'd13,5'd10,5'd12,5'd2,5'd12,5'd6,5'd10,5'd5,5'd16,5'd5,5'd3,5'd3,5'd0,5'd0,5'd1,5'd9,5'd13,5'd2,5'd4,5'd3,5'd12,5'd10,5'd6,5'd7,5'd12,5'd6,5'd15,5'd9,5'd6,5'd4,5'd12,5'd5,5'd16,5'd1,5'd15,5'd11,5'd11,5'd7,5'd15,5'd8,5'd13,5'd2,5'd14,5'd0,5'd10,5'd11,5'd7,5'd0,5'd22,5'd0,5'd19,5'd3,5'd12,5'd8,5'd9,5'd8,5'd13,5'd8,5'd15,5'd11,5'd12,5'd7,5'd22,5'd3,5'd14,5'd7,5'd13,5'd11,5'd15,5'd1,5'd21,5'd0,5'd6,5'd2,5'd13,5'd0,5'd14,5'd4,5'd17,5'd6,5'd12,5'd5,5'd14,5'd6,5'd9,5'd2,5'd12,5'd3,5'd13,5'd0,5'd7,5'd6,5'd8,5'd0,5'd13,5'd7,5'd17,5'd12,5'd17,5'd0,5'd11,5'd1,5'd7,5'd0,5'd11,5'd10,5'd5,5'd2,5'd20,5'd3,5'd19,5'd6,5'd8,5'd4,5'd7,5'd20,5'd5,5'd10,5'd3,5'd11,5'd5,5'd14,5'd10,5'd12,5'd2,5'd19,5'd6,5'd15,5'd10,5'd15,5'd9,5'd9,5'd8,5'd0,5'd9,5'd10,5'd9,5'd12,5'd0,5'd13,5'd9,5'd17,5'd7,5'd12,5'd10,5'd14,5'd5,5'd12,5'd2,5'd8,5'd6,5'd12,5'd9,5'd3,5'd0,5'd0,5'd6,5'd10,5'd0,5'd4,5'd7,5'd14,5'd6,5'd16,5'd3,5'd4,5'd4,5'd3,5'd5,5'd16,5'd5,5'd17,5'd12,5'd10,5'd11,5'd0,5'd4,5'd16,5'd3,5'd10,5'd7,5'd12,5'd7,5'd10,5'd6,5'd16,5'd3,5'd12,5'd9,5'd13,5'd8,5'd13,5'd2,5'd13,5'd0,5'd6,5'd0,5'd10,5'd1,5'd15,5'd2,5'd11,5'd0,5'd5,5'd10,5'd13,5'd10,5'd13,5'd10,5'd13,5'd7,5'd13,5'd1,5'd15,5'd0,5'd9,5'd7,5'd21,5'd3,5'd21,5'd7,5'd11,5'd7,5'd10,5'd0,5'd6,5'd12,5'd12,5'd2,5'd4,5'd0,5'd13,5'd0,5'd5,5'd5,5'd20,5'd2,5'd0,5'd7,5'd5,5'd2,5'd7,5'd7,5'd14,5'd5,5'd10,5'd4,5'd12,5'd1,5'd16,5'd2,5'd18,5'd9,5'd12,5'd5,5'd2,5'd9,5'd6,5'd10,5'd1,5'd12,5'd5,5'd0,5'd21,5'd2,5'd10,5'd11,5'd9,5'd9,5'd6,5'd4,5'd12,5'd10,5'd11,5'd5,5'd10,5'd2,5'd9,5'd3,5'd18,5'd7,5'd18,5'd3,5'd7,5'd9,5'd11,5'd0,5'd18,5'd2,5'd6,5'd0,5'd11,5'd3,5'd8,5'd4,5'd1,5'd4,5'd0,5'd14,5'd0,5'd14,5'd6,5'd12,5'd8,5'd12,5'd0,5'd13,5'd7,5'd11,5'd2,5'd13,5'd8,5'd12,5'd10,5'd16,5'd10,5'd1,5'd0,5'd14,5'd9,5'd13,5'd0,5'd10,5'd8,5'd14,5'd9,5'd13,5'd10,5'd12,5'd4,5'd9,5'd0,5'd15,5'd0,5'd16,5'd5,5'd17,5'd7,5'd3,5'd2,5'd13,5'd2,5'd13,5'd1,5'd13,5'd12,5'd13,5'd2,5'd20,5'd4,5'd9,5'd6,5'd12,5'd7,5'd6,5'd0,5'd4,5'd3,5'd15,5'd1,5'd6,5'd1,5'd1,5'd7,5'd0,5'd5,5'd17,5'd6,5'd16,5'd1,5'd19,5'd0,5'd7,5'd12,5'd14,5'd7,5'd15,5'd3,5'd14,5'd1,5'd15,5'd4,5'd18,5'd11,5'd11,5'd9,5'd9,5'd1,5'd1,5'd0,5'd9,5'd1,5'd11,5'd12,5'd12,5'd7,5'd14,5'd6,5'd11,5'd1,5'd11,5'd0,5'd4,5'd10,5'd12,5'd10,5'd11,5'd8,5'd10,5'd11,5'd12,5'd0,5'd13,5'd3,5'd11,5'd8,5'd14,5'd9,5'd10,5'd11,5'd10,5'd8,5'd14,5'd1,5'd14,5'd0,5'd0,5'd8,5'd6,5'd1,5'd13,5'd1,5'd9,5'd3,5'd15,5'd0,5'd14,5'd1,5'd14,5'd3,5'd15,5'd6,5'd12,5'd9,5'd15,5'd4,5'd6,5'd4,5'd9,5'd1,5'd3,5'd4,5'd19,5'd1,5'd9,5'd6,5'd7,5'd1,5'd20,5'd11,5'd12,5'd12,5'd13,5'd9,5'd13,5'd5,5'd17,5'd3,5'd14,5'd2,5'd12,5'd8,5'd7,5'd1,5'd12,5'd2,5'd14,5'd2,5'd20,5'd7,5'd15,5'd0,5'd1,5'd8,5'd11,5'd8,5'd15,5'd6,5'd10,5'd10,5'd6,5'd7,5'd9,5'd11,5'd13,5'd8,5'd12,5'd7,5'd14,5'd1,5'd0,5'd1,5'd13,5'd0,5'd11,5'd1,5'd14,5'd5,5'd6,5'd1,5'd5,5'd1,5'd12,5'd0,5'd21,5'd0,5'd17,5'd0,5'd8,5'd9,5'd13,5'd8,5'd7,5'd4,5'd14,5'd6,5'd15,5'd8,5'd14,5'd6,5'd6,5'd8,5'd18,5'd4,5'd2,5'd2,5'd17,5'd4,5'd6,5'd3,5'd16,5'd0,5'd14,5'd11,5'd10,5'd6,5'd8,5'd6,5'd16,5'd3,5'd6,5'd8,5'd10,5'd5,5'd12,5'd0,5'd5,5'd0,5'd12,5'd9,5'd16,5'd2,5'd20,5'd0,5'd15,5'd4,5'd18,5'd4,5'd16,5'd5,5'd17,5'd12,5'd18,5'd10,5'd13,5'd4,5'd17,5'd7,5'd13,5'd7,5'd11,5'd2,5'd14,5'd0,5'd13,5'd9,5'd12,5'd4,5'd9,5'd3,5'd14,5'd2,5'd5,5'd0,5'd8,5'd2,5'd16,5'd11,5'd7,5'd1,5'd12,5'd0,5'd14,5'd0,5'd9,5'd9,5'd13,5'd10,5'd7,5'd9,5'd12,5'd7,5'd8,5'd5,5'd15,5'd9,5'd12,5'd7,5'd15,5'd3,5'd15,5'd10,5'd7,5'd11,5'd10,5'd1,5'd15,5'd1,5'd11,5'd2,5'd17,5'd7,5'd10,5'd10,5'd6,5'd6,5'd13,5'd3,5'd6,5'd0,5'd15,5'd0,5'd4,5'd0,5'd6,5'd8,5'd12,5'd3,5'd12,5'd12,5'd15,5'd10,5'd13,5'd4,5'd16,5'd4,5'd3,5'd11,5'd4,5'd5,5'd14,5'd12,5'd14,5'd9,5'd7,5'd4,5'd14,5'd6,5'd9,5'd0,5'd14,5'd3,5'd19,5'd6,5'd16,5'd7,5'd16,5'd11,5'd11,5'd9,5'd2,5'd3,5'd9,5'd8,5'd5,5'd4,5'd10,5'd3,5'd10,5'd3,5'd7,5'd3,5'd10,5'd9,5'd7,5'd10,5'd1,5'd9,5'd6,5'd0,5'd1,5'd10,5'd6,5'd12,5'd0,5'd13,5'd0,5'd8,5'd4,5'd16,5'd0,5'd14,5'd5,5'd14,5'd5,5'd12,5'd11,5'd6,5'd11,5'd11,5'd0,5'd4,5'd9,5'd7,5'd9,5'd5,5'd10,5'd12,5'd5,5'd2,5'd3,5'd12,5'd0,5'd18,5'd9,5'd9,5'd0,5'd2,5'd0,5'd15,5'd9,5'd11,5'd11,5'd10,5'd10,5'd1,5'd11,5'd17,5'd5,5'd6,5'd4,5'd11,5'd9,5'd5,5'd8,5'd3,5'd1,5'd12,5'd1,5'd19,5'd0,5'd15,5'd7,5'd20,5'd3,5'd13,5'd9,5'd7,5'd5,5'd16,5'd8,5'd11,5'd10,5'd13,5'd0,5'd18,5'd3,5'd18,5'd8,5'd14,5'd12,5'd9,5'd11,5'd9,5'd9,5'd9,5'd9,5'd14,5'd6,5'd4,5'd10,5'd13,5'd9,5'd1,5'd8,5'd4,5'd2,5'd14,5'd4,5'd11,5'd8,5'd10,5'd4,5'd11,5'd5,5'd0,5'd0,5'd13,5'd8,5'd20,5'd3,5'd15,5'd0,5'd15,5'd0,5'd17,5'd4,5'd15,5'd2,5'd9,5'd0,5'd15,5'd2,5'd9,5'd1,5'd13,5'd8,5'd14,5'd7,5'd9,5'd0,5'd12,5'd12,5'd12,5'd10,5'd12,5'd10,5'd12,5'd2,5'd17,5'd5,5'd13,5'd3,5'd3,5'd2,5'd12,5'd8,5'd20,5'd4,5'd13,5'd2,5'd15,5'd3,5'd11,5'd0,5'd9,5'd7,5'd7,5'd13,5'd10,5'd14,5'd10,5'd12,5'd12,5'd12,5'd3,5'd12,5'd1,5'd19,5'd0,5'd17,5'd9,5'd7,5'd10,5'd12,5'd2,5'd0,5'd0,5'd8,5'd2,5'd11,5'd12,5'd8,5'd6,5'd4,5'd3,5'd15,5'd10,5'd12,5'd7,5'd12,5'd7,5'd9,5'd7,5'd12,5'd0,5'd18,5'd2,5'd1,5'd1,5'd6,5'd4,5'd18,5'd1,5'd6,5'd0,5'd14,5'd8,5'd0,5'd4,5'd10,5'd5,5'd15,5'd1,5'd19,5'd10,5'd19,5'd4,5'd3,5'd2,5'd14,5'd3,5'd17,5'd4,5'd7,5'd8,5'd13,5'd9,5'd13,5'd6,5'd14,5'd0,5'd19,5'd8,5'd12,5'd12,5'd15,5'd1,5'd10,5'd4,5'd16,5'd5,5'd14,5'd12,5'd12,5'd9,5'd17,5'd1,5'd20,5'd10,5'd11,5'd10,5'd14,5'd7,5'd10,5'd12,5'd13,5'd1,5'd2,5'd11,5'd13,5'd8,5'd10,5'd10,5'd0,5'd2,5'd9,5'd0,5'd12,5'd0,5'd3,5'd5,5'd8,5'd8,5'd17,5'd4,5'd14,5'd6,5'd5,5'd0,5'd18,5'd1,5'd3,5'd1,5'd14,5'd3,5'd14,5'd10,5'd14,5'd2,5'd12,5'd12,5'd12,5'd7,5'd15,5'd11,5'd5,5'd4,5'd18,5'd3,5'd18,5'd8,5'd10,5'd7,5'd9,5'd6,5'd2,5'd4,5'd17,5'd6,5'd7,5'd8,5'd1,5'd2,5'd7,5'd12,5'd8,5'd14,5'd9,5'd11,5'd10,5'd5,5'd12,5'd7,5'd11,5'd10,5'd5,5'd14,5'd2,5'd3,5'd0,5'd18,5'd1,5'd17,5'd0,5'd19,5'd6,5'd8,5'd4,5'd14,5'd10,5'd12,5'd6,5'd9,5'd1,5'd19,5'd1,5'd9,5'd8,5'd12,5'd6,5'd3,5'd5,5'd9,5'd5,5'd13,5'd2,5'd11,5'd0,5'd12,5'd10,5'd13,5'd7,5'd13,5'd2,5'd18,5'd3,5'd4,5'd9,5'd4,5'd11,5'd7,5'd6,5'd3,5'd2,5'd20,5'd1,5'd22,5'd8,5'd15,5'd0,5'd17,5'd1,5'd18,5'd3,5'd16,5'd4,5'd17,5'd3,5'd8,5'd0,5'd19,5'd5,5'd4,5'd0,5'd11,5'd10,5'd14,5'd3,5'd16,5'd5,5'd17,5'd4,5'd13,5'd1,5'd14,5'd0,5'd6,5'd0,5'd13,5'd0,5'd14,5'd0,5'd20,5'd1,5'd12,5'd12,5'd14,5'd7,5'd13,5'd11,5'd12,5'd10,5'd13,5'd8,5'd13,5'd8,5'd13,5'd0,5'd5,5'd0,5'd15,5'd0,5'd15,5'd5,5'd17,5'd9,5'd12,5'd2,5'd0,5'd0,5'd17,5'd0,5'd18,5'd1,5'd2,5'd0,5'd13,5'd2,5'd20,5'd0,5'd15,5'd6,5'd10,5'd0,5'd3,5'd9,5'd13,5'd7,5'd15,5'd1,5'd7,5'd8,5'd4,5'd8,5'd11,5'd6,5'd9,5'd9,5'd8,5'd4,5'd10,5'd10,5'd0,5'd0,5'd0,5'd16,5'd3,5'd12,5'd11,5'd10,5'd7,5'd16,5'd0,5'd7,5'd12,5'd8,5'd10,5'd7,5'd3,5'd14,5'd0,5'd15,5'd0,5'd15,5'd4,5'd15,5'd3,5'd15,5'd4,5'd12,5'd8,5'd12,5'd9,5'd12,5'd1,5'd16,5'd0,5'd18,5'd0,5'd12,5'd7,5'd8,5'd10,5'd4,5'd11,5'd9,5'd12,5'd8,5'd8,5'd14,5'd2,5'd20,5'd2,5'd6,5'd8,5'd13,5'd9,5'd6,5'd12,5'd9,5'd5,5'd13,5'd0,5'd18,5'd5,5'd12,5'd5,5'd13,5'd0,5'd2,5'd0,5'd3,5'd3,5'd17,5'd8,5'd15,5'd11,5'd11,5'd3,5'd16,5'd3,5'd14,5'd0,5'd9,5'd1,5'd18,5'd6,5'd16,5'd9,5'd16,5'd1,5'd5,5'd1,5'd5,5'd2,5'd13,5'd0,5'd15,5'd9,5'd16,5'd3,5'd10,5'd9,5'd15,5'd1,5'd13,5'd6,5'd18,5'd5,5'd14,5'd10,5'd12,5'd12,5'd11,5'd12,5'd16,5'd9,5'd8,5'd2,5'd20,5'd3,5'd8,5'd4,5'd14,5'd8,5'd14,5'd4,5'd14,5'd1,5'd19,5'd2,5'd3,5'd8,5'd15,5'd11,5'd6,5'd6,5'd2,5'd0,5'd7,5'd2,5'd4,5'd5,5'd2,5'd9,5'd12,5'd5,5'd12,5'd0,5'd12,5'd2,5'd17,5'd9,5'd11,5'd5,5'd13,5'd3,5'd12,5'd3,5'd12,5'd12,5'd7,5'd3,5'd11,5'd1,5'd16,5'd9,5'd12,5'd4,5'd8,5'd8,5'd17,5'd6,5'd11,5'd8,5'd9,5'd5,5'd14,5'd6,5'd5,5'd0,5'd12,5'd1,5'd12,5'd2,5'd12,5'd0,5'd12,5'd7,5'd10,5'd10,5'd5,5'd9,5'd11,5'd11,5'd5,5'd8,5'd10,5'd0,5'd14,5'd5,5'd12,5'd2,5'd3,5'd11,5'd12,5'd11,5'd11,5'd7,5'd10,5'd12,5'd16,5'd3,5'd16,5'd3,5'd15,5'd10,5'd12,5'd11,5'd7,5'd12,5'd16,5'd0,5'd9,5'd1,5'd15,5'd0,5'd14,5'd1,5'd20,5'd2,5'd2,5'd1,5'd12,5'd0,5'd13,5'd5,5'd14,5'd7,5'd11,5'd1,5'd10,5'd9,5'd6,5'd9,5'd5,5'd8,5'd13,5'd3,5'd18,5'd2,5'd20,5'd0,5'd6,5'd0,5'd12,5'd10,5'd20,5'd0,5'd6,5'd8,5'd4,5'd5,5'd8,5'd0,5'd20,5'd8,5'd20,5'd3,5'd11,5'd8,5'd1,5'd7,5'd2,5'd17,5'd7,5'd9,5'd1,5'd11,5'd6,5'd14,5'd12,5'd6,5'd1,5'd18,5'd2,5'd12,5'd7,5'd14,5'd10,5'd12,5'd9,5'd20,5'd0,5'd12,5'd5,5'd14,5'd11,5'd12,5'd5,5'd13,5'd4,5'd6,5'd0,5'd9,5'd8,5'd5,5'd3,5'd8,5'd1,5'd9,5'd9,5'd13,5'd2,5'd4,5'd9,5'd13,5'd11,5'd12,5'd9,5'd18,5'd9,5'd10,5'd5,5'd7,5'd2,5'd3,5'd0,5'd0,5'd10,5'd6,5'd4,5'd5,5'd3,5'd12,5'd4,5'd12,5'd11,5'd8,5'd10,5'd1,5'd5,5'd2,5'd0,5'd5,5'd3,5'd19,5'd5,5'd13,5'd9,5'd9,5'd5,5'd5,5'd5,5'd16,5'd0,5'd16,5'd6,5'd12,5'd7,5'd14,5'd7,5'd13,5'd4,5'd15,5'd0,5'd10,5'd11,5'd18,5'd7,5'd11,5'd6,5'd13,5'd2,5'd10,5'd5,5'd18,5'd0,5'd12,5'd6,5'd12,5'd9,5'd5,5'd2,5'd14,5'd2,5'd14,5'd10,5'd4,5'd8,5'd12,5'd0,5'd14,5'd0,5'd12,5'd2,5'd20,5'd2,5'd10,5'd0,5'd11,5'd3,5'd8,5'd2,5'd11,5'd7,5'd9,5'd4,5'd7,5'd14,5'd9,5'd14,5'd7,5'd11,5'd2,5'd8,5'd1,5'd6,5'd1,5'd12,5'd9,5'd11,5'd1,5'd9,5'd8,5'd14,5'd3,5'd11,5'd7,5'd12,5'd12,5'd15,5'd8,5'd5,5'd11,5'd4,5'd10,5'd9,5'd8,5'd12,5'd11,5'd11,5'd0,5'd12,5'd11,5'd18,5'd6,5'd15,5'd1,5'd13,5'd8,5'd12,5'd8,5'd12,5'd10,5'd6,5'd0,5'd15,5'd1,5'd12,5'd2,5'd12,5'd8,5'd13,5'd0,5'd15,5'd0,5'd17,5'd0,5'd12,5'd7,5'd10,5'd5,5'd16,5'd5,5'd13,5'd1,5'd15,5'd4,5'd12,5'd4,5'd13,5'd1,5'd1,5'd0,5'd11,5'd9,5'd18,5'd0,5'd20,5'd0,5'd19,5'd1,5'd12,5'd5,5'd13,5'd8,5'd9,5'd0,5'd4,5'd11,5'd12,5'd10,5'd12,5'd2,5'd3,5'd10,5'd3,5'd3,5'd14,5'd1,5'd10,5'd2,5'd16,5'd0,5'd15,5'd3,5'd20,5'd2,5'd16,5'd2,5'd15,5'd9,5'd20,5'd8,5'd19,5'd1,5'd8,5'd5,5'd15,5'd0,5'd12,5'd5,5'd10,5'd2,5'd4,5'd10,5'd6,5'd17,5'd3,5'd14,5'd2,5'd4,5'd8,5'd10,5'd0,5'd13,5'd0,5'd20,5'd3,5'd19,5'd0,5'd1,5'd2,5'd22,5'd3,5'd18,5'd2,5'd12,5'd3,5'd11,5'd1,5'd13,5'd12,5'd2,5'd2,5'd18,5'd0,5'd2,5'd8,5'd18,5'd9,5'd9,5'd1,5'd8,5'd9,5'd11,5'd11,5'd12,5'd4,5'd17,5'd8,5'd13,5'd6,5'd13,5'd8,5'd14,5'd0,5'd15,5'd10,5'd17,5'd7,5'd5,5'd0,5'd15,5'd6,5'd15,5'd5,5'd15,5'd9,5'd13,5'd12,5'd13,5'd1,5'd14,5'd7,5'd6,5'd3,5'd1,5'd1,5'd5,5'd1,5'd3,5'd8,5'd5,5'd5,5'd3,5'd5,5'd8,5'd7,5'd12,5'd6,5'd14,5'd10,5'd10,5'd5,5'd13,5'd0,5'd11,5'd6,5'd16,5'd6,5'd7,5'd8,5'd13,5'd4,5'd13,5'd8,5'd13,5'd3,5'd9,5'd3,5'd18,5'd3,5'd11,5'd5,5'd10,5'd3,5'd8,5'd7,5'd2,5'd17,5'd1,5'd12,5'd3,5'd3,5'd0,5'd12,5'd6,5'd11,5'd3,5'd15,5'd8,5'd14,5'd11,5'd14,5'd0,5'd15,5'd0,5'd10,5'd10,5'd5,5'd6,5'd8,5'd5,5'd17,5'd0,5'd15,5'd6,5'd4,5'd3,5'd19,5'd3,5'd19,5'd3,5'd15,5'd2,5'd8,5'd3,5'd6,5'd0,5'd13,5'd9,5'd13,5'd8,5'd10,5'd0,5'd20,5'd3,5'd20,5'd8,5'd13,5'd12,5'd12,5'd3,5'd3,5'd6,5'd14,5'd6,5'd14,5'd9,5'd13,5'd0,5'd15,5'd12,5'd22,5'd7,5'd11,5'd8,5'd22,5'd5,5'd18,5'd5,5'd14,5'd2,5'd12,5'd0,5'd18,5'd9,5'd3,5'd2,5'd19,5'd0,5'd15,5'd1,5'd14,5'd9,5'd14,5'd0,5'd10,5'd8,5'd10,5'd2,5'd3,5'd9,5'd1,5'd8,5'd10,5'd6,5'd8,5'd10,5'd5,5'd9,5'd6,5'd16,5'd10,5'd12,5'd11,5'd6,5'd6,5'd14,5'd10,5'd14,5'd12,5'd17,5'd2,5'd18,5'd2,5'd14,5'd5,5'd8,5'd6,5'd19,5'd7,5'd15,5'd1,5'd12,5'd9,5'd15,5'd0,5'd6,5'd3,5'd13,5'd0,5'd12,5'd0,5'd19,5'd0,5'd14,5'd6,5'd2,5'd3,5'd12,5'd12,5'd12,5'd4,5'd6,5'd10,5'd8,5'd0,5'd5,5'd5,5'd10,5'd1,5'd6,5'd8,5'd14,5'd9,5'd9,5'd8,5'd14,5'd1,5'd17,5'd0,5'd9,5'd0,5'd18,5'd7,5'd18,5'd6,5'd20,5'd8,5'd14,5'd9,5'd13,5'd10,5'd9,5'd8,5'd12,5'd6,5'd13,5'd5,5'd20,5'd3,5'd3,5'd3,5'd11,5'd5,5'd14,5'd8,5'd10,5'd6,5'd12,5'd11,5'd11,5'd12,5'd6,5'd16,5'd4,5'd5,5'd7,5'd14,5'd0,5'd16,5'd8,5'd12,5'd9,5'd13,5'd0,5'd6,5'd1,5'd6,5'd7,5'd15,5'd8,5'd12,5'd4,5'd12,5'd7,5'd16,5'd1,5'd20,5'd6,5'd14,5'd2,5'd4,5'd0,5'd15,5'd3,5'd18,5'd5,5'd17,5'd0,5'd14,5'd1,5'd12,5'd1,5'd14,5'd1,5'd18,5'd9,5'd13,5'd9,5'd15,5'd8,5'd11,5'd5,5'd15,5'd3,5'd15,5'd10,5'd12,5'd6,5'd5,5'd0,5'd18,5'd3,5'd18,5'd0,5'd21,5'd9,5'd16,5'd10,5'd3,5'd2,5'd9,5'd7,5'd11,5'd4,5'd5,5'd10,5'd6,5'd8,5'd12,5'd3,5'd10,5'd1,5'd15,5'd1,5'd12,5'd8,5'd9,5'd10,5'd13,5'd11,5'd5,5'd2,5'd14,5'd7,5'd9,5'd8,5'd15,5'd8,5'd14,5'd9,5'd13,5'd10,5'd8,5'd0,5'd18,5'd0,5'd9,5'd4,5'd0,5'd2,5'd16,5'd6,5'd12,5'd12,5'd9,5'd8,5'd9,5'd0,5'd8,5'd0,5'd15,5'd8,5'd15,5'd0,5'd15,5'd0,5'd7,5'd8,5'd7,5'd9,5'd6,5'd9,5'd12,5'd10,5'd13,5'd1,5'd14,5'd6,5'd12,5'd3,5'd15,5'd8,5'd10,5'd4,5'd7,5'd3,5'd17,5'd11,5'd15,5'd3,5'd14,5'd1,5'd20,5'd10,5'd9,5'd11,5'd8,5'd4,5'd12,5'd0,5'd10,5'd8,5'd10,5'd10,5'd13,5'd4,5'd12,5'd0,5'd3,5'd9,5'd12,5'd5,5'd7,5'd4,5'd14,5'd5,5'd12,5'd2,5'd13,5'd10,5'd13,5'd9,5'd13,5'd0,5'd13,5'd1,5'd18,5'd3,5'd18,5'd6,5'd11,5'd10,5'd11,5'd0,5'd13,5'd2,5'd1,5'd0,5'd13,5'd2,5'd5,5'd2,5'd5,5'd2,5'd20,5'd9,5'd5,5'd4,5'd10,5'd10,5'd6,5'd6,5'd0,5'd13,5'd3,5'd13,5'd6,5'd18,5'd9,5'd14,5'd9,5'd14,5'd12,5'd13,5'd0,5'd7,5'd9,5'd12,5'd9,5'd1,5'd0,5'd7,5'd8,5'd8,5'd8,5'd13,5'd1,5'd13,5'd12,5'd13,5'd7,5'd14,5'd10,5'd8,5'd7,5'd8,5'd3,5'd18,5'd5,5'd14,5'd2,5'd9,5'd2,5'd16,5'd3,5'd18,5'd3,5'd18,5'd9,5'd4,5'd0,5'd9,5'd10,5'd6,5'd8,5'd19,5'd4,5'd16,5'd5,5'd8,5'd12,5'd3,5'd8,5'd10,5'd3,5'd3,5'd6,5'd4,5'd4,5'd14,5'd5,5'd3,5'd2,5'd2,5'd9,5'd12,5'd0,5'd8,5'd8,5'd14,5'd0,5'd17,5'd8,5'd14,5'd4,5'd12,5'd2,5'd20,5'd5,5'd6,5'd1,5'd6,5'd0,5'd7,5'd6,5'd10,5'd1,5'd9,5'd11,5'd11,5'd9,5'd11,5'd8,5'd11,5'd4,5'd8,5'd6,5'd9,5'd10,5'd12,5'd9,5'd11,5'd9,5'd10,5'd5,5'd15,5'd1,5'd14,5'd3,5'd5,5'd1,5'd3,5'd2,5'd4,5'd1,5'd15,5'd8,5'd6,5'd3,5'd14,5'd1,5'd8,5'd3,5'd19,5'd2,5'd4,5'd8,5'd10,5'd6,5'd0,5'd17,5'd1,5'd12,5'd10,5'd12,5'd0,5'd12,5'd2,5'd20,5'd11,5'd20,5'd2,5'd2,5'd10,5'd2,5'd5,5'd8,5'd4,5'd18,5'd5,5'd9,5'd6,5'd11,5'd9,5'd5,5'd8,5'd5,5'd7,5'd11,5'd8,5'd20,5'd4,5'd12,5'd9,5'd16,5'd5,5'd5,5'd9,5'd8,5'd1,5'd10,5'd6,5'd4,5'd11,5'd5,5'd6,5'd5,5'd8,5'd3,5'd10,5'd6}
`define RECTANGLE2_Y1 {5'd1,5'd17,5'd2,5'd19,5'd19,5'd19,5'd19,5'd14,5'd16,5'd19,5'd19,5'd6,5'd19,5'd12,5'd12,5'd20,5'd16,5'd18,5'd14,5'd13,5'd13,5'd13,5'd13,5'd8,5'd15,5'd15,5'd15,5'd13,5'd13,5'd13,5'd13,5'd8,5'd8,5'd0,5'd20,5'd1,5'd1,5'd0,5'd14,5'd13,5'd9,5'd11,5'd1,5'd0,5'd0,5'd9,5'd9,5'd2,5'd13,5'd1,5'd2,5'd14,5'd14,5'd5,5'd6,5'd6,5'd8,5'd8,5'd5,5'd11,5'd17,5'd20,5'd19,5'd17,5'd18,5'd17,5'd4,5'd8,5'd8,5'd9,5'd7,5'd7,5'd7,5'd5,5'd9,5'd16,5'd4,5'd3,5'd4,5'd0,5'd6,5'd5,5'd0,5'd1,5'd9,5'd10,5'd9,5'd13,5'd12,5'd2,5'd2,5'd13,5'd13,5'd10,5'd13,5'd10,5'd10,5'd14,5'd12,5'd13,5'd12,5'd3,5'd3,5'd0,5'd6,5'd6,5'd15,5'd12,5'd12,5'd15,5'd12,5'd8,5'd8,5'd4,5'd5,5'd11,5'd12,5'd14,5'd14,5'd4,5'd4,5'd3,5'd12,5'd2,5'd5,5'd6,5'd5,5'd19,5'd19,5'd16,5'd16,5'd16,5'd16,5'd0,5'd0,5'd16,5'd16,5'd20,5'd18,5'd21,5'd22,5'd6,5'd6,5'd6,5'd0,5'd2,5'd8,5'd7,5'd7,5'd11,5'd11,5'd11,5'd7,5'd9,5'd4,5'd6,5'd9,5'd11,5'd17,5'd17,5'd12,5'd11,5'd11,5'd7,5'd7,5'd4,5'd3,5'd5,5'd5,5'd3,5'd3,5'd0,5'd1,5'd8,5'd12,5'd15,5'd19,5'd13,5'd2,5'd6,5'd11,5'd20,5'd16,5'd13,5'd6,5'd14,5'd14,5'd6,5'd6,5'd2,5'd4,5'd9,5'd12,5'd16,5'd18,5'd14,5'd16,5'd1,5'd5,5'd7,5'd7,5'd1,5'd2,5'd16,5'd15,5'd5,5'd4,5'd7,5'd0,5'd6,5'd2,5'd2,5'd0,5'd0,5'd0,5'd0,5'd8,5'd8,5'd4,5'd9,5'd2,5'd8,5'd8,5'd7,5'd8,5'd9,5'd19,5'd19,5'd0,5'd0,5'd0,5'd7,5'd7,5'd7,5'd0,5'd0,5'd1,5'd11,5'd7,5'd19,5'd6,5'd6,5'd3,5'd2,5'd17,5'd2,5'd8,5'd6,5'd3,5'd6,5'd6,5'd20,5'd8,5'd8,5'd3,5'd2,5'd1,5'd2,5'd2,5'd9,5'd10,5'd10,5'd13,5'd13,5'd2,5'd10,5'd8,5'd8,5'd7,5'd6,5'd6,5'd6,5'd13,5'd0,5'd19,5'd6,5'd1,5'd9,5'd15,5'd7,5'd14,5'd10,5'd12,5'd12,5'd16,5'd19,5'd14,5'd15,5'd13,5'd13,5'd4,5'd10,5'd1,5'd1,5'd4,5'd12,5'd6,5'd10,5'd15,5'd0,5'd1,5'd7,5'd8,5'd8,5'd9,5'd14,5'd4,5'd0,5'd0,5'd0,5'd4,5'd18,5'd18,5'd6,5'd7,5'd7,5'd16,5'd4,5'd0,5'd19,5'd12,5'd8,5'd9,5'd5,5'd6,5'd8,5'd12,5'd1,5'd0,5'd0,5'd14,5'd14,5'd6,5'd7,5'd11,5'd0,5'd0,5'd6,5'd0,5'd7,5'd9,5'd0,5'd16,5'd2,5'd3,5'd19,5'd13,5'd9,5'd17,5'd13,5'd0,5'd0,5'd7,5'd7,5'd6,5'd0,5'd1,5'd11,5'd2,5'd6,5'd1,5'd1,5'd2,5'd1,5'd15,5'd15,5'd15,5'd15,5'd4,5'd4,5'd9,5'd0,5'd3,5'd9,5'd6,5'd3,5'd1,5'd1,5'd20,5'd20,5'd6,5'd7,5'd8,5'd20,5'd17,5'd8,5'd2,5'd15,5'd20,5'd17,5'd17,5'd15,5'd18,5'd18,5'd5,5'd11,5'd11,5'd11,5'd1,5'd9,5'd14,5'd7,5'd0,5'd12,5'd0,5'd1,5'd20,5'd14,5'd1,5'd6,5'd3,5'd0,5'd4,5'd9,5'd6,5'd6,5'd9,5'd22,5'd1,5'd0,5'd0,5'd1,5'd15,5'd10,5'd10,5'd15,5'd15,5'd6,5'd17,5'd7,5'd7,5'd11,5'd0,5'd5,5'd1,5'd4,5'd7,5'd8,5'd17,5'd4,5'd17,5'd3,5'd17,5'd14,5'd17,5'd15,5'd12,5'd7,5'd7,5'd9,5'd9,5'd10,5'd0,5'd17,5'd17,5'd13,5'd13,5'd1,5'd13,5'd13,5'd13,5'd5,5'd10,5'd8,5'd4,5'd4,5'd5,5'd10,5'd14,5'd14,5'd12,5'd5,5'd10,5'd8,5'd9,5'd6,5'd6,5'd11,5'd11,5'd8,5'd10,5'd1,5'd16,5'd1,5'd1,5'd18,5'd19,5'd12,5'd11,5'd17,5'd4,5'd22,5'd20,5'd14,5'd9,5'd11,5'd8,5'd8,5'd8,5'd12,5'd2,5'd5,5'd7,5'd0,5'd0,5'd1,5'd8,5'd6,5'd9,5'd2,5'd5,5'd0,5'd0,5'd17,5'd15,5'd20,5'd8,5'd6,5'd2,5'd4,5'd13,5'd5,5'd2,5'd7,5'd7,5'd12,5'd6,5'd10,5'd10,5'd1,5'd1,5'd10,5'd19,5'd10,5'd1,5'd11,5'd0,5'd13,5'd2,5'd2,5'd11,5'd19,5'd7,5'd4,5'd4,5'd13,5'd13,5'd16,5'd5,5'd6,5'd5,5'd12,5'd12,5'd0,5'd0,5'd1,5'd0,5'd9,5'd4,5'd9,5'd9,5'd9,5'd6,5'd20,5'd0,5'd2,5'd2,5'd17,5'd17,5'd20,5'd20,5'd20,5'd17,5'd9,5'd9,5'd6,5'd8,5'd17,5'd9,5'd10,5'd14,5'd19,5'd17,5'd18,5'd18,5'd6,5'd10,5'd12,5'd18,5'd1,5'd13,5'd11,5'd9,5'd5,5'd9,5'd17,5'd2,5'd8,5'd8,5'd22,5'd6,5'd12,5'd16,5'd0,5'd0,5'd6,5'd3,5'd10,5'd1,5'd11,5'd12,5'd2,5'd15,5'd3,5'd4,5'd19,5'd20,5'd20,5'd15,5'd15,5'd12,5'd12,5'd10,5'd10,5'd6,5'd16,5'd12,5'd3,5'd11,5'd8,5'd8,5'd0,5'd6,5'd12,5'd12,5'd16,5'd0,5'd2,5'd14,5'd9,5'd8,5'd11,5'd10,5'd10,5'd8,5'd10,5'd20,5'd5,5'd11,5'd9,5'd9,5'd10,5'd0,5'd15,5'd15,5'd14,5'd16,5'd16,5'd16,5'd18,5'd10,5'd14,5'd14,5'd10,5'd1,5'd1,5'd0,5'd10,5'd0,5'd8,5'd7,5'd9,5'd0,5'd0,5'd4,5'd0,5'd2,5'd2,5'd6,5'd5,5'd0,5'd0,5'd4,5'd0,5'd5,5'd5,5'd1,5'd1,5'd17,5'd17,5'd18,5'd19,5'd19,5'd4,5'd11,5'd18,5'd19,5'd10,5'd3,5'd11,5'd11,5'd8,5'd6,5'd8,5'd8,5'd8,5'd8,5'd8,5'd5,5'd18,5'd11,5'd16,5'd17,5'd4,5'd8,5'd4,5'd21,5'd21,5'd14,5'd14,5'd9,5'd7,5'd3,5'd0,5'd17,5'd17,5'd0,5'd4,5'd2,5'd7,5'd4,5'd0,5'd2,5'd11,5'd10,5'd5,5'd6,5'd8,5'd8,5'd16,5'd9,5'd5,5'd6,5'd3,5'd6,5'd18,5'd14,5'd14,5'd12,5'd6,5'd8,5'd1,5'd12,5'd18,5'd15,5'd2,5'd2,5'd2,5'd2,5'd4,5'd4,5'd2,5'd6,5'd20,5'd7,5'd7,5'd1,5'd6,5'd0,5'd0,5'd6,5'd6,5'd3,5'd14,5'd2,5'd2,5'd1,5'd1,5'd3,5'd12,5'd14,5'd19,5'd15,5'd15,5'd15,5'd23,5'd18,5'd6,5'd11,5'd1,5'd3,5'd7,5'd7,5'd14,5'd14,5'd8,5'd8,5'd12,5'd12,5'd12,5'd12,5'd20,5'd4,5'd19,5'd19,5'd16,5'd1,5'd1,5'd8,5'd6,5'd2,5'd9,5'd11,5'd16,5'd14,5'd3,5'd5,5'd0,5'd16,5'd4,5'd9,5'd1,5'd1,5'd6,5'd5,5'd11,5'd7,5'd16,5'd0,5'd4,5'd4,5'd4,5'd4,5'd16,5'd9,5'd1,5'd1,5'd0,5'd1,5'd16,5'd1,5'd21,5'd1,5'd14,5'd14,5'd6,5'd2,5'd10,5'd10,5'd12,5'd19,5'd10,5'd17,5'd18,5'd18,5'd19,5'd19,5'd18,5'd4,5'd3,5'd3,5'd0,5'd0,5'd5,5'd5,5'd0,5'd0,5'd8,5'd7,5'd10,5'd7,5'd1,5'd1,5'd12,5'd10,5'd14,5'd1,5'd0,5'd0,5'd6,5'd14,5'd19,5'd8,5'd10,5'd7,5'd7,5'd14,5'd13,5'd3,5'd6,5'd1,5'd8,5'd5,5'd0,5'd19,5'd10,5'd3,5'd16,5'd22,5'd7,5'd2,5'd2,5'd3,5'd3,5'd17,5'd1,5'd1,5'd0,5'd4,5'd6,5'd7,5'd4,5'd4,5'd5,5'd5,5'd8,5'd10,5'd10,5'd2,5'd19,5'd9,5'd4,5'd2,5'd19,5'd20,5'd21,5'd21,5'd18,5'd5,5'd16,5'd16,5'd17,5'd17,5'd15,5'd9,5'd11,5'd11,5'd15,5'd18,5'd18,5'd11,5'd11,5'd1,5'd5,5'd1,5'd5,5'd6,5'd0,5'd8,5'd1,5'd16,5'd20,5'd17,5'd18,5'd1,5'd13,5'd1,5'd5,5'd5,5'd0,5'd0,5'd6,5'd6,5'd5,5'd18,5'd19,5'd6,5'd8,5'd8,5'd15,5'd16,5'd1,5'd7,5'd2,5'd2,5'd0,5'd0,5'd18,5'd11,5'd20,5'd4,5'd10,5'd0,5'd16,5'd12,5'd5,5'd7,5'd1,5'd10,5'd15,5'd10,5'd12,5'd12,5'd12,5'd12,5'd12,5'd9,5'd10,5'd10,5'd8,5'd17,5'd17,5'd12,5'd12,5'd14,5'd14,5'd8,5'd9,5'd8,5'd13,5'd2,5'd13,5'd13,5'd3,5'd4,5'd0,5'd0,5'd0,5'd7,5'd4,5'd5,5'd9,5'd9,5'd0,5'd9,5'd6,5'd13,5'd15,5'd8,5'd3,5'd4,5'd12,5'd3,5'd0,5'd19,5'd20,5'd20,5'd6,5'd2,5'd3,5'd0,5'd1,5'd14,5'd15,5'd0,5'd6,5'd11,5'd0,5'd8,5'd7,5'd10,5'd16,5'd10,5'd11,5'd11,5'd10,5'd0,5'd1,5'd1,5'd8,5'd8,5'd0,5'd0,5'd2,5'd2,5'd0,5'd0,5'd12,5'd0,5'd3,5'd9,5'd10,5'd10,5'd13,5'd6,5'd6,5'd17,5'd10,5'd14,5'd12,5'd0,5'd8,5'd5,5'd10,5'd4,5'd7,5'd5,5'd9,5'd6,5'd7,5'd6,5'd18,5'd18,5'd15,5'd8,5'd18,5'd19,5'd20,5'd18,5'd0,5'd8,5'd1,5'd6,5'd3,5'd7,5'd2,5'd2,5'd2,5'd4,5'd8,5'd3,5'd3,5'd6,5'd15,5'd15,5'd22,5'd15,5'd19,5'd19,5'd0,5'd5,5'd2,5'd3,5'd4,5'd7,5'd3,5'd9,5'd12,5'd12,5'd0,5'd17,5'd3,5'd0,5'd18,5'd16,5'd16,5'd16,5'd4,5'd4,5'd17,5'd19,5'd0,5'd0,5'd6,5'd6,5'd7,5'd15,5'd10,5'd6,5'd0,5'd20,5'd16,5'd2,5'd6,5'd10,5'd22,5'd16,5'd6,5'd16,5'd2,5'd8,5'd10,5'd15,5'd10,5'd5,5'd3,5'd16,5'd1,5'd1,5'd0,5'd0,5'd18,5'd0,5'd0,5'd6,5'd6,5'd1,5'd0,5'd21,5'd14,5'd11,5'd0,5'd0,5'd3,5'd0,5'd12,5'd7,5'd15,5'd1,5'd12,5'd12,5'd19,5'd18,5'd11,5'd15,5'd2,5'd2,5'd18,5'd20,5'd9,5'd13,5'd13,5'd18,5'd20,5'd18,5'd6,5'd7,5'd13,5'd13,5'd13,5'd6,5'd0,5'd4,5'd18,5'd10,5'd15,5'd12,5'd2,5'd2,5'd4,5'd0,5'd19,5'd14,5'd14,5'd3,5'd7,5'd2,5'd1,5'd0,5'd0,5'd7,5'd11,5'd4,5'd9,5'd8,5'd4,5'd2,5'd2,5'd7,5'd11,5'd9,5'd10,5'd15,5'd18,5'd1,5'd1,5'd3,5'd7,5'd7,5'd11,5'd3,5'd22,5'd13,5'd7,5'd0,5'd13,5'd15,5'd0,5'd2,5'd0,5'd10,5'd5,5'd21,5'd21,5'd6,5'd4,5'd9,5'd9,5'd7,5'd13,5'd5,5'd5,5'd6,5'd5,5'd1,5'd1,5'd0,5'd7,5'd1,5'd21,5'd13,5'd2,5'd0,5'd0,5'd10,5'd23,5'd1,5'd3,5'd0,5'd10,5'd10,5'd12,5'd8,5'd9,5'd9,5'd9,5'd8,5'd7,5'd5,5'd9,5'd2,5'd17,5'd13,5'd18,5'd14,5'd13,5'd18,5'd18,5'd19,5'd19,5'd6,5'd5,5'd2,5'd19,5'd18,5'd17,5'd8,5'd19,5'd17,5'd9,5'd6,5'd11,5'd0,5'd0,5'd8,5'd16,5'd3,5'd2,5'd1,5'd3,5'd3,5'd3,5'd6,5'd2,5'd3,5'd5,5'd6,5'd9,5'd19,5'd7,5'd4,5'd1,5'd13,5'd4,5'd11,5'd4,5'd8,5'd18,5'd3,5'd6,5'd11,5'd0,5'd7,5'd5,5'd5,5'd4,5'd5,5'd1,5'd1,5'd4,5'd4,5'd4,5'd4,5'd4,5'd1,5'd5,5'd5,5'd19,5'd5,5'd7,5'd5,5'd12,5'd13,5'd2,5'd18,5'd12,5'd11,5'd7,5'd4,5'd9,5'd6,5'd8,5'd11,5'd15,5'd15,5'd4,5'd15,5'd13,5'd14,5'd15,5'd15,5'd8,5'd8,5'd11,5'd11,5'd11,5'd22,5'd3,5'd8,5'd2,5'd3,5'd2,5'd2,5'd2,5'd18,5'd16,5'd17,5'd8,5'd8,5'd4,5'd4,5'd2,5'd4,5'd14,5'd10,5'd5,5'd1,5'd10,5'd10,5'd8,5'd10,5'd9,5'd9,5'd6,5'd6,5'd16,5'd12,5'd16,5'd16,5'd10,5'd0,5'd1,5'd2,5'd19,5'd14,5'd6,5'd6,5'd3,5'd3,5'd20,5'd17,5'd4,5'd0,5'd0,5'd0,5'd3,5'd10,5'd15,5'd3,5'd0,5'd1,5'd7,5'd2,5'd18,5'd2,5'd7,5'd0,5'd6,5'd13,5'd7,5'd7,5'd18,5'd10,5'd18,5'd16,5'd17,5'd18,5'd1,5'd20,5'd21,5'd1,5'd18,5'd18,5'd18,5'd14,5'd7,5'd7,5'd9,5'd8,5'd14,5'd14,5'd14,5'd18,5'd7,5'd18,5'd9,5'd0,5'd6,5'd11,5'd13,5'd13,5'd9,5'd19,5'd4,5'd4,5'd0,5'd4,5'd11,5'd5,5'd12,5'd20,5'd7,5'd3,5'd15,5'd0,5'd7,5'd10,5'd2,5'd4,5'd21,5'd12,5'd0,5'd12,5'd12,5'd11,5'd1,5'd4,5'd19,5'd6,5'd8,5'd11,5'd11,5'd3,5'd3,5'd5,5'd5,5'd5,5'd5,5'd6,5'd6,5'd12,5'd12,5'd7,5'd6,5'd9,5'd4,5'd8,5'd15,5'd9,5'd16,5'd9,5'd10,5'd15,5'd18,5'd16,5'd0,5'd5,5'd3,5'd19,5'd17,5'd13,5'd13,5'd12,5'd0,5'd7,5'd12,5'd7,5'd13,5'd7,5'd14,5'd14,5'd7,5'd7,5'd7,5'd12,5'd22,5'd18,5'd13,5'd14,5'd13,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd2,5'd15,5'd12,5'd7,5'd10,5'd10,5'd8,5'd8,5'd1,5'd2,5'd0,5'd0,5'd9,5'd18,5'd18,5'd1,5'd0,5'd16,5'd16,5'd17,5'd12,5'd10,5'd10,5'd10,5'd7,5'd9,5'd12,5'd17,5'd16,5'd6,5'd6,5'd18,5'd9,5'd14,5'd9,5'd12,5'd5,5'd10,5'd8,5'd8,5'd7,5'd6,5'd5,5'd8,5'd0,5'd8,5'd7,5'd8,5'd16,5'd16,5'd17,5'd16,5'd18,5'd19,5'd0,5'd0,5'd0,5'd6,5'd2,5'd8,5'd10,5'd6,5'd3,5'd10,5'd11,5'd3,5'd1,5'd0,5'd2,5'd2,5'd0,5'd0,5'd5,5'd8,5'd10,5'd1,5'd7,5'd0,5'd0,5'd0,5'd4,5'd17,5'd10,5'd4,5'd6,5'd6,5'd11,5'd21,5'd14,5'd1,5'd7,5'd9,5'd19,5'd13,5'd3,5'd5,5'd5,5'd12,5'd2,5'd10,5'd7,5'd18,5'd1,5'd0,5'd9,5'd22,5'd6,5'd17,5'd8,5'd0,5'd0,5'd17,5'd17,5'd14,5'd14,5'd11,5'd14,5'd8,5'd8,5'd0,5'd6,5'd5,5'd5,5'd8,5'd8,5'd20,5'd18,5'd18,5'd8,5'd13,5'd4,5'd9,5'd17,5'd10,5'd15,5'd8,5'd7,5'd13,5'd2,5'd0,5'd0,5'd0,5'd0,5'd2,5'd5,5'd11,5'd11,5'd5,5'd7,5'd12,5'd1,5'd13,5'd4,5'd5,5'd5,5'd16,5'd6,5'd5,5'd19,5'd3,5'd8,5'd6,5'd19,5'd20,5'd6,5'd0,5'd0,5'd8,5'd11,5'd8,5'd6,5'd11,5'd2,5'd13,5'd0,5'd2,5'd5,5'd2,5'd2,5'd15,5'd2,5'd2,5'd1,5'd17,5'd17,5'd18,5'd18,5'd15,5'd15,5'd13,5'd6,5'd6,5'd8,5'd3,5'd15,5'd10,5'd13,5'd6,5'd8,5'd5,5'd16,5'd5,5'd6,5'd5,5'd5,5'd21,5'd15,5'd0,5'd18,5'd4,5'd0,5'd2,5'd2,5'd8,5'd8,5'd5,5'd5,5'd17,5'd17,5'd11,5'd0,5'd16,5'd23,5'd7,5'd11,5'd1,5'd7,5'd0,5'd11,5'd14,5'd3,5'd4,5'd5,5'd9,5'd11,5'd15,5'd1,5'd2,5'd4,5'd8,5'd0,5'd16,5'd16,5'd4,5'd5,5'd12,5'd1,5'd19,5'd19,5'd8,5'd15,5'd7,5'd8,5'd4,5'd7,5'd9,5'd9,5'd15,5'd19,5'd16,5'd7,5'd15,5'd10,5'd10,5'd8,5'd10,5'd13,5'd22,5'd16,5'd16,5'd2,5'd1,5'd19,5'd18,5'd19,5'd19,5'd19,5'd8,5'd5,5'd9,5'd11,5'd7,5'd2,5'd12,5'd12,5'd15,5'd6,5'd2,5'd15,5'd1,5'd1,5'd5,5'd13,5'd8,5'd8,5'd3,5'd3,5'd7,5'd7,5'd0,5'd5,5'd3,5'd0,5'd3,5'd1,5'd18,5'd18,5'd1,5'd1,5'd6,5'd6,5'd3,5'd17,5'd16,5'd13,5'd1,5'd17,5'd14,5'd6,5'd10,5'd10,5'd3,5'd3,5'd0,5'd1,5'd14,5'd14,5'd5,5'd0,5'd0,5'd12,5'd11,5'd10,5'd0,5'd8,5'd20,5'd12,5'd11,5'd11,5'd0,5'd0,5'd3,5'd3,5'd16,5'd18,5'd8,5'd11,5'd6,5'd3,5'd1,5'd4,5'd12,5'd2,5'd11,5'd17,5'd8,5'd8,5'd19,5'd8,5'd18,5'd6,5'd1,5'd9,5'd7,5'd16,5'd16,5'd0,5'd9,5'd5,5'd9,5'd4,5'd4,5'd12,5'd11,5'd11,5'd16,5'd12,5'd6,5'd12,5'd4,5'd0,5'd10,5'd18,5'd10,5'd10,5'd6,5'd5,5'd5,5'd0,5'd16,5'd8,5'd15,5'd16,5'd5,5'd11,5'd16,5'd14,5'd11,5'd11,5'd20,5'd14,5'd1,5'd0,5'd0,5'd12,5'd11,5'd14,5'd14,5'd9,5'd5,5'd7,5'd11,5'd6,5'd12,5'd13,5'd8,5'd5,5'd19,5'd19,5'd2,5'd6,5'd4,5'd5,5'd9,5'd6,5'd3,5'd12,5'd4,5'd7,5'd7,5'd4,5'd9,5'd5,5'd17,5'd5,5'd17,5'd1,5'd1,5'd0,5'd5,5'd0,5'd18,5'd6,5'd11,5'd14,5'd16,5'd7,5'd16,5'd11,5'd11,5'd6,5'd6,5'd0,5'd4,5'd10,5'd0,5'd13,5'd11,5'd14,5'd16,5'd8,5'd7,5'd11,5'd9,5'd3,5'd21,5'd12,5'd11,5'd0,5'd7,5'd6,5'd2,5'd7,5'd20,5'd12,5'd8,5'd16,5'd12,5'd14,5'd3,5'd13,5'd5,5'd16,5'd15,5'd18,5'd1,5'd2,5'd2,5'd3,5'd7,5'd18,5'd0,5'd1,5'd20,5'd3,5'd0,5'd8,5'd0,5'd11,5'd10,5'd9,5'd11,5'd10,5'd2,5'd7,5'd21,5'd4,5'd6,5'd18,5'd16,5'd6,5'd18,5'd19,5'd17,5'd20,5'd21,5'd12,5'd10,5'd11,5'd10,5'd10,5'd4,5'd0,5'd5,5'd2,5'd4,5'd13,5'd7,5'd10,5'd3,5'd0,5'd0,5'd6,5'd11,5'd11,5'd8,5'd8,5'd13,5'd11,5'd9,5'd9,5'd5,5'd12,5'd12,5'd6,5'd8,5'd18,5'd17,5'd17,5'd17,5'd0,5'd5,5'd3,5'd11,5'd11,5'd18,5'd18,5'd17,5'd10,5'd8,5'd19,5'd0,5'd4,5'd2,5'd11,5'd0,5'd10,5'd14,5'd16,5'd9,5'd10,5'd13,5'd19,5'd16,5'd3,5'd5,5'd13,5'd6,5'd5,5'd6,5'd6,5'd9,5'd9,5'd12,5'd0,5'd9,5'd16,5'd17,5'd13,5'd17,5'd17,5'd4,5'd5,5'd5,5'd5,5'd0,5'd9,5'd6,5'd7,5'd11,5'd8,5'd6,5'd7,5'd12,5'd12,5'd16,5'd17,5'd3,5'd0,5'd1,5'd10,5'd23,5'd11,5'd0,5'd0,5'd11,5'd3,5'd4,5'd20,5'd11,5'd11,5'd14,5'd11,5'd1,5'd3,5'd3,5'd12,5'd12,5'd5,5'd5,5'd6,5'd6,5'd5,5'd14,5'd14,5'd19,5'd3,5'd0,5'd7,5'd2,5'd3,5'd0,5'd2,5'd10,5'd19,5'd2,5'd8,5'd13,5'd7,5'd4,5'd5,5'd5,5'd21,5'd6,5'd9,5'd11,5'd14,5'd14,5'd5,5'd9,5'd11,5'd5,5'd2,5'd2,5'd20,5'd20,5'd4,5'd4,5'd4,5'd4,5'd2,5'd2,5'd10,5'd10,5'd4,5'd4,5'd5,5'd6,5'd10,5'd9,5'd8,5'd4,5'd10,5'd22,5'd6,5'd5,5'd8,5'd5,5'd11,5'd10,5'd0,5'd0,5'd6,5'd3,5'd20,5'd19,5'd2,5'd8,5'd8,5'd14,5'd15,5'd18,5'd17,5'd3,5'd11,5'd2,5'd0,5'd20,5'd5,5'd10,5'd12,5'd8,5'd6,5'd3,5'd2,5'd17,5'd7,5'd20,5'd1,5'd7,5'd0,5'd0,5'd17,5'd8,5'd11,5'd11,5'd14,5'd11,5'd20,5'd11,5'd0,5'd12,5'd2,5'd0,5'd6,5'd19,5'd16,5'd5,5'd10,5'd0,5'd3,5'd16,5'd16,5'd2,5'd12,5'd14,5'd15,5'd3,5'd6,5'd7,5'd13,5'd0,5'd3,5'd6,5'd6,5'd7,5'd6,5'd2,5'd2,5'd12,5'd12,5'd8,5'd8,5'd11,5'd19,5'd0,5'd0,5'd4,5'd4,5'd11,5'd15,5'd1,5'd1,5'd5,5'd5,5'd6,5'd11,5'd13,5'd16,5'd15,5'd17,5'd12,5'd5,5'd1,5'd1,5'd7,5'd17,5'd10,5'd10,5'd9,5'd10,5'd2,5'd1,5'd5,5'd13,5'd1,5'd4,5'd5,5'd3,5'd10,5'd1,5'd6,5'd7,5'd3,5'd2,5'd6,5'd0,5'd12,5'd8,5'd0,5'd0,5'd11,5'd3,5'd0,5'd0,5'd0,5'd0,5'd6,5'd6,5'd20,5'd17,5'd18,5'd3,5'd11,5'd11,5'd20,5'd20,5'd14,5'd20,5'd19,5'd7,5'd12,5'd7,5'd5,5'd8,5'd21,5'd12,5'd0,5'd6,5'd3,5'd8,5'd8,5'd8,5'd2,5'd0,5'd17,5'd6,5'd13,5'd7,5'd7,5'd3,5'd0,5'd6,5'd5,5'd6,5'd2,5'd2,5'd2,5'd7,5'd0,5'd15,5'd5,5'd7,5'd7,5'd0,5'd0,5'd14,5'd5,5'd4,5'd0,5'd18,5'd17,5'd15,5'd15,5'd18,5'd1,5'd0,5'd0,5'd9,5'd8,5'd7,5'd11,5'd13,5'd0,5'd20,5'd2,5'd16,5'd11,5'd15,5'd0,5'd1,5'd6,5'd6,5'd12,5'd18,5'd18,5'd0,5'd0,5'd17,5'd9,5'd11,5'd11,5'd17,5'd17,5'd23,5'd6,5'd7,5'd7,5'd8,5'd7,5'd12,5'd3,5'd8,5'd17,5'd0,5'd0,5'd2,5'd14,5'd20,5'd2,5'd7,5'd7,5'd16,5'd4,5'd18,5'd4,5'd1,5'd6,5'd11,5'd11,5'd2,5'd5,5'd8,5'd1,5'd15,5'd8,5'd6,5'd7,5'd11,5'd6,5'd3,5'd13,5'd19,5'd4,5'd16,5'd14,5'd8,5'd15,5'd7,5'd17,5'd17,5'd6,5'd11,5'd1,5'd17,5'd10,5'd6,5'd4,5'd7,5'd9,5'd17,5'd1,5'd1,5'd0,5'd17,5'd14,5'd15,5'd14,5'd14,5'd12,5'd12,5'd0,5'd0,5'd4,5'd7,5'd0,5'd6,5'd13,5'd16,5'd22,5'd12,5'd1,5'd1,5'd12,5'd14,5'd13,5'd8,5'd5,5'd14,5'd8,5'd14,5'd0,5'd0,5'd2,5'd11,5'd5,5'd5,5'd20,5'd5,5'd6,5'd6,5'd9,5'd6,5'd6,5'd14,5'd4,5'd7,5'd14,5'd13,5'd14,5'd12,5'd6,5'd7,5'd2,5'd14,5'd22,5'd19,5'd2,5'd5,5'd3,5'd19,5'd1,5'd3,5'd4,5'd4,5'd0,5'd19,5'd18,5'd13,5'd17,5'd19,5'd10,5'd4,5'd3,5'd3,5'd0,5'd0,5'd7,5'd7,5'd15,5'd15,5'd14,5'd11,5'd11,5'd12,5'd0,5'd0,5'd0,5'd9,5'd6,5'd7,5'd0,5'd10,5'd16,5'd16,5'd10,5'd10,5'd0,5'd3,5'd6,5'd2,5'd4,5'd8,5'd10,5'd7,5'd6,5'd20,5'd2,5'd2,5'd0,5'd1,5'd14,5'd14,5'd16,5'd16,5'd1,5'd11,5'd17,5'd8,5'd2,5'd8,5'd14,5'd2,5'd1,5'd11,5'd3,5'd17,5'd15,5'd8,5'd7,5'd7,5'd21,5'd0,5'd3,5'd1,5'd2,5'd14,5'd20,5'd7,5'd0,5'd0,5'd6,5'd16,5'd11,5'd7,5'd6,5'd9,5'd14,5'd8,5'd6,5'd15,5'd20,5'd18,5'd18,5'd19,5'd7,5'd6,5'd0,5'd0,5'd4,5'd0,5'd5,5'd8,5'd16,5'd6,5'd10,5'd7,5'd1,5'd7,5'd12,5'd12,5'd11,5'd3,5'd2,5'd5,5'd1,5'd12,5'd0,5'd23,5'd1,5'd0,5'd19,5'd3,5'd4,5'd13,5'd5,5'd11,5'd2,5'd18,5'd4,5'd19,5'd16,5'd16,5'd6,5'd1,5'd1,5'd0,5'd0,5'd0,5'd4,5'd13,5'd12,5'd11,5'd11,5'd11,5'd11,5'd11,5'd5,5'd3,5'd20,5'd0,5'd0,5'd1,5'd0,5'd3,5'd0,5'd0,5'd15,5'd10,5'd14,5'd14,5'd15,5'd8,5'd8,5'd6,5'd14,5'd17,5'd13,5'd12,5'd7,5'd0,5'd0,5'd1,5'd1,5'd5,5'd4,5'd12,5'd20,5'd5,5'd10,5'd2,5'd5,5'd16,5'd16,5'd12,5'd11,5'd8,5'd3,5'd1,5'd6,5'd0,5'd19,5'd17,5'd15,5'd5,5'd5,5'd6,5'd0,5'd9,5'd11,5'd19,5'd8,5'd18,5'd16,5'd0,5'd0,5'd8,5'd8,5'd10,5'd0,5'd12,5'd16,5'd4,5'd4,5'd4,5'd17,5'd2,5'd19,5'd16,5'd8,5'd12,5'd12,5'd23,5'd18,5'd6,5'd6,5'd13,5'd6,5'd20,5'd6,5'd11,5'd0,5'd3,5'd8,5'd6,5'd6,5'd0,5'd6,5'd3,5'd0,5'd5,5'd6,5'd17,5'd17,5'd17,5'd12,5'd5,5'd1,5'd1,5'd10,5'd18,5'd17,5'd13,5'd8,5'd12,5'd14,5'd11,5'd1,5'd3,5'd3,5'd17,5'd12,5'd1,5'd5,5'd7,5'd7,5'd13,5'd11,5'd5,5'd1,5'd1,5'd7,5'd1,5'd3,5'd4,5'd5,5'd2,5'd1,5'd13,5'd1,5'd16,5'd6,5'd8,5'd1,5'd1,5'd8,5'd21,5'd12,5'd5,5'd13,5'd11,5'd3,5'd13,5'd20,5'd6,5'd6,5'd0,5'd5,5'd8,5'd5,5'd11,5'd3,5'd11,5'd14,5'd2,5'd12,5'd4,5'd8,5'd3,5'd19,5'd11,5'd13,5'd5,5'd20,5'd12,5'd4,5'd7}
`define RECTANGLE2_X2 {5'd15,5'd24,5'd18,5'd12,5'd21,5'd9,5'd24,5'd18,5'd22,5'd18,5'd24,5'd12,5'd24,5'd3,5'd24,5'd18,5'd12,5'd11,5'd21,5'd11,5'd21,5'd20,5'd22,5'd13,5'd21,5'd18,5'd22,5'd9,5'd19,5'd6,5'd23,5'd4,5'd24,5'd7,5'd21,5'd6,5'd21,5'd5,5'd15,5'd15,5'd24,5'd18,5'd13,5'd10,5'd16,5'd14,5'd22,5'd16,5'd22,5'd21,5'd14,5'd10,5'd16,5'd13,5'd14,5'd11,5'd12,5'd14,5'd23,5'd16,5'd16,5'd12,5'd18,5'd18,5'd23,5'd11,5'd24,5'd14,5'd23,5'd17,5'd17,5'd18,5'd20,5'd18,5'd16,5'd15,5'd24,5'd19,5'd15,5'd12,5'd14,5'd15,5'd14,5'd18,5'd23,5'd10,5'd22,5'd7,5'd13,5'd12,5'd13,5'd9,5'd21,5'd15,5'd24,5'd6,5'd21,5'd14,5'd18,5'd20,5'd16,5'd12,5'd18,5'd14,5'd24,5'd18,5'd24,5'd12,5'd15,5'd18,5'd15,5'd9,5'd24,5'd12,5'd18,5'd11,5'd15,5'd7,5'd21,5'd8,5'd17,5'd16,5'd12,5'd19,5'd23,5'd12,5'd21,5'd18,5'd23,5'd10,5'd24,5'd9,5'd24,5'd5,5'd24,5'd7,5'd22,5'd16,5'd24,5'd9,5'd21,5'd3,5'd23,5'd10,5'd21,5'd10,5'd24,5'd10,5'd24,5'd6,5'd24,5'd23,5'd24,5'd10,5'd18,5'd11,5'd24,5'd13,5'd24,5'd18,5'd14,5'd15,5'd14,5'd7,5'd24,5'd18,5'd23,5'd14,5'd14,5'd4,5'd22,5'd7,5'd24,5'd17,5'd23,5'd15,5'd15,5'd13,5'd22,5'd4,5'd23,5'd20,5'd16,5'd11,5'd20,5'd8,5'd21,5'd12,5'd13,5'd10,5'd24,5'd15,5'd18,5'd10,5'd21,5'd15,5'd18,5'd9,5'd14,5'd18,5'd12,5'd24,5'd12,5'd17,5'd10,5'd21,5'd12,5'd15,5'd15,5'd13,5'd8,5'd20,5'd7,5'd19,5'd4,5'd22,5'd6,5'd21,5'd10,5'd17,5'd14,5'd24,5'd21,5'd22,5'd16,5'd22,5'd20,5'd15,5'd7,5'd18,5'd18,5'd15,5'd14,5'd22,5'd9,5'd16,5'd13,5'd16,5'd10,5'd23,5'd7,5'd17,5'd12,5'd14,5'd14,5'd14,5'd15,5'd13,5'd12,5'd15,5'd12,5'd19,5'd4,5'd22,5'd3,5'd22,5'd9,5'd16,5'd13,5'd24,5'd8,5'd24,5'd18,5'd23,5'd6,5'd22,5'd10,5'd21,5'd13,5'd13,5'd5,5'd19,5'd10,5'd20,5'd19,5'd13,5'd12,5'd23,5'd12,5'd15,5'd14,5'd18,5'd9,5'd24,5'd8,5'd14,5'd8,5'd14,5'd17,5'd14,5'd14,5'd15,5'd4,5'd21,5'd2,5'd19,5'd10,5'd18,5'd3,5'd20,5'd8,5'd22,5'd6,5'd24,5'd12,5'd24,5'd13,5'd20,5'd12,5'd20,5'd6,5'd21,5'd18,5'd16,5'd11,5'd18,5'd15,5'd23,5'd13,5'd19,5'd12,5'd12,5'd11,5'd18,5'd13,5'd22,5'd19,5'd12,5'd9,5'd19,5'd5,5'd23,5'd12,5'd14,5'd14,5'd16,5'd9,5'd14,5'd12,5'd15,5'd17,5'd13,5'd18,5'd24,5'd9,5'd21,5'd13,5'd23,5'd16,5'd16,5'd11,5'd15,5'd11,5'd15,5'd19,5'd16,5'd15,5'd18,5'd12,5'd19,5'd12,5'd15,5'd14,5'd23,5'd14,5'd15,5'd10,5'd23,5'd6,5'd22,5'd6,5'd18,5'd9,5'd24,5'd6,5'd17,5'd3,5'd24,5'd13,5'd17,5'd14,5'd13,5'd9,5'd16,5'd16,5'd17,5'd10,5'd23,5'd9,5'd24,5'd18,5'd23,5'd10,5'd24,5'd6,5'd22,5'd11,5'd16,5'd16,5'd17,5'd14,5'd22,5'd12,5'd21,5'd6,5'd21,5'd14,5'd24,5'd8,5'd14,5'd12,5'd7,5'd19,5'd11,5'd15,5'd12,5'd24,5'd19,5'd12,5'd12,5'd16,5'd3,5'd23,5'd9,5'd18,5'd6,5'd21,5'd12,5'd21,5'd8,5'd20,5'd10,5'd13,5'd12,5'd16,5'd22,5'd20,5'd17,5'd21,5'd17,5'd21,5'd12,5'd21,5'd11,5'd21,5'd21,5'd14,5'd13,5'd24,5'd10,5'd18,5'd12,5'd24,5'd9,5'd24,5'd11,5'd22,5'd2,5'd17,5'd12,5'd16,5'd12,5'd18,5'd20,5'd23,5'd11,5'd15,5'd12,5'd22,5'd12,5'd20,5'd6,5'd18,5'd12,5'd19,5'd9,5'd18,5'd9,5'd20,5'd11,5'd14,5'd10,5'd19,5'd7,5'd19,5'd16,5'd24,5'd12,5'd23,5'd14,5'd15,5'd21,5'd22,5'd4,5'd15,5'd9,5'd15,5'd12,5'd14,5'd21,5'd22,5'd13,5'd14,5'd8,5'd19,5'd7,5'd21,5'd19,5'd24,5'd9,5'd23,5'd11,5'd15,5'd11,5'd24,5'd13,5'd14,5'd12,5'd19,5'd16,5'd16,5'd17,5'd24,5'd14,5'd18,5'd10,5'd17,5'd8,5'd19,5'd9,5'd23,5'd14,5'd16,5'd14,5'd23,5'd15,5'd15,5'd4,5'd21,5'd24,5'd16,5'd18,5'd12,5'd2,5'd24,5'd5,5'd24,5'd8,5'd15,5'd11,5'd15,5'd11,5'd16,5'd9,5'd16,5'd20,5'd17,5'd13,5'd24,5'd10,5'd20,5'd12,5'd15,5'd19,5'd16,5'd3,5'd23,5'd18,5'd24,5'd11,5'd22,5'd9,5'd23,5'd7,5'd20,5'd8,5'd14,5'd11,5'd20,5'd13,5'd15,5'd17,5'd18,5'd9,5'd20,5'd6,5'd17,5'd14,5'd16,5'd19,5'd22,5'd12,5'd21,5'd14,5'd21,5'd24,5'd14,5'd19,5'd17,5'd18,5'd13,5'd14,5'd24,5'd4,5'd22,5'd6,5'd21,5'd18,5'd16,5'd9,5'd10,5'd21,5'd10,5'd20,5'd17,5'd20,5'd10,5'd19,5'd12,5'd14,5'd5,5'd22,5'd9,5'd18,5'd12,5'd20,5'd11,5'd15,5'd16,5'd24,5'd15,5'd12,5'd12,5'd23,5'd11,5'd22,5'd11,5'd23,5'd10,5'd18,5'd15,5'd16,5'd12,5'd19,5'd22,5'd18,5'd15,5'd24,5'd12,5'd22,5'd5,5'd24,5'd7,5'd19,5'd19,5'd20,5'd16,5'd23,5'd10,5'd24,5'd7,5'd20,5'd20,5'd21,5'd8,5'd19,5'd7,5'd21,5'd17,5'd14,5'd18,5'd24,5'd8,5'd20,5'd6,5'd12,5'd12,5'd17,5'd9,5'd16,5'd8,5'd18,5'd5,5'd14,5'd11,5'd15,5'd11,5'd16,5'd11,5'd22,5'd9,5'd24,5'd18,5'd14,5'd19,5'd24,5'd13,5'd13,5'd11,5'd19,5'd14,5'd17,5'd13,5'd17,5'd13,5'd17,5'd11,5'd17,5'd3,5'd24,5'd4,5'd20,5'd17,5'd23,5'd21,5'd23,5'd13,5'd17,5'd14,5'd17,5'd6,5'd13,5'd22,5'd21,5'd20,5'd22,5'd4,5'd15,5'd24,5'd23,5'd15,5'd24,5'd4,5'd24,5'd15,5'd20,5'd20,5'd17,5'd10,5'd19,5'd9,5'd14,5'd11,5'd13,5'd7,5'd22,5'd6,5'd22,5'd12,5'd16,5'd10,5'd22,5'd12,5'd24,5'd12,5'd12,5'd19,5'd20,5'd19,5'd23,5'd20,5'd14,5'd13,5'd15,5'd18,5'd15,5'd10,5'd14,5'd13,5'd13,5'd11,5'd12,5'd22,5'd24,5'd6,5'd21,5'd9,5'd21,5'd5,5'd17,5'd15,5'd15,5'd6,5'd24,5'd8,5'd24,5'd18,5'd13,5'd9,5'd16,5'd20,5'd20,5'd23,5'd10,5'd24,5'd24,5'd20,5'd12,5'd18,5'd16,5'd18,5'd19,5'd15,5'd13,5'd17,5'd14,5'd19,5'd12,5'd17,5'd12,5'd19,5'd12,5'd23,5'd4,5'd24,5'd14,5'd20,5'd9,5'd14,5'd10,5'd23,5'd11,5'd15,5'd12,5'd14,5'd6,5'd15,5'd9,5'd24,5'd8,5'd24,5'd19,5'd24,5'd16,5'd22,5'd4,5'd15,5'd3,5'd15,5'd6,5'd15,5'd18,5'd15,5'd4,5'd22,5'd9,5'd15,5'd12,5'd18,5'd10,5'd24,5'd3,5'd24,5'd9,5'd21,5'd10,5'd24,5'd20,5'd24,5'd17,5'd24,5'd7,5'd19,5'd8,5'd18,5'd5,5'd23,5'd4,5'd12,5'd15,5'd24,5'd9,5'd17,5'd12,5'd21,5'd9,5'd17,5'd6,5'd20,5'd13,5'd13,5'd15,5'd15,5'd20,5'd24,5'd9,5'd21,5'd12,5'd15,5'd24,5'd15,5'd12,5'd21,5'd11,5'd17,5'd5,5'd15,5'd12,5'd14,5'd13,5'd13,5'd12,5'd15,5'd12,5'd17,5'd18,5'd15,5'd12,5'd21,5'd11,5'd14,5'd10,5'd16,5'd11,5'd12,5'd16,5'd14,5'd15,5'd24,5'd20,5'd24,5'd6,5'd24,5'd12,5'd24,5'd11,5'd23,5'd7,5'd13,5'd9,5'd21,5'd10,5'd24,5'd13,5'd23,5'd9,5'd21,5'd9,5'd16,5'd15,5'd19,5'd14,5'd24,5'd20,5'd16,5'd7,5'd22,5'd8,5'd24,5'd4,5'd18,5'd16,5'd17,5'd19,5'd23,5'd13,5'd20,5'd15,5'd15,5'd11,5'd15,5'd7,5'd19,5'd12,5'd20,5'd12,5'd18,5'd11,5'd22,5'd10,5'd21,5'd4,5'd17,5'd4,5'd22,5'd9,5'd17,5'd18,5'd23,5'd15,5'd20,5'd14,5'd17,5'd11,5'd20,5'd14,5'd19,5'd14,5'd12,5'd21,5'd15,5'd12,5'd16,5'd10,5'd17,5'd11,5'd12,5'd11,5'd23,5'd9,5'd17,5'd19,5'd17,5'd19,5'd20,5'd10,5'd24,5'd21,5'd24,5'd5,5'd22,5'd7,5'd24,5'd18,5'd18,5'd11,5'd15,5'd11,5'd13,5'd12,5'd19,5'd9,5'd18,5'd13,5'd17,5'd11,5'd15,5'd16,5'd24,5'd7,5'd23,5'd4,5'd20,5'd8,5'd24,5'd8,5'd21,5'd17,5'd20,5'd13,5'd12,5'd7,5'd16,5'd12,5'd20,5'd18,5'd18,5'd10,5'd16,5'd18,5'd16,5'd20,5'd19,5'd12,5'd24,5'd13,5'd18,5'd4,5'd22,5'd9,5'd24,5'd6,5'd20,5'd8,5'd20,5'd7,5'd19,5'd20,5'd19,5'd12,5'd17,5'd7,5'd20,5'd10,5'd20,5'd12,5'd21,5'd20,5'd24,5'd3,5'd15,5'd11,5'd24,5'd19,5'd24,5'd21,5'd24,5'd11,5'd23,5'd10,5'd24,5'd8,5'd22,5'd13,5'd12,5'd10,5'd23,5'd24,5'd23,5'd12,5'd15,5'd15,5'd21,5'd14,5'd13,5'd12,5'd15,5'd11,5'd23,5'd19,5'd24,5'd11,5'd14,5'd9,5'd17,5'd21,5'd17,5'd14,5'd17,5'd18,5'd15,5'd5,5'd24,5'd7,5'd16,5'd12,5'd20,5'd17,5'd14,5'd11,5'd24,5'd14,5'd14,5'd21,5'd24,5'd9,5'd24,5'd24,5'd23,5'd9,5'd24,5'd16,5'd18,5'd12,5'd19,5'd18,5'd21,5'd14,5'd20,5'd12,5'd21,5'd10,5'd24,5'd13,5'd20,5'd19,5'd20,5'd14,5'd20,5'd11,5'd19,5'd11,5'd17,5'd9,5'd12,5'd6,5'd20,5'd5,5'd21,5'd8,5'd18,5'd16,5'd18,5'd13,5'd13,5'd14,5'd22,5'd6,5'd15,5'd13,5'd21,5'd7,5'd14,5'd20,5'd12,5'd12,5'd12,5'd22,5'd13,5'd15,5'd11,5'd14,5'd7,5'd16,5'd10,5'd12,5'd22,5'd24,5'd14,5'd24,5'd11,5'd24,5'd18,5'd17,5'd10,5'd24,5'd23,5'd23,5'd10,5'd19,5'd10,5'd14,5'd13,5'd24,5'd13,5'd13,5'd6,5'd22,5'd13,5'd13,5'd12,5'd23,5'd12,5'd14,5'd11,5'd24,5'd21,5'd23,5'd6,5'd24,5'd12,5'd15,5'd11,5'd23,5'd10,5'd24,5'd13,5'd15,5'd16,5'd14,5'd13,5'd12,5'd17,5'd23,5'd10,5'd24,5'd20,5'd15,5'd14,5'd23,5'd10,5'd22,5'd5,5'd15,5'd4,5'd23,5'd7,5'd17,5'd9,5'd23,5'd7,5'd24,5'd17,5'd15,5'd10,5'd19,5'd13,5'd16,5'd15,5'd24,5'd6,5'd24,5'd21,5'd24,5'd10,5'd16,5'd17,5'd14,5'd13,5'd15,5'd14,5'd15,5'd10,5'd15,5'd9,5'd22,5'd12,5'd15,5'd11,5'd24,5'd15,5'd21,5'd22,5'd20,5'd13,5'd20,5'd13,5'd14,5'd20,5'd14,5'd11,5'd24,5'd4,5'd16,5'd16,5'd24,5'd9,5'd21,5'd9,5'd24,5'd6,5'd23,5'd19,5'd24,5'd22,5'd16,5'd6,5'd24,5'd20,5'd23,5'd19,5'd17,5'd10,5'd16,5'd13,5'd18,5'd19,5'd15,5'd13,5'd16,5'd12,5'd14,5'd12,5'd15,5'd22,5'd21,5'd12,5'd19,5'd19,5'd21,5'd4,5'd24,5'd16,5'd22,5'd9,5'd23,5'd12,5'd21,5'd6,5'd13,5'd9,5'd16,5'd17,5'd13,5'd16,5'd14,5'd18,5'd12,5'd14,5'd21,5'd22,5'd12,5'd21,5'd20,5'd22,5'd7,5'd24,5'd15,5'd17,5'd14,5'd20,5'd22,5'd24,5'd9,5'd17,5'd20,5'd20,5'd24,5'd17,5'd18,5'd21,5'd17,5'd21,5'd12,5'd14,5'd9,5'd18,5'd10,5'd16,5'd16,5'd14,5'd6,5'd24,5'd14,5'd23,5'd19,5'd24,5'd8,5'd24,5'd7,5'd18,5'd12,5'd18,5'd12,5'd24,5'd11,5'd15,5'd9,5'd19,5'd5,5'd23,5'd13,5'd23,5'd20,5'd21,5'd10,5'd18,5'd7,5'd21,5'd7,5'd18,5'd11,5'd16,5'd11,5'd19,5'd11,5'd18,5'd5,5'd24,5'd12,5'd18,5'd18,5'd24,5'd22,5'd15,5'd8,5'd20,5'd10,5'd19,5'd23,5'd21,5'd11,5'd20,5'd4,5'd23,5'd12,5'd13,5'd14,5'd19,5'd8,5'd12,5'd18,5'd15,5'd7,5'd22,5'd13,5'd15,5'd10,5'd16,5'd14,5'd24,5'd8,5'd16,5'd9,5'd23,5'd18,5'd21,5'd7,5'd16,5'd16,5'd19,5'd10,5'd20,5'd15,5'd21,5'd6,5'd24,5'd23,5'd21,5'd10,5'd23,5'd15,5'd20,5'd12,5'd20,5'd10,5'd14,5'd14,5'd17,5'd9,5'd17,5'd13,5'd24,5'd6,5'd20,5'd6,5'd20,5'd11,5'd14,5'd17,5'd15,5'd12,5'd22,5'd9,5'd20,5'd10,5'd17,5'd16,5'd2,5'd24,5'd12,5'd16,5'd10,5'd16,5'd12,5'd14,5'd12,5'd23,5'd15,5'd12,5'd14,5'd13,5'd10,5'd19,5'd11,5'd21,5'd6,5'd24,5'd7,5'd23,5'd5,5'd24,5'd9,5'd16,5'd10,5'd18,5'd13,5'd14,5'd18,5'd18,5'd5,5'd23,5'd7,5'd15,5'd13,5'd13,5'd10,5'd23,5'd17,5'd18,5'd11,5'd19,5'd14,5'd14,5'd4,5'd15,5'd14,5'd19,5'd10,5'd22,5'd11,5'd24,5'd21,5'd22,5'd12,5'd24,5'd20,5'd19,5'd13,5'd21,5'd4,5'd22,5'd2,5'd23,5'd9,5'd16,5'd12,5'd23,5'd7,5'd24,5'd8,5'd21,5'd7,5'd20,5'd5,5'd12,5'd4,5'd23,5'd18,5'd22,5'd9,5'd13,5'd12,5'd20,5'd9,5'd22,5'd8,5'd22,5'd15,5'd20,5'd12,5'd20,5'd19,5'd24,5'd5,5'd23,5'd10,5'd20,5'd11,5'd24,5'd10,5'd18,5'd15,5'd17,5'd11,5'd17,5'd17,5'd14,5'd12,5'd17,5'd11,5'd17,5'd13,5'd17,5'd9,5'd23,5'd23,5'd24,5'd18,5'd24,5'd7,5'd19,5'd11,5'd14,5'd4,5'd24,5'd6,5'd23,5'd22,5'd24,5'd19,5'd22,5'd20,5'd15,5'd4,5'd22,5'd9,5'd24,5'd9,5'd14,5'd10,5'd21,5'd12,5'd15,5'd9,5'd17,5'd3,5'd17,5'd14,5'd24,5'd11,5'd13,5'd9,5'd15,5'd14,5'd16,5'd19,5'd14,5'd14,5'd4,5'd12,5'd8,5'd24,5'd15,5'd18,5'd17,5'd15,5'd16,5'd22,5'd6,5'd18,5'd21,5'd18,5'd14,5'd17,5'd5,5'd18,5'd9,5'd24,5'd9,5'd24,5'd19,5'd24,5'd9,5'd21,5'd6,5'd14,5'd12,5'd16,5'd11,5'd22,5'd11,5'd23,5'd8,5'd24,5'd6,5'd16,5'd12,5'd17,5'd14,5'd23,5'd17,5'd14,5'd21,5'd16,5'd10,5'd16,5'd4,5'd22,5'd4,5'd24,5'd11,5'd16,5'd12,5'd12,5'd19,5'd16,5'd8,5'd23,5'd6,5'd24,5'd12,5'd19,5'd11,5'd22,5'd12,5'd24,5'd7,5'd24,5'd12,5'd24,5'd9,5'd16,5'd13,5'd13,5'd21,5'd24,5'd21,5'd16,5'd18,5'd16,5'd12,5'd24,5'd8,5'd18,5'd14,5'd18,5'd20,5'd23,5'd19,5'd23,5'd11,5'd22,5'd9,5'd24,5'd11,5'd24,5'd19,5'd15,5'd15,5'd24,5'd11,5'd15,5'd12,5'd24,5'd12,5'd24,5'd13,5'd14,5'd14,5'd14,5'd19,5'd23,5'd11,5'd17,5'd4,5'd22,5'd5,5'd16,5'd10,5'd20,5'd10,5'd16,5'd10,5'd20,5'd9,5'd21,5'd22,5'd22,5'd12,5'd24,5'd13,5'd20,5'd9,5'd23,5'd4,5'd17,5'd21,5'd20,5'd19,5'd22,5'd15,5'd23,5'd16,5'd24,5'd9,5'd24,5'd7,5'd22,5'd12,5'd15,5'd9,5'd16,5'd12,5'd21,5'd6,5'd14,5'd14,5'd12,5'd6,5'd14,5'd8,5'd23,5'd15,5'd21,5'd10,5'd17,5'd16,5'd22,5'd9,5'd14,5'd15,5'd15,5'd18,5'd20,5'd15,5'd19,5'd24,5'd21,5'd19,5'd21,5'd21,5'd21,5'd6,5'd23,5'd11,5'd15,5'd14,5'd19,5'd13,5'd15,5'd14,5'd23,5'd16,5'd13,5'd10,5'd24,5'd7,5'd21,5'd20,5'd22,5'd13,5'd13,5'd16,5'd14,5'd8,5'd12,5'd18,5'd17,5'd5,5'd17,5'd9,5'd21,5'd12,5'd14,5'd13,5'd13,5'd20,5'd23,5'd18,5'd18,5'd12,5'd23,5'd9,5'd21,5'd4,5'd23,5'd21,5'd23,5'd4,5'd16,5'd21,5'd24,5'd11,5'd16,5'd9,5'd15,5'd16,5'd14,5'd12,5'd22,5'd15,5'd24,5'd11,5'd16,5'd6,5'd21,5'd4,5'd22,5'd9,5'd24,5'd6,5'd18,5'd12,5'd22,5'd24,5'd19,5'd16,5'd23,5'd10,5'd16,5'd4,5'd24,5'd16,5'd24,5'd9,5'd13,5'd15,5'd24,5'd17,5'd7,5'd22,5'd8,5'd12,5'd9,5'd14,5'd10,5'd18,5'd15,5'd18,5'd7,5'd22,5'd22,5'd19,5'd17,5'd18,5'd12,5'd16,5'd15,5'd24,5'd6,5'd20,5'd10,5'd19,5'd13,5'd23,5'd12,5'd22,5'd8,5'd24,5'd8,5'd18,5'd15,5'd24,5'd18,5'd17,5'd7,5'd15,5'd11,5'd15,5'd22,5'd20,5'd11,5'd15,5'd13,5'd14,5'd14,5'd24,5'd13,5'd14,5'd17,5'd18,5'd5,5'd21,5'd10,5'd24,5'd13,5'd24,5'd13,5'd19,5'd11,5'd16,5'd7,5'd14,5'd16,5'd13,5'd17,5'd12,5'd18,5'd22,5'd11,5'd23,5'd5,5'd21,5'd8,5'd24,5'd11,5'd15,5'd19,5'd24,5'd11,5'd20,5'd21,5'd20,5'd12,5'd18,5'd10,5'd17,5'd9,5'd23,5'd8,5'd17,5'd23,5'd14,5'd13,5'd22,5'd10,5'd13,5'd10,5'd20,5'd18,5'd17,5'd8,5'd24,5'd4,5'd14,5'd12,5'd16,5'd13,5'd21,5'd10,5'd17,5'd10,5'd22,5'd12,5'd24,5'd11,5'd23,5'd19,5'd23,5'd9,5'd24,5'd4,5'd22,5'd4,5'd14,5'd18,5'd14,5'd21,5'd16,5'd20,5'd13,5'd17,5'd16,5'd9,5'd9,5'd17,5'd13,5'd17,5'd11,5'd15,5'd11,5'd17,5'd21,5'd18,5'd7,5'd15,5'd13,5'd21,5'd10,5'd15,5'd16,5'd17,5'd7,5'd15,5'd12,5'd17,5'd16,5'd17,5'd14,5'd21,5'd13,5'd20,5'd13,5'd15,5'd11,5'd14,5'd13,5'd17,5'd22,5'd18,5'd17,5'd23,5'd17,5'd18,5'd22,5'd21,5'd10,5'd18,5'd13,5'd14,5'd12,5'd24,5'd9,5'd24,5'd19,5'd24,5'd20,5'd24,5'd11,5'd16,5'd9,5'd24,5'd18,5'd21,5'd23,5'd24,5'd12,5'd17,5'd9,5'd19,5'd8,5'd23,5'd10,5'd24,5'd13,5'd17,5'd8,5'd24,5'd20,5'd24,5'd6,5'd13,5'd11,5'd24,5'd4,5'd24,5'd5,5'd24,5'd19,5'd24,5'd12,5'd16,5'd16,5'd15,5'd20,5'd22,5'd13,5'd14,5'd12,5'd14,5'd4,5'd12,5'd14,5'd21,5'd15,5'd17,5'd20,5'd14,5'd8,5'd22,5'd8,5'd24,5'd5,5'd22,5'd4,5'd22,5'd20,5'd24,5'd11,5'd23,5'd16,5'd21,5'd23,5'd17,5'd12,5'd19,5'd22,5'd19,5'd9,5'd14,5'd20,5'd13,5'd24,5'd7,5'd18,5'd10,5'd21,5'd11,5'd21,5'd12,5'd14,5'd12,5'd19,5'd10,5'd22,5'd6,5'd21,5'd2,5'd23,5'd22,5'd24,5'd21,5'd24,5'd21,5'd15,5'd10,5'd15,5'd10,5'd21,5'd18,5'd12,5'd6,5'd22,5'd6,5'd22,5'd14,5'd24,5'd15,5'd15,5'd22,5'd18,5'd13,5'd15,5'd13,5'd15,5'd7,5'd20,5'd11,5'd16,5'd11,5'd18,5'd9,5'd21,5'd5,5'd18,5'd13,5'd21,5'd13,5'd23,5'd6,5'd16,5'd15,5'd16,5'd8,5'd18,5'd11,5'd15,5'd14,5'd15,5'd11,5'd24,5'd8,5'd12,5'd21,5'd24,5'd10,5'd23,5'd19,5'd12,5'd16,5'd13,5'd10,5'd22,5'd19,5'd17,5'd11,5'd16,5'd12,5'd19,5'd12,5'd20,5'd8,5'd23,5'd20,5'd15,5'd8,5'd18,5'd16,5'd18,5'd11,5'd16,5'd14,5'd16,5'd16,5'd16,5'd6,5'd23,5'd21,5'd21,5'd6,5'd15,5'd19,5'd14,5'd18,5'd16,5'd17,5'd7,5'd22,5'd2,5'd24,5'd7,5'd21,5'd6,5'd14,5'd11,5'd19,5'd6,5'd19,5'd10,5'd16,5'd13,5'd16,5'd9,5'd24,5'd14,5'd24,5'd13,5'd19,5'd9,5'd17,5'd7,5'd19,5'd9,5'd24,5'd18,5'd13,5'd5,5'd21,5'd5,5'd21,5'd21,5'd18,5'd6,5'd17,5'd9,5'd24,5'd6,5'd21,5'd11,5'd15,5'd16,5'd21,5'd4,5'd24,5'd19,5'd24,5'd10,5'd15,5'd14,5'd24,5'd21,5'd21,5'd18,5'd15,5'd18,5'd16,5'd11,5'd15,5'd24,5'd24,5'd14,5'd23,5'd11,5'd14,5'd10,5'd23,5'd11,5'd21,5'd10,5'd19,5'd7,5'd20,5'd6,5'd24,5'd15,5'd24,5'd20,5'd21,5'd9,5'd24,5'd10,5'd23,5'd15,5'd23,5'd10,5'd15,5'd16,5'd14,5'd4,5'd24,5'd15,5'd24,5'd16,5'd14,5'd17,5'd13,5'd14,5'd10,5'd16,5'd8,5'd22,5'd12,5'd19,5'd15,5'd13,5'd9,5'd16,5'd12,5'd19,5'd13,5'd22,5'd4,5'd21,5'd5,5'd16,5'd15,5'd16,5'd8,5'd22,5'd9,5'd17,5'd3,5'd15,5'd11,5'd17,5'd21,5'd24,5'd11,5'd21,5'd18,5'd24,5'd5,5'd24,5'd24,5'd20,5'd17,5'd24,5'd12,5'd24,5'd19,5'd23,5'd11,5'd18,5'd19,5'd16,5'd22,5'd20,5'd12,5'd21,5'd19,5'd24,5'd10,5'd16,5'd15,5'd15,5'd10,5'd16,5'd7,5'd23,5'd19,5'd18,5'd6,5'd24,5'd16,5'd24,5'd17,5'd22,5'd14,5'd23,5'd11,5'd15,5'd13,5'd18,5'd15,5'd15,5'd11,5'd18,5'd10,5'd22,5'd9,5'd22,5'd6,5'd13,5'd10,5'd19,5'd16,5'd12,5'd12,5'd21,5'd13,5'd13,5'd14,5'd12,5'd19,5'd20,5'd23,5'd13,5'd24,5'd24,5'd19,5'd16,5'd18,5'd15,5'd18,5'd9,5'd19,5'd12,5'd23,5'd14,5'd24,5'd14,5'd14,5'd18,5'd16,5'd16,5'd22,5'd4,5'd23,5'd11,5'd24,5'd21,5'd23,5'd9,5'd24,5'd6,5'd21,5'd7,5'd19,5'd3,5'd18,5'd10,5'd20,5'd12,5'd24,5'd19,5'd24,5'd11,5'd15,5'd14,5'd24,5'd11,5'd14,5'd8,5'd24,5'd16,5'd24,5'd12,5'd14,5'd18,5'd23,5'd6,5'd24,5'd18,5'd24,5'd3,5'd24,5'd11,5'd19,5'd12,5'd22,5'd22,5'd15,5'd10,5'd16,5'd8,5'd19,5'd14,5'd18,5'd16,5'd14,5'd21,5'd15,5'd12,5'd18,5'd11,5'd21,5'd10,5'd15,5'd11,5'd14,5'd13,5'd24,5'd20,5'd17,5'd12,5'd15,5'd11,5'd24,5'd10,5'd16,5'd11,5'd15,5'd12,5'd13,5'd6,5'd24,5'd16,5'd15,5'd17,5'd24,5'd5,5'd18,5'd7,5'd17,5'd14,5'd17,5'd16,5'd15,5'd9,5'd17,5'd9,5'd24,5'd9,5'd16,5'd6,5'd16,5'd6,5'd17,5'd16,5'd13,5'd11,5'd18,5'd12,5'd15,5'd13,5'd15,5'd14,5'd17,5'd12,5'd18,5'd6,5'd20,5'd16,5'd15,5'd7,5'd17,5'd9,5'd20,5'd13,5'd22,5'd19,5'd24,5'd11,5'd23,5'd15,5'd14,5'd20,5'd16,5'd19,5'd23,5'd12,5'd15,5'd15,5'd15,5'd11,5'd14,5'd11,5'd21,5'd18,5'd21,5'd11,5'd17,5'd10,5'd17,5'd20,5'd19,5'd10,5'd21,5'd9,5'd22,5'd12,5'd15,5'd11,5'd15,5'd12,5'd15,5'd9,5'd24,5'd21,5'd24,5'd18,5'd15,5'd13,5'd13,5'd11,5'd24,5'd9,5'd23,5'd20,5'd20,5'd4,5'd24,5'd4,5'd24,5'd20,5'd22,5'd14,5'd23,5'd7,5'd16,5'd13,5'd20,5'd12,5'd18,5'd17,5'd21,5'd22,5'd15,5'd19,5'd10,5'd15,5'd10,5'd15,5'd22,5'd24,5'd12,5'd18,5'd12,5'd15,5'd13,5'd23,5'd18,5'd19,5'd10,5'd18,5'd11,5'd16,5'd11,5'd16,5'd20,5'd16,5'd12,5'd20,5'd19,5'd16,5'd10,5'd18,5'd6,5'd21,5'd9,5'd17,5'd19,5'd15,5'd21,5'd20,5'd6,5'd21,5'd6,5'd21,5'd11,5'd21,5'd22,5'd15,5'd13,5'd18,5'd16,5'd24,5'd8,5'd20,5'd10,5'd19,5'd23,5'd22,5'd10,5'd14,5'd6,5'd21,5'd14,5'd22,5'd10,5'd19,5'd12,5'd12,5'd11,5'd22,5'd15,5'd14,5'd9,5'd17,5'd10,5'd16,5'd6,5'd23,5'd11,5'd16,5'd8,5'd22,5'd4,5'd22,5'd8,5'd24,5'd23,5'd24,5'd10,5'd17,5'd14,5'd14,5'd19,5'd15,5'd13,5'd13,5'd14,5'd13,5'd16,5'd14,5'd20,5'd16,5'd18,5'd15,5'd12,5'd14,5'd11,5'd13,5'd15,5'd14,5'd12,5'd19,5'd10,5'd23,5'd10,5'd19,5'd11,5'd21,5'd4,5'd20,5'd19,5'd24,5'd14,5'd18,5'd11,5'd17,5'd9,5'd16,5'd5,5'd21,5'd8,5'd22,5'd16,5'd14,5'd18,5'd6,5'd19,5'd19,5'd19,5'd12,5'd14,5'd19,5'd14,5'd4,5'd22,5'd22,5'd22,5'd4,5'd12,5'd12,5'd23,5'd12,5'd16,5'd7,5'd21,5'd18,5'd15,5'd9,5'd13,5'd14,5'd20,5'd16,5'd19,5'd17,5'd13,5'd16,5'd22,5'd6,5'd14,5'd11,5'd19,5'd19,5'd19,5'd15,5'd16,5'd20,5'd14,5'd18,5'd11,5'd15,5'd17,5'd18,5'd7,5'd17,5'd21,5'd14,5'd18}
`define RECTANGLE2_Y2 {5'd12,5'd21,5'd22,5'd21,5'd21,5'd21,5'd21,5'd15,5'd17,5'd20,5'd21,5'd11,5'd21,5'd18,5'd18,5'd23,5'd20,5'd21,5'd18,5'd18,5'd18,5'd16,5'd15,5'd15,5'd18,5'd19,5'd19,5'd18,5'd18,5'd17,5'd17,5'd14,5'd14,5'd10,5'd22,5'd8,5'd8,5'd7,5'd19,5'd17,5'd10,5'd13,5'd13,5'd9,5'd9,5'd18,5'd12,5'd4,5'd24,5'd13,5'd8,5'd23,5'd23,5'd11,5'd15,5'd9,5'd11,5'd13,5'd6,5'd16,5'd20,5'd22,5'd21,5'd18,5'd19,5'd20,5'd7,5'd11,5'd11,5'd11,5'd9,5'd10,5'd10,5'd8,5'd14,5'd18,5'd5,5'd6,5'd7,5'd9,5'd15,5'd11,5'd9,5'd2,5'd11,5'd12,5'd12,5'd16,5'd22,5'd20,5'd20,5'd15,5'd15,5'd12,5'd14,5'd17,5'd17,5'd21,5'd16,5'd16,5'd23,5'd20,5'd20,5'd10,5'd7,5'd7,5'd16,5'd18,5'd18,5'd16,5'd18,5'd13,5'd13,5'd9,5'd10,5'd14,5'd18,5'd19,5'd19,5'd23,5'd23,5'd18,5'd24,5'd4,5'd10,5'd9,5'd11,5'd20,5'd20,5'd18,5'd18,5'd18,5'd18,5'd6,5'd6,5'd20,5'd20,5'd22,5'd21,5'd23,5'd23,5'd15,5'd15,5'd14,5'd19,5'd4,5'd9,5'd9,5'd8,5'd14,5'd14,5'd24,5'd9,5'd15,5'd7,5'd9,5'd11,5'd16,5'd18,5'd18,5'd18,5'd17,5'd17,5'd14,5'd14,5'd6,5'd4,5'd14,5'd14,5'd13,5'd13,5'd18,5'd2,5'd10,5'd13,5'd18,5'd23,5'd24,5'd3,5'd16,5'd12,5'd23,5'd21,5'd20,5'd9,5'd19,5'd19,5'd15,5'd15,5'd5,5'd5,5'd12,5'd21,5'd19,5'd21,5'd16,5'd20,5'd6,5'd11,5'd10,5'd13,5'd5,5'd8,5'd18,5'd17,5'd9,5'd7,5'd13,5'd16,5'd15,5'd22,5'd22,5'd22,5'd22,5'd14,5'd14,5'd24,5'd24,5'd20,5'd13,5'd10,5'd10,5'd9,5'd12,5'd10,5'd10,5'd20,5'd23,5'd24,5'd24,5'd13,5'd13,5'd12,5'd9,5'd22,5'd22,5'd10,5'd16,5'd11,5'd21,5'd10,5'd12,5'd13,5'd8,5'd20,5'd8,5'd15,5'd11,5'd9,5'd11,5'd11,5'd22,5'd24,5'd24,5'd22,5'd20,5'd3,5'd10,5'd10,5'd14,5'd13,5'd13,5'd16,5'd16,5'd8,5'd12,5'd15,5'd15,5'd13,5'd11,5'd11,5'd13,5'd19,5'd24,5'd20,5'd9,5'd23,5'd12,5'd24,5'd13,5'd18,5'd13,5'd14,5'd14,5'd24,5'd24,5'd19,5'd21,5'd20,5'd20,5'd13,5'd13,5'd19,5'd19,5'd23,5'd17,5'd9,5'd12,5'd24,5'd23,5'd11,5'd9,5'd11,5'd11,5'd12,5'd16,5'd13,5'd24,5'd15,5'd24,5'd14,5'd19,5'd19,5'd13,5'd13,5'd13,5'd20,5'd8,5'd9,5'd23,5'd16,5'd12,5'd13,5'd13,5'd13,5'd11,5'd14,5'd6,5'd5,5'd5,5'd19,5'd19,5'd15,5'd15,5'd16,5'd7,5'd9,5'd16,5'd9,5'd13,5'd15,5'd9,5'd17,5'd3,5'd10,5'd21,5'd17,5'd11,5'd19,5'd17,5'd24,5'd24,5'd16,5'd13,5'd9,5'd7,5'd16,5'd14,5'd15,5'd9,5'd7,5'd7,5'd9,5'd2,5'd17,5'd18,5'd17,5'd17,5'd14,5'd14,5'd12,5'd9,5'd12,5'd12,5'd10,5'd12,5'd11,5'd11,5'd23,5'd23,5'd15,5'd10,5'd20,5'd23,5'd21,5'd20,5'd11,5'd17,5'd22,5'd18,5'd18,5'd17,5'd20,5'd20,5'd8,5'd12,5'd17,5'd17,5'd4,5'd15,5'd16,5'd9,5'd3,5'd18,5'd6,5'd8,5'd23,5'd16,5'd15,5'd11,5'd6,5'd10,5'd7,5'd15,5'd11,5'd8,5'd11,5'd23,5'd9,5'd6,5'd6,5'd7,5'd19,5'd17,5'd17,5'd24,5'd24,5'd11,5'd24,5'd12,5'd12,5'd16,5'd9,5'd12,5'd7,5'd23,5'd12,5'd11,5'd24,5'd7,5'd24,5'd22,5'd24,5'd16,5'd24,5'd16,5'd24,5'd15,5'd8,5'd12,5'd11,5'd14,5'd12,5'd19,5'd19,5'd15,5'd15,5'd21,5'd24,5'd19,5'd19,5'd12,5'd14,5'd9,5'd11,5'd22,5'd11,5'd17,5'd20,5'd24,5'd18,5'd14,5'd14,5'd15,5'd13,5'd12,5'd12,5'd15,5'd15,5'd11,5'd16,5'd10,5'd19,5'd12,5'd12,5'd20,5'd21,5'd14,5'd14,5'd19,5'd10,5'd23,5'd23,5'd24,5'd14,5'd20,5'd17,5'd17,5'd17,5'd13,5'd4,5'd10,5'd12,5'd6,5'd6,5'd11,5'd10,5'd10,5'd18,5'd4,5'd6,5'd19,5'd19,5'd19,5'd16,5'd22,5'd17,5'd15,5'd4,5'd6,5'd19,5'd10,5'd4,5'd12,5'd9,5'd15,5'd10,5'd16,5'd16,5'd11,5'd11,5'd16,5'd24,5'd19,5'd11,5'd14,5'd19,5'd22,5'd12,5'd3,5'd14,5'd23,5'd11,5'd14,5'd14,5'd18,5'd18,5'd20,5'd11,5'd12,5'd24,5'd19,5'd19,5'd24,5'd24,5'd7,5'd7,5'd12,5'd14,5'd12,5'd12,5'd16,5'd15,5'd24,5'd24,5'd13,5'd13,5'd18,5'd18,5'd22,5'd22,5'd22,5'd19,5'd15,5'd15,5'd15,5'd17,5'd20,5'd12,5'd14,5'd22,5'd23,5'd20,5'd21,5'd21,5'd9,5'd12,5'd20,5'd24,5'd2,5'd15,5'd16,5'd14,5'd14,5'd14,5'd24,5'd8,5'd9,5'd13,5'd23,5'd15,5'd17,5'd17,5'd22,5'd22,5'd12,5'd13,5'd12,5'd4,5'd15,5'd20,5'd21,5'd19,5'd5,5'd6,5'd21,5'd24,5'd24,5'd24,5'd24,5'd18,5'd18,5'd16,5'd16,5'd15,5'd20,5'd22,5'd24,5'd21,5'd10,5'd15,5'd9,5'd12,5'd15,5'd14,5'd18,5'd9,5'd10,5'd21,5'd13,5'd20,5'd20,5'd20,5'd20,5'd9,5'd12,5'd22,5'd9,5'd17,5'd18,5'd13,5'd12,5'd23,5'd17,5'd17,5'd18,5'd18,5'd18,5'd21,5'd21,5'd15,5'd19,5'd16,5'd14,5'd9,5'd9,5'd9,5'd15,5'd14,5'd23,5'd10,5'd11,5'd18,5'd18,5'd10,5'd9,5'd10,5'd10,5'd15,5'd10,5'd9,5'd9,5'd14,5'd24,5'd15,5'd15,5'd17,5'd17,5'd19,5'd19,5'd20,5'd20,5'd20,5'd17,5'd12,5'd20,5'd21,5'd20,5'd5,5'd17,5'd17,5'd13,5'd13,5'd13,5'd15,5'd13,5'd13,5'd13,5'd14,5'd20,5'd16,5'd19,5'd19,5'd13,5'd9,5'd13,5'd24,5'd24,5'd18,5'd18,5'd12,5'd10,5'd24,5'd5,5'd18,5'd18,5'd5,5'd15,5'd3,5'd8,5'd7,5'd5,5'd15,5'd12,5'd19,5'd9,5'd7,5'd10,5'd15,5'd20,5'd14,5'd18,5'd9,5'd23,5'd9,5'd21,5'd19,5'd19,5'd18,5'd11,5'd12,5'd2,5'd18,5'd19,5'd24,5'd16,5'd7,5'd4,5'd3,5'd13,5'd5,5'd17,5'd15,5'd23,5'd10,5'd10,5'd11,5'd15,5'd6,5'd9,5'd13,5'd15,5'd4,5'd16,5'd13,5'd13,5'd10,5'd14,5'd16,5'd17,5'd22,5'd24,5'd18,5'd18,5'd18,5'd24,5'd19,5'd15,5'd16,5'd6,5'd6,5'd8,5'd8,5'd16,5'd16,5'd10,5'd11,5'd16,5'd16,5'd23,5'd16,5'd21,5'd14,5'd22,5'd22,5'd18,5'd8,5'd7,5'd16,5'd15,5'd8,5'd19,5'd12,5'd21,5'd16,5'd10,5'd11,5'd4,5'd22,5'd13,5'd12,5'd11,5'd11,5'd15,5'd14,5'd20,5'd15,5'd18,5'd2,5'd7,5'd7,5'd8,5'd7,5'd18,5'd11,5'd10,5'd11,5'd19,5'd11,5'd20,5'd11,5'd24,5'd11,5'd23,5'd23,5'd11,5'd11,5'd15,5'd15,5'd19,5'd20,5'd17,5'd20,5'd21,5'd21,5'd21,5'd20,5'd19,5'd8,5'd5,5'd4,5'd16,5'd16,5'd21,5'd21,5'd6,5'd6,5'd13,5'd11,5'd17,5'd9,5'd12,5'd12,5'd14,5'd13,5'd20,5'd12,5'd9,5'd9,5'd18,5'd23,5'd22,5'd15,5'd14,5'd9,5'd9,5'd16,5'd15,5'd8,5'd9,5'd7,5'd12,5'd12,5'd12,5'd22,5'd17,5'd8,5'd18,5'd24,5'd13,5'd21,5'd15,5'd8,5'd8,5'd20,5'd5,5'd7,5'd2,5'd11,5'd9,5'd13,5'd17,5'd17,5'd15,5'd14,5'd12,5'd18,5'd24,5'd4,5'd23,5'd12,5'd7,5'd4,5'd24,5'd21,5'd23,5'd23,5'd21,5'd13,5'd19,5'd19,5'd19,5'd19,5'd17,5'd12,5'd15,5'd15,5'd24,5'd24,5'd21,5'd16,5'd18,5'd2,5'd9,5'd9,5'd8,5'd7,5'd8,5'd12,5'd7,5'd18,5'd22,5'd21,5'd19,5'd7,5'd24,5'd4,5'd11,5'd14,5'd9,5'd9,5'd15,5'd15,5'd12,5'd21,5'd21,5'd9,5'd14,5'd10,5'd17,5'd18,5'd10,5'd14,5'd22,5'd22,5'd9,5'd9,5'd19,5'd12,5'd23,5'd6,5'd16,5'd9,5'd20,5'd14,5'd10,5'd10,5'd4,5'd16,5'd17,5'd20,5'd17,5'd17,5'd19,5'd19,5'd16,5'd11,5'd13,5'd13,5'd10,5'd20,5'd19,5'd19,5'd18,5'd18,5'd16,5'd9,5'd10,5'd10,5'd17,5'd23,5'd16,5'd16,5'd4,5'd7,5'd9,5'd9,5'd13,5'd10,5'd8,5'd9,5'd15,5'd15,5'd11,5'd15,5'd12,5'd18,5'd24,5'd11,5'd9,5'd5,5'd24,5'd9,5'd5,5'd20,5'd24,5'd24,5'd8,5'd5,5'd12,5'd14,5'd19,5'd19,5'd18,5'd5,5'd10,5'd13,5'd9,5'd14,5'd10,5'd15,5'd17,5'd13,5'd13,5'd13,5'd17,5'd9,5'd14,5'd14,5'd10,5'd10,5'd17,5'd17,5'd22,5'd22,5'd14,5'd14,5'd24,5'd18,5'd17,5'd15,5'd16,5'd16,5'd20,5'd9,5'd10,5'd20,5'd13,5'd16,5'd18,5'd9,5'd20,5'd7,5'd12,5'd6,5'd8,5'd8,5'd12,5'd7,5'd9,5'd9,5'd21,5'd21,5'd24,5'd12,5'd20,5'd21,5'd24,5'd20,5'd11,5'd13,5'd10,5'd9,5'd13,5'd11,5'd14,5'd14,5'd7,5'd7,5'd12,5'd5,5'd14,5'd15,5'd24,5'd24,5'd23,5'd24,5'd24,5'd21,5'd24,5'd9,5'd7,5'd5,5'd9,5'd13,5'd6,5'd16,5'd16,5'd17,5'd23,5'd18,5'd6,5'd23,5'd19,5'd17,5'd18,5'd18,5'd5,5'd5,5'd19,5'd20,5'd21,5'd21,5'd11,5'd9,5'd11,5'd19,5'd15,5'd9,5'd8,5'd24,5'd19,5'd4,5'd15,5'd16,5'd24,5'd19,5'd15,5'd19,5'd22,5'd10,5'd16,5'd23,5'd16,5'd11,5'd6,5'd19,5'd17,5'd17,5'd9,5'd9,5'd20,5'd9,5'd9,5'd15,5'd16,5'd2,5'd6,5'd24,5'd20,5'd14,5'd13,5'd11,5'd6,5'd12,5'd24,5'd12,5'd16,5'd7,5'd16,5'd17,5'd24,5'd21,5'd14,5'd20,5'd5,5'd3,5'd20,5'd24,5'd12,5'd15,5'd15,5'd19,5'd22,5'd21,5'd12,5'd12,5'd15,5'd17,5'd17,5'd10,5'd9,5'd13,5'd19,5'd23,5'd24,5'd16,5'd3,5'd8,5'd8,5'd13,5'd20,5'd23,5'd23,5'd6,5'd9,5'd4,5'd3,5'd9,5'd9,5'd13,5'd22,5'd12,5'd11,5'd11,5'd7,5'd12,5'd12,5'd14,5'd16,5'd15,5'd14,5'd18,5'd21,5'd5,5'd2,5'd5,5'd12,5'd11,5'd12,5'd16,5'd23,5'd18,5'd13,5'd6,5'd18,5'd18,5'd9,5'd20,5'd6,5'd15,5'd12,5'd24,5'd24,5'd10,5'd10,5'd16,5'd16,5'd11,5'd15,5'd8,5'd8,5'd7,5'd8,5'd17,5'd17,5'd18,5'd11,5'd12,5'd24,5'd19,5'd12,5'd24,5'd24,5'd16,5'd24,5'd14,5'd12,5'd9,5'd11,5'd13,5'd20,5'd12,5'd12,5'd13,5'd13,5'd12,5'd12,5'd7,5'd15,5'd6,5'd20,5'd18,5'd24,5'd18,5'd18,5'd21,5'd21,5'd21,5'd21,5'd9,5'd8,5'd4,5'd21,5'd19,5'd21,5'd11,5'd21,5'd18,5'd11,5'd7,5'd16,5'd9,5'd9,5'd13,5'd18,5'd4,5'd8,5'd19,5'd8,5'd14,5'd14,5'd15,5'd8,5'd4,5'd10,5'd9,5'd12,5'd21,5'd8,5'd13,5'd4,5'd20,5'd13,5'd17,5'd6,5'd11,5'd21,5'd10,5'd15,5'd14,5'd5,5'd9,5'd8,5'd11,5'd17,5'd10,5'd10,5'd10,5'd6,5'd6,5'd6,5'd6,5'd8,5'd7,5'd10,5'd10,5'd23,5'd7,5'd12,5'd11,5'd15,5'd15,5'd4,5'd20,5'd13,5'd16,5'd10,5'd7,5'd16,5'd10,5'd10,5'd16,5'd24,5'd24,5'd20,5'd19,5'd19,5'd20,5'd17,5'd24,5'd11,5'd11,5'd14,5'd12,5'd12,5'd23,5'd8,5'd11,5'd8,5'd6,5'd5,5'd10,5'd13,5'd23,5'd19,5'd21,5'd15,5'd15,5'd14,5'd14,5'd8,5'd14,5'd18,5'd14,5'd9,5'd10,5'd17,5'd17,5'd16,5'd16,5'd16,5'd16,5'd15,5'd9,5'd20,5'd17,5'd20,5'd20,5'd16,5'd6,5'd5,5'd4,5'd20,5'd19,5'd22,5'd22,5'd8,5'd8,5'd24,5'd20,5'd14,5'd8,5'd7,5'd7,5'd12,5'd19,5'd23,5'd8,5'd18,5'd14,5'd11,5'd15,5'd21,5'd3,5'd16,5'd9,5'd15,5'd19,5'd12,5'd9,5'd21,5'd13,5'd20,5'd18,5'd18,5'd19,5'd24,5'd24,5'd24,5'd24,5'd21,5'd21,5'd20,5'd17,5'd10,5'd10,5'd11,5'd9,5'd16,5'd16,5'd16,5'd21,5'd16,5'd21,5'd13,5'd9,5'd15,5'd15,5'd22,5'd22,5'd18,5'd20,5'd21,5'd21,5'd6,5'd21,5'd19,5'd14,5'd14,5'd23,5'd11,5'd6,5'd19,5'd7,5'd12,5'd12,5'd6,5'd24,5'd22,5'd17,5'd18,5'd23,5'd23,5'd17,5'd8,5'd13,5'd20,5'd13,5'd12,5'd22,5'd23,5'd7,5'd7,5'd7,5'd7,5'd8,5'd8,5'd9,5'd9,5'd16,5'd16,5'd21,5'd18,5'd12,5'd9,5'd15,5'd24,5'd11,5'd21,5'd16,5'd17,5'd19,5'd24,5'd20,5'd24,5'd11,5'd4,5'd22,5'd19,5'd16,5'd16,5'd15,5'd6,5'd12,5'd18,5'd16,5'd16,5'd14,5'd16,5'd16,5'd10,5'd8,5'd8,5'd18,5'd23,5'd23,5'd17,5'd18,5'd20,5'd23,5'd23,5'd21,5'd21,5'd20,5'd20,5'd4,5'd19,5'd17,5'd10,5'd15,5'd15,5'd14,5'd14,5'd10,5'd9,5'd6,5'd6,5'd16,5'd19,5'd20,5'd24,5'd9,5'd19,5'd20,5'd20,5'd19,5'd14,5'd13,5'd14,5'd9,5'd12,5'd13,5'd18,5'd20,5'd12,5'd15,5'd21,5'd13,5'd19,5'd12,5'd15,5'd24,5'd17,5'd13,5'd13,5'd11,5'd15,5'd14,5'd13,5'd12,5'd13,5'd13,5'd13,5'd18,5'd17,5'd19,5'd18,5'd19,5'd21,5'd9,5'd9,5'd9,5'd15,5'd12,5'd10,5'd13,5'd9,5'd6,5'd13,5'd12,5'd4,5'd2,5'd9,5'd13,5'd13,5'd11,5'd11,5'd11,5'd14,5'd12,5'd2,5'd13,5'd9,5'd9,5'd9,5'd13,5'd19,5'd13,5'd5,5'd14,5'd15,5'd17,5'd24,5'd22,5'd7,5'd10,5'd16,5'd24,5'd18,5'd14,5'd8,5'd8,5'd15,5'd5,5'd23,5'd23,5'd20,5'd4,5'd5,5'd11,5'd24,5'd8,5'd22,5'd10,5'd16,5'd5,5'd19,5'd19,5'd16,5'd16,5'd22,5'd16,5'd12,5'd12,5'd16,5'd15,5'd13,5'd13,5'd17,5'd11,5'd22,5'd21,5'd21,5'd11,5'd16,5'd11,5'd13,5'd19,5'd20,5'd16,5'd11,5'd11,5'd17,5'd6,5'd9,5'd9,5'd13,5'd15,5'd13,5'd6,5'd17,5'd17,5'd11,5'd11,5'd20,5'd16,5'd21,5'd9,5'd8,5'd8,5'd19,5'd9,5'd9,5'd21,5'd11,5'd9,5'd9,5'd20,5'd22,5'd9,5'd18,5'd18,5'd17,5'd20,5'd9,5'd9,5'd12,5'd11,5'd14,5'd12,5'd4,5'd8,5'd13,5'd13,5'd21,5'd13,5'd3,5'd2,5'd18,5'd18,5'd20,5'd20,5'd17,5'd17,5'd23,5'd9,5'd8,5'd15,5'd6,5'd17,5'd14,5'd23,5'd12,5'd11,5'd12,5'd18,5'd14,5'd15,5'd15,5'd14,5'd24,5'd18,5'd9,5'd20,5'd24,5'd21,5'd15,5'd23,5'd11,5'd11,5'd15,5'd15,5'd20,5'd20,5'd15,5'd13,5'd17,5'd24,5'd14,5'd14,5'd10,5'd10,5'd6,5'd12,5'd19,5'd5,5'd5,5'd8,5'd16,5'd13,5'd24,5'd3,5'd4,5'd7,5'd10,5'd2,5'd20,5'd20,5'd12,5'd11,5'd17,5'd7,5'd21,5'd21,5'd16,5'd24,5'd16,5'd12,5'd14,5'd24,5'd14,5'd14,5'd18,5'd21,5'd19,5'd9,5'd18,5'd14,5'd17,5'd14,5'd13,5'd17,5'd24,5'd19,5'd18,5'd4,5'd2,5'd21,5'd19,5'd21,5'd20,5'd21,5'd11,5'd8,5'd16,5'd15,5'd12,5'd4,5'd17,5'd17,5'd21,5'd7,5'd10,5'd21,5'd3,5'd3,5'd14,5'd15,5'd9,5'd9,5'd15,5'd21,5'd12,5'd13,5'd19,5'd14,5'd7,5'd19,5'd12,5'd20,5'd21,5'd21,5'd11,5'd11,5'd15,5'd11,5'd7,5'd20,5'd17,5'd15,5'd3,5'd20,5'd16,5'd13,5'd17,5'd17,5'd4,5'd4,5'd6,5'd7,5'd15,5'd16,5'd9,5'd9,5'd9,5'd17,5'd17,5'd17,5'd6,5'd10,5'd24,5'd13,5'd19,5'd19,5'd19,5'd19,5'd12,5'd12,5'd18,5'd19,5'd11,5'd15,5'd15,5'd14,5'd2,5'd8,5'd21,5'd3,5'd15,5'd22,5'd16,5'd16,5'd23,5'd16,5'd21,5'd15,5'd4,5'd15,5'd10,5'd23,5'd23,5'd18,5'd17,5'd11,5'd15,5'd12,5'd12,5'd19,5'd13,5'd16,5'd24,5'd13,5'd13,5'd14,5'd12,5'd9,5'd16,5'd24,5'd17,5'd13,5'd9,5'd10,5'd10,5'd9,5'd19,5'd15,5'd17,5'd22,5'd6,5'd15,5'd18,5'd22,5'd12,5'd13,5'd22,5'd17,5'd8,5'd13,5'd13,5'd13,5'd14,5'd24,5'd24,5'd19,5'd14,5'd17,5'd14,5'd12,5'd17,5'd24,5'd10,5'd13,5'd20,5'd21,5'd3,5'd12,5'd5,5'd7,5'd12,5'd9,5'd8,5'd18,5'd13,5'd11,5'd11,5'd7,5'd24,5'd7,5'd18,5'd7,5'd18,5'd24,5'd24,5'd6,5'd7,5'd9,5'd22,5'd8,5'd12,5'd21,5'd22,5'd8,5'd22,5'd24,5'd24,5'd12,5'd12,5'd12,5'd6,5'd15,5'd12,5'd14,5'd16,5'd24,5'd24,5'd15,5'd16,5'd18,5'd12,5'd6,5'd24,5'd18,5'd14,5'd6,5'd16,5'd9,5'd7,5'd13,5'd24,5'd15,5'd15,5'd19,5'd15,5'd24,5'd4,5'd19,5'd11,5'd17,5'd17,5'd20,5'd3,5'd11,5'd11,5'd12,5'd12,5'd19,5'd6,5'd2,5'd23,5'd4,5'd15,5'd10,5'd6,5'd15,5'd19,5'd15,5'd16,5'd18,5'd8,5'd13,5'd23,5'd7,5'd7,5'd20,5'd19,5'd12,5'd24,5'd21,5'd19,5'd24,5'd24,5'd20,5'd15,5'd16,5'd14,5'd14,5'd9,5'd9,5'd9,5'd4,5'd14,5'd23,5'd14,5'd18,5'd10,5'd9,5'd9,5'd10,5'd22,5'd15,5'd11,5'd12,5'd17,5'd17,5'd11,5'd12,5'd16,5'd16,5'd16,5'd15,5'd18,5'd19,5'd19,5'd19,5'd18,5'd2,5'd6,5'd6,5'd17,5'd17,5'd20,5'd20,5'd18,5'd15,5'd10,5'd21,5'd7,5'd10,5'd7,5'd21,5'd18,5'd14,5'd16,5'd18,5'd12,5'd14,5'd18,5'd21,5'd17,5'd4,5'd11,5'd24,5'd15,5'd11,5'd15,5'd15,5'd13,5'd13,5'd13,5'd5,5'd16,5'd22,5'd21,5'd17,5'd18,5'd18,5'd15,5'd15,5'd23,5'd23,5'd9,5'd23,5'd12,5'd8,5'd14,5'd15,5'd7,5'd12,5'd16,5'd16,5'd19,5'd19,5'd20,5'd10,5'd12,5'd13,5'd24,5'd17,5'd9,5'd6,5'd20,5'd20,5'd6,5'd22,5'd15,5'd16,5'd16,5'd15,5'd6,5'd11,5'd6,5'd14,5'd14,5'd23,5'd23,5'd9,5'd9,5'd9,5'd17,5'd19,5'd24,5'd6,5'd6,5'd9,5'd11,5'd22,5'd23,5'd11,5'd11,5'd20,5'd11,5'd9,5'd16,5'd8,5'd10,5'd11,5'd10,5'd23,5'd9,5'd14,5'd24,5'd19,5'd19,5'd8,5'd11,5'd14,5'd8,5'd8,5'd8,5'd22,5'd22,5'd14,5'd14,5'd13,5'd11,5'd9,5'd9,5'd16,5'd16,5'd24,5'd24,5'd24,5'd9,5'd14,5'd17,5'd14,5'd9,5'd14,5'd23,5'd9,5'd24,5'd10,5'd24,5'd20,5'd16,5'd9,5'd9,5'd15,5'd15,5'd22,5'd21,5'd24,5'd11,5'd9,5'd19,5'd17,5'd19,5'd18,5'd8,5'd22,5'd20,5'd8,5'd24,5'd8,5'd12,5'd20,5'd13,5'd9,5'd7,5'd11,5'd20,5'd18,5'd22,5'd2,5'd12,5'd9,5'd9,5'd19,5'd12,5'd18,5'd17,5'd16,5'd18,5'd23,5'd17,5'd6,5'd18,5'd3,5'd6,5'd13,5'd24,5'd19,5'd11,5'd12,5'd3,5'd6,5'd20,5'd20,5'd22,5'd14,5'd19,5'd16,5'd6,5'd15,5'd13,5'd17,5'd21,5'd12,5'd21,5'd21,5'd16,5'd20,5'd4,5'd4,5'd17,5'd17,5'd14,5'd14,5'd17,5'd21,5'd17,5'd17,5'd6,5'd6,5'd13,5'd24,5'd10,5'd10,5'd16,5'd16,5'd7,5'd17,5'd18,5'd18,5'd18,5'd18,5'd15,5'd9,5'd17,5'd17,5'd16,5'd20,5'd17,5'd17,5'd14,5'd17,5'd24,5'd10,5'd14,5'd15,5'd2,5'd8,5'd9,5'd24,5'd16,5'd13,5'd16,5'd16,5'd4,5'd4,5'd15,5'd18,5'd17,5'd15,5'd9,5'd18,5'd14,5'd13,5'd5,5'd5,5'd8,5'd5,5'd9,5'd9,5'd23,5'd19,5'd19,5'd12,5'd13,5'd13,5'd22,5'd22,5'd22,5'd22,5'd21,5'd19,5'd17,5'd12,5'd17,5'd10,5'd24,5'd14,5'd5,5'd11,5'd6,5'd12,5'd13,5'd12,5'd5,5'd13,5'd20,5'd15,5'd19,5'd13,5'd10,5'd10,5'd9,5'd16,5'd11,5'd24,5'd9,5'd11,5'd17,5'd14,5'd9,5'd17,5'd19,5'd19,5'd14,5'd24,5'd24,5'd24,5'd11,5'd15,5'd24,5'd23,5'd18,5'd18,5'd18,5'd19,5'd3,5'd5,5'd5,5'd11,5'd11,5'd11,5'd12,5'd15,5'd8,5'd23,5'd5,5'd20,5'd14,5'd19,5'd24,5'd2,5'd8,5'd9,5'd18,5'd19,5'd19,5'd9,5'd9,5'd22,5'd16,5'd20,5'd20,5'd20,5'd20,5'd24,5'd8,5'd10,5'd10,5'd10,5'd10,5'd19,5'd14,5'd13,5'd19,5'd14,5'd14,5'd8,5'd16,5'd24,5'd8,5'd13,5'd13,5'd23,5'd23,5'd21,5'd7,5'd18,5'd15,5'd15,5'd15,5'd6,5'd14,5'd15,5'd22,5'd24,5'd18,5'd15,5'd11,5'd17,5'd9,5'd6,5'd16,5'd21,5'd5,5'd22,5'd18,5'd11,5'd18,5'd11,5'd19,5'd19,5'd12,5'd13,5'd24,5'd19,5'd13,5'd15,5'd8,5'd13,5'd15,5'd20,5'd7,5'd7,5'd6,5'd19,5'd15,5'd16,5'd16,5'd16,5'd18,5'd18,5'd9,5'd9,5'd14,5'd14,5'd11,5'd9,5'd15,5'd19,5'd23,5'd15,5'd20,5'd20,5'd16,5'd16,5'd20,5'd14,5'd20,5'd16,5'd10,5'd16,5'd9,5'd9,5'd4,5'd12,5'd8,5'd8,5'd22,5'd8,5'd15,5'd15,5'd21,5'd20,5'd15,5'd16,5'd5,5'd15,5'd22,5'd20,5'd19,5'd16,5'd11,5'd10,5'd6,5'd24,5'd23,5'd24,5'd10,5'd11,5'd11,5'd22,5'd15,5'd12,5'd22,5'd22,5'd9,5'd20,5'd19,5'd21,5'd21,5'd24,5'd17,5'd6,5'd18,5'd18,5'd9,5'd9,5'd16,5'd11,5'd18,5'd18,5'd16,5'd14,5'd13,5'd13,5'd6,5'd10,5'd19,5'd15,5'd16,5'd13,5'd19,5'd14,5'd18,5'd18,5'd12,5'd12,5'd23,5'd24,5'd9,5'd22,5'd7,5'd12,5'd17,5'd10,5'd15,5'd22,5'd11,5'd11,5'd6,5'd10,5'd16,5'd22,5'd19,5'd19,5'd7,5'd15,5'd22,5'd12,5'd16,5'd10,5'd19,5'd16,5'd14,5'd16,5'd6,5'd19,5'd17,5'd16,5'd11,5'd11,5'd24,5'd19,5'd6,5'd5,5'd5,5'd23,5'd24,5'd17,5'd18,5'd18,5'd9,5'd18,5'd12,5'd8,5'd15,5'd16,5'd24,5'd10,5'd8,5'd24,5'd24,5'd20,5'd21,5'd21,5'd16,5'd15,5'd13,5'd13,5'd11,5'd9,5'd8,5'd11,5'd17,5'd11,5'd16,5'd12,5'd7,5'd18,5'd14,5'd14,5'd14,5'd4,5'd3,5'd11,5'd10,5'd18,5'd9,5'd24,5'd2,5'd9,5'd23,5'd6,5'd20,5'd21,5'd11,5'd14,5'd6,5'd19,5'd13,5'd20,5'd18,5'd18,5'd24,5'd23,5'd23,5'd24,5'd24,5'd17,5'd10,5'd15,5'd14,5'd17,5'd17,5'd19,5'd12,5'd12,5'd7,5'd12,5'd22,5'd6,5'd6,5'd3,5'd6,5'd7,5'd6,5'd8,5'd18,5'd24,5'd22,5'd21,5'd24,5'd19,5'd19,5'd11,5'd21,5'd19,5'd17,5'd14,5'd23,5'd22,5'd22,5'd8,5'd9,5'd15,5'd7,5'd17,5'd23,5'd11,5'd12,5'd6,5'd9,5'd22,5'd22,5'd22,5'd13,5'd21,5'd4,5'd15,5'd24,5'd6,5'd22,5'd21,5'd16,5'd11,5'd11,5'd11,5'd24,5'd15,5'd12,5'd22,5'd18,5'd20,5'd18,5'd9,5'd9,5'd11,5'd11,5'd16,5'd9,5'd21,5'd19,5'd14,5'd14,5'd19,5'd18,5'd3,5'd20,5'd18,5'd10,5'd17,5'd17,5'd24,5'd24,5'd15,5'd15,5'd17,5'd15,5'd23,5'd12,5'd15,5'd6,5'd6,5'd12,5'd15,5'd15,5'd9,5'd15,5'd6,5'd5,5'd12,5'd11,5'd19,5'd19,5'd20,5'd16,5'd12,5'd2,5'd21,5'd16,5'd19,5'd19,5'd19,5'd10,5'd15,5'd21,5'd15,5'd24,5'd16,5'd16,5'd20,5'd14,5'd6,5'd11,5'd10,5'd10,5'd24,5'd12,5'd12,5'd10,5'd10,5'd8,5'd10,5'd14,5'd13,5'd24,5'd15,5'd14,5'd23,5'd11,5'd20,5'd12,5'd23,5'd16,5'd16,5'd10,5'd24,5'd18,5'd15,5'd20,5'd14,5'd6,5'd19,5'd22,5'd15,5'd19,5'd11,5'd14,5'd18,5'd15,5'd17,5'd6,5'd16,5'd19,5'd5,5'd16,5'd11,5'd10,5'd6,5'd24,5'd14,5'd21,5'd24,5'd22,5'd15,5'd11,5'd10}
`define RECTANGLE2_WEIGHTS {32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384}
`define RECTANGLE3_X1 {5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd3,5'd18,5'd0,5'd0,5'd11,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd13,5'd4,5'd16,5'd7,5'd3,5'd6,5'd15,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd6,5'd12,5'd10,5'd11,5'd0,5'd7,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd14,5'd7,5'd12,5'd0,5'd12,5'd0,5'd0,5'd3,5'd19,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd5,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd8,5'd10,5'd0,5'd0,5'd7,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd10,5'd7,5'd0,5'd0,5'd5,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd8,5'd4,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd8,5'd0,5'd13,5'd0,5'd0,5'd12,5'd0,5'd11,5'd10,5'd0,5'd2,5'd0,5'd0,5'd9,5'd11,5'd5,5'd15,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd14,5'd6,5'd0,5'd9,5'd12,5'd0,5'd13,5'd3,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd4,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd12,5'd10,5'd3,5'd13,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd6,5'd0,5'd0,5'd11,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd1,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd5,5'd9,5'd12,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd7,5'd15,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd2,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd9,5'd7,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd2,5'd20,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd20,5'd0,5'd0,5'd12,5'd11,5'd0,5'd0,5'd3,5'd19,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd7,5'd14,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd12,5'd13,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd16,5'd9,5'd12,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd1,5'd11,5'd0,5'd0,5'd11,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd9,5'd3,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd3,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd10,5'd6,5'd14,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd12,5'd7,5'd12,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd9,5'd0,5'd0,5'd5,5'd11,5'd11,5'd12,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd11,5'd6,5'd11,5'd0,5'd11,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd15,5'd0,5'd0,5'd0,5'd4,5'd9,5'd13,5'd12,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd12,5'd7,5'd11,5'd0,5'd5,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd12,5'd5,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd7,5'd15,5'd12,5'd0,5'd12,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd11,5'd3,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd7,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd14,5'd0,5'd6,5'd12,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd10,5'd0,5'd0,5'd0,5'd1,5'd0,5'd0,5'd12,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd7,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd5,5'd0,5'd9,5'd0,5'd6,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd1,5'd6,5'd12,5'd0,5'd0,5'd11,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd4,5'd15,5'd0,5'd0,5'd0,5'd17,5'd7,5'd2,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd4,5'd0,5'd0,5'd16,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd12,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd7,5'd0,5'd12,5'd10,5'd0,5'd0,5'd0,5'd0,5'd9,5'd11,5'd5,5'd15,5'd0,5'd15,5'd0,5'd0,5'd10,5'd10,5'd0,5'd0,5'd7,5'd0,5'd11,5'd10,5'd11,5'd7,5'd11,5'd0,5'd5,5'd14,5'd12,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd14,5'd4,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd1,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd14,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd5,5'd15,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd10,5'd4,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd11,5'd0,5'd0,5'd0,5'd0,5'd7,5'd14,5'd0,5'd0,5'd4,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd5,5'd3,5'd10,5'd8,5'd11,5'd16,5'd10,5'd6,5'd0,5'd11,5'd11,5'd9,5'd0,5'd10,5'd0,5'd9,5'd0,5'd9,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd6,5'd9,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd10,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd2,5'd11,5'd9,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd12,5'd5,5'd11,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd1,5'd0,5'd0,5'd0,5'd0,5'd7,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd6,5'd0,5'd8,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd1,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd4,5'd0,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd7,5'd4,5'd17,5'd0,5'd0,5'd4,5'd8,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd16,5'd0,5'd16,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd10,5'd10,5'd0,5'd0,5'd7,5'd0,5'd0,5'd5,5'd0,5'd10,5'd0,5'd8,5'd0,5'd16,5'd0,5'd4,5'd10,5'd9,5'd0,5'd1,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd12,5'd8,5'd0,5'd0,5'd10,5'd11,5'd0,5'd6,5'd0,5'd0,5'd0,5'd1,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd12,5'd4,5'd16,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd7,5'd11,5'd0,5'd0,5'd0,5'd12,5'd7,5'd0,5'd0,5'd0,5'd0,5'd2,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd5,5'd0,5'd0,5'd6,5'd14,5'd6,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd12,5'd0,5'd0,5'd7,5'd0,5'd0,5'd10,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd4,5'd16,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd7,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd5,5'd0,5'd0,5'd5,5'd14,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd1,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd8,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd17,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd15,5'd0,5'd0,5'd3,5'd10,5'd10,5'd4,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd1,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd3,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd2,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd2,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd9,5'd12,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd11,5'd0,5'd0,5'd0,5'd2,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd11,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0}
`define RECTANGLE3_Y1 {5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd18,5'd18,5'd0,5'd0,5'd21,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd17,5'd14,5'd14,5'd10,5'd22,5'd8,5'd8,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd13,5'd9,5'd10,5'd14,5'd0,5'd19,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd6,5'd20,5'd20,5'd0,5'd21,5'd0,5'd0,5'd15,5'd15,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd9,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd16,5'd11,5'd0,5'd0,5'd12,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd15,5'd15,5'd0,5'd0,5'd11,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd11,5'd9,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd13,5'd0,5'd8,5'd0,5'd0,5'd16,5'd0,5'd13,5'd13,5'd0,5'd11,5'd0,5'd0,5'd5,5'd5,5'd19,5'd19,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd12,5'd0,5'd12,5'd12,5'd0,5'd12,5'd11,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd9,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd6,5'd6,5'd7,5'd19,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd12,5'd0,5'd0,5'd15,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd13,5'd12,5'd12,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd11,5'd11,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd14,5'd0,5'd0,5'd16,5'd15,5'd0,5'd0,5'd13,5'd13,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd15,5'd15,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd16,5'd14,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd18,5'd16,5'd16,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd14,5'd0,5'd0,5'd10,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd13,5'd14,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd5,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd21,5'd19,5'd19,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd7,5'd16,5'd15,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd4,5'd0,5'd0,5'd12,5'd11,5'd11,5'd15,5'd0,5'd0,5'd0,5'd0,5'd2,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd11,5'd20,5'd11,5'd0,5'd11,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd6,5'd0,5'd0,5'd0,5'd9,5'd12,5'd12,5'd14,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd17,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd2,5'd11,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd15,5'd15,5'd12,5'd0,5'd21,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd13,5'd13,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd9,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd16,5'd0,5'd9,5'd10,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd21,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd11,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd9,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd9,5'd0,5'd19,5'd0,5'd9,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd9,5'd9,5'd0,5'd0,5'd12,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd6,5'd18,5'd0,5'd0,5'd0,5'd6,5'd15,5'd12,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd18,5'd0,5'd0,5'd18,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd9,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd11,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd11,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd8,5'd0,5'd5,5'd10,5'd0,5'd0,5'd0,5'd0,5'd15,5'd15,5'd14,5'd14,5'd0,5'd14,5'd0,5'd0,5'd9,5'd10,5'd0,5'd0,5'd16,5'd0,5'd16,5'd16,5'd15,5'd9,5'd20,5'd0,5'd20,5'd20,5'd16,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd8,5'd7,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd7,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd16,5'd17,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd14,5'd16,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd19,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd6,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd20,5'd12,5'd15,5'd21,5'd13,5'd19,5'd12,5'd15,5'd0,5'd17,5'd13,5'd13,5'd0,5'd15,5'd0,5'd13,5'd0,5'd13,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd11,5'd11,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd4,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd22,5'd21,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd19,5'd9,5'd9,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd12,5'd11,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd7,5'd0,5'd2,5'd20,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd14,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd3,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd13,5'd17,5'd17,5'd0,5'd0,5'd6,5'd7,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd16,5'd0,5'd16,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd12,5'd12,5'd0,5'd0,5'd16,5'd0,5'd0,5'd13,5'd0,5'd12,5'd0,5'd16,5'd0,5'd17,5'd0,5'd9,5'd10,5'd10,5'd0,5'd19,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd9,5'd7,5'd0,5'd0,5'd15,5'd15,5'd0,5'd15,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd2,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd11,5'd15,5'd15,5'd0,5'd0,5'd0,5'd5,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd9,5'd9,5'd0,5'd0,5'd0,5'd6,5'd6,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd9,5'd0,5'd0,5'd19,5'd19,5'd8,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd20,5'd0,5'd14,5'd19,5'd0,5'd0,5'd15,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd17,5'd17,5'd0,5'd17,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd8,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd18,5'd0,5'd3,5'd5,5'd5,5'd0,5'd0,5'd0,5'd0,5'd15,5'd8,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd13,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd7,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd18,5'd0,5'd0,5'd14,5'd14,5'd11,5'd9,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd11,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd18,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd3,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd11,5'd11,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd11,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd11,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0}
`define RECTANGLE3_X2 {5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd6,5'd21,5'd0,5'd0,5'd22,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd18,5'd8,5'd20,5'd9,5'd12,5'd9,5'd18,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd15,5'd18,5'd14,5'd17,5'd0,5'd11,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd19,5'd12,5'd17,5'd0,5'd18,5'd0,5'd0,5'd5,5'd21,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd13,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd12,5'd16,5'd0,5'd0,5'd12,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd17,5'd14,5'd0,5'd0,5'd9,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd14,5'd13,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd13,5'd0,5'd18,5'd0,5'd0,5'd17,5'd0,5'd19,5'd14,5'd0,5'd12,5'd0,5'd0,5'd13,5'd15,5'd9,5'd19,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd18,5'd12,5'd0,5'd11,5'd18,5'd0,5'd15,5'd6,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd13,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd17,5'd13,5'd6,5'd18,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd15,5'd0,5'd0,5'd20,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd12,5'd12,5'd15,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd9,5'd17,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd17,5'd15,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd4,5'd22,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd22,5'd0,5'd0,5'd17,5'd13,5'd0,5'd0,5'd5,5'd21,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd10,5'd17,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd17,5'd17,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd19,5'd12,5'd15,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd22,5'd0,5'd0,5'd17,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd13,5'd5,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd12,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd16,5'd10,5'd18,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd16,5'd12,5'd14,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd18,5'd0,5'd0,5'd14,5'd13,5'd13,5'd14,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd13,5'd11,5'd13,5'd0,5'd13,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd19,5'd0,5'd0,5'd0,5'd14,5'd11,5'd15,5'd21,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd17,5'd14,5'd16,5'd0,5'd9,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd24,5'd13,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd9,5'd17,5'd21,5'd0,5'd22,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd21,5'd13,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd10,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd17,5'd0,5'd13,5'd17,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd16,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd24,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd13,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd12,5'd0,5'd15,5'd0,5'd13,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd18,5'd0,5'd0,5'd22,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd7,5'd19,5'd0,5'd0,5'd0,5'd20,5'd11,5'd13,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd8,5'd0,5'd0,5'd20,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd19,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd22,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd18,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd13,5'd0,5'd24,5'd14,5'd0,5'd0,5'd0,5'd0,5'd13,5'd15,5'd9,5'd19,5'd0,5'd19,5'd0,5'd0,5'd18,5'd14,5'd0,5'd0,5'd10,5'd0,5'd14,5'd13,5'd13,5'd13,5'd16,5'd0,5'd10,5'd19,5'd16,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd17,5'd7,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd17,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd9,5'd19,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd13,5'd13,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd17,5'd0,5'd0,5'd0,5'd0,5'd10,5'd17,5'd0,5'd0,5'd8,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd10,5'd13,5'd20,5'd14,5'd22,5'd20,5'd19,5'd12,5'd0,5'd14,5'd15,5'd13,5'd0,5'd12,5'd0,5'd13,5'd0,5'd13,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd15,5'd12,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd16,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd21,5'd16,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd19,5'd12,5'd17,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd18,5'd18,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd12,5'd0,5'd12,5'd12,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd9,5'd0,5'd15,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd14,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd14,5'd7,5'd20,5'd0,5'd0,5'd7,5'd12,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd20,5'd0,5'd20,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd14,5'd14,5'd0,5'd0,5'd13,5'd0,5'd0,5'd12,5'd0,5'd14,5'd0,5'd12,5'd0,5'd20,5'd0,5'd12,5'd15,5'd14,5'd0,5'd12,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd18,5'd12,5'd0,5'd0,5'd18,5'd14,5'd0,5'd14,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd18,5'd8,5'd20,5'd0,5'd0,5'd0,5'd12,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd14,5'd20,5'd0,5'd0,5'd0,5'd24,5'd13,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd13,5'd0,5'd0,5'd10,5'd18,5'd12,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd17,5'd0,5'd12,5'd11,5'd0,5'd0,5'd12,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd8,5'd20,5'd0,5'd20,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd13,5'd0,5'd12,5'd10,5'd19,5'd0,5'd0,5'd0,5'd0,5'd21,5'd12,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd13,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd20,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd18,5'd0,5'd0,5'd6,5'd14,5'd19,5'd12,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd15,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd12,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd13,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd14,5'd19,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd17,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd15,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0}
`define RECTANGLE3_Y2 {5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd24,5'd24,5'd0,5'd0,5'd24,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd21,5'd20,5'd20,5'd20,5'd24,5'd15,5'd15,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd18,5'd14,5'd15,5'd17,5'd0,5'd24,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd24,5'd24,5'd0,5'd24,5'd0,5'd0,5'd24,5'd24,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd13,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd21,5'd15,5'd0,5'd0,5'd18,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd22,5'd22,5'd0,5'd0,5'd16,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd21,5'd11,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd19,5'd0,5'd12,5'd0,5'd0,5'd20,5'd0,5'd17,5'd21,5'd0,5'd14,5'd0,5'd0,5'd10,5'd10,5'd24,5'd24,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd15,5'd0,5'd21,5'd15,5'd0,5'd21,5'd21,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd11,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd12,5'd12,5'd13,5'd23,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd24,5'd0,5'd0,5'd17,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd17,5'd18,5'd18,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd23,5'd23,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd21,5'd21,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd24,5'd0,5'd0,5'd23,5'd24,5'd0,5'd0,5'd24,5'd24,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd21,5'd21,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd21,5'd19,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd22,5'd22,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd16,5'd0,5'd0,5'd18,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd18,5'd23,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd10,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd24,5'd24,5'd24,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd13,5'd24,5'd24,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd8,5'd0,5'd0,5'd15,5'd21,5'd21,5'd24,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd21,5'd24,5'd21,5'd0,5'd21,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0,5'd11,5'd23,5'd23,5'd16,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd16,5'd19,5'd24,5'd0,5'd24,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd4,5'd18,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd19,5'd0,5'd23,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd16,5'd16,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd15,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd22,5'd0,5'd12,5'd14,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd22,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd14,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd12,5'd0,5'd23,5'd0,5'd12,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd18,5'd18,5'd0,5'd0,5'd20,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd12,5'd23,5'd0,5'd0,5'd0,5'd12,5'd20,5'd19,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd23,5'd0,5'd0,5'd23,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd12,5'd0,5'd0,5'd0,5'd0,5'd7,5'd0,5'd0,5'd0,5'd0,5'd14,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd14,5'd0,5'd8,5'd18,5'd0,5'd0,5'd0,5'd0,5'd22,5'd22,5'd24,5'd24,5'd0,5'd24,5'd0,5'd0,5'd13,5'd19,5'd0,5'd0,5'd24,5'd0,5'd23,5'd23,5'd24,5'd12,5'd24,5'd0,5'd24,5'd24,5'd22,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd16,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd14,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd23,5'd24,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd21,5'd18,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd23,5'd0,5'd0,5'd0,5'd0,5'd20,5'd20,5'd0,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd24,5'd18,5'd24,5'd24,5'd17,5'd24,5'd15,5'd18,5'd0,5'd24,5'd18,5'd18,5'd0,5'd24,5'd0,5'd18,5'd0,5'd18,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd22,5'd17,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd7,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd24,5'd24,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd22,5'd12,5'd13,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd18,5'd14,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd10,5'd0,5'd4,5'd24,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd24,5'd0,5'd19,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd11,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd5,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd20,5'd24,5'd24,5'd0,5'd0,5'd12,5'd13,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd0,5'd24,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd20,5'd20,5'd0,5'd0,5'd21,5'd0,5'd0,5'd20,5'd0,5'd20,5'd0,5'd22,5'd0,5'd24,5'd0,5'd12,5'd15,5'd15,5'd0,5'd22,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd12,5'd12,5'd0,5'd0,5'd18,5'd22,5'd0,5'd18,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd9,5'd0,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd17,5'd24,5'd24,5'd0,5'd0,5'd0,5'd10,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd13,5'd0,5'd0,5'd0,5'd9,5'd12,5'd0,5'd0,5'd0,5'd0,5'd20,5'd0,5'd0,5'd20,5'd0,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd12,5'd0,5'd0,5'd24,5'd24,5'd11,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd0,5'd16,5'd24,5'd0,5'd0,5'd24,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd0,5'd24,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd16,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd21,5'd0,5'd5,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd17,5'd16,5'd0,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd19,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd13,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd0,5'd0,5'd24,5'd21,5'd22,5'd12,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd17,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd8,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd20,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd24,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd16,5'd0,5'd0,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd17,5'd17,5'd16,5'd0,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd16,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd23,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd18,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0}
`define RECTANGLE3_WEIGHTS {32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0}
`define FEATURE_THRESHOLD {32'd4294967293,32'd10,32'd0,32'd4294967294,32'd7,32'd3,32'd4294967291,32'd2,32'd0,32'd4294967295,32'd4294967294,32'd9,32'd2,32'd4294967289,32'd4,32'd4294967291,32'd14,32'd6,32'd0,32'd6,32'd4294967292,32'd4294967294,32'd0,32'd10,32'd3,32'd1,32'd4294967276,32'd4294967293,32'd4294967291,32'd5,32'd4294967287,32'd5,32'd4294967291,32'd6,32'd4294967292,32'd1,32'd4294967295,32'd3,32'd1,32'd4294967295,32'd1,32'd0,32'd4294967294,32'd3,32'd4294967293,32'd4294967289,32'd4294967289,32'd1,32'd18,32'd4294967266,32'd10,32'd2,32'd4294967291,32'd0,32'd2,32'd4,32'd4294967293,32'd4294967288,32'd2,32'd4294967292,32'd0,32'd0,32'd1,32'd1,32'd1,32'd2,32'd9,32'd2,32'd4294967282,32'd3,32'd0,32'd4294967283,32'd4294967266,32'd4294967286,32'd4294967294,32'd0,32'd4294967294,32'd4294967285,32'd1,32'd4,32'd4294967295,32'd3,32'd4,32'd4294967295,32'd4294967293,32'd1,32'd7,32'd4294967294,32'd5,32'd1,32'd2,32'd4,32'd4294967293,32'd3,32'd1,32'd4294967290,32'd4,32'd0,32'd2,32'd4294967288,32'd16,32'd4294967282,32'd4294967266,32'd36,32'd4294967294,32'd2,32'd1,32'd4294967292,32'd1,32'd4294967295,32'd4294967293,32'd4294967285,32'd4294967281,32'd4294967294,32'd4294967293,32'd3,32'd4294967291,32'd2,32'd4294967292,32'd4294967295,32'd2,32'd4294967281,32'd4294967282,32'd5,32'd14,32'd1,32'd4294967287,32'd1,32'd4294967294,32'd1,32'd4294967291,32'd4294967293,32'd1,32'd4294967286,32'd8,32'd4294967293,32'd3,32'd1,32'd4294967294,32'd1,32'd0,32'd6,32'd4294967293,32'd4294967285,32'd0,32'd6,32'd4294967294,32'd4294967289,32'd4294967295,32'd4294967294,32'd8,32'd54,32'd4294967285,32'd4294967292,32'd4294967291,32'd4294967292,32'd4294967291,32'd7,32'd2,32'd4294967294,32'd4294967293,32'd0,32'd0,32'd21,32'd2,32'd6,32'd4294967295,32'd1,32'd4294967295,32'd1,32'd4294967291,32'd4294967295,32'd4294967295,32'd4294967294,32'd4294967295,32'd0,32'd4294967293,32'd4294967292,32'd4294967295,32'd4294967293,32'd0,32'd4294967295,32'd20,32'd3,32'd6,32'd1,32'd7,32'd4294967294,32'd5,32'd2,32'd0,32'd6,32'd4294967286,32'd0,32'd2,32'd4294967295,32'd0,32'd3,32'd2,32'd4294967284,32'd0,32'd4,32'd4294967292,32'd1,32'd3,32'd6,32'd4294967293,32'd7,32'd2,32'd1,32'd7,32'd11,32'd11,32'd16,32'd4294967291,32'd1,32'd4294967274,32'd4294967288,32'd12,32'd1,32'd4294967292,32'd4294967287,32'd1,32'd25,32'd1,32'd1,32'd4294967295,32'd4294967292,32'd4294967295,32'd4294967294,32'd41,32'd4294967295,32'd4294967292,32'd4294967295,32'd4294967294,32'd4,32'd3,32'd2,32'd4,32'd8,32'd10,32'd6,32'd4294967287,32'd3,32'd5,32'd10,32'd4294967291,32'd11,32'd0,32'd4,32'd4294967294,32'd0,32'd7,32'd4294967293,32'd2,32'd0,32'd4294967295,32'd4294967291,32'd12,32'd4294967286,32'd9,32'd4294967285,32'd2,32'd10,32'd2,32'd11,32'd9,32'd4294967280,32'd4294967294,32'd4294967291,32'd1,32'd4294967295,32'd4294967293,32'd4294967266,32'd1,32'd3,32'd4294967293,32'd6,32'd3,32'd4294967292,32'd4294967295,32'd15,32'd4294967295,32'd0,32'd10,32'd5,32'd1,32'd0,32'd11,32'd20,32'd4294967292,32'd4294967292,32'd0,32'd0,32'd2,32'd4294967292,32'd4294967293,32'd0,32'd6,32'd4,32'd17,32'd4294967295,32'd4294967292,32'd2,32'd4294967290,32'd4294967294,32'd28,32'd47,32'd0,32'd4294967285,32'd4294967295,32'd1,32'd4294967294,32'd14,32'd2,32'd4,32'd3,32'd4294967295,32'd4294967293,32'd4,32'd1,32'd4294967293,32'd4294967289,32'd4294967295,32'd4294967293,32'd4294967293,32'd5,32'd4,32'd8,32'd4294967293,32'd5,32'd4294967292,32'd4,32'd6,32'd4294967294,32'd4294967287,32'd4294967292,32'd4,32'd4294967294,32'd1,32'd4294967286,32'd6,32'd1,32'd0,32'd4294967280,32'd5,32'd7,32'd4,32'd4294967294,32'd4294967287,32'd4294967293,32'd7,32'd4294967294,32'd4294967295,32'd7,32'd1,32'd4294967285,32'd4294967294,32'd4,32'd4,32'd4,32'd0,32'd4294967294,32'd4294967295,32'd4294967294,32'd4294967286,32'd4294967292,32'd8,32'd4294967285,32'd4294967280,32'd4294967295,32'd4294967294,32'd4294967295,32'd4294967294,32'd3,32'd0,32'd4294967291,32'd8,32'd6,32'd4294967293,32'd3,32'd4294967290,32'd4294967295,32'd6,32'd0,32'd0,32'd4294967292,32'd2,32'd4294967294,32'd1,32'd4294967294,32'd4294967294,32'd4294967292,32'd3,32'd4294967291,32'd4294967295,32'd1,32'd0,32'd19,32'd3,32'd4294967293,32'd4294967294,32'd4294967294,32'd10,32'd4294967292,32'd3,32'd0,32'd4294967295,32'd5,32'd4,32'd3,32'd14,32'd4294967289,32'd1,32'd9,32'd3,32'd6,32'd1,32'd4294967276,32'd4294967292,32'd0,32'd7,32'd1,32'd4,32'd4294967281,32'd4294967280,32'd4294967283,32'd4294967291,32'd4294967290,32'd7,32'd1,32'd9,32'd5,32'd4294967292,32'd30,32'd4294967280,32'd4294967292,32'd4294967291,32'd4294967281,32'd14,32'd1,32'd4294967295,32'd4294967292,32'd4,32'd10,32'd1,32'd4294967291,32'd12,32'd1,32'd5,32'd4294967294,32'd4294967291,32'd29,32'd1,32'd4294967293,32'd2,32'd3,32'd4294967294,32'd4294967287,32'd4294967294,32'd3,32'd2,32'd4294967295,32'd1,32'd4294967287,32'd0,32'd4294967295,32'd5,32'd4294967289,32'd4294967285,32'd38,32'd0,32'd4294967289,32'd4294967289,32'd5,32'd2,32'd4294967295,32'd1,32'd4294967292,32'd4294967293,32'd4294967295,32'd2,32'd4294967294,32'd2,32'd4294967294,32'd4294967294,32'd4294967285,32'd4294967294,32'd0,32'd3,32'd4294967292,32'd0,32'd1,32'd7,32'd19,32'd8,32'd4294967293,32'd3,32'd4,32'd3,32'd4294967294,32'd4294967290,32'd4294967293,32'd4294967289,32'd4294967286,32'd4294967293,32'd2,32'd14,32'd85,32'd4294967294,32'd0,32'd4294967293,32'd5,32'd0,32'd4294967295,32'd4,32'd4294967291,32'd4294967295,32'd0,32'd4294967295,32'd4294967294,32'd4294967284,32'd4,32'd4294967286,32'd4294967290,32'd4294967294,32'd4294967292,32'd1,32'd8,32'd4294967266,32'd37,32'd1,32'd1,32'd4294967280,32'd4294967267,32'd4294967294,32'd4294967294,32'd4294967290,32'd0,32'd2,32'd4294967294,32'd4294967290,32'd3,32'd4294967290,32'd6,32'd4294967293,32'd4294967293,32'd4294967293,32'd4294967294,32'd4294967294,32'd26,32'd0,32'd1,32'd4294967295,32'd2,32'd4294967287,32'd4294967288,32'd4294967295,32'd4294967290,32'd2,32'd4,32'd4,32'd4294967294,32'd12,32'd4294967294,32'd7,32'd7,32'd4294967295,32'd1,32'd4294967294,32'd3,32'd4294967293,32'd0,32'd5,32'd4294967295,32'd0,32'd4294967294,32'd4294967291,32'd4294967291,32'd4294967293,32'd2,32'd4294967290,32'd4294967289,32'd2,32'd4294967288,32'd4294967291,32'd1,32'd4294967286,32'd4294967287,32'd0,32'd4294967292,32'd4294967292,32'd5,32'd4,32'd4294967288,32'd4294967287,32'd5,32'd2,32'd4294967295,32'd0,32'd3,32'd5,32'd0,32'd4294967291,32'd4294967290,32'd5,32'd4,32'd3,32'd13,32'd3,32'd4294967294,32'd4294967292,32'd9,32'd4294967288,32'd4,32'd2,32'd11,32'd4294967283,32'd5,32'd3,32'd3,32'd4294967289,32'd1,32'd7,32'd5,32'd4294967293,32'd0,32'd20,32'd4294967259,32'd5,32'd4294967283,32'd4294967292,32'd4294967294,32'd4294967294,32'd2,32'd2,32'd4294967292,32'd0,32'd4294967293,32'd4294967292,32'd14,32'd1,32'd23,32'd4294967278,32'd1,32'd4294967294,32'd1,32'd4294967291,32'd4294967292,32'd66,32'd4294967291,32'd9,32'd2,32'd4294967295,32'd4294967284,32'd4294967278,32'd2,32'd0,32'd12,32'd4294967292,32'd1,32'd2,32'd0,32'd4294967291,32'd4294967287,32'd4294967290,32'd1,32'd5,32'd8,32'd4294967287,32'd5,32'd4294967287,32'd26,32'd4294967255,32'd4294967294,32'd3,32'd13,32'd4294967289,32'd4294967295,32'd14,32'd4294967293,32'd4294967294,32'd1,32'd11,32'd4294967295,32'd4,32'd4294967295,32'd5,32'd0,32'd1,32'd4294967295,32'd1,32'd4294967295,32'd11,32'd1,32'd4294967293,32'd4,32'd1,32'd4294967294,32'd4294967289,32'd2,32'd3,32'd4294967294,32'd7,32'd9,32'd4294967284,32'd2,32'd6,32'd4294967290,32'd2,32'd4294967293,32'd4294967287,32'd4294967295,32'd4294967289,32'd4294967294,32'd4294967294,32'd5,32'd4294967284,32'd4294967290,32'd6,32'd0,32'd4294967294,32'd68,32'd9,32'd2,32'd4294967295,32'd4,32'd4294967291,32'd4294967294,32'd4294967294,32'd4294967290,32'd2,32'd5,32'd4,32'd4294967295,32'd10,32'd4294967295,32'd4294967295,32'd4,32'd4294967289,32'd4294967295,32'd4294967294,32'd4294967294,32'd4294967295,32'd4294967287,32'd1,32'd4294967291,32'd2,32'd3,32'd4294967292,32'd4,32'd4294967295,32'd4294967292,32'd1,32'd4,32'd4294967256,32'd4294967287,32'd6,32'd1,32'd4294967292,32'd0,32'd19,32'd8,32'd5,32'd11,32'd13,32'd4294967291,32'd4294967294,32'd5,32'd0,32'd4294967288,32'd4294967293,32'd1,32'd4294967294,32'd7,32'd4294967289,32'd1,32'd7,32'd4294967290,32'd0,32'd1,32'd4294967294,32'd4294967293,32'd3,32'd2,32'd4294967295,32'd4294967295,32'd2,32'd4,32'd24,32'd6,32'd2,32'd4294967293,32'd4,32'd4,32'd4294967288,32'd4294967289,32'd0,32'd4294967292,32'd4294967294,32'd0,32'd4294967295,32'd3,32'd0,32'd5,32'd0,32'd13,32'd4294967292,32'd6,32'd4294967295,32'd0,32'd2,32'd0,32'd9,32'd4294967294,32'd4294967292,32'd2,32'd8,32'd6,32'd4294967291,32'd4294967287,32'd5,32'd4294967292,32'd3,32'd4,32'd0,32'd4294967281,32'd2,32'd4294967292,32'd4294967294,32'd15,32'd4294967283,32'd4294967294,32'd3,32'd7,32'd4294967288,32'd2,32'd2,32'd0,32'd4294967293,32'd4294967295,32'd4294967291,32'd5,32'd1,32'd4294967288,32'd4294967294,32'd4294967286,32'd4294967281,32'd4294967274,32'd4294967294,32'd3,32'd6,32'd4294967294,32'd4294967295,32'd4294967294,32'd3,32'd0,32'd2,32'd25,32'd6,32'd2,32'd6,32'd4294967295,32'd0,32'd4,32'd4294967288,32'd8,32'd6,32'd6,32'd4294967291,32'd5,32'd4294967288,32'd4294967295,32'd4294967295,32'd2,32'd13,32'd4294967287,32'd0,32'd4294967288,32'd1,32'd4,32'd6,32'd4294967280,32'd4294967295,32'd4294967294,32'd4294967291,32'd4294967294,32'd4294967294,32'd9,32'd7,32'd4294967295,32'd4294967294,32'd4294967281,32'd4294967290,32'd0,32'd4294967289,32'd4294967295,32'd4294967294,32'd9,32'd4294967294,32'd1,32'd4294967294,32'd13,32'd4294967290,32'd4294967295,32'd4294967290,32'd0,32'd4294967291,32'd6,32'd4294967290,32'd4294967294,32'd4294967295,32'd2,32'd4294967295,32'd2,32'd4294967295,32'd4294967291,32'd53,32'd3,32'd4294967294,32'd4,32'd3,32'd1,32'd4294967295,32'd4294967295,32'd2,32'd4294967294,32'd4294967294,32'd0,32'd4294967294,32'd2,32'd2,32'd2,32'd0,32'd4294967289,32'd4294967295,32'd4294967294,32'd0,32'd4294967292,32'd4294967292,32'd1,32'd6,32'd4294967294,32'd10,32'd41,32'd4294967289,32'd1,32'd4294967290,32'd4294967288,32'd4294967293,32'd4294967295,32'd2,32'd3,32'd1,32'd4294967293,32'd4294967293,32'd4294967290,32'd2,32'd4294967295,32'd4294967294,32'd4294967294,32'd4294967295,32'd0,32'd9,32'd4294967292,32'd2,32'd4294967293,32'd4294967290,32'd4294967293,32'd4294967293,32'd4294967291,32'd2,32'd4294967295,32'd4294967291,32'd4294967289,32'd4294967293,32'd4,32'd4294967295,32'd1,32'd10,32'd4294967295,32'd11,32'd4294967293,32'd0,32'd0,32'd3,32'd4294967282,32'd7,32'd1,32'd4294967294,32'd0,32'd4294967293,32'd1,32'd4294967294,32'd4294967286,32'd3,32'd8,32'd4294967287,32'd4294967286,32'd5,32'd1,32'd1,32'd4,32'd2,32'd4294967280,32'd4294967294,32'd4294967294,32'd4294967294,32'd4294967283,32'd3,32'd4294967294,32'd4294967292,32'd2,32'd4294967295,32'd4294967291,32'd3,32'd2,32'd3,32'd3,32'd4294967288,32'd4294967294,32'd13,32'd5,32'd4294967279,32'd4294967295,32'd4294967285,32'd0,32'd33,32'd6,32'd4294967292,32'd5,32'd4294967286,32'd4294967292,32'd4294967291,32'd0,32'd4294967295,32'd4294967287,32'd0,32'd4294967294,32'd1,32'd1,32'd4294967295,32'd11,32'd4294967291,32'd4294967289,32'd8,32'd0,32'd4294967294,32'd4294967282,32'd4294967271,32'd4294967292,32'd1,32'd4294967293,32'd4294967295,32'd4,32'd4294967285,32'd0,32'd2,32'd2,32'd4294967289,32'd4294967294,32'd4294967295,32'd0,32'd4294967285,32'd4294967278,32'd4294967293,32'd4294967295,32'd4294967278,32'd0,32'd4294967294,32'd2,32'd5,32'd5,32'd6,32'd3,32'd2,32'd4294967291,32'd14,32'd4294967293,32'd4294967289,32'd4294967293,32'd6,32'd4,32'd4,32'd0,32'd1,32'd8,32'd4,32'd1,32'd4294967288,32'd4294967290,32'd2,32'd4294967289,32'd4294967290,32'd4,32'd1,32'd3,32'd10,32'd4294967293,32'd4294967255,32'd7,32'd22,32'd2,32'd7,32'd4294967295,32'd1,32'd0,32'd0,32'd2,32'd4294967290,32'd4294967295,32'd4294967295,32'd4294967294,32'd4294967295,32'd7,32'd0,32'd0,32'd4,32'd1,32'd44,32'd1,32'd4294967293,32'd3,32'd4294967289,32'd0,32'd4294967291,32'd11,32'd2,32'd4,32'd4294967293,32'd2,32'd10,32'd4294967293,32'd1,32'd0,32'd0,32'd4294967293,32'd1,32'd4294967295,32'd4294967295,32'd1,32'd4294967295,32'd24,32'd5,32'd4294967292,32'd6,32'd2,32'd4294967293,32'd6,32'd4294967282,32'd4294967295,32'd2,32'd1,32'd6,32'd4294967287,32'd3,32'd4294967295,32'd3,32'd4294967291,32'd4294967294,32'd4294967293,32'd9,32'd4294967289,32'd1,32'd3,32'd4,32'd2,32'd1,32'd2,32'd4294967294,32'd4294967295,32'd4294967295,32'd4294967293,32'd4,32'd2,32'd14,32'd4294967295,32'd4294967291,32'd8,32'd1,32'd8,32'd5,32'd7,32'd9,32'd4294967294,32'd28,32'd4294967291,32'd4294967295,32'd4294967293,32'd3,32'd0,32'd4294967289,32'd4294967294,32'd4294967286,32'd4294967294,32'd17,32'd4294967295,32'd0,32'd5,32'd4294967293,32'd4294967292,32'd11,32'd1,32'd0,32'd4294967291,32'd1,32'd8,32'd4,32'd4294967291,32'd4294967294,32'd4294967294,32'd4,32'd4294967295,32'd4294967294,32'd1,32'd2,32'd12,32'd1,32'd4294967295,32'd4,32'd0,32'd2,32'd4294967291,32'd4294967291,32'd4294967291,32'd6,32'd7,32'd4294967290,32'd20,32'd25,32'd0,32'd9,32'd14,32'd0,32'd1,32'd4294967292,32'd4294967292,32'd6,32'd4294967294,32'd0,32'd6,32'd4294967285,32'd0,32'd4294967295,32'd4294967295,32'd0,32'd6,32'd1,32'd4294967291,32'd0,32'd3,32'd4294967293,32'd4,32'd4294967295,32'd5,32'd1,32'd2,32'd2,32'd5,32'd2,32'd2,32'd4294967280,32'd6,32'd4294967286,32'd3,32'd0,32'd2,32'd4294967290,32'd4294967295,32'd4294967292,32'd4294967293,32'd4294967290,32'd4294967294,32'd4294967293,32'd4294967290,32'd4,32'd9,32'd4294967295,32'd4294967293,32'd4294967293,32'd4294967284,32'd4294967291,32'd4294967295,32'd2,32'd3,32'd4294967295,32'd4,32'd0,32'd3,32'd1,32'd9,32'd4294967281,32'd4294967281,32'd4294967290,32'd4294967291,32'd13,32'd4294967292,32'd0,32'd5,32'd7,32'd4294967290,32'd4294967294,32'd4294967292,32'd1,32'd4294967287,32'd4294967290,32'd4294967294,32'd3,32'd3,32'd4294967289,32'd3,32'd3,32'd1,32'd4294967295,32'd4294967295,32'd4294967290,32'd0,32'd3,32'd4294967294,32'd4294967286,32'd2,32'd2,32'd4294967294,32'd4294967292,32'd12,32'd1,32'd1,32'd4294967292,32'd4294967295,32'd4294967292,32'd0,32'd0,32'd4294967294,32'd6,32'd4294967295,32'd4294967290,32'd2,32'd4294967293,32'd4294967293,32'd2,32'd4294967291,32'd4294967291,32'd4,32'd4294967290,32'd5,32'd0,32'd4294967294,32'd1,32'd3,32'd4,32'd1,32'd16,32'd4294967292,32'd6,32'd4294967292,32'd8,32'd1,32'd0,32'd0,32'd4294967292,32'd3,32'd2,32'd4294967295,32'd6,32'd4294967295,32'd13,32'd0,32'd7,32'd4294967293,32'd4294967288,32'd4294967289,32'd11,32'd11,32'd3,32'd3,32'd4,32'd4294967294,32'd14,32'd4294967290,32'd22,32'd12,32'd1,32'd3,32'd6,32'd6,32'd4294967292,32'd4294967293,32'd4294967295,32'd4,32'd1,32'd4294967290,32'd0,32'd4294967295,32'd4294967293,32'd2,32'd0,32'd0,32'd4294967295,32'd4294967293,32'd4294967286,32'd13,32'd5,32'd4294967293,32'd4294967287,32'd4294967291,32'd2,32'd4294967292,32'd4294967291,32'd4294967279,32'd4294967291,32'd3,32'd5,32'd4294967281,32'd1,32'd29,32'd4294967289,32'd4294967293,32'd15,32'd22,32'd1,32'd4294967291,32'd1,32'd9,32'd4294967294,32'd4294967294,32'd4294967295,32'd4,32'd2,32'd4294967293,32'd4294967292,32'd8,32'd3,32'd2,32'd4294967294,32'd1,32'd23,32'd4294967287,32'd1,32'd15,32'd4294967281,32'd4,32'd4294967294,32'd4294967286,32'd5,32'd4294967294,32'd3,32'd0,32'd6,32'd2,32'd1,32'd4,32'd4294967291,32'd4294967294,32'd4294967293,32'd4294967295,32'd4294967292,32'd4,32'd4294967294,32'd4294967293,32'd4294967291,32'd0,32'd4,32'd12,32'd3,32'd4294967292,32'd4294967294,32'd4294967295,32'd9,32'd20,32'd4294967293,32'd4294967294,32'd4294967293,32'd0,32'd4294967295,32'd4294967288,32'd4294967293,32'd5,32'd4,32'd4294967294,32'd4294967294,32'd4294967293,32'd1,32'd4294967295,32'd4294967293,32'd4294967290,32'd4294967288,32'd4294967294,32'd4294967293,32'd4294967292,32'd3,32'd4294967293,32'd4294967292,32'd0,32'd3,32'd12,32'd4294967289,32'd2,32'd1,32'd0,32'd0,32'd0,32'd4294967294,32'd4,32'd0,32'd4294967295,32'd4294967295,32'd2,32'd18,32'd2,32'd5,32'd12,32'd21,32'd1,32'd4294967291,32'd4294967293,32'd4294967292,32'd4294967295,32'd4294967295,32'd4294967293,32'd2,32'd4294967288,32'd12,32'd4294967295,32'd0,32'd4294967293,32'd2,32'd7,32'd2,32'd4294967293,32'd4294967293,32'd4294967294,32'd3,32'd7,32'd4294967278,32'd3,32'd4294967292,32'd7,32'd4294967290,32'd0,32'd4294967281,32'd4294967287,32'd4294967288,32'd1,32'd4,32'd10,32'd5,32'd6,32'd3,32'd4294967291,32'd3,32'd4294967295,32'd4294967287,32'd4294967293,32'd4294967294,32'd10,32'd4294967293,32'd3,32'd5,32'd4294967293,32'd6,32'd3,32'd4294967294,32'd4294967294,32'd1,32'd4,32'd0,32'd14,32'd0,32'd4294967291,32'd4294967284,32'd4294967283,32'd4294967294,32'd4294967295,32'd2,32'd0,32'd4294967294,32'd2,32'd3,32'd11,32'd4294967290,32'd2,32'd4294967292,32'd4,32'd4294967289,32'd1,32'd3,32'd3,32'd4294967292,32'd6,32'd1,32'd4,32'd1,32'd4,32'd0,32'd4294967292,32'd3,32'd4294967295,32'd4,32'd4294967294,32'd3,32'd4294967294,32'd3,32'd4294967295,32'd1,32'd4294967292,32'd4294967284,32'd10,32'd1,32'd4294967285,32'd4294967293,32'd5,32'd3,32'd7,32'd4294967290,32'd2,32'd1,32'd8,32'd1,32'd3,32'd4294967291,32'd1,32'd6,32'd12,32'd2,32'd1,32'd1,32'd4294967290,32'd2,32'd4294967294,32'd3,32'd4294967295,32'd4294967295,32'd4294967294,32'd3,32'd1,32'd0,32'd5,32'd12,32'd4294967280,32'd7,32'd0,32'd4294967295,32'd4294967295,32'd4,32'd4294967289,32'd4294967291,32'd4294967258,32'd4294967292,32'd4294967294,32'd4294967289,32'd1,32'd0,32'd7,32'd4294967293,32'd4294967294,32'd4294967293,32'd4294967291,32'd4294967295,32'd7,32'd0,32'd4294967293,32'd1,32'd1,32'd7,32'd2,32'd28,32'd4294967286,32'd4294967291,32'd6,32'd1,32'd42,32'd4294967294,32'd3,32'd11,32'd0,32'd14,32'd29,32'd4294967294,32'd1,32'd7,32'd4,32'd4294967294,32'd4294967293,32'd4294967293,32'd4294967294,32'd12,32'd0,32'd4294967294,32'd4294967294,32'd4294967294,32'd1,32'd54,32'd4294967293,32'd5,32'd9,32'd0,32'd6,32'd6,32'd14,32'd0,32'd4294967293,32'd4294967293,32'd3,32'd4294967293,32'd5,32'd4,32'd4294967293,32'd8,32'd4294967293,32'd4294967283,32'd0,32'd4294967294,32'd4294967290,32'd4294967286,32'd24,32'd3,32'd4294967293,32'd4294967290,32'd3,32'd2,32'd0,32'd4294967293,32'd0,32'd4294967292,32'd4294967290,32'd17,32'd4294967287,32'd2,32'd4294967286,32'd3,32'd8,32'd4294967292,32'd3,32'd5,32'd2,32'd27,32'd4294967295,32'd4294967289,32'd0,32'd4294967294,32'd9,32'd4294967295,32'd4294967294,32'd4294967293,32'd1,32'd2,32'd4294967282,32'd0,32'd4294967292,32'd1,32'd4294967285,32'd4294967294,32'd2,32'd4294967292,32'd4294967295,32'd4294967294,32'd4294967292,32'd0,32'd4294967295,32'd4294967295,32'd1,32'd4294967294,32'd4294967291,32'd4294967293,32'd3,32'd4294967291,32'd4294967284,32'd4294967288,32'd8,32'd1,32'd4294967292,32'd2,32'd4294967292,32'd4,32'd4294967295,32'd4294967292,32'd0,32'd0,32'd4294967293,32'd2,32'd0,32'd4294967293,32'd3,32'd4294967293,32'd4294967294,32'd4294967290,32'd4294967293,32'd2,32'd58,32'd4294967294,32'd4294967293,32'd2,32'd3,32'd4294967291,32'd3,32'd1,32'd3,32'd0,32'd0,32'd4294967288,32'd1,32'd1,32'd4294967279,32'd1,32'd3,32'd4294967291,32'd4294967291,32'd4294967294,32'd6,32'd5,32'd1,32'd4294967284,32'd2,32'd7,32'd6,32'd4294967291,32'd4294967290,32'd1,32'd4294967292,32'd3,32'd5,32'd4294967294,32'd13,32'd2,32'd4294967293,32'd4294967290,32'd2,32'd5,32'd4294967292,32'd1,32'd4294967293,32'd7,32'd10,32'd1,32'd0,32'd4,32'd4294967295,32'd4294967289,32'd4294967292,32'd2,32'd7,32'd13,32'd4294967295,32'd4294967295,32'd1,32'd1,32'd4294967293,32'd2,32'd5,32'd1,32'd4294967293,32'd1,32'd2,32'd4294967295,32'd4294967293,32'd4294967291,32'd7,32'd4294967292,32'd1,32'd4294967291,32'd4294967295,32'd4294967295,32'd2,32'd4294967282,32'd4294967290,32'd4294967293,32'd4294967287,32'd4294967293,32'd3,32'd4294967295,32'd1,32'd4294967294,32'd4294967291,32'd4294967293,32'd4294967295,32'd4294967295,32'd1,32'd4,32'd2,32'd1,32'd4294967293,32'd3,32'd4294967292,32'd4,32'd0,32'd0,32'd1,32'd10,32'd3,32'd1,32'd1,32'd3,32'd4294967292,32'd3,32'd4294967295,32'd5,32'd14,32'd2,32'd0,32'd3,32'd7,32'd4294967295,32'd4294967291,32'd3,32'd4294967293,32'd1,32'd4294967293,32'd4294967291,32'd0,32'd5,32'd4294967294,32'd4,32'd0,32'd0,32'd4,32'd4294967287,32'd4,32'd3,32'd4294967290,32'd1,32'd4294967295,32'd4294967294,32'd4294967292,32'd5,32'd4,32'd4294967295,32'd7,32'd4294967279,32'd4294967295,32'd1,32'd4294967288,32'd4294967292,32'd4294967287,32'd20,32'd4294967291,32'd1,32'd3,32'd7,32'd2,32'd4294967292,32'd10,32'd11,32'd4294967294,32'd6,32'd4294967284,32'd10,32'd4294967295,32'd4294967282,32'd7,32'd0,32'd4,32'd4294967294,32'd3,32'd4294967285,32'd3,32'd4294967295,32'd3,32'd6,32'd4294967285,32'd4294967291,32'd8,32'd2,32'd2,32'd4294967293,32'd0,32'd6,32'd4,32'd4294967293,32'd4294967290,32'd1,32'd0,32'd1,32'd6,32'd1,32'd4294967294,32'd1,32'd5,32'd4294967290,32'd0,32'd4294967294,32'd4294967294,32'd4294967293,32'd4294967292,32'd4294967290,32'd2,32'd4294967295,32'd16,32'd4294967295,32'd7,32'd2,32'd15,32'd0,32'd4294967290,32'd1,32'd3,32'd4294967295,32'd4294967295,32'd0,32'd4294967292,32'd14,32'd8,32'd4294967293,32'd2,32'd3,32'd4294967294,32'd4294967294,32'd4294967293,32'd4294967245,32'd5,32'd4294967295,32'd2,32'd1,32'd4294967289,32'd3,32'd0,32'd4294967288,32'd0,32'd4294967292,32'd4,32'd0,32'd2,32'd12,32'd4294967295,32'd4294967290,32'd20,32'd15,32'd4294967294,32'd4294967286,32'd4294967291,32'd3,32'd11,32'd3,32'd4294967294,32'd1,32'd4294967293,32'd1,32'd4294967293,32'd4294967294,32'd4294967294,32'd4294967294,32'd13,32'd10,32'd4294967294,32'd6,32'd5,32'd6,32'd4,32'd4294967291,32'd0,32'd4294967293,32'd3,32'd4294967295,32'd2,32'd4294967293,32'd4294967291,32'd1,32'd0,32'd13,32'd0,32'd2,32'd4294967294,32'd4,32'd3,32'd4294967292,32'd4294967291,32'd0,32'd4294967294,32'd5,32'd0,32'd0,32'd0,32'd2,32'd4294967293,32'd15,32'd4,32'd4294967293,32'd4294967291,32'd0,32'd4294967293,32'd7,32'd4294967289,32'd4294967294,32'd4294967289,32'd0,32'd2,32'd4294967295,32'd4,32'd4,32'd6,32'd0,32'd6,32'd4294967294,32'd8,32'd4294967290,32'd4294967295,32'd4294967294,32'd4294967289,32'd4294967295,32'd4294967292,32'd4294967293,32'd1,32'd5,32'd15,32'd0,32'd4294967280,32'd4294967294,32'd7,32'd3,32'd5,32'd70,32'd12,32'd4294967295,32'd4294967294,32'd4294967285,32'd0,32'd3,32'd10,32'd4294967290,32'd0,32'd4,32'd4,32'd2,32'd4294967294,32'd4294967293,32'd7,32'd4294967295,32'd4,32'd1,32'd3,32'd0,32'd4294967291,32'd4294967294,32'd3,32'd1,32'd6,32'd4294967289,32'd4294967295,32'd7,32'd4294967290,32'd1,32'd2,32'd17,32'd4294967285,32'd4294967293,32'd1,32'd4294967289,32'd4294967293,32'd4294967293,32'd3,32'd1,32'd4294967293,32'd4294967287,32'd7,32'd4294967295,32'd4294967289,32'd4294967285,32'd4294967289,32'd4294967293,32'd4294967294,32'd4294967295,32'd4294967279,32'd11,32'd4294967292,32'd0,32'd6,32'd0,32'd4294967295,32'd4294967293,32'd6,32'd4294967295,32'd8,32'd4294967293,32'd27,32'd4294967295,32'd1,32'd2,32'd4294967294,32'd1,32'd4294967288,32'd4294967295,32'd16,32'd4294967291,32'd4294967292,32'd4294967288,32'd4294967289,32'd3,32'd1,32'd0,32'd4294967293,32'd3,32'd1,32'd1,32'd4,32'd4294967294,32'd0,32'd1,32'd2,32'd4294967295,32'd1,32'd4,32'd4,32'd6,32'd0,32'd4,32'd1,32'd2,32'd4294967294,32'd5,32'd4,32'd6,32'd2,32'd4,32'd5,32'd10,32'd4294967294,32'd2,32'd21,32'd2,32'd6,32'd3,32'd4294967294,32'd4294967289,32'd1,32'd4,32'd2,32'd4294967294,32'd4294967284,32'd3,32'd1,32'd3,32'd4294967290,32'd24,32'd4294967290,32'd3,32'd4294967293,32'd4294967287,32'd9,32'd4294967295,32'd4294967287,32'd4294967289,32'd4,32'd1,32'd1,32'd12,32'd4294967294,32'd1,32'd4294967289,32'd10,32'd0,32'd1,32'd9,32'd4294967275,32'd4294967293,32'd8,32'd5,32'd5,32'd6,32'd4294967288,32'd11,32'd0,32'd4,32'd2,32'd0,32'd4294967294,32'd5,32'd4294967294,32'd4294967292,32'd4294967292,32'd2,32'd4294967295,32'd4294967293,32'd4294967293,32'd2,32'd4294967291,32'd2,32'd2,32'd4294967294,32'd1,32'd2,32'd4294967287,32'd4294967273,32'd29,32'd2,32'd4294967284,32'd7,32'd0,32'd4294967292,32'd3,32'd3,32'd3,32'd0,32'd4294967288,32'd4294967290,32'd4294967294,32'd4294967295,32'd4294967291,32'd4294967294,32'd4294967293,32'd4294967295,32'd4294967294,32'd2,32'd0,32'd4294967294,32'd4294967292,32'd12,32'd2,32'd4294967293,32'd4294967293,32'd4294967295,32'd4294967291,32'd3,32'd4294967295,32'd0,32'd2,32'd3,32'd12,32'd4,32'd4294967294,32'd2,32'd4294967293,32'd4294967294,32'd1,32'd4294967295,32'd7,32'd4294967294,32'd3,32'd1,32'd4294967281,32'd6,32'd4294967295,32'd4294967283,32'd4294967294,32'd4294967295,32'd4294967294,32'd2,32'd18,32'd1,32'd4,32'd2,32'd2,32'd0,32'd7,32'd1,32'd4294967293,32'd3,32'd1,32'd24,32'd0,32'd4294967292,32'd4294967291,32'd4294967292,32'd1,32'd1,32'd1,32'd1,32'd2,32'd4294967295,32'd7,32'd4294967290,32'd4294967294,32'd4294967293,32'd4294967280,32'd4294967290,32'd4294967290,32'd4294967280,32'd4294967282,32'd4294967290,32'd4294967290,32'd0,32'd2,32'd4,32'd0,32'd3,32'd4294967284,32'd1,32'd4294967292,32'd4294967291,32'd0,32'd4294967295,32'd4294967295,32'd4,32'd4294967293,32'd3,32'd4294967292,32'd7,32'd4,32'd4294967293,32'd4,32'd2,32'd4294967290,32'd8,32'd4294967295,32'd6,32'd4294967292,32'd4,32'd1,32'd4294967289,32'd4294967295,32'd4294967292,32'd4294967295,32'd1,32'd4,32'd5,32'd0,32'd4294967293,32'd4294967293,32'd9,32'd4294967294,32'd4294967288,32'd4294967291,32'd4294967292,32'd5,32'd2,32'd26,32'd3,32'd5,32'd4294967292,32'd4294967295,32'd5,32'd4294967293,32'd4294967293,32'd4294967294,32'd2,32'd8,32'd4294967293,32'd4294967293,32'd6,32'd4294967293,32'd4294967292,32'd2,32'd4294967295,32'd4294967284,32'd4294967291,32'd4,32'd1,32'd5,32'd4294967293,32'd35,32'd0,32'd1,32'd4294967288,32'd4294967278,32'd6,32'd4294967291,32'd4294967295,32'd4294967285,32'd4294967293,32'd4294967294,32'd4294967291,32'd4294967291,32'd4294967295,32'd4294967294,32'd3,32'd4294967288,32'd4294967287,32'd4294967293,32'd1,32'd1,32'd4294967294,32'd23,32'd4294967290,32'd4294967292,32'd4294967287,32'd15,32'd12,32'd4294967259,32'd0,32'd3,32'd4294967291,32'd13,32'd1,32'd4294967294,32'd4294967293,32'd2,32'd4294967286,32'd4294967284,32'd0,32'd0,32'd2,32'd4294967292,32'd0,32'd4294967293,32'd4294967291,32'd6,32'd4294967295,32'd4294967291,32'd4294967288,32'd4294967292,32'd12,32'd1,32'd4294967295,32'd4294967295,32'd5,32'd4294967295,32'd11,32'd4294967290,32'd1,32'd2,32'd4294967290,32'd4,32'd1,32'd2,32'd7,32'd3,32'd2,32'd4,32'd18,32'd4294967294,32'd4294967290,32'd36,32'd3,32'd1,32'd4294967295,32'd13,32'd1,32'd4,32'd0,32'd4294967286,32'd4294967292,32'd4,32'd4294967295,32'd4294967287,32'd4294967286,32'd2,32'd10,32'd4294967294,32'd4294967295,32'd21,32'd1,32'd42,32'd4294967293,32'd7,32'd5,32'd12,32'd0,32'd4294967286,32'd4294967292,32'd4294967294,32'd4,32'd7,32'd1,32'd4294967295,32'd4294967295,32'd4294967292,32'd4294967290,32'd4294967292,32'd4294967290,32'd4294967294,32'd0,32'd5,32'd4294967294,32'd4294967270,32'd5,32'd2,32'd4294967285,32'd0,32'd6,32'd4294967294,32'd3,32'd1,32'd4294967292,32'd3,32'd5,32'd8,32'd3,32'd4294967295,32'd4294967294,32'd3,32'd5,32'd0,32'd1,32'd4,32'd4,32'd0,32'd4294967291,32'd4294967292,32'd5,32'd4294967295,32'd6,32'd3,32'd2,32'd4294967295,32'd18,32'd4294967292,32'd2,32'd2,32'd4,32'd2,32'd4294967284,32'd17,32'd4294967290,32'd0,32'd7,32'd19,32'd4294967294,32'd4294967277,32'd4294967292,32'd4294967288,32'd4294967290,32'd4294967295,32'd0,32'd4294967295,32'd1,32'd2,32'd4294967292,32'd0,32'd4294967293,32'd4294967292,32'd4294967293,32'd4294967294,32'd4294967288,32'd4294967294,32'd4294967292,32'd4294967293,32'd0,32'd4294967293,32'd4294967291,32'd4294967295,32'd4294967293,32'd1,32'd3,32'd4,32'd4294967294,32'd4294967295,32'd4294967291,32'd4294967294,32'd4294967294,32'd4294967267,32'd4294967289,32'd1,32'd1,32'd0,32'd5,32'd4294967295,32'd3,32'd4294967290,32'd4294967294,32'd5,32'd4294967295,32'd4294967283,32'd4294967293,32'd4294967295,32'd0,32'd0,32'd8,32'd5,32'd0,32'd0,32'd4294967293,32'd0,32'd4294967291,32'd4294967295,32'd2,32'd4294967287,32'd4294967289,32'd5,32'd4294967294,32'd2,32'd6,32'd2,32'd2,32'd6,32'd2,32'd4294967294,32'd4294967292,32'd4294967293,32'd8,32'd4294967288,32'd4294967269,32'd17,32'd4294967287,32'd4294967291,32'd7,32'd6,32'd16,32'd4294967295,32'd4294967295,32'd2,32'd4294967293,32'd3,32'd4294967294,32'd4294967295,32'd7,32'd6,32'd0,32'd3,32'd4294967288,32'd4294967291,32'd4294967293,32'd2,32'd4294967293,32'd4294967294,32'd4294967295,32'd4294967295,32'd4294967295,32'd4294967282,32'd4,32'd4294967295,32'd4294967289,32'd0,32'd4294967291,32'd4294967291,32'd0,32'd4,32'd1,32'd3,32'd4,32'd1,32'd1,32'd0,32'd1,32'd1,32'd8,32'd4294967292,32'd0,32'd4294967295,32'd4294967291,32'd4294967294,32'd3,32'd2,32'd3,32'd1,32'd4,32'd4,32'd1,32'd4294967282,32'd0,32'd2,32'd1,32'd1,32'd4294967295,32'd2,32'd1,32'd4294967294,32'd30,32'd9,32'd4294967292,32'd2,32'd0,32'd3,32'd4294967290,32'd2,32'd4294967295,32'd3,32'd0,32'd1,32'd4294967292,32'd4294967288,32'd4294967293,32'd5,32'd4294967290,32'd4294967292,32'd8,32'd4294967295,32'd23,32'd4294967273,32'd4294967294,32'd7,32'd3,32'd5,32'd4294967294,32'd4294967292,32'd0,32'd5,32'd1,32'd8,32'd4294967287,32'd4294967290,32'd4,32'd3,32'd4294967294,32'd0,32'd4,32'd0,32'd2,32'd2,32'd12,32'd4,32'd4294967290,32'd4294967290,32'd9,32'd0,32'd15,32'd0,32'd3,32'd4294967286,32'd4294967293,32'd4294967290,32'd0,32'd4294967295,32'd0,32'd4294967294,32'd4294967291,32'd33,32'd11,32'd0,32'd2,32'd4294967292,32'd4294967294,32'd2,32'd4294967293,32'd4294967293,32'd4294967294,32'd4294967291,32'd1,32'd3,32'd4294967292,32'd4294967292,32'd3,32'd4,32'd10,32'd4294967295,32'd4294967294,32'd0,32'd4294967293,32'd4294967295,32'd4294967295,32'd4,32'd0,32'd4,32'd1,32'd4294967293,32'd1,32'd1,32'd11,32'd0,32'd10,32'd24,32'd5,32'd4294967287,32'd4294967294,32'd4294967295,32'd4294967293,32'd2,32'd0,32'd7,32'd6,32'd4294967295,32'd3,32'd3,32'd4294967292,32'd3,32'd4294967279,32'd0,32'd4294967291,32'd4294967288,32'd4294967295,32'd4294967291,32'd4,32'd4294967295,32'd2,32'd4294967291,32'd1,32'd4294967260,32'd3,32'd2,32'd1,32'd1,32'd19,32'd2,32'd4294967288,32'd4294967290,32'd3,32'd0,32'd4294967286,32'd4,32'd0,32'd4294967295,32'd5,32'd2,32'd2,32'd48,32'd4294967291,32'd4294967289,32'd15,32'd0,32'd11,32'd4294967290,32'd4294967287,32'd6,32'd6,32'd4294967295,32'd4,32'd0,32'd2,32'd2,32'd4,32'd9,32'd12,32'd1,32'd2,32'd4294967278,32'd4294967293,32'd2,32'd4294967295,32'd4294967295,32'd2,32'd1,32'd4294967294,32'd5,32'd12,32'd3,32'd3,32'd4294967293,32'd1,32'd4294967294,32'd0,32'd13,32'd2,32'd1,32'd3,32'd2,32'd4294967292}
`define FEATURE_ABOVE {32'd0,32'd215,32'd28,32'd4294967292,32'd4294967157,32'd4294967181,32'd15,32'd111,32'd44,32'd4294967275,32'd23,32'd4294967183,32'd4294967265,32'd4294967276,32'd88,32'd4294967273,32'd4294967230,32'd81,32'd27,32'd4294967243,32'd18,32'd4294967293,32'd4294967291,32'd75,32'd4294967241,32'd35,32'd16,32'd4294967273,32'd10,32'd4294967189,32'd15,32'd60,32'd10,32'd202,32'd19,32'd4294967237,32'd4294967284,32'd51,32'd4294967264,32'd8,32'd85,32'd4294967288,32'd7,32'd4294967159,32'd20,32'd4294967272,32'd11,32'd15,32'd51,32'd4294967277,32'd4294967268,32'd4294967231,32'd15,32'd0,32'd86,32'd38,32'd25,32'd4294967288,32'd71,32'd4294967278,32'd4294967258,32'd23,32'd40,32'd43,32'd62,32'd4294967220,32'd4294967184,32'd92,32'd10,32'd4294967178,32'd4294967249,32'd10,32'd10,32'd4294967276,32'd26,32'd37,32'd22,32'd4294967278,32'd33,32'd4294967122,32'd4294967289,32'd76,32'd4294967184,32'd4294967291,32'd0,32'd19,32'd200,32'd4294967293,32'd4294967163,32'd34,32'd54,32'd4294967167,32'd9,32'd4294967237,32'd4294967212,32'd4294967274,32'd53,32'd4294967249,32'd36,32'd4294967276,32'd46,32'd4294967269,32'd9,32'd56,32'd4,32'd51,32'd59,32'd4294967293,32'd4294967293,32'd4294967266,32'd18,32'd4294967273,32'd11,32'd4294967256,32'd4294967295,32'd4294967121,32'd17,32'd19,32'd8,32'd0,32'd4294967229,32'd4294967275,32'd0,32'd53,32'd4294967201,32'd45,32'd22,32'd40,32'd8,32'd4294967215,32'd16,32'd4294967292,32'd4294967230,32'd4294967271,32'd116,32'd4294967270,32'd50,32'd16,32'd4294967295,32'd4294967208,32'd40,32'd140,32'd4294967294,32'd4294967292,32'd41,32'd4294967113,32'd4294967284,32'd4294967290,32'd4294967283,32'd4294967289,32'd4294967054,32'd229,32'd18,32'd4294967268,32'd7,32'd4294967270,32'd18,32'd4294967237,32'd105,32'd4294967272,32'd26,32'd4294967250,32'd4294967284,32'd4294967086,32'd32,32'd122,32'd25,32'd7,32'd24,32'd27,32'd4294967292,32'd4294967294,32'd25,32'd4294967216,32'd21,32'd40,32'd24,32'd4294967290,32'd28,32'd4294967263,32'd25,32'd4294967258,32'd109,32'd4294967186,32'd115,32'd18,32'd4294967279,32'd4294967265,32'd95,32'd4294967205,32'd33,32'd4294967194,32'd21,32'd4294967196,32'd52,32'd4294967257,32'd4294967215,32'd54,32'd28,32'd4294967237,32'd4294967245,32'd82,32'd4294967288,32'd44,32'd4294967177,32'd62,32'd3,32'd4294967218,32'd34,32'd36,32'd24,32'd41,32'd4294967106,32'd4294967024,32'd4294967269,32'd54,32'd4294967288,32'd5,32'd122,32'd24,32'd4294967272,32'd14,32'd49,32'd150,32'd4294967158,32'd71,32'd4294967275,32'd17,32'd1,32'd21,32'd4294967188,32'd4294967288,32'd3,32'd4294967294,32'd4294967291,32'd4294967094,32'd57,32'd4294967245,32'd90,32'd4294967090,32'd4294967025,32'd4294967174,32'd4294967270,32'd4294967290,32'd167,32'd4294967041,32'd4294967276,32'd4294966934,32'd6,32'd34,32'd4294967266,32'd26,32'd4294967178,32'd4294967290,32'd56,32'd46,32'd0,32'd6,32'd43,32'd5,32'd4294967115,32'd14,32'd4294967231,32'd314,32'd4294967214,32'd4294966679,32'd4294967154,32'd16,32'd4294967274,32'd21,32'd10,32'd4294967283,32'd4294967267,32'd15,32'd27,32'd36,32'd4294967289,32'd4294967251,32'd4294967172,32'd7,32'd35,32'd134,32'd0,32'd25,32'd191,32'd4294967179,32'd14,32'd4294967288,32'd80,32'd306,32'd4294967273,32'd22,32'd9,32'd33,32'd60,32'd7,32'd4294967264,32'd35,32'd84,32'd37,32'd325,32'd4294967295,32'd4294967294,32'd4294967260,32'd4294967275,32'd23,32'd4294967113,32'd4294967053,32'd9,32'd1,32'd6,32'd66,32'd4294967267,32'd4294967255,32'd4294967197,32'd4294967232,32'd34,32'd4294967259,32'd4294967268,32'd45,32'd4294967230,32'd29,32'd4294967272,32'd4294967273,32'd4294967277,32'd31,32'd57,32'd79,32'd4294967049,32'd23,32'd79,32'd0,32'd66,32'd46,32'd4294967262,32'd7,32'd4294967291,32'd77,32'd4294967291,32'd4294967277,32'd4294967290,32'd4294967104,32'd38,32'd42,32'd4294967291,32'd4294967218,32'd4294967125,32'd4294967188,32'd4294967256,32'd11,32'd4294967293,32'd4294967176,32'd4294967257,32'd4294967288,32'd128,32'd39,32'd4294967273,32'd27,32'd45,32'd83,32'd4294967211,32'd29,32'd4294967271,32'd24,32'd4294967264,32'd20,32'd4294967290,32'd4294963456,32'd4294967272,32'd10,32'd4,32'd31,32'd4294967237,32'd24,32'd4294967203,32'd4294967268,32'd4294967267,32'd88,32'd53,32'd6,32'd69,32'd16,32'd4294967254,32'd62,32'd4294967226,32'd4294967289,32'd4294967291,32'd4294967261,32'd4294967294,32'd78,32'd4294967268,32'd20,32'd4294967291,32'd4294967227,32'd4294967292,32'd24,32'd4294967191,32'd4294967252,32'd92,32'd4294967234,32'd4294967265,32'd4294967288,32'd4,32'd44,32'd4294967264,32'd57,32'd36,32'd4294967211,32'd55,32'd58,32'd50,32'd394,32'd8,32'd4294967231,32'd4294967128,32'd67,32'd4294967096,32'd27,32'd7,32'd3,32'd26,32'd138,32'd35,32'd47,32'd14,32'd4294967288,32'd16,32'd4294967277,32'd8,32'd4294967183,32'd28,32'd175,32'd4294967173,32'd1,32'd116,32'd4294967263,32'd4,32'd3,32'd14,32'd83,32'd41,32'd4294967267,32'd4,32'd4294967114,32'd4294967195,32'd76,32'd18,32'd160,32'd54,32'd79,32'd22,32'd4294967277,32'd89,32'd4294967217,32'd20,32'd4294967151,32'd4294967186,32'd4294967271,32'd4294967287,32'd7,32'd4294967273,32'd20,32'd9,32'd65,32'd29,32'd4294967255,32'd2,32'd4294967138,32'd18,32'd4294967270,32'd4294967155,32'd11,32'd12,32'd4294967288,32'd98,32'd145,32'd4294967285,32'd1,32'd14,32'd4294967293,32'd4294967295,32'd4294967175,32'd4294967290,32'd4294967225,32'd20,32'd4294967271,32'd17,32'd3,32'd26,32'd118,32'd7,32'd4294967255,32'd39,32'd89,32'd4294966893,32'd75,32'd17,32'd53,32'd64,32'd4294967160,32'd26,32'd4294967265,32'd32,32'd4294967274,32'd11,32'd4294967295,32'd4294967129,32'd188,32'd4294966845,32'd4294967295,32'd37,32'd4294967290,32'd4294967236,32'd4294967238,32'd4294967290,32'd4294967186,32'd9,32'd4294967262,32'd39,32'd4,32'd23,32'd4294967270,32'd4294967242,32'd4294967294,32'd0,32'd4294967278,32'd0,32'd8,32'd4294967206,32'd4294967288,32'd4294963456,32'd4294967246,32'd31,32'd4294967271,32'd16,32'd1,32'd24,32'd4294967291,32'd4294967281,32'd4294967198,32'd21,32'd4294967271,32'd4294967218,32'd4294967274,32'd112,32'd1,32'd26,32'd4294967275,32'd3,32'd4294967257,32'd91,32'd4294967243,32'd4294967275,32'd4294967294,32'd4294967233,32'd4294967270,32'd22,32'd4294967251,32'd4,32'd52,32'd70,32'd4294967176,32'd4294967289,32'd129,32'd22,32'd140,32'd94,32'd4294967266,32'd76,32'd4294967295,32'd4294967254,32'd4294967271,32'd4294967272,32'd4294967130,32'd30,32'd18,32'd4294967294,32'd4294967294,32'd5,32'd4294967274,32'd4294967225,32'd0,32'd20,32'd33,32'd16,32'd4294967292,32'd29,32'd4294967292,32'd4294967291,32'd12,32'd17,32'd4294967295,32'd4294967224,32'd126,32'd17,32'd4294967242,32'd4294967228,32'd205,32'd4294967258,32'd23,32'd57,32'd4294967182,32'd67,32'd4294967259,32'd4294967277,32'd82,32'd75,32'd50,32'd78,32'd38,32'd4294967260,32'd7,32'd111,32'd12,32'd73,32'd4294967282,32'd4294967108,32'd15,32'd4294967099,32'd4294967232,32'd59,32'd10,32'd25,32'd4294967127,32'd59,32'd8,32'd4294967243,32'd53,32'd4294967277,32'd4294967006,32'd4294967287,32'd18,32'd4294967269,32'd4294967293,32'd4294967201,32'd4294967210,32'd4294967287,32'd4294967281,32'd4294967295,32'd4,32'd130,32'd4294967275,32'd119,32'd15,32'd72,32'd21,32'd22,32'd4294967292,32'd4294967290,32'd4294967094,32'd4294967291,32'd4294967215,32'd4294967194,32'd4294967290,32'd4294967287,32'd6,32'd48,32'd4294967219,32'd293,32'd5,32'd4294967227,32'd50,32'd4294967227,32'd8,32'd4294967278,32'd8,32'd15,32'd4294967218,32'd61,32'd18,32'd4294967190,32'd24,32'd4294967165,32'd15,32'd3,32'd4294967110,32'd65,32'd8,32'd4294967260,32'd68,32'd4294967293,32'd21,32'd24,32'd4294967150,32'd4294967255,32'd97,32'd9,32'd4294967269,32'd4294967225,32'd4294967260,32'd10,32'd58,32'd4294967269,32'd4294967248,32'd9,32'd23,32'd4294967189,32'd42,32'd4294967292,32'd19,32'd4294967253,32'd4294967280,32'd4294967274,32'd4294967239,32'd95,32'd16,32'd4294967164,32'd4294967044,32'd4294967274,32'd4294967193,32'd4294967291,32'd22,32'd4294967244,32'd11,32'd4294967264,32'd2,32'd32,32'd11,32'd4294967260,32'd38,32'd7,32'd26,32'd197,32'd4294967201,32'd97,32'd4294967294,32'd70,32'd21,32'd4294967292,32'd1,32'd4294967276,32'd50,32'd75,32'd4294967114,32'd4294967254,32'd103,32'd4294967266,32'd4294967239,32'd210,32'd8,32'd4294967263,32'd30,32'd4294967259,32'd3,32'd4294967288,32'd41,32'd4294967273,32'd66,32'd4294967172,32'd4,32'd110,32'd30,32'd4294967293,32'd85,32'd4294967132,32'd4,32'd4294967272,32'd95,32'd4294967197,32'd0,32'd4294967254,32'd4294967148,32'd122,32'd66,32'd4294967079,32'd4294967087,32'd4294967250,32'd1,32'd4294967176,32'd32,32'd0,32'd1,32'd4294967166,32'd4294967288,32'd60,32'd2,32'd4294967193,32'd86,32'd4294967269,32'd30,32'd4294967209,32'd27,32'd3,32'd4294967226,32'd4294967183,32'd4294967261,32'd4294967261,32'd40,32'd33,32'd88,32'd51,32'd63,32'd5,32'd4294967143,32'd4294967230,32'd4294967290,32'd3,32'd0,32'd12,32'd4294967252,32'd25,32'd4294967267,32'd4294967225,32'd18,32'd4294967223,32'd25,32'd139,32'd4294967294,32'd4294967209,32'd4294967259,32'd4294967279,32'd38,32'd30,32'd420,32'd24,32'd4294967273,32'd4294967270,32'd89,32'd94,32'd4294967289,32'd11,32'd4294966996,32'd18,32'd83,32'd54,32'd10,32'd18,32'd4294967202,32'd17,32'd2,32'd4294966721,32'd4294967276,32'd21,32'd85,32'd4294967195,32'd4294967275,32'd4294967282,32'd70,32'd36,32'd4294967269,32'd5,32'd4294967273,32'd4294967203,32'd4294967240,32'd15,32'd4294967252,32'd6,32'd4294967289,32'd15,32'd4294967264,32'd89,32'd142,32'd4294967273,32'd8,32'd26,32'd4294967196,32'd37,32'd105,32'd4294967155,32'd124,32'd4294967224,32'd4294967187,32'd34,32'd13,32'd4294967286,32'd4294967274,32'd211,32'd4294967205,32'd4294966969,32'd4294967276,32'd110,32'd4294967287,32'd4294967291,32'd6,32'd33,32'd243,32'd15,32'd11,32'd8,32'd11,32'd4294967167,32'd44,32'd19,32'd4294967273,32'd4294967264,32'd4294967291,32'd0,32'd2,32'd4294967258,32'd4294967224,32'd18,32'd2,32'd17,32'd4294967263,32'd29,32'd4294967270,32'd7,32'd0,32'd104,32'd4294967272,32'd57,32'd4294967289,32'd4294967115,32'd4294967288,32'd4294967288,32'd4294967273,32'd24,32'd4294967290,32'd4294967258,32'd4294967273,32'd6,32'd6,32'd4294967241,32'd4294967248,32'd71,32'd2,32'd19,32'd4294967090,32'd4294967266,32'd4294967255,32'd75,32'd4294967212,32'd44,32'd7,32'd3,32'd4294967184,32'd23,32'd4294967268,32'd28,32'd6,32'd4294967254,32'd4294967191,32'd4294967244,32'd4294967253,32'd7,32'd4294967292,32'd11,32'd18,32'd5,32'd4294967265,32'd29,32'd4294967238,32'd20,32'd77,32'd159,32'd4294967289,32'd51,32'd4294967270,32'd18,32'd4294967265,32'd38,32'd27,32'd4294967170,32'd54,32'd4294967291,32'd4294967294,32'd23,32'd94,32'd4294967276,32'd4294967293,32'd21,32'd9,32'd32,32'd4294967177,32'd21,32'd4294967202,32'd4294967289,32'd4294967295,32'd4294967269,32'd0,32'd17,32'd53,32'd4294967248,32'd4294967262,32'd4294967292,32'd3,32'd4294967168,32'd4294967258,32'd40,32'd62,32'd27,32'd4294967165,32'd16,32'd4294967208,32'd18,32'd38,32'd4294967243,32'd78,32'd4294967260,32'd4294967260,32'd4294967278,32'd0,32'd4294967258,32'd4294967265,32'd15,32'd43,32'd110,32'd4294967277,32'd11,32'd4294967151,32'd4294967275,32'd65,32'd63,32'd0,32'd8,32'd4294967293,32'd4294967293,32'd4294967271,32'd15,32'd4294967243,32'd2,32'd4294967294,32'd4294967272,32'd4294967294,32'd9,32'd4294967151,32'd4294967273,32'd42,32'd4294967256,32'd4294967273,32'd2,32'd4294966862,32'd48,32'd4294967278,32'd4294967292,32'd4294967293,32'd2,32'd4294967134,32'd4294967210,32'd4294967295,32'd4294966998,32'd4294967289,32'd20,32'd4294967266,32'd32,32'd4294967258,32'd14,32'd4294967243,32'd28,32'd16,32'd54,32'd0,32'd69,32'd4294967270,32'd5,32'd144,32'd21,32'd4294967293,32'd16,32'd4294967277,32'd22,32'd41,32'd6,32'd4294967294,32'd4294967292,32'd4294967278,32'd41,32'd34,32'd64,32'd4294967291,32'd4294967293,32'd10,32'd35,32'd4294967266,32'd6,32'd4294967295,32'd27,32'd4294967269,32'd30,32'd4294967291,32'd4294967288,32'd4294967123,32'd4294967253,32'd89,32'd55,32'd34,32'd19,32'd54,32'd19,32'd4294967275,32'd20,32'd182,32'd4294967216,32'd4294967228,32'd26,32'd50,32'd4294967232,32'd39,32'd65,32'd4294967288,32'd4294967288,32'd35,32'd11,32'd4294967287,32'd4294967205,32'd4294967217,32'd4294967219,32'd99,32'd20,32'd4294967287,32'd4294967262,32'd51,32'd49,32'd4294967240,32'd28,32'd8,32'd29,32'd10,32'd24,32'd4,32'd19,32'd4294967252,32'd0,32'd4,32'd4294967164,32'd15,32'd33,32'd4294967169,32'd52,32'd119,32'd54,32'd4294967256,32'd4294967263,32'd4294967294,32'd4294967272,32'd4294967276,32'd4294967080,32'd4294967295,32'd4294967168,32'd4294967289,32'd117,32'd151,32'd18,32'd66,32'd48,32'd4294967219,32'd20,32'd4294967208,32'd24,32'd6,32'd74,32'd4294967257,32'd42,32'd4294967206,32'd4294967293,32'd4294967068,32'd35,32'd4294967274,32'd124,32'd4294967293,32'd4294967290,32'd4294967182,32'd37,32'd65,32'd19,32'd4294967148,32'd4294967287,32'd107,32'd21,32'd0,32'd4294967254,32'd4294967051,32'd18,32'd29,32'd103,32'd4294967184,32'd4294967165,32'd34,32'd70,32'd3,32'd26,32'd4294967251,32'd26,32'd4294967137,32'd66,32'd4294967158,32'd32,32'd4294967268,32'd91,32'd4294967170,32'd59,32'd70,32'd56,32'd78,32'd4294967272,32'd105,32'd4294967291,32'd4294967287,32'd4294967290,32'd4294967278,32'd4,32'd18,32'd4294967271,32'd16,32'd4294967265,32'd4294967011,32'd4294967293,32'd4294967285,32'd4294967198,32'd4294967292,32'd4294967288,32'd4294966687,32'd56,32'd42,32'd4294967292,32'd39,32'd4294967202,32'd4294967209,32'd4294967279,32'd7,32'd4294967262,32'd4294967235,32'd4294967272,32'd4,32'd20,32'd4294967237,32'd4294967079,32'd4294967244,32'd4294967267,32'd48,32'd3,32'd74,32'd4294967289,32'd17,32'd4294967277,32'd4294967096,32'd69,32'd18,32'd267,32'd369,32'd4294967242,32'd73,32'd4294967165,32'd4294967262,32'd61,32'd4294967295,32'd4294967274,32'd41,32'd1,32'd4294967274,32'd62,32'd1,32'd4294967253,32'd0,32'd5,32'd32,32'd79,32'd4294967269,32'd7,32'd29,32'd4294967156,32'd19,32'd79,32'd4294967279,32'd95,32'd53,32'd4294967218,32'd4294967235,32'd101,32'd69,32'd4294967209,32'd18,32'd43,32'd12,32'd86,32'd36,32'd4294967238,32'd19,32'd1,32'd18,32'd4294967295,32'd11,32'd4294967270,32'd20,32'd4294967291,32'd4294967251,32'd61,32'd22,32'd4294967277,32'd1,32'd4294967290,32'd4,32'd4294967292,32'd4294967218,32'd41,32'd4294967280,32'd69,32'd29,32'd4294967178,32'd49,32'd4294967042,32'd21,32'd4,32'd4,32'd4294967266,32'd82,32'd3,32'd4294967261,32'd115,32'd77,32'd4294967291,32'd4294967270,32'd4294967266,32'd32,32'd4294967265,32'd6,32'd4,32'd49,32'd4294967186,32'd12,32'd4294967175,32'd4294967265,32'd18,32'd31,32'd4294967261,32'd22,32'd4,32'd4294967217,32'd4294967265,32'd17,32'd60,32'd32,32'd4,32'd19,32'd4294967157,32'd66,32'd4294967203,32'd18,32'd4294967262,32'd29,32'd13,32'd34,32'd4294967263,32'd4294967180,32'd1,32'd20,32'd54,32'd4294967286,32'd3,32'd103,32'd4294967271,32'd29,32'd4294967191,32'd5,32'd23,32'd30,32'd12,32'd53,32'd65,32'd78,32'd28,32'd77,32'd4294967221,32'd64,32'd10,32'd4294967233,32'd67,32'd9,32'd27,32'd4294967267,32'd39,32'd4294967218,32'd22,32'd33,32'd4294967281,32'd4294967115,32'd27,32'd4294967063,32'd0,32'd4294967291,32'd25,32'd93,32'd4294967121,32'd4294967204,32'd100,32'd4294967022,32'd19,32'd4294966976,32'd9,32'd4294967207,32'd126,32'd4294967154,32'd50,32'd4294967058,32'd4294967145,32'd4294967295,32'd0,32'd4294967259,32'd4294967205,32'd51,32'd17,32'd6,32'd27,32'd4294967277,32'd4294967210,32'd4,32'd33,32'd4294967250,32'd28,32'd4294967295,32'd98,32'd4294967199,32'd2,32'd4294967277,32'd4294967274,32'd4294967189,32'd22,32'd4294967266,32'd14,32'd4294967261,32'd47,32'd4294967188,32'd9,32'd25,32'd139,32'd4294967270,32'd2,32'd4294967168,32'd4294967099,32'd21,32'd23,32'd43,32'd1280,32'd4294967255,32'd4294967289,32'd5,32'd45,32'd44,32'd0,32'd4294967293,32'd4294967179,32'd45,32'd4294967247,32'd4294967274,32'd4294967247,32'd4294967155,32'd2,32'd11,32'd4294967024,32'd4294967273,32'd4294967215,32'd4294967289,32'd16,32'd74,32'd4294967288,32'd4294967197,32'd41,32'd4294967204,32'd48,32'd4294967219,32'd129,32'd4294967292,32'd22,32'd4294967269,32'd31,32'd4294967274,32'd4294967165,32'd4294967255,32'd30,32'd2,32'd4294967248,32'd58,32'd4294967125,32'd4294967159,32'd22,32'd4294967265,32'd4294967289,32'd4294967145,32'd133,32'd4294967262,32'd19,32'd6,32'd26,32'd4294967258,32'd0,32'd4294967294,32'd4294967233,32'd4294967117,32'd4294967284,32'd2,32'd20,32'd4294967219,32'd28,32'd4294967266,32'd19,32'd4294967272,32'd28,32'd4294967269,32'd23,32'd4294967193,32'd22,32'd0,32'd57,32'd50,32'd4294967179,32'd4294967272,32'd54,32'd4294967211,32'd31,32'd15,32'd35,32'd31,32'd35,32'd4294967208,32'd4294967222,32'd4294967215,32'd51,32'd98,32'd63,32'd4294967025,32'd250,32'd4294967236,32'd4294967215,32'd16,32'd4294967294,32'd18,32'd4294967268,32'd4,32'd4294967270,32'd4294967242,32'd4294967277,32'd4294967156,32'd11,32'd35,32'd4294967270,32'd52,32'd4294967010,32'd4294967259,32'd4294967295,32'd9,32'd2,32'd4294967268,32'd64,32'd4294967293,32'd69,32'd1,32'd62,32'd17,32'd4294967229,32'd17,32'd4294967274,32'd4,32'd14,32'd4294967209,32'd200,32'd4294967104,32'd4294967176,32'd4294967145,32'd4294967290,32'd126,32'd3,32'd14,32'd4294967276,32'd24,32'd4294967047,32'd25,32'd4294967249,32'd4294967216,32'd4294967261,32'd4294966921,32'd4294967155,32'd24,32'd4294967262,32'd85,32'd4294967153,32'd37,32'd93,32'd32,32'd4294967267,32'd26,32'd4294967288,32'd4294967295,32'd4294967267,32'd101,32'd4294967252,32'd20,32'd4294967213,32'd54,32'd4294967187,32'd21,32'd15,32'd10,32'd4294967156,32'd15,32'd31,32'd90,32'd56,32'd4294967288,32'd4294967238,32'd90,32'd4294967126,32'd38,32'd4294967149,32'd4294967262,32'd4,32'd4294967259,32'd4294967263,32'd4294967199,32'd4294967270,32'd32,32'd4294967261,32'd73,32'd4294967293,32'd77,32'd4294967269,32'd23,32'd76,32'd37,32'd4294967272,32'd4294967292,32'd128,32'd4294967200,32'd79,32'd18,32'd4294967147,32'd4294967282,32'd4294967039,32'd62,32'd44,32'd18,32'd20,32'd348,32'd4294967133,32'd4294967231,32'd4294967187,32'd79,32'd0,32'd4294967162,32'd4294967269,32'd4294967210,32'd10,32'd30,32'd4294967295,32'd67,32'd39,32'd4294967200,32'd4294967170,32'd4294966789,32'd4294967277,32'd4294967153,32'd5,32'd29,32'd2,32'd4294967151,32'd4294967270,32'd4294967290,32'd4294967291,32'd4294967282,32'd4294967239,32'd23,32'd53,32'd42,32'd151,32'd20,32'd5,32'd26,32'd4294967270,32'd4294967256,32'd4294967141,32'd35,32'd4294967247,32'd40,32'd29,32'd97,32'd4294967132,32'd116,32'd4294967210,32'd4294967270,32'd4294967087,32'd41,32'd4294967164,32'd5,32'd4294967274,32'd68,32'd4294967275,32'd70,32'd4294967131,32'd4294967268,32'd4294967285,32'd102,32'd4294967116,32'd4294967260,32'd4294967294,32'd3,32'd4294967247,32'd4294967061,32'd32,32'd1,32'd22,32'd0,32'd4294967276,32'd4294967060,32'd20,32'd99,32'd160,32'd15,32'd102,32'd52,32'd4294967194,32'd4294967247,32'd29,32'd0,32'd55,32'd4294967269,32'd4294967194,32'd4294967188,32'd0,32'd4294967158,32'd4294967291,32'd4294967289,32'd4294967281,32'd1,32'd16,32'd4294967272,32'd159,32'd4294967151,32'd20,32'd4294967268,32'd75,32'd33,32'd33,32'd0,32'd4294967265,32'd4294967273,32'd22,32'd144,32'd2,32'd22,32'd4,32'd4294967205,32'd4294967158,32'd4294967293,32'd79,32'd90,32'd4294967240,32'd4294966979,32'd4294967277,32'd4294967292,32'd45,32'd0,32'd4294967155,32'd1,32'd18,32'd4294967272,32'd59,32'd142,32'd15,32'd9,32'd22,32'd35,32'd4,32'd2,32'd4294967238,32'd4294967294,32'd27,32'd4294967251,32'd24,32'd17,32'd25,32'd4294967264,32'd103,32'd5,32'd19,32'd4294967293,32'd4294967207,32'd4294967292,32'd19,32'd4294967274,32'd105,32'd16,32'd20,32'd54,32'd20,32'd4294967183,32'd36,32'd8,32'd4294967269,32'd8,32'd4,32'd71,32'd34,32'd4294967261,32'd4294967247,32'd4294967293,32'd4294967276,32'd4294967268,32'd4294967283,32'd39,32'd93,32'd4294967254,32'd0,32'd4294967172,32'd4294967207,32'd5,32'd4294967207,32'd13,32'd110,32'd46,32'd4294967243,32'd3,32'd22,32'd53,32'd4294967258,32'd75,32'd4294967195,32'd4294967272,32'd8,32'd4294967292,32'd100,32'd4294967242,32'd25,32'd4294967294,32'd4294967243,32'd156,32'd4294967208,32'd4294967295,32'd20,32'd28,32'd3,32'd39,32'd44,32'd4294967277,32'd4294966697,32'd4294967148,32'd16,32'd4294967273,32'd4294967251,32'd214,32'd26,32'd26,32'd26,32'd4294967076,32'd4294967136,32'd132,32'd4294967293,32'd4294967070,32'd4294967259,32'd4294967263,32'd22,32'd34,32'd95,32'd4294967045,32'd33,32'd4294967257,32'd4294967265,32'd56,32'd4,32'd4294967158,32'd4294966947,32'd80,32'd18,32'd66,32'd4294967245,32'd11,32'd4294967288,32'd1,32'd81,32'd5,32'd54,32'd4294967294,32'd4294967289,32'd4294967256,32'd68,32'd4294967269,32'd15,32'd4294967293,32'd15,32'd0,32'd4294967118,32'd4294967252,32'd105,32'd4294967272,32'd14,32'd1,32'd4294967274,32'd2,32'd71,32'd59,32'd4294967231,32'd28,32'd17,32'd4294967184,32'd22,32'd4294967135,32'd31,32'd12,32'd43,32'd119,32'd4294967250,32'd50,32'd53,32'd4294967168,32'd25,32'd4294967167,32'd4294967263,32'd123,32'd4294966977,32'd4294967147,32'd43,32'd69,32'd4294967069,32'd4294967263,32'd18,32'd58,32'd30,32'd4294967206,32'd20,32'd4294967294,32'd4294967262,32'd4294967151,32'd4294967236,32'd32,32'd38,32'd4294967229,32'd4294967224,32'd4294967263,32'd42,32'd76,32'd5,32'd4294967198,32'd4294967281,32'd4294967294,32'd27,32'd93,32'd116,32'd10,32'd91,32'd4294967263,32'd24,32'd8,32'd29,32'd4294967253,32'd7,32'd141,32'd4294967270,32'd55,32'd74,32'd73,32'd39,32'd4294967207,32'd248,32'd122,32'd4294967295,32'd206,32'd4294967292,32'd158,32'd4294967230,32'd17,32'd275,32'd24,32'd78,32'd3,32'd4294967053,32'd20,32'd30,32'd4294967249,32'd4294967157,32'd4294967139,32'd4294967289,32'd4294967295,32'd4294967052,32'd73,32'd60,32'd0,32'd4,32'd4294967169,32'd4294967213,32'd23,32'd4294967269,32'd48,32'd4,32'd51,32'd4294967162,32'd33,32'd4294967277,32'd48,32'd4294967125,32'd1,32'd7,32'd20,32'd4294967290,32'd8,32'd4294967294,32'd20,32'd31,32'd2,32'd4294967128,32'd22,32'd4294967173,32'd4294967231,32'd70,32'd4294967200,32'd4294967274,32'd63,32'd4294967168,32'd28,32'd4294967271,32'd27,32'd4294967275,32'd4294967020,32'd163,32'd31,32'd25,32'd46,32'd5,32'd26,32'd4294967268,32'd6,32'd149,32'd4294967286,32'd4294967210,32'd75,32'd4294967271,32'd48,32'd29,32'd14,32'd17,32'd4294967291,32'd184,32'd27,32'd4294967230,32'd4294967237,32'd4294967258,32'd2,32'd71,32'd53,32'd4294967243,32'd19,32'd4294967293,32'd4294967246,32'd4294967102,32'd4294967205,32'd4294967292,32'd4294967258,32'd4294967295,32'd4294967275,32'd4294967259,32'd2,32'd1,32'd6,32'd129,32'd79,32'd4294967266,32'd4294967157,32'd99,32'd118,32'd80,32'd23,32'd4294967234,32'd4294967285,32'd4294967136,32'd4294967265,32'd4294967184,32'd25,32'd4294967293,32'd4294967203,32'd4294967230,32'd4294967124,32'd44,32'd4294967239,32'd6,32'd4294967112,32'd91,32'd1,32'd4294967264,32'd31,32'd4294967260,32'd4294967158,32'd34,32'd34,32'd24,32'd46,32'd4294967210,32'd90,32'd66,32'd4294967271,32'd2,32'd4294967243,32'd0,32'd4294967118,32'd22,32'd4294967295,32'd7,32'd27,32'd112,32'd16,32'd73,32'd4294967154,32'd4294966968,32'd4294967239,32'd68,32'd4294967259,32'd117,32'd4294967293,32'd4294967289,32'd4,32'd12,32'd4294967252,32'd20,32'd4294967266,32'd52,32'd71,32'd76,32'd4294967248,32'd21,32'd4294967258,32'd4294966981,32'd4294967183,32'd98,32'd4294967082,32'd4294967200,32'd6,32'd23,32'd4294967276,32'd27,32'd4294967153,32'd149,32'd4294967292,32'd27,32'd4294967175,32'd75,32'd50,32'd4294967292,32'd4294967295,32'd4294967043,32'd4294967257,32'd4294967174,32'd56,32'd4294967243,32'd4294967236,32'd19,32'd0,32'd4294967205,32'd66,32'd4294967137,32'd4294967294,32'd0,32'd4294967139,32'd4294967294,32'd18,32'd48,32'd4294967099,32'd8,32'd4294967293,32'd4294967219,32'd4294967269,32'd24,32'd4294967267,32'd4294967234,32'd42,32'd21,32'd4294967294,32'd4294966967,32'd4294967245,32'd24,32'd4294967269,32'd4294967294,32'd7,32'd30,32'd4294967294,32'd21,32'd4294967098,32'd23,32'd4294967205,32'd4294967140,32'd51,32'd4294967287,32'd4294967274,32'd137,32'd6,32'd4294967144,32'd4294967267,32'd132,32'd4294967248,32'd77,32'd4294967260,32'd4294967277,32'd49,32'd25,32'd3,32'd4294967170,32'd2,32'd19,32'd4294967267,32'd4,32'd67,32'd4294967269,32'd4294967239,32'd24,32'd4294967097,32'd61,32'd4294967229,32'd74,32'd16,32'd47,32'd26,32'd15,32'd4294967205,32'd25,32'd87,32'd57,32'd73,32'd10,32'd4294967270,32'd4294967184,32'd4294967257,32'd4294967260,32'd67,32'd49,32'd201,32'd4294967216,32'd4294967189,32'd4294967195,32'd4294967164,32'd4294967255,32'd69,32'd4294967090,32'd50,32'd152,32'd4294967091,32'd4294967272,32'd9,32'd99,32'd4294967233,32'd93,32'd2,32'd4294967291,32'd43,32'd4294967200,32'd69,32'd0,32'd89,32'd4294967274,32'd52,32'd4294967258,32'd26,32'd94,32'd4294967275,32'd4294967275,32'd8,32'd4294967204,32'd50,32'd18,32'd4294967130,32'd4294967273,32'd46,32'd4294967291,32'd269,32'd4294967228,32'd4294967247,32'd38,32'd4,32'd4294967292,32'd190,32'd4294967194,32'd72,32'd69,32'd18,32'd4294967143,32'd55,32'd4294967139,32'd4294967212,32'd4294967200,32'd21,32'd68,32'd2,32'd4294967292,32'd17,32'd76,32'd4294967285,32'd4294967294,32'd21,32'd4294967147,32'd25,32'd143,32'd4294967248,32'd6,32'd92,32'd141,32'd4294967291,32'd4294967264,32'd99,32'd27,32'd25,32'd74,32'd33,32'd6,32'd4294967206,32'd72,32'd67,32'd7,32'd23,32'd4294967268,32'd22,32'd6,32'd28,32'd8,32'd28,32'd4294967229,32'd4294967236,32'd4294967173,32'd4294967279,32'd4294967252,32'd20,32'd94,32'd4294967206,32'd4294967260,32'd27,32'd15,32'd4294967292,32'd67,32'd42,32'd4294967153,32'd40,32'd72,32'd129,32'd74,32'd4294967262,32'd48,32'd4294967272,32'd28,32'd24,32'd4294967287,32'd4294967049,32'd4294967284,32'd4294967165,32'd26,32'd4294967270,32'd50,32'd4294967238,32'd15,32'd4294967270,32'd4294967274,32'd3,32'd4294967261,32'd4294967182,32'd25,32'd91,32'd4294967256,32'd17,32'd43,32'd4294967113,32'd32,32'd0,32'd4294967252,32'd3,32'd105,32'd22,32'd5,32'd4294967269,32'd2,32'd53,32'd33,32'd40,32'd86,32'd4294967197,32'd4294967289,32'd4294967074,32'd4294967294,32'd3,32'd25,32'd4294967266,32'd20,32'd4294967261,32'd12,32'd4294967272,32'd4294967295,32'd6,32'd4294967287,32'd104,32'd4294967104,32'd14,32'd61,32'd4294967269,32'd4294967217,32'd0,32'd19,32'd4294967229,32'd4294967279,32'd4,32'd4294967218,32'd4294967264,32'd127,32'd1,32'd96,32'd4294967018,32'd3,32'd4294966955,32'd59,32'd4294967266,32'd125,32'd4294967228,32'd4294967204,32'd5,32'd4294967159,32'd29,32'd26,32'd4294967254,32'd4294967294,32'd8,32'd33,32'd4294967121,32'd4294967188,32'd4294967208,32'd24,32'd6,32'd4294967229,32'd9,32'd26,32'd4294967261,32'd4294967239,32'd68,32'd37,32'd168,32'd74,32'd82,32'd3,32'd4294967268,32'd195,32'd0,32'd3,32'd32,32'd56,32'd4294967238,32'd4294967295,32'd31,32'd4294967086,32'd20,32'd4294967272,32'd35,32'd4294967270,32'd19,32'd4294967268,32'd62,32'd33,32'd4294967110,32'd4294967267,32'd98,32'd4294967247,32'd52,32'd4294967295,32'd15,32'd102,32'd8,32'd4294967247,32'd18,32'd4294967239,32'd4294967290,32'd4294967293,32'd20,32'd4294967253,32'd34,32'd76,32'd4,32'd3,32'd2,32'd4294967210,32'd37,32'd7,32'd4294967140,32'd4294967270,32'd31,32'd4294967295,32'd146,32'd138,32'd4294967294,32'd19,32'd160,32'd4294967268,32'd4294967208,32'd102,32'd4294967288,32'd2,32'd4294967205,32'd4294967291,32'd27,32'd4294967228,32'd4294967261,32'd4294967167,32'd26,32'd4294967227,32'd4294967283,32'd3,32'd4294967085,32'd4294967204,32'd33,32'd1,32'd4294967279,32'd4294967090,32'd4294967245,32'd13,32'd26,32'd4294967108,32'd4294967269,32'd77,32'd17,32'd4294967160,32'd4294967172,32'd4294967254,32'd102,32'd47,32'd49,32'd94,32'd95,32'd52,32'd68,32'd140,32'd4294967263,32'd36,32'd98,32'd4294967162,32'd29,32'd4294967292,32'd4294966949,32'd40,32'd118,32'd30,32'd4294967292,32'd20,32'd4294966996,32'd4294967253,32'd4294967259,32'd19,32'd130,32'd4294967075,32'd9,32'd4294967254,32'd4294967000,32'd32,32'd66,32'd22,32'd4294967160,32'd156,32'd139,32'd4294967258,32'd4294967293,32'd26,32'd4294967250,32'd130,32'd4294967137,32'd4294967213,32'd4294967262,32'd4294967281,32'd4294967293,32'd16,32'd4294967265,32'd6,32'd10,32'd43,32'd90,32'd4294967276,32'd2,32'd156,32'd4294967158,32'd19,32'd34,32'd4294967204,32'd9,32'd4294967244,32'd4294967206,32'd20,32'd4294967169,32'd110,32'd104,32'd4294967200,32'd4294967192,32'd35,32'd4294967122,32'd4294967111,32'd32,32'd48,32'd4294967091,32'd4294967241,32'd32,32'd23,32'd4294967256,32'd121,32'd4294967235,32'd108,32'd86,32'd4294967192,32'd16,32'd4294967075,32'd8,32'd4294967209,32'd58,32'd37,32'd51,32'd4294967217,32'd142,32'd19,32'd42,32'd4294967102,32'd4294967132,32'd4294967273,32'd0,32'd21,32'd4294967292,32'd4294967294,32'd4294967252,32'd4294967283,32'd5,32'd83,32'd196,32'd20,32'd4294967213,32'd40,32'd0,32'd24,32'd4294967242,32'd20,32'd5,32'd19,32'd4294967262,32'd41,32'd5,32'd21,32'd4294967234,32'd4,32'd8,32'd4294967076,32'd135,32'd25,32'd7,32'd31,32'd4294967260,32'd4294967269,32'd4294967264,32'd25,32'd4294967161,32'd91,32'd16,32'd4294967144,32'd8,32'd4294967012,32'd0,32'd24,32'd4294967103,32'd4294967229,32'd4294967295,32'd29,32'd4294967239,32'd56,32'd25,32'd4294967159,32'd4294967118,32'd49,32'd4294967224,32'd30,32'd4294967184,32'd22,32'd4294967221,32'd33,32'd4294967247,32'd34,32'd91,32'd4294967206,32'd65,32'd115,32'd74,32'd38,32'd105,32'd4294967198,32'd8,32'd4294967285,32'd1,32'd4294967053,32'd4294967268,32'd4294967290,32'd157,32'd29,32'd7,32'd4294967137,32'd48,32'd4294967098,32'd9,32'd23,32'd60,32'd31,32'd4294967081,32'd4294967282,32'd4294967247,32'd4294967104,32'd58,32'd4294967189,32'd133,32'd4294967294,32'd4294967255,32'd30,32'd65,32'd25,32'd4294967247,32'd4294967272,32'd13,32'd30,32'd5,32'd4294967082,32'd4294967236,32'd21,32'd55,32'd44,32'd6,32'd4294967237,32'd4294967132,32'd66,32'd4294967028,32'd4294967126,32'd23,32'd4294967171,32'd18,32'd4294967237,32'd76,32'd53,32'd4294967262,32'd4294967236,32'd24,32'd4294967283,32'd29,32'd39,32'd76,32'd4294967136,32'd64,32'd63,32'd122,32'd87,32'd16,32'd48,32'd4294967103,32'd72,32'd81,32'd8,32'd4294967186,32'd4294967161,32'd27,32'd103,32'd4294967213,32'd0,32'd57,32'd4294967227,32'd4294967163,32'd5,32'd4294967168,32'd8,32'd82,32'd4294967223,32'd63,32'd5,32'd17,32'd7,32'd4294967190,32'd4294967255,32'd31,32'd4294967098,32'd4294967273,32'd106,32'd4294967289,32'd15,32'd4294967208,32'd61,32'd79,32'd4294967230,32'd29,32'd4294967206,32'd4294967126,32'd25,32'd134,32'd4294967256,32'd4294967273,32'd146,32'd109,32'd4294967232,32'd46,32'd46,32'd68,32'd82,32'd71,32'd134,32'd4294967220,32'd4294967263,32'd4294967294,32'd66,32'd31,32'd68,32'd39,32'd4294967134,32'd30,32'd4294967261,32'd32,32'd4294967214,32'd4294967274,32'd4294967222,32'd4294967277,32'd12,32'd126,32'd4294967025,32'd50,32'd68,32'd2,32'd16,32'd100,32'd9,32'd25,32'd10,32'd18,32'd4294967210,32'd4294967189,32'd4294967254,32'd38,32'd109,32'd156,32'd168,32'd4294967268,32'd10,32'd87,32'd9,32'd4294967204,32'd20,32'd4294967091,32'd4294967229,32'd4294967105,32'd69,32'd6,32'd4294967173,32'd59,32'd162,32'd48,32'd95,32'd180,32'd139,32'd27,32'd4294967251,32'd4294967290,32'd5,32'd91,32'd35,32'd4294967134,32'd4294967150,32'd4294967261,32'd4294966991,32'd4294967135,32'd13,32'd50,32'd7,32'd81,32'd4294967258,32'd32,32'd4294967247,32'd23,32'd4294967087,32'd4294967181,32'd4294967124,32'd30,32'd35,32'd4294967278,32'd122,32'd150,32'd75,32'd66,32'd177,32'd98,32'd4294967159,32'd13,32'd138,32'd30,32'd36,32'd4294966957,32'd51,32'd4294967240,32'd4294966917,32'd123,32'd120,32'd197,32'd4294967289,32'd4294967257,32'd164,32'd30,32'd4294967096,32'd20,32'd4294967237,32'd155,32'd186,32'd4294967124,32'd135,32'd54,32'd106,32'd4294967092,32'd128,32'd188,32'd4294967102,32'd99,32'd146,32'd4294967228,32'd4294967271,32'd174,32'd4294967258,32'd4294967211,32'd119,32'd69,32'd58,32'd4294967017,32'd221,32'd90,32'd151,32'd4294967095,32'd109,32'd57,32'd56,32'd4294967056,32'd161,32'd151,32'd136,32'd170,32'd4294967012}
`define FEATURE_BELOW {32'd62,32'd4294967279,32'd4294967272,32'd4294967194,32'd14,32'd4294967290,32'd4294967218,32'd4294967276,32'd4294967289,32'd83,32'd4294967239,32'd4294967290,32'd25,32'd96,32'd9,32'd90,32'd24,32'd4294967273,32'd4294967291,32'd10,32'd4294967261,32'd4294967198,32'd33,32'd4294967274,32'd21,32'd4294967268,32'd4294967266,32'd82,32'd149,32'd4294967292,32'd4294967170,32'd4294967273,32'd43,32'd4294967279,32'd4294967169,32'd4,32'd33,32'd4294967272,32'd27,32'd4294967250,32'd5,32'd4294967146,32'd101,32'd4294967288,32'd4294967229,32'd47,32'd108,32'd4294967255,32'd4,32'd151,32'd17,32'd3,32'd4294967242,32'd4294967216,32'd0,32'd4294967269,32'd4294967247,32'd4294967105,32'd2,32'd156,32'd28,32'd4294967258,32'd4294967288,32'd4294967267,32'd4294967292,32'd4294967295,32'd20,32'd4294967275,32'd54,32'd4294967291,32'd28,32'd4294967236,32'd151,32'd100,32'd4294967250,32'd4294967266,32'd4294967196,32'd210,32'd4294967256,32'd4294967289,32'd57,32'd4294967272,32'd19,32'd4294967188,32'd36,32'd4294967251,32'd11,32'd4294967202,32'd20,32'd4294967263,32'd4,32'd4294967290,32'd69,32'd5,32'd18,32'd92,32'd7,32'd10,32'd4294967289,32'd122,32'd4294967287,32'd50,32'd89,32'd4294967271,32'd95,32'd4294967269,32'd3,32'd4294967176,32'd25,32'd42,32'd4294967272,32'd105,32'd150,32'd36,32'd44,32'd4294967288,32'd4294967225,32'd4294967253,32'd103,32'd4294967211,32'd18,32'd116,32'd65,32'd4294967265,32'd21,32'd4294967268,32'd4294967203,32'd4294967266,32'd129,32'd2,32'd4294967209,32'd4294967177,32'd25,32'd84,32'd7,32'd83,32'd4294967292,32'd4294967253,32'd81,32'd4294967295,32'd4294967274,32'd4294967275,32'd67,32'd4294967185,32'd4294967286,32'd4294967289,32'd66,32'd4294967118,32'd57,32'd4294967115,32'd15,32'd4294967278,32'd4294967202,32'd50,32'd149,32'd68,32'd4294967135,32'd9,32'd4,32'd74,32'd4294967241,32'd23,32'd30,32'd4294967289,32'd4294967284,32'd4294967274,32'd4294967224,32'd4294967228,32'd4294967261,32'd4294967254,32'd102,32'd4294967195,32'd4294967232,32'd3,32'd4294967226,32'd4294967262,32'd4294967195,32'd4294967111,32'd4294967228,32'd42,32'd4294967244,32'd37,32'd2,32'd2,32'd4,32'd4294967239,32'd17,32'd62,32'd4294967288,32'd5,32'd4294967232,32'd4,32'd4294967232,32'd5,32'd4294967266,32'd48,32'd12,32'd4294967244,32'd4294967177,32'd80,32'd13,32'd5,32'd4294967100,32'd0,32'd4294967291,32'd6,32'd4294967232,32'd16,32'd4294967255,32'd4294967273,32'd4294967261,32'd2,32'd4294967288,32'd16,32'd44,32'd4294967291,32'd4294967085,32'd59,32'd4294967277,32'd4294967294,32'd57,32'd4294966600,32'd4294967271,32'd9,32'd4294967290,32'd2,32'd103,32'd4294967182,32'd4294967227,32'd4294967231,32'd4294967292,32'd30,32'd4294967237,32'd46,32'd4294967181,32'd15,32'd4294967271,32'd29,32'd4294967275,32'd15,32'd4294967286,32'd20,32'd42,32'd26,32'd4294967278,32'd14,32'd117,32'd15,32'd4294967240,32'd4294967293,32'd42,32'd4294967281,32'd4294967292,32'd53,32'd4294967270,32'd4294967286,32'd4294967227,32'd74,32'd4294967268,32'd114,32'd4294967288,32'd4294967053,32'd5,32'd11,32'd4294967294,32'd15,32'd4294967290,32'd4294967215,32'd100,32'd4294967231,32'd4294967241,32'd25,32'd38,32'd4294967069,32'd4294967263,32'd3,32'd4294967158,32'd17,32'd4294967290,32'd46,32'd4294967261,32'd4,32'd4294967205,32'd4294967269,32'd4294967277,32'd21,32'd4294967251,32'd32,32'd4294967272,32'd13,32'd107,32'd4294967187,32'd4294967242,32'd4294967295,32'd4294967271,32'd57,32'd37,32'd4294967276,32'd4294967273,32'd4294967287,32'd4294967279,32'd36,32'd4294967192,32'd23,32'd125,32'd4294967222,32'd4294967289,32'd17,32'd4294967233,32'd85,32'd4294967241,32'd4294967291,32'd45,32'd24,32'd4294967294,32'd18,32'd4294967264,32'd42,32'd44,32'd2,32'd4,32'd4294967240,32'd66,32'd27,32'd139,32'd4294967250,32'd4294967269,32'd4294967294,32'd4294967287,32'd4294967259,32'd4294967272,32'd83,32'd4294967270,32'd1,32'd36,32'd94,32'd4294967168,32'd4294967292,32'd4294967180,32'd25,32'd4294967163,32'd18,32'd4294967265,32'd4294967275,32'd4294967170,32'd23,32'd4294967290,32'd19,32'd24,32'd302,32'd4294967189,32'd17,32'd32,32'd30,32'd4294967274,32'd4294967275,32'd96,32'd4294967227,32'd4294967265,32'd4294967294,32'd2,32'd4294967275,32'd75,32'd4294967262,32'd52,32'd4294967123,32'd4294967123,32'd14,32'd107,32'd165,32'd4294967215,32'd4294967229,32'd11,32'd4294967232,32'd1,32'd32,32'd68,32'd5,32'd4294967264,32'd43,32'd4294967269,32'd4294967116,32'd37,32'd4294967291,32'd5,32'd34,32'd4294967146,32'd21,32'd4294967186,32'd4294967288,32'd61,32'd4294967260,32'd4294967114,32'd19,32'd4294967143,32'd4294967168,32'd7,32'd36,32'd4294967268,32'd32,32'd86,32'd60,32'd4294967195,32'd4294967251,32'd97,32'd4294967265,32'd4294967234,32'd33,32'd4294967236,32'd4294967235,32'd4294967208,32'd4294967280,32'd162,32'd4,32'd19,32'd4294967269,32'd18,32'd4294967263,32'd139,32'd4294967213,32'd4294967288,32'd4294967276,32'd4294967292,32'd4294967265,32'd4294963456,32'd4294967062,32'd4294967217,32'd153,32'd46,32'd4294967294,32'd2,32'd4294967277,32'd20,32'd4294967219,32'd5,32'd34,32'd62,32'd4294967227,32'd4294967167,32'd4294967273,32'd4294967291,32'd40,32'd44,32'd4294967288,32'd19,32'd4294967273,32'd4294967245,32'd4294967277,32'd0,32'd4294967273,32'd4294967255,32'd149,32'd10,32'd1,32'd4294967252,32'd4294967291,32'd17,32'd58,32'd61,32'd4294967231,32'd18,32'd4294967256,32'd40,32'd4294967270,32'd4294967240,32'd24,32'd56,32'd4294967290,32'd4294967265,32'd63,32'd20,32'd4294967244,32'd152,32'd4294967079,32'd3,32'd4294967275,32'd25,32'd4294967214,32'd4294966817,32'd4294967198,32'd59,32'd4294967291,32'd30,32'd4,32'd4294967285,32'd66,32'd4294966834,32'd4294967225,32'd4294967252,32'd4294967276,32'd91,32'd20,32'd7,32'd4294967274,32'd17,32'd4294967270,32'd4294967183,32'd4294967266,32'd7,32'd4294967290,32'd4294967230,32'd54,32'd4294967271,32'd119,32'd142,32'd4294967205,32'd19,32'd4294967276,32'd17,32'd4294967197,32'd4294967271,32'd4294967164,32'd18,32'd9,32'd45,32'd4294967292,32'd119,32'd32,32'd4294967274,32'd4294967226,32'd4294967276,32'd65,32'd18,32'd4294967166,32'd102,32'd216,32'd89,32'd4294967236,32'd17,32'd4294967074,32'd14,32'd16,32'd4294967289,32'd74,32'd4294967234,32'd4294967211,32'd4294967222,32'd4294967159,32'd26,32'd4294967294,32'd4294967263,32'd75,32'd24,32'd102,32'd8,32'd4294967211,32'd4294967256,32'd116,32'd78,32'd31,32'd4294967288,32'd12,32'd25,32'd4294967181,32'd18,32'd66,32'd4294967177,32'd20,32'd108,32'd4294967261,32'd6,32'd2,32'd50,32'd4294967275,32'd4294967205,32'd4294967276,32'd9,32'd54,32'd4294967292,32'd4294967189,32'd22,32'd86,32'd26,32'd4294967292,32'd4294967262,32'd4294967248,32'd74,32'd4294967187,32'd58,32'd132,32'd29,32'd4294967204,32'd4294967207,32'd4294967256,32'd4294967085,32'd4294967150,32'd4294967218,32'd4294967145,32'd76,32'd4294967233,32'd4294967220,32'd4294967157,32'd17,32'd4294967271,32'd4294967106,32'd19,32'd29,32'd4294967275,32'd43,32'd4294967237,32'd4294967266,32'd5,32'd4294967272,32'd61,32'd91,32'd4294967267,32'd4294967273,32'd4294967247,32'd4294967248,32'd4294967181,32'd28,32'd117,32'd4294967274,32'd595,32'd4294967273,32'd21,32'd4294967288,32'd4294967090,32'd4294967289,32'd20,32'd4294967271,32'd93,32'd4294967260,32'd15,32'd4294967272,32'd77,32'd14,32'd4294967284,32'd131,32'd17,32'd4294967050,32'd4294967096,32'd51,32'd60,32'd4294967293,32'd17,32'd4294967056,32'd31,32'd4294967183,32'd97,32'd4294967276,32'd41,32'd4294967276,32'd4294967220,32'd4294967272,32'd4294967247,32'd4294967256,32'd63,32'd4294967150,32'd17,32'd4294967176,32'd22,32'd4294967293,32'd48,32'd4294966790,32'd165,32'd4294967268,32'd29,32'd4294967279,32'd122,32'd5,32'd4294967284,32'd7,32'd178,32'd223,32'd123,32'd4294967252,32'd18,32'd4294967268,32'd4294967228,32'd4294967292,32'd4294967224,32'd4294967291,32'd4294966840,32'd4294967224,32'd21,32'd4294967269,32'd60,32'd30,32'd6,32'd4294967170,32'd4294967257,32'd4294967259,32'd18,32'd19,32'd7,32'd4294967237,32'd22,32'd6,32'd23,32'd4294967232,32'd4294967293,32'd51,32'd27,32'd4294967238,32'd4294967202,32'd4294967293,32'd4294967278,32'd4294967193,32'd4294967060,32'd20,32'd21,32'd103,32'd16,32'd4294967273,32'd4294967123,32'd4294967291,32'd15,32'd107,32'd29,32'd4294967170,32'd4294967239,32'd10,32'd82,32'd37,32'd44,32'd4294967260,32'd282,32'd51,32'd5,32'd4294967239,32'd4294967260,32'd4294967277,32'd23,32'd4294967269,32'd66,32'd4294967269,32'd4294967235,32'd4294967164,32'd83,32'd162,32'd0,32'd4294967271,32'd19,32'd23,32'd3,32'd55,32'd31,32'd4294967277,32'd72,32'd44,32'd4294967223,32'd37,32'd56,32'd4294967031,32'd4294967285,32'd125,32'd4294967278,32'd4294967293,32'd74,32'd4294967273,32'd4294967240,32'd4294967175,32'd2,32'd4294967290,32'd128,32'd93,32'd0,32'd0,32'd120,32'd26,32'd21,32'd4294967273,32'd4294967282,32'd4294967289,32'd15,32'd25,32'd92,32'd4294967295,32'd4294967226,32'd4294967178,32'd109,32'd0,32'd49,32'd4294967260,32'd122,32'd9,32'd4294967280,32'd87,32'd4294967200,32'd9,32'd4294967205,32'd4294967173,32'd22,32'd3,32'd47,32'd59,32'd4294967237,32'd4294967214,32'd4294967255,32'd4294967193,32'd4294967268,32'd82,32'd4294967290,32'd18,32'd4294967125,32'd53,32'd4294967205,32'd147,32'd20,32'd4294967262,32'd40,32'd21,32'd4294967244,32'd17,32'd4294967262,32'd11,32'd4294967199,32'd25,32'd37,32'd32,32'd4294967267,32'd4294967257,32'd4294967280,32'd4294967237,32'd79,32'd28,32'd4294967273,32'd9,32'd4294967147,32'd165,32'd4294967287,32'd4294967268,32'd4294967274,32'd3,32'd4294967242,32'd4294967034,32'd4294967294,32'd4294967218,32'd4294967195,32'd14,32'd134,32'd4294967278,32'd4294967273,32'd22,32'd108,32'd17,32'd4294967271,32'd5,32'd57,32'd27,32'd86,32'd15,32'd10,32'd4294967164,32'd18,32'd113,32'd4294967109,32'd4294966902,32'd35,32'd9,32'd4294967276,32'd34,32'd4294967238,32'd4294967273,32'd4294967293,32'd4294967287,32'd4294967275,32'd19,32'd4294967276,32'd24,32'd4294967292,32'd4294967266,32'd4294967248,32'd19,32'd91,32'd8,32'd4294967294,32'd18,32'd120,32'd8,32'd4294966961,32'd32,32'd4294967224,32'd4294967288,32'd4294967278,32'd4294966900,32'd4294967247,32'd220,32'd4294967246,32'd20,32'd4294967267,32'd4294967045,32'd84,32'd37,32'd4294967157,32'd52,32'd4294967220,32'd17,32'd4,32'd4294967287,32'd4294967210,32'd4294967190,32'd34,32'd4294967290,32'd58,32'd43,32'd4294967210,32'd9,32'd84,32'd0,32'd4294967128,32'd15,32'd4294967092,32'd29,32'd98,32'd4294967288,32'd4294967126,32'd21,32'd109,32'd96,32'd4294967223,32'd26,32'd25,32'd4294967292,32'd4294967216,32'd4294967254,32'd4294967288,32'd24,32'd26,32'd2,32'd0,32'd4294967274,32'd4294967235,32'd101,32'd4294967293,32'd4294967263,32'd50,32'd4294967282,32'd4294967228,32'd23,32'd4294967294,32'd17,32'd18,32'd140,32'd4294967147,32'd112,32'd4294967246,32'd68,32'd51,32'd4294967241,32'd11,32'd4294967214,32'd4294967271,32'd10,32'd4294967101,32'd4294967289,32'd69,32'd4294967182,32'd49,32'd4294967281,32'd4294967254,32'd23,32'd4294967267,32'd84,32'd4294967185,32'd4294967153,32'd4294967257,32'd65,32'd4294967160,32'd4294967236,32'd4294967212,32'd4294967284,32'd0,32'd4294967224,32'd3,32'd81,32'd4294967169,32'd33,32'd4294967184,32'd4294967127,32'd4294967259,32'd45,32'd54,32'd83,32'd4294967155,32'd21,32'd53,32'd4294967233,32'd4294967261,32'd4294967238,32'd3,32'd4294967158,32'd23,32'd4294967201,32'd4294967221,32'd92,32'd4294967227,32'd34,32'd32,32'd40,32'd4294967186,32'd29,32'd33,32'd4294967136,32'd4294967269,32'd6,32'd169,32'd181,32'd4294967290,32'd24,32'd4294967271,32'd5,32'd4294967224,32'd111,32'd4294967198,32'd51,32'd64,32'd4294967042,32'd5,32'd73,32'd4294967203,32'd19,32'd4294967191,32'd103,32'd4294967290,32'd22,32'd4294967266,32'd24,32'd98,32'd41,32'd4294967286,32'd2,32'd221,32'd37,32'd4294967195,32'd26,32'd4294967289,32'd21,32'd4294967211,32'd17,32'd4294967141,32'd4294967258,32'd42,32'd4294967288,32'd24,32'd4294967171,32'd10,32'd4294967257,32'd4294967252,32'd4294967288,32'd4294967217,32'd4294967292,32'd47,32'd70,32'd4294967277,32'd4294967187,32'd4294967196,32'd4294967111,32'd160,32'd4294967203,32'd4294967267,32'd118,32'd4294967205,32'd20,32'd249,32'd4294967279,32'd4294967262,32'd4294967290,32'd4294967141,32'd37,32'd4294967236,32'd4294967285,32'd57,32'd83,32'd4294967209,32'd4294967277,32'd58,32'd4294967267,32'd4294967151,32'd22,32'd4294967290,32'd17,32'd4294967273,32'd1,32'd4294967264,32'd4294967287,32'd4294967269,32'd4294967234,32'd113,32'd4294967229,32'd4294967277,32'd23,32'd3,32'd4294967281,32'd4294967268,32'd18,32'd4294967266,32'd4294967294,32'd4294967110,32'd40,32'd4294967261,32'd308,32'd4294967007,32'd22,32'd1,32'd24,32'd4294967274,32'd4294967205,32'd4294967052,32'd32,32'd4294967269,32'd2,32'd23,32'd4294967270,32'd4294967232,32'd4294967269,32'd4294967244,32'd4294967287,32'd4294967231,32'd4294967271,32'd22,32'd83,32'd4294967229,32'd15,32'd4294967249,32'd4294967288,32'd4294967292,32'd4294967280,32'd4294967275,32'd4294967290,32'd25,32'd18,32'd4294967193,32'd35,32'd142,32'd14,32'd4294967197,32'd21,32'd4294967098,32'd6,32'd4294967276,32'd4294967157,32'd4294967268,32'd4294967277,32'd5,32'd4294967249,32'd3,32'd4294967221,32'd4294967229,32'd4294967295,32'd44,32'd4294967295,32'd3,32'd84,32'd4294967289,32'd4294967293,32'd125,32'd4,32'd4294967174,32'd39,32'd4294967295,32'd4294967273,32'd4294967268,32'd4294967068,32'd4294967291,32'd30,32'd4294967272,32'd4294967233,32'd4294967189,32'd34,32'd4294967291,32'd4294967113,32'd4294967249,32'd4294967295,32'd0,32'd26,32'd4294967244,32'd4294967283,32'd4294967195,32'd4294967284,32'd31,32'd4294967198,32'd4294967295,32'd4294967256,32'd2,32'd4294967226,32'd121,32'd4294967278,32'd14,32'd4294967255,32'd4294967254,32'd4294967232,32'd4294967227,32'd68,32'd4,32'd4294967163,32'd57,32'd4294967154,32'd43,32'd4294967219,32'd4294966921,32'd65,32'd4294966976,32'd43,32'd18,32'd4294967185,32'd25,32'd4294967295,32'd83,32'd4294967076,32'd14,32'd4294967269,32'd4294967270,32'd4294967161,32'd4294967281,32'd0,32'd20,32'd306,32'd69,32'd31,32'd22,32'd82,32'd111,32'd4294967255,32'd26,32'd4294967288,32'd23,32'd57,32'd3,32'd4294967225,32'd4,32'd4294967118,32'd4294967192,32'd206,32'd18,32'd4294967272,32'd4294967058,32'd4294967278,32'd10,32'd10,32'd4294967295,32'd4294967292,32'd31,32'd4294967268,32'd38,32'd135,32'd2,32'd4294967214,32'd45,32'd4294967272,32'd96,32'd19,32'd53,32'd4294967237,32'd4294967261,32'd4294967273,32'd30,32'd4294967238,32'd4294967270,32'd4294967292,32'd4294967079,32'd4294967270,32'd52,32'd4294967272,32'd4294967294,32'd3,32'd27,32'd4294967273,32'd4294967294,32'd2,32'd4294967227,32'd4294967262,32'd118,32'd4294967270,32'd4294967286,32'd15,32'd4294967235,32'd4294967210,32'd4294967147,32'd4294967182,32'd240,32'd63,32'd4294967245,32'd4294967147,32'd18,32'd4294967263,32'd4294967253,32'd169,32'd81,32'd4294967144,32'd92,32'd4294967157,32'd22,32'd4294967262,32'd50,32'd4294967266,32'd4294967265,32'd4294967292,32'd4294967273,32'd4294967288,32'd4294967188,32'd4294967217,32'd80,32'd67,32'd7,32'd4294967187,32'd43,32'd4294967275,32'd6,32'd4294967139,32'd41,32'd60,32'd4294967293,32'd50,32'd90,32'd4294967217,32'd0,32'd4294967295,32'd212,32'd4294967295,32'd23,32'd4294967239,32'd4294967259,32'd44,32'd4294967164,32'd4294967215,32'd23,32'd59,32'd4294967207,32'd4294967264,32'd4294967260,32'd4294967206,32'd4294967173,32'd4294967293,32'd4294967290,32'd6,32'd4294967198,32'd58,32'd4294967198,32'd4294967214,32'd4294967260,32'd80,32'd21,32'd4294967182,32'd4294967143,32'd4294967253,32'd69,32'd4294967191,32'd4294967294,32'd129,32'd4294967205,32'd6,32'd172,32'd4294967233,32'd4294967269,32'd4294967208,32'd4294967255,32'd4294967252,32'd4294967261,32'd4294967186,32'd4294967249,32'd91,32'd4294967270,32'd87,32'd9,32'd4294967294,32'd4294967227,32'd4294967271,32'd58,32'd3,32'd4,32'd4294967279,32'd4294967262,32'd44,32'd4294967289,32'd4294967294,32'd4294967288,32'd100,32'd4294967158,32'd4294967220,32'd4294967273,32'd19,32'd4294967295,32'd7,32'd4294967288,32'd4294967220,32'd4294967287,32'd132,32'd4,32'd5,32'd4294967290,32'd5,32'd4294967288,32'd16,32'd4294967174,32'd40,32'd28,32'd21,32'd4294967264,32'd4294966968,32'd4294967226,32'd4294967262,32'd248,32'd24,32'd4294967225,32'd4294967284,32'd25,32'd4294967269,32'd4294967180,32'd4294967294,32'd4294967295,32'd31,32'd182,32'd45,32'd4294967295,32'd4294967222,32'd61,32'd4294966944,32'd48,32'd4294967294,32'd0,32'd176,32'd4294967254,32'd2,32'd74,32'd26,32'd4294967295,32'd15,32'd4294967251,32'd4294967203,32'd4294967262,32'd12,32'd29,32'd54,32'd4294967219,32'd1,32'd4294967263,32'd72,32'd4294967186,32'd22,32'd4294967263,32'd26,32'd125,32'd31,32'd4294967292,32'd66,32'd4294967236,32'd16,32'd108,32'd25,32'd4294967115,32'd4294967198,32'd4294967270,32'd57,32'd4294967295,32'd4294967268,32'd0,32'd4294967269,32'd4,32'd3,32'd4294967144,32'd4294967232,32'd81,32'd4294967227,32'd164,32'd21,32'd25,32'd4294967267,32'd4294967199,32'd35,32'd4294967267,32'd21,32'd4294967294,32'd4294967146,32'd76,32'd76,32'd4294967292,32'd0,32'd46,32'd4294967288,32'd4294967187,32'd3,32'd38,32'd97,32'd4294967151,32'd17,32'd4294967292,32'd78,32'd4294967188,32'd4294967176,32'd8,32'd4294967285,32'd79,32'd4294967166,32'd115,32'd4294967163,32'd122,32'd4294967157,32'd5,32'd4294967234,32'd4294967169,32'd4294967281,32'd4294967253,32'd17,32'd185,32'd4294967275,32'd18,32'd4294967192,32'd4294967193,32'd4294967224,32'd4294967218,32'd4294967222,32'd30,32'd35,32'd42,32'd4294967175,32'd4294967236,32'd4294967270,32'd18,32'd4294967278,32'd18,32'd5,32'd4294967210,32'd4294967195,32'd4294967187,32'd51,32'd78,32'd63,32'd30,32'd232,32'd15,32'd4294967238,32'd4294967288,32'd124,32'd4294967271,32'd4294967288,32'd30,32'd4294967184,32'd44,32'd4294967207,32'd23,32'd4294967266,32'd81,32'd4294967268,32'd77,32'd4294967269,32'd4294967047,32'd6,32'd4294967175,32'd107,32'd104,32'd4294967248,32'd25,32'd4294967277,32'd17,32'd4294967292,32'd17,32'd4294967139,32'd9,32'd4294967204,32'd4294967001,32'd155,32'd4294967238,32'd4294967288,32'd4294967227,32'd19,32'd15,32'd37,32'd14,32'd4294967292,32'd4294967293,32'd54,32'd1,32'd4294967292,32'd4294967293,32'd4294967272,32'd4294967262,32'd59,32'd4294967211,32'd4294966997,32'd43,32'd58,32'd6,32'd23,32'd4294967216,32'd2,32'd4294967289,32'd0,32'd4294967196,32'd4294967229,32'd84,32'd4294967294,32'd4294967139,32'd4294967254,32'd4294967293,32'd4294967260,32'd60,32'd14,32'd4294967293,32'd4294967291,32'd4294967251,32'd4294967292,32'd33,32'd4294967209,32'd19,32'd49,32'd20,32'd86,32'd4294967283,32'd48,32'd4294967295,32'd4294967149,32'd4294967291,32'd78,32'd4294967191,32'd4294967266,32'd4294967288,32'd150,32'd64,32'd4294967273,32'd26,32'd4294967269,32'd4294967193,32'd4294967293,32'd19,32'd4294967290,32'd4294967282,32'd4294967261,32'd4294967267,32'd4294967245,32'd12,32'd4294967292,32'd22,32'd5,32'd4294967286,32'd4294967176,32'd31,32'd80,32'd23,32'd4294967227,32'd4294967261,32'd4294967147,32'd4294967290,32'd4294967256,32'd30,32'd4294967295,32'd15,32'd354,32'd22,32'd4294967203,32'd4294967205,32'd4294967192,32'd19,32'd103,32'd113,32'd4294966986,32'd37,32'd30,32'd4294967129,32'd4294967258,32'd4294967244,32'd4294967271,32'd4294967155,32'd4294967187,32'd4294967209,32'd152,32'd50,32'd2,32'd4294967230,32'd58,32'd4294967259,32'd4294967213,32'd4294967259,32'd28,32'd4294967247,32'd73,32'd73,32'd20,32'd4294967264,32'd21,32'd4294967216,32'd20,32'd4294967270,32'd41,32'd4294967269,32'd17,32'd58,32'd24,32'd4294967272,32'd19,32'd39,32'd86,32'd4294967210,32'd34,32'd4294967289,32'd4294967266,32'd4294967194,32'd4294967272,32'd4294967188,32'd23,32'd4294967290,32'd4294967217,32'd4294967273,32'd11,32'd4294967246,32'd3,32'd4294967264,32'd17,32'd17,32'd4294967238,32'd4294967186,32'd4294967293,32'd66,32'd19,32'd4294967294,32'd75,32'd4294967291,32'd70,32'd4294967075,32'd49,32'd4294967186,32'd4294967030,32'd109,32'd4294967295,32'd4294967292,32'd4294967213,32'd89,32'd4294967292,32'd4294967259,32'd4294967278,32'd4294967183,32'd45,32'd107,32'd4294967144,32'd4294967274,32'd67,32'd4294967250,32'd79,32'd2,32'd16,32'd4294967133,32'd4294967287,32'd4294967270,32'd22,32'd4294967288,32'd61,32'd4294967131,32'd4294967287,32'd4294967192,32'd15,32'd4294967183,32'd4294967196,32'd131,32'd4294967282,32'd4294967274,32'd4294967131,32'd4294967228,32'd4294967218,32'd4294967258,32'd79,32'd4294967192,32'd30,32'd4294967142,32'd4294967286,32'd30,32'd4294967219,32'd4294967233,32'd4294967233,32'd74,32'd4294967291,32'd4294967205,32'd4294967119,32'd4294967129,32'd22,32'd4294967097,32'd4294967094,32'd200,32'd1,32'd4294967224,32'd4294967120,32'd4294967257,32'd4294967217,32'd6,32'd4294967220,32'd4294967208,32'd32,32'd4294967204,32'd135,32'd4294967256,32'd4294967241,32'd65,32'd22,32'd4294967093,32'd77,32'd110,32'd114,32'd4294967247,32'd4294967284,32'd56,32'd56,32'd5,32'd20,32'd4294967149,32'd20,32'd4294967184,32'd4294967265,32'd4294967244,32'd49,32'd4294967115,32'd4294967195,32'd4294967224,32'd119,32'd4294967192,32'd20,32'd92,32'd311,32'd4294967144,32'd1,32'd18,32'd4294967202,32'd4294967177,32'd30,32'd4294967275,32'd27,32'd4294967171,32'd4294967081,32'd4294967246,32'd147,32'd4294967254,32'd4294967290,32'd279,32'd14,32'd4294967292,32'd4294967241,32'd105,32'd25,32'd4294967276,32'd4294967203,32'd4294967254,32'd4294967244,32'd4294967290,32'd15,32'd4294967274,32'd27,32'd4294967290,32'd49,32'd60,32'd4294967265,32'd4294967257,32'd0,32'd4294967289,32'd4294967254,32'd32,32'd29,32'd4294967264,32'd156,32'd4294967294,32'd15,32'd4294967268,32'd4294967231,32'd4294967265,32'd20,32'd4294967226,32'd69,32'd4294967178,32'd4294967289,32'd4294967213,32'd4294967274,32'd4294967112,32'd33,32'd39,32'd1,32'd84,32'd4294967192,32'd4294967130,32'd4294966935,32'd4294967185,32'd21,32'd29,32'd1,32'd122,32'd4294966591,32'd4294967163,32'd49,32'd4294967171,32'd4294967282,32'd4294967264,32'd19,32'd4294967253,32'd4294967213,32'd3,32'd4294967222,32'd4294967295,32'd4294967247,32'd4294967229,32'd4294967277,32'd4294967272,32'd23,32'd4294967262,32'd4294967286,32'd4294967294,32'd4294967237,32'd4294967295,32'd40,32'd4294967271,32'd14,32'd4294967295,32'd4294967259,32'd4294967264,32'd21,32'd81,32'd4294967164,32'd4294967261,32'd4294967176,32'd6,32'd4294967264,32'd4294967113,32'd53,32'd0,32'd36,32'd4294967245,32'd4294967277,32'd22,32'd20,32'd75,32'd4294967291,32'd4294967264,32'd146,32'd9,32'd69,32'd4294967110,32'd4294967152,32'd4294967264,32'd4294967286,32'd4294967185,32'd4294967289,32'd75,32'd4294967132,32'd4294967177,32'd4294967187,32'd58,32'd52,32'd4294967266,32'd65,32'd4294967235,32'd4294967242,32'd4294967232,32'd4294967180,32'd84,32'd4294967277,32'd11,32'd4294967165,32'd6,32'd4294967124,32'd8,32'd13,32'd4294967156,32'd4294967278,32'd4294967174,32'd4294967270,32'd27,32'd4294967289,32'd4294967066,32'd4294967256,32'd39,32'd4294967293,32'd22,32'd4294967036,32'd58,32'd4294967289,32'd4294967282,32'd4294967260,32'd38,32'd4294967210,32'd22,32'd7,32'd4294967223,32'd78,32'd4294967289,32'd4294967211,32'd4294967291,32'd4294967294,32'd4294967281,32'd264,32'd4294967271,32'd4294967292,32'd109,32'd4294967215,32'd4294967198,32'd4294967057,32'd283,32'd4294967145,32'd4294967112,32'd4294967251,32'd42,32'd4294967291,32'd4294967259,32'd4294967295,32'd33,32'd4294967268,32'd24,32'd137,32'd4294967283,32'd4294967294,32'd4294967207,32'd98,32'd4294967253,32'd176,32'd19,32'd4294967275,32'd4294967242,32'd4294967248,32'd0,32'd4294967179,32'd4294967243,32'd86,32'd162,32'd4294967274,32'd72,32'd5,32'd4294967293,32'd147,32'd4294967285,32'd4294967246,32'd4294966781,32'd4294967234,32'd78,32'd4294967274,32'd4294967252,32'd15,32'd17,32'd49,32'd77,32'd4294967262,32'd4294967290,32'd36,32'd4294967156,32'd4294967143,32'd22,32'd4294967293,32'd26,32'd4294967099,32'd45,32'd4294967148,32'd27,32'd53,32'd130,32'd4294967154,32'd61,32'd4294967270,32'd4294967295,32'd88,32'd26,32'd4294967267,32'd4,32'd4294967265,32'd4294967129,32'd20,32'd58,32'd1,32'd43,32'd5,32'd4294967274,32'd4294967107,32'd28,32'd20,32'd24,32'd4294967245,32'd29,32'd4294967180,32'd27,32'd4294967257,32'd158,32'd104,32'd4294967174,32'd86,32'd27,32'd4294967236,32'd4294967204,32'd4294967159,32'd4294967225,32'd46,32'd4294967224,32'd4294967181,32'd87,32'd70,32'd23,32'd51,32'd4294967292,32'd4294967222,32'd4294967169,32'd192,32'd4294967252,32'd4294967295,32'd4294967236,32'd0,32'd4294967295,32'd14,32'd17,32'd4294967276,32'd46,32'd8,32'd4294967120,32'd42,32'd4294967194,32'd118,32'd38,32'd4294967207,32'd70,32'd4294967273,32'd4294967263,32'd4294967290,32'd28,32'd4294967097,32'd50,32'd19,32'd1,32'd8,32'd4294967292,32'd23,32'd4294967207,32'd4294967264,32'd245,32'd4294967265,32'd4294967295,32'd10,32'd4294967090,32'd4294967257,32'd2,32'd2,32'd4294967262,32'd103,32'd4294967154,32'd15,32'd42,32'd24,32'd4294967261,32'd37,32'd18,32'd4294967102,32'd4294967162,32'd17,32'd4294967265,32'd19,32'd4294967160,32'd43,32'd4294967294,32'd87,32'd4294967239,32'd4294967272,32'd4294967291,32'd177,32'd4294967135,32'd42,32'd104,32'd4294967244,32'd95,32'd19,32'd4294967256,32'd4294967077,32'd4294967121,32'd21,32'd31,32'd4294967230,32'd117,32'd74,32'd4294967203,32'd4294967244,32'd4294967132,32'd4294967050,32'd4294967293,32'd4294967246,32'd9,32'd25,32'd4294967255,32'd73,32'd228,32'd1,32'd4294967180,32'd17,32'd105,32'd4294967295,32'd35,32'd4294967286,32'd75,32'd63,32'd4294967250,32'd4294967159,32'd4294967146,32'd15,32'd4294967140,32'd4294967191,32'd156,32'd175,32'd4294967259,32'd20,32'd36,32'd4294967212,32'd0,32'd4294967283,32'd30,32'd4294967284,32'd4294967169,32'd4294967231,32'd4294967162,32'd4294967231,32'd42,32'd4294967144,32'd4294967249,32'd4294967192,32'd4294967187,32'd4294967217,32'd21,32'd3,32'd20,32'd49,32'd7,32'd4294967261,32'd6,32'd9,32'd24,32'd3,32'd16,32'd36,32'd4294967289,32'd4294967291,32'd4294967283,32'd4294967275,32'd20,32'd100,32'd232,32'd4294967271,32'd25,32'd4294967271,32'd62,32'd4294967050,32'd4294967286,32'd5,32'd4294967292,32'd4294967160,32'd4294967293,32'd155,32'd4294967294,32'd48,32'd4294967194,32'd4294967269,32'd39,32'd223,32'd88,32'd8,32'd4294967268,32'd4294967226,32'd18,32'd151,32'd4294967265,32'd4294967073,32'd12,32'd25,32'd29,32'd4294967253,32'd81,32'd4294967079,32'd10,32'd5,32'd1,32'd4294967265,32'd4294967074,32'd4294967294,32'd4294967278,32'd4294967294,32'd19,32'd6,32'd4294967168,32'd4294967258,32'd48,32'd4294967007,32'd4294967112,32'd4294967258,32'd48,32'd4294967140,32'd4294967233,32'd0,32'd4294967117,32'd4294967271,32'd45,32'd4294967180,32'd4294967290,32'd4294967270,32'd103,32'd101,32'd3,32'd4294967240,32'd4294967179,32'd4294967261,32'd4294967226,32'd4294967145,32'd34,32'd4294967257,32'd4294967267,32'd4294967185,32'd4294967205,32'd118,32'd4294967228,32'd4294967176,32'd4294967252,32'd4294967180,32'd4294967201,32'd30,32'd44,32'd11,32'd42,32'd74,32'd4294967217,32'd4294967260,32'd34,32'd118,32'd4294967200,32'd4294967186,32'd151,32'd4294967247,32'd4294967222,32'd15,32'd4294967177,32'd4294967221,32'd4294967243,32'd4294967166,32'd78,32'd4294967283,32'd125,32'd4294967213,32'd4294967244,32'd89,32'd4294967291,32'd83,32'd1,32'd4294967283,32'd122,32'd0,32'd29,32'd4294966903,32'd123,32'd47,32'd4294967175,32'd24,32'd8,32'd4294967267,32'd4294967264,32'd53,32'd4294967230,32'd4294967262,32'd4294967294,32'd4294967290,32'd4294967131,32'd23,32'd4294967176,32'd6,32'd4294967219,32'd117,32'd124,32'd76,32'd4294967257,32'd4294967221,32'd4294967248,32'd4294967279,32'd7,32'd87,32'd4294967293,32'd104,32'd4294967158,32'd4294967152,32'd85,32'd4294967217,32'd77,32'd382,32'd207,32'd66,32'd4294967163,32'd32,32'd4294967266,32'd24,32'd4294967209,32'd4294967272,32'd125,32'd26,32'd4294967128,32'd4294967193,32'd33,32'd59,32'd4294967171,32'd21,32'd98,32'd4,32'd4294967100,32'd0,32'd4294967292,32'd128,32'd4294967292,32'd4294967272,32'd136,32'd4294967289,32'd25,32'd33,32'd4294967151,32'd22,32'd4294967229,32'd4294967173,32'd61,32'd126,32'd4294967171,32'd4294967275,32'd3,32'd20,32'd21,32'd4294967186,32'd4294967131,32'd37,32'd4294967162,32'd4294967108,32'd117,32'd59,32'd4294967242,32'd4294967181,32'd4294967257,32'd4294967195,32'd4294967180,32'd4294967171,32'd56,32'd4294967275,32'd89,32'd4294967186,32'd4294967265,32'd4294967260,32'd19,32'd4294967139,32'd4294967226,32'd4294967293,32'd4294967222,32'd145,32'd2,32'd106,32'd4294967181,32'd100,32'd4294967286,32'd4294967249,32'd16,32'd96,32'd4294967285,32'd33,32'd4294967276,32'd4294967143,32'd4294967093,32'd4294967267,32'd177,32'd37,32'd4294967104,32'd22,32'd99,32'd4294967034,32'd4294967129,32'd48,32'd4294967214,32'd4294967260,32'd126,32'd4294967151,32'd60,32'd7,32'd4294967250,32'd4294967203,32'd25,32'd108,32'd4294967213,32'd4294967122,32'd4294967293,32'd4294967271,32'd105,32'd4294967228,32'd1,32'd123,32'd23,32'd4294967260,32'd107,32'd4294967149,32'd27,32'd4294966902,32'd4294967081,32'd25,32'd47,32'd5,32'd4294967177,32'd24,32'd81,32'd4294967145,32'd17,32'd15,32'd4294967192,32'd4294967108,32'd129,32'd2,32'd27,32'd4294967182,32'd4294967240,32'd3,32'd76,32'd4294967255,32'd4294967041,32'd20,32'd34,32'd108,32'd4294967283,32'd4294967226,32'd4294967206,32'd4294967247,32'd4294967244,32'd4294967153,32'd4294967205,32'd4294967224,32'd91,32'd4294967219,32'd4294967263,32'd29,32'd4294967235,32'd76,32'd4294967292,32'd4294967259,32'd4294967267,32'd4294967263,32'd4294967008,32'd4294967195,32'd4294967292,32'd54,32'd63,32'd4294967127,32'd4294967269,32'd18,32'd4294967168,32'd48,32'd4294967292,32'd4294967219,32'd4294967258,32'd4294967233,32'd6,32'd4294967289,32'd4294967264,32'd51,32'd4294967038,32'd4294967174,32'd58,32'd4294967295,32'd2,32'd32,32'd87,32'd73,32'd4294967023,32'd4294967105,32'd99,32'd218,32'd4294967195,32'd4294967286,32'd4294967263,32'd47,32'd4294967127,32'd4294967292,32'd6,32'd4294967019,32'd4294967235,32'd22,32'd4294967150,32'd25,32'd17,32'd4294967177,32'd8,32'd4294967283,32'd4294967261,32'd27,32'd12,32'd4294967179,32'd6,32'd26,32'd4294967228,32'd4294967229,32'd4,32'd20,32'd4294967220,32'd4294967190,32'd96,32'd0,32'd51,32'd4294967282,32'd4294967255,32'd42,32'd4294967140,32'd30,32'd4294967076,32'd39,32'd4294967223,32'd4294967150,32'd4294967165,32'd130,32'd4294967216,32'd4294967041,32'd4294967244,32'd20,32'd3,32'd54,32'd4294967107,32'd4294967214,32'd4294967018,32'd125,32'd61,32'd44,32'd4294967158,32'd4294967282,32'd4294967272,32'd4294967215,32'd25,32'd4294967211,32'd4294967092,32'd4294967178,32'd54,32'd4294967156,32'd4294967162,32'd4294967148,32'd106,32'd4294967274,32'd4294967152,32'd4294967146,32'd27,32'd251,32'd4294967177,32'd24,32'd4294967268,32'd4294967262,32'd4294967156,32'd4294967155,32'd91,32'd60,32'd123,32'd4294967071,32'd9,32'd4294967281,32'd4294967197,32'd20,32'd4294967166,32'd19,32'd4294967055,32'd4294967157,32'd4,32'd50,32'd4294967004,32'd4294967195,32'd43,32'd4294967238,32'd4294967181,32'd18,32'd5,32'd4294967231,32'd32,32'd4294967208,32'd21,32'd4294967162,32'd40,32'd4294967263,32'd107,32'd4294967156,32'd4294967239,32'd71,32'd4294967204,32'd4294967246,32'd4294967199,32'd4294967138,32'd4294967163,32'd25,32'd4294967173,32'd102,32'd4294967083,32'd18,32'd134,32'd113,32'd4294967269,32'd4294967164,32'd4294967165,32'd27,32'd4294967247,32'd26,32'd4294967161,32'd4294967193,32'd4294967248,32'd4294967166,32'd1,32'd120,32'd56,32'd27,32'd4294967245,32'd37,32'd4294967263,32'd75,32'd81,32'd4294967100,32'd4294967244,32'd4294967187,32'd103,32'd72,32'd4294967177,32'd4294967192,32'd4294967136,32'd24,32'd45,32'd4294967188,32'd4294967238,32'd4294967234,32'd4294967059,32'd71,32'd11,32'd4294967246,32'd4,32'd20,32'd4294967194,32'd38,32'd4294967182,32'd46,32'd4294967243,32'd4294967237,32'd167,32'd73,32'd4294967161,32'd223,32'd4294967131,32'd4294967225,32'd4294967223,32'd33,32'd4294967167,32'd4294967153,32'd4294967182,32'd4294967259,32'd4294967011,32'd4294967244,32'd26,32'd4294967252,32'd2,32'd4294967155,32'd18,32'd10,32'd4294967100,32'd4294967261,32'd37,32'd4294967000,32'd4294967260,32'd42,32'd27,32'd4294967121,32'd31,32'd4294967141,32'd4294967266,32'd37,32'd4294967265,32'd4294967107,32'd4294967164,32'd4294967092,32'd28,32'd132,32'd4294967165,32'd7,32'd45,32'd4294967254,32'd159,32'd4294967176,32'd32,32'd4294967243,32'd4294967284,32'd52,32'd4294967138,32'd33,32'd39,32'd4294967156,32'd4294967261,32'd201,32'd141,32'd4294967252,32'd4294967265,32'd82,32'd4294967170,32'd4294967134,32'd4294967200,32'd4294967186,32'd4294967135,32'd4294967182,32'd25,32'd110,32'd89,32'd4294967253,32'd4294967221,32'd4294967251,32'd4294967227,32'd8,32'd4294967118,32'd111,32'd4294967134,32'd29,32'd97,32'd34,32'd48,32'd4294967149,32'd4294967286,32'd2,32'd4294967222,32'd4294967248,32'd185,32'd4294967168,32'd4294967291,32'd4294967120,32'd4294967161,32'd4294967128,32'd4294967130,32'd26,32'd26,32'd106,32'd4294967162,32'd4294967251,32'd4294967288,32'd4294967262,32'd95,32'd4294967090,32'd4294967271,32'd4294967074,32'd58,32'd4294967128,32'd34,32'd62,32'd36,32'd4294967220,32'd160,32'd39,32'd4294967272,32'd4294967240,32'd4294967142,32'd4294967158,32'd4294967234,32'd4294967140,32'd4294966870,32'd142,32'd54,32'd4294966999,32'd4294967249,32'd4294967199,32'd32,32'd19,32'd50,32'd9,32'd23,32'd4294967111,32'd4294967188,32'd4294966998,32'd4294967233,32'd184,32'd4294966966,32'd127,32'd4294967045,32'd23,32'd62,32'd22,32'd4294966983,32'd4294967173,32'd191,32'd4294967240,32'd4294967256,32'd4294967189,32'd4294967109,32'd4294967222,32'd4294967096,32'd148,32'd4294967062,32'd4294967289,32'd4294967176,32'd4294967072,32'd8,32'd4294967248,32'd114,32'd22,32'd4294967244,32'd4294967283,32'd4294967256,32'd226,32'd194,32'd4294967275,32'd4294967166,32'd36,32'd4294967088,32'd135,32'd4294967244,32'd4294967257,32'd47,32'd4294967231,32'd4294967117,32'd4294967212,32'd59,32'd4294967085,32'd4294967166,32'd50,32'd4294967218,32'd4294967251,32'd143,32'd187,32'd4294967242,32'd148,32'd119,32'd4294967251,32'd4294967157,32'd4294966954,32'd34,32'd4294967225,32'd4294967047,32'd4294967089,32'd159,32'd4294967186,32'd4294967107,32'd4294967080,32'd71,32'd4294967196,32'd4294967184,32'd4294967103,32'd4294967057,32'd267}
