localparam int[13] pyramid_widths = {320, 266, 222, 185, 154, 128, 107, 89, 74, 62, 51, 43, 35};
localparam int[13] pyramid_heights = {240, 199, 166, 138, 115, 96, 80, 66, 55, 46, 38, 32, 26};

/*
320 x 240 - 63936 windows
266 x 199 - 42350 windows
222 x 166
185 x 138
154 x 115
128 x 96
107 x 80
89 x 66
74 x 55
62 x 46
51 x 38
43 x 32
35 x 26
*/