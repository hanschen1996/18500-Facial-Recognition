/** @file vj_weights.vh
 *  @brief Viola-Jones weights data structure
 */

// assume we use haarcascade_frontalface_default.xml
#define NUM_STAGE 25
#define NUM_FEATURE 2913
#define WINDOW_SIZE 24

localparam logic [24:0][31:0] stage_num_feature = {9, 25, 52, 84, 136, 189, 251, 323, 406, 497, 596, 711, 838, 973, 1109, 1246, 1405, 1560, 1729, 1925, 2122, 2303, 2502, 2713, 2913};

localparam logic [24:0][31:0] stage_threshold = {-258, -255, -238, -228, -225, -211, -206, -199, -197, -187, -198, -190, -183, -190, -175, -180, -184, -174, -166, -164, -168, -170, -167, -173, -153};

localparam logic [2912:0][31:0] rectangle1_xs = {6, 6, 3, 8, 3, 6, 5, 11, 4, 6, 6, 1, 0, 9, 5, 5, 13, 7, 10, 2, 18, 0, 9, 7, 5, 0, 5, 9, 9, 6, 3, 5, 18, 1, 0, 5, 2, 8, 2, 0, 20, 0, 18, 0, 12, 0, 12, 8, 5, 1, 17, 0, 6, 6, 0, 4, 2, 19, 1, 0, 1, 14, 3, 6, 8, 15, 1, 4, 0, 3, 1, 5, 3, 14, 1, 11, 5, 6, 9, 9, 7, 10, 8, 3, 6, 0, 4, 11, 0, 11, 4, 11, 9, 9, 1, 10, 6, 7, 0, 6, 1, 6, 2, 20, 0, 2, 0, 12, 5, 11, 0, 12, 6, 8, 0, 10, 3, 2, 2, 3, 5, 9, 4, 4, 6, 3, 0, 6, 6, 3, 1, 8, 0, 12, 0, 19, 0, 6, 7, 9, 0, 4, 7, 18, 0, 18, 0, 16, 2, 9, 2, 14, 5, 15, 0, 8, 7, 0, 1, 14, 7, 10, 4, 10, 1, 10, 5, 8, 6, 7, 0, 1, 5, 12, 6, 7, 0, 2, 2, 14, 8, 14, 8, 17, 6, 13, 3, 9, 0, 0, 6, 7, 10, 1, 5, 9, 20, 2, 5, 0, 5, 0, 6, 0, 1, 2, 2, 0, 9, 7, 11, 6, 18, 3, 18, 1, 11, 0, 13, 7, 11, 8, 13, 2, 3, 0, 9, 4, 7, 0, 7, 7, 3, 0, 3, 4, 13, 9, 5, 1, 10, 0, 1, 4, 0, 2, 9, 5, 17, 1, 14, 3, 15, 9, 17, 3, 7, 1, 10, 0, 15, 3, 12, 6, 14, 1, 13, 7, 12, 6, 6, 7, 7, 8, 7, 0, 15, 0, 15, 7, 15, 0, 8, 0, 3, 0, 9, 10, 7, 5, 14, 2, 0, 4, 9, 0, 18, 0, 8, 8, 11, 7, 12, 6, 15, 5, 9, 7, 14, 2, 5, 9, 12, 9, 3, 6, 12, 1, 12, 1, 10, 3, 10, 0, 6, 6, 5, 4, 11, 7, 3, 2, 3, 8, 16, 7, 18, 0, 18, 3, 18, 0, 5, 6, 10, 8, 15, 3, 15, 2, 8, 8, 15, 4, 13, 7, 18, 1, 14, 1, 4, 1, 10, 0, 15, 3, 15, 3, 15, 0, 4, 2, 14, 6, 17, 1, 16, 7, 12, 4, 10, 2, 15, 0, 6, 1, 6, 0, 8, 9, 6, 0, 16, 0, 14, 1, 5, 4, 16, 0, 10, 9, 9, 3, 6, 8, 0, 14, 5, 9, 0, 3, 3, 20, 0, 8, 6, 9, 1, 9, 7, 13, 7, 14, 2, 18, 6, 18, 7, 18, 0, 9, 0, 17, 1, 14, 6, 3, 9, 12, 6, 6, 1, 10, 5, 5, 0, 0, 1, 6, 4, 1, 5, 0, 3, 2, 6, 14, 0, 14, 0, 0, 0, 5, 3, 6, 0, 13, 7, 9, 1, 13, 5, 16, 4, 0, 5, 12, 2, 15, 0, 12, 11, 9, 8, 12, 3, 6, 7, 12, 10, 16, 4, 2, 5, 10, 8, 6, 6, 0, 1, 3, 3, 0, 10, 8, 5, 0, 14, 9, 14, 1, 15, 0, 17, 2, 3, 9, 18, 0, 4, 2, 14, 0, 18, 5, 21, 6, 8, 7, 21, 10, 15, 0, 11, 7, 12, 6, 14, 6, 3, 3, 0, 10, 11, 6, 16, 3, 16, 0, 10, 0, 13, 7, 5, 0, 6, 3, 8, 2, 15, 3, 17, 1, 19, 1, 4, 6, 15, 0, 15, 3, 8, 6, 5, 10, 10, 0, 15, 0, 12, 9, 12, 6, 15, 0, 11, 6, 10, 0, 3, 3, 0, 0, 12, 2, 7, 0, 3, 6, 5, 11, 0, 18, 3, 9, 0, 13, 0, 13, 4, 13, 5, 7, 6, 14, 4, 11, 0, 13, 2, 10, 8, 14, 6, 8, 7, 8, 5, 3, 0, 5, 0, 3, 1, 5, 1, 1, 3, 6, 6, 14, 1, 11, 10, 11, 7, 12, 2, 14, 6, 14, 0, 5, 1, 13, 7, 12, 0, 7, 7, 8, 1, 13, 5, 14, 4, 12, 9, 11, 5, 8, 1, 9, 3, 12, 8, 2, 0, 14, 2, 2, 6, 5, 1, 7, 3, 9, 2, 18, 3, 20, 2, 1, 0, 19, 0, 18, 0, 7, 0, 10, 8, 4, 2, 7, 3, 16, 5, 10, 4, 2, 6, 1, 12, 0, 15, 5, 8, 1, 17, 8, 17, 7, 15, 2, 10, 0, 20, 1, 15, 0, 16, 2, 10, 1, 11, 3, 3, 10, 3, 0, 12, 8, 10, 9, 4, 0, 9, 8, 13, 5, 0, 1, 19, 0, 16, 0, 12, 7, 9, 0, 1, 1, 13, 0, 12, 4, 15, 1, 3, 2, 13, 1, 3, 7, 12, 0, 13, 0, 15, 0, 13, 5, 0, 2, 0, 1, 15, 0, 6, 8, 10, 8, 12, 6, 13, 1, 15, 6, 13, 5, 6, 0, 11, 9, 10, 8, 3, 10, 4, 9, 5, 2, 13, 8, 12, 2, 7, 3, 11, 0, 3, 1, 11, 9, 9, 1, 6, 1, 8, 2, 11, 7, 11, 5, 11, 5, 4, 2, 7, 9, 2, 8, 3, 8, 0, 6, 0, 20, 0, 0, 0, 14, 0, 1, 5, 4, 8, 6, 2, 11, 2, 5, 9, 8, 6, 10, 0, 18, 2, 3, 2, 13, 6, 9, 7, 18, 9, 6, 0, 13, 0, 13, 5, 11, 4, 6, 0, 12, 0, 12, 5, 5, 5, 3, 7, 13, 2, 19, 1, 5, 0, 2, 5, 1, 3, 8, 6, 10, 1, 8, 3, 5, 4, 6, 7, 0, 0, 3, 2, 7, 5, 10, 9, 18, 4, 10, 9, 11, 7, 4, 2, 13, 7, 3, 1, 8, 3, 5, 8, 9, 0, 6, 0, 13, 5, 1, 9, 9, 5, 4, 0, 16, 9, 8, 8, 10, 7, 5, 2, 18, 1, 6, 9, 10, 6, 8, 1, 9, 6, 17, 2, 7, 1, 1, 9, 3, 16, 0, 16, 0, 8, 5, 4, 0, 6, 0, 20, 8, 6, 0, 6, 0, 20, 0, 15, 0, 13, 5, 5, 3, 6, 6, 10, 1, 11, 5, 12, 5, 13, 0, 8, 1, 2, 2, 17, 1, 7, 0, 15, 1, 9, 0, 16, 4, 7, 9, 12, 8, 15, 3, 15, 1, 15, 6, 10, 6, 11, 6, 11, 9, 3, 2, 3, 3, 4, 0, 10, 0, 5, 8, 11, 5, 5, 10, 10, 7, 1, 0, 12, 2, 12, 1, 12, 0, 5, 6, 14, 5, 9, 1, 8, 3, 12, 0, 8, 4, 12, 9, 9, 1, 8, 3, 7, 10, 10, 3, 12, 3, 10, 5, 7, 6, 12, 2, 0, 0, 0, 5, 1, 9, 2, 5, 4, 2, 7, 0, 2, 3, 6, 9, 15, 8, 3, 2, 19, 1, 14, 4, 14, 6, 14, 4, 0, 1, 20, 0, 8, 7, 16, 5, 11, 10, 10, 7, 14, 5, 12, 6, 11, 1, 15, 9, 10, 3, 16, 7, 15, 0, 13, 2, 5, 1, 5, 1, 14, 4, 14, 4, 18, 1, 2, 0, 12, 3, 16, 3, 9, 9, 15, 7, 17, 3, 3, 0, 2, 0, 13, 5, 5, 5, 18, 0, 3, 2, 2, 5, 6, 6, 13, 5, 6, 0, 18, 0, 12, 6, 0, 3, 9, 5, 4, 10, 8, 2, 8, 0, 18, 0, 9, 1, 2, 7, 8, 4, 10, 2, 15, 3, 15, 4, 15, 0, 15, 0, 10, 1, 7, 10, 8, 3, 7, 0, 10, 7, 5, 5, 6, 3, 16, 0, 0, 0, 10, 10, 4, 0, 9, 3, 6, 11, 5, 4, 2, 7, 1, 13, 5, 11, 6, 3, 0, 10, 6, 6, 0, 18, 0, 11, 0, 2, 1, 18, 0, 17, 0, 0, 0, 10, 7, 15, 3, 15, 0, 15, 0, 5, 0, 9, 3, 9, 5, 9, 8, 10, 5, 9, 7, 11, 9, 6, 1, 16, 0, 8, 0, 3, 0, 6, 0, 14, 1, 13, 4, 12, 2, 16, 3, 14, 8, 9, 0, 4, 5, 15, 0, 8, 1, 14, 4, 16, 3, 18, 1, 11, 0, 15, 7, 22, 0, 18, 0, 3, 6, 7, 2, 4, 9, 4, 3, 18, 2, 4, 7, 7, 6, 12, 0, 8, 2, 13, 5, 9, 5, 3, 2, 11, 3, 9, 1, 15, 1, 9, 6, 10, 7, 10, 4, 0, 3, 19, 0, 17, 1, 18, 0, 3, 2, 9, 5, 10, 8, 7, 9, 5, 8, 8, 6, 14, 6, 8, 2, 2, 0, 0, 7, 6, 14, 4, 2, 6, 9, 7, 6, 5, 18, 0, 18, 2, 5, 11, 15, 7, 7, 10, 10, 2, 14, 8, 14, 3, 14, 1, 3, 1, 18, 0, 5, 6, 14, 4, 15, 0, 0, 3, 3, 0, 1, 0, 2, 2, 0, 10, 10, 6, 11, 9, 2, 1, 13, 6, 10, 6, 14, 6, 9, 8, 17, 1, 14, 7, 3, 1, 14, 0, 12, 0, 10, 1, 15, 6, 6, 8, 14, 0, 10, 6, 7, 9, 10, 8, 7, 4, 17, 3, 10, 2, 3, 4, 15, 7, 15, 1, 11, 5, 10, 4, 0, 4, 10, 0, 6, 1, 18, 4, 6, 1, 1, 2, 12, 0, 10, 7, 9, 4, 6, 5, 10, 8, 9, 3, 4, 6, 8, 0, 11, 2, 8, 0, 0, 2, 4, 10, 7, 9, 17, 0, 16, 1, 12, 3, 12, 3, 12, 8, 10, 6, 13, 1, 7, 2, 0, 9, 0, 9, 2, 13, 4, 20, 8, 0, 0, 3, 3, 13, 5, 13, 2, 9, 8, 12, 8, 8, 11, 9, 0, 9, 1, 12, 6, 13, 1, 9, 2, 15, 0, 9, 2, 15, 4, 17, 0, 15, 0, 9, 3, 16, 0, 13, 0, 0, 5, 8, 4, 10, 8, 11, 4, 14, 2, 4, 8, 1, 7, 13, 8, 4, 3, 14, 8, 3, 4, 3, 9, 9, 7, 12, 6, 18, 3, 18, 0, 13, 5, 11, 3, 16, 5, 7, 1, 2, 3, 17, 5, 13, 0, 15, 1, 12, 1, 3, 6, 5, 9, 11, 4, 6, 5, 11, 5, 1, 7, 6, 6, 11, 5, 6, 0, 2, 0, 9, 9, 12, 0, 1, 3, 2, 5, 10, 8, 5, 6, 7, 5, 4, 0, 9, 9, 6, 9, 10, 5, 14, 5, 14, 0, 16, 4, 8, 0, 13, 0, 0, 6, 10, 1, 0, 2, 2, 1, 10, 7, 9, 7, 3, 7, 3, 8, 3, 6, 1, 5, 8, 3, 0, 2, 4, 9, 9, 14, 7, 14, 4, 17, 1, 14, 0, 9, 3, 14, 4, 7, 7, 14, 10, 14, 5, 4, 9, 3, 4, 16, 4, 6, 10, 9, 6, 5, 3, 6, 0, 6, 0, 4, 0, 15, 0, 6, 3, 12, 6, 6, 9, 10, 7, 14, 2, 11, 1, 15, 1, 10, 4, 7, 10, 13, 3, 13, 5, 10, 7, 15, 5, 8, 7, 12, 6, 7, 6, 5, 3, 3, 0, 14, 0, 1, 1, 7, 9, 10, 2, 8, 0, 5, 2, 14, 3, 9, 4, 0, 7, 11, 0, 14, 2, 11, 7, 6, 4, 14, 4, 13, 8, 17, 4, 15, 3, 12, 0, 16, 2, 15, 0, 18, 0, 16, 5, 12, 0, 5, 0, 8, 5, 10, 6, 6, 3, 12, 0, 0, 5, 10, 9, 8, 0, 16, 3, 6, 0, 14, 0, 2, 4, 12, 0, 6, 1, 11, 3, 15, 6, 9, 4, 7, 5, 11, 7, 8, 0, 10, 0, 20, 0, 12, 1, 5, 1, 6, 5, 11, 1, 11, 0, 3, 1, 0, 1, 11, 4, 12, 4, 13, 1, 9, 0, 6, 6, 10, 6, 13, 2, 11, 1, 1, 0, 13, 5, 18, 0, 11, 0, 12, 1, 7, 8, 6, 2, 14, 3, 15, 5, 11, 7, 11, 9, 4, 9, 17, 1, 7, 6, 9, 1, 19, 0, 3, 1, 2, 4, 6, 4, 15, 3, 8, 3, 15, 3, 5, 1, 14, 0, 15, 3, 9, 1, 13, 1, 6, 8, 0, 0, 4, 1, 14, 1, 10, 6, 10, 7, 14, 6, 8, 3, 5, 0, 9, 4, 10, 8, 7, 8, 11, 7, 4, 0, 7, 1, 11, 6, 7, 7, 9, 0, 7, 1, 9, 0, 1, 1, 9, 3, 9, 9, 16, 2, 13, 1, 14, 3, 13, 7, 4, 9, 7, 0, 15, 1, 14, 4, 15, 3, 0, 7, 1, 1, 6, 1, 15, 3, 4, 0, 6, 4, 6, 0, 3, 4, 20, 0, 11, 6, 11, 1, 11, 1, 11, 0, 3, 7, 17, 5, 16, 0, 6, 0, 3, 2, 10, 10, 11, 9, 5, 6, 10, 0, 6, 4, 14, 0, 1, 8, 13, 10, 7, 8, 7, 2, 11, 7, 13, 0, 12, 8, 12, 6, 14, 0, 14, 0, 4, 1, 4, 0, 3, 9, 0, 6, 2, 18, 0, 11, 9, 7, 1, 18, 5, 18, 0, 9, 2, 10, 5, 9, 7, 10, 4, 6, 0, 3, 9, 6, 2, 19, 0, 5, 5, 1, 8, 6, 9, 2, 5, 8, 9, 14, 2, 10, 1, 11, 4, 6, 5, 9, 7, 7, 2, 5, 7, 0, 0, 16, 5, 5, 0, 11, 0, 4, 2, 3, 2, 6, 0, 3, 0, 5, 1, 19, 3, 19, 7, 9, 0, 15, 1, 9, 7, 9, 7, 9, 7, 9, 10, 5, 0, 9, 2, 15, 1, 6, 0, 6, 0, 13, 2, 13, 5, 11, 7, 10, 3, 14, 4, 4, 5, 7, 2, 10, 3, 16, 0, 0, 4, 10, 7, 13, 3, 16, 2, 3, 4, 4, 3, 8, 2, 14, 7, 4, 0, 10, 5, 0, 0, 3, 9, 0, 6, 8, 2, 12, 5, 14, 5, 6, 7, 11, 7, 13, 0, 1, 6, 10, 3, 0, 0, 3, 7, 10, 8, 12, 6, 16, 2, 10, 8, 14, 0, 11, 3, 10, 0, 19, 4, 4, 0, 6, 19, 0, 18, 0, 5, 10, 9, 0, 7, 1, 8, 0, 13, 10, 13, 7, 4, 0, 0, 6, 7, 0, 13, 3, 12, 2, 9, 6, 14, 5, 10, 6, 14, 4, 14, 0, 13, 2, 6, 0, 19, 1, 15, 3, 11, 7, 14, 3, 20, 7, 7, 2, 15, 7, 13, 5, 3, 5, 9, 3, 19, 0, 20, 0, 7, 4, 10, 0, 7, 0, 13, 1, 7, 0, 6, 8, 7, 1, 16, 5, 7, 4, 6, 9, 15, 6, 12, 7, 6, 10, 10, 3, 4, 2, 13, 7, 1, 0, 0, 3, 3, 3, 13, 2, 10, 6, 2, 2, 10, 8, 13, 3, 3, 2, 14, 3, 5, 2, 17, 2, 0, 7, 15, 5, 11, 6, 11, 5, 15, 4, 12, 6, 5, 9, 12, 4, 4, 5, 14, 9, 9, 9, 1, 2, 12, 6, 12, 8, 7, 0, 4, 2, 15, 0, 6, 6, 8, 1, 6, 7, 10, 3, 15, 1, 15, 10, 15, 6, 15, 6, 16, 2, 2, 6, 9, 2, 16, 0, 15, 8, 15, 0, 12, 3, 13, 0, 10, 7, 4, 0, 6, 3, 9, 5, 5, 3, 5, 6, 0, 2, 8, 18, 0, 4, 6, 4, 4, 7, 0, 13, 5, 3, 0, 14, 0, 14, 0, 6, 0, 14, 6, 15, 8, 4, 5, 7, 10, 5, 1, 18, 0, 13, 0, 12, 7, 14, 0, 14, 2, 14, 1, 3, 5, 5, 8, 9, 6, 5, 8, 6, 3, 13, 3, 12, 7, 13, 7, 11, 7, 5, 8, 4, 0, 0, 0, 9, 3, 12, 8, 10, 5, 2, 6, 8, 9, 15, 1, 11, 5, 6, 1, 2, 7, 10, 3, 7, 7, 9, 1, 13, 3, 8, 6, 4, 0, 3, 2, 16, 4, 16, 1, 15, 3, 18, 0, 4, 2, 17, 1, 8, 0, 11, 0, 19, 2, 3, 4, 7, 3, 8, 4, 10, 3, 15, 0, 6, 9, 12, 8, 16, 8, 6, 0, 17, 0, 9, 1, 7, 7, 7, 3, 9, 3, 6, 1, 16, 0, 0, 3, 4, 0, 20, 1, 18, 0, 8, 4, 7, 6, 7, 9, 8, 8, 8, 4, 7, 0, 12, 4, 8, 9, 14, 7, 4, 10, 12, 0, 16, 5, 10, 2, 2, 7, 3, 2, 15, 2, 10, 4, 15, 0, 18, 0, 15, 3, 12, 0, 11, 9, 12, 3, 5, 0, 8, 6, 14, 9, 6, 6, 1, 12, 3, 9, 4, 11, 3, 5, 4, 9, 8, 16, 3, 6, 8, 0, 0, 5, 0, 2, 9, 9, 9, 5, 2, 6, 5, 18, 0, 10, 6, 3, 5, 17, 0, 9, 5, 11, 0, 6, 4, 9, 5, 6, 7, 11, 1, 18, 0, 0, 0, 6, 0, 19, 4, 19, 1, 3, 0, 12, 7, 12, 2, 14, 0, 15, 0, 14, 0, 5, 0, 3, 5, 4, 3, 4, 4, 16, 6, 13, 3, 12, 5, 10, 6, 6, 0, 12, 0, 12, 9, 6, 0, 2, 0, 6, 0, 0, 4, 12, 6, 15, 3, 6, 5, 12, 0, 11, 10, 9, 1, 6, 1, 7, 0, 10, 9, 10, 8, 9, 1, 0, 6, 8, 5, 4, 4, 8, 1, 10, 1, 0, 1, 5, 0, 9, 1, 8, 8, 5, 9, 6, 2, 10, 7, 14, 8, 9, 3, 5, 4, 6, 9, 12, 6, 9, 5, 5, 9, 11, 2, 15, 3, 3, 5, 16, 0, 13, 1, 15, 5, 6, 2, 14, 10, 13, 3, 13, 3, 11, 0, 0, 6, 18, 0, 15, 1, 15, 0, 3, 0, 15, 0, 12, 3, 16, 0, 9};

localparam logic [2912:0][31:0] rectangle1_ys = {4, 4, 9, 18, 5, 5, 8, 14, 0, 6, 4, 8, 2, 9, 6, 0, 11, 5, 8, 5, 0, 6, 6, 18, 7, 3, 8, 6, 5, 6, 21, 6, 1, 1, 8, 6, 12, 1, 13, 1, 2, 5, 4, 3, 1, 6, 1, 1, 5, 10, 13, 4, 4, 5, 1, 10, 17, 3, 3, 1, 7, 7, 12, 6, 7, 15, 17, 4, 1, 0, 5, 8, 14, 15, 15, 6, 5, 0, 0, 6, 0, 6, 6, 8, 0, 0, 7, 6, 20, 6, 13, 6, 6, 12, 22, 7, 7, 6, 14, 18, 1, 16, 4, 4, 4, 16, 12, 0, 10, 8, 8, 0, 0, 14, 16, 8, 19, 10, 9, 0, 6, 5, 5, 14, 13, 16, 0, 6, 1, 2, 8, 9, 12, 16, 16, 1, 2, 8, 5, 17, 7, 1, 5, 1, 1, 0, 0, 7, 10, 9, 15, 7, 6, 8, 8, 6, 7, 14, 10, 12, 0, 0, 3, 0, 1, 0, 0, 18, 3, 3, 10, 10, 11, 11, 11, 10, 13, 4, 0, 0, 0, 1, 1, 6, 14, 14, 18, 4, 17, 2, 8, 5, 5, 4, 0, 15, 0, 0, 22, 0, 6, 1, 5, 1, 2, 8, 12, 12, 7, 1, 2, 4, 1, 15, 5, 5, 0, 4, 0, 0, 6, 7, 17, 18, 18, 20, 15, 4, 6, 14, 9, 6, 6, 10, 16, 6, 0, 0, 7, 20, 5, 2, 1, 0, 0, 21, 7, 7, 8, 15, 15, 0, 6, 1, 2, 14, 6, 2, 4, 17, 7, 1, 13, 13, 6, 12, 1, 0, 2, 2, 18, 6, 7, 3, 4, 1, 2, 3, 3, 0, 8, 8, 14, 14, 10, 0, 1, 6, 9, 0, 0, 0, 11, 9, 8, 12, 12, 12, 7, 7, 0, 0, 3, 3, 2, 10, 14, 13, 5, 17, 18, 0, 4, 4, 3, 1, 16, 3, 5, 2, 14, 21, 14, 2, 4, 6, 8, 14, 6, 6, 7, 3, 12, 6, 6, 9, 6, 6, 2, 18, 2, 2, 10, 0, 0, 0, 12, 6, 12, 5, 8, 6, 12, 12, 1, 1, 9, 21, 13, 13, 6, 0, 7, 4, 0, 0, 12, 12, 12, 12, 14, 13, 15, 0, 1, 1, 14, 3, 1, 0, 6, 10, 15, 1, 9, 0, 15, 15, 7, 12, 8, 14, 10, 3, 17, 13, 0, 3, 5, 7, 6, 8, 15, 1, 8, 5, 2, 7, 7, 6, 1, 1, 18, 4, 16, 7, 7, 2, 20, 12, 2, 0, 0, 15, 8, 3, 5, 4, 6, 4, 4, 4, 22, 14, 14, 11, 11, 9, 12, 0, 0, 17, 17, 6, 6, 4, 0, 0, 15, 8, 12, 2, 20, 0, 13, 10, 3, 5, 7, 0, 0, 1, 17, 15, 15, 16, 13, 0, 4, 5, 4, 0, 0, 7, 7, 5, 13, 0, 7, 2, 2, 2, 6, 5, 6, 0, 3, 7, 7, 7, 6, 14, 0, 2, 4, 3, 4, 0, 6, 0, 10, 21, 6, 5, 2, 7, 7, 17, 18, 6, 18, 18, 9, 9, 3, 17, 15, 17, 3, 3, 0, 0, 0, 0, 3, 11, 0, 0, 8, 12, 0, 6, 0, 2, 7, 6, 1, 4, 3, 1, 0, 0, 13, 5, 1, 2, 10, 4, 10, 10, 14, 7, 1, 1, 5, 9, 16, 12, 14, 13, 5, 5, 5, 5, 1, 1, 15, 9, 2, 2, 0, 0, 17, 5, 2, 2, 7, 7, 0, 0, 6, 7, 6, 6, 3, 0, 9, 7, 6, 0, 14, 14, 12, 2, 16, 16, 0, 0, 8, 5, 13, 14, 6, 0, 1, 6, 0, 11, 20, 11, 12, 11, 11, 4, 15, 0, 0, 2, 0, 18, 7, 14, 2, 3, 6, 8, 4, 8, 2, 16, 0, 2, 11, 3, 16, 17, 13, 9, 7, 8, 2, 17, 18, 3, 6, 0, 0, 10, 11, 5, 6, 5, 3, 21, 10, 4, 8, 9, 6, 6, 5, 4, 4, 10, 10, 2, 2, 4, 4, 4, 4, 18, 18, 2, 2, 5, 8, 7, 5, 14, 14, 11, 9, 6, 19, 5, 5, 4, 6, 10, 7, 2, 18, 9, 2, 0, 3, 2, 5, 0, 3, 14, 9, 11, 5, 6, 6, 5, 5, 10, 10, 0, 3, 1, 7, 12, 6, 7, 18, 2, 3, 2, 0, 0, 5, 22, 10, 1, 0, 3, 15, 13, 8, 8, 2, 5, 8, 8, 6, 0, 9, 0, 5, 5, 5, 4, 16, 16, 9, 13, 10, 9, 0, 11, 5, 5, 6, 6, 5, 6, 13, 5, 2, 15, 17, 13, 10, 6, 14, 12, 10, 0, 11, 2, 4, 0, 17, 6, 10, 16, 16, 16, 11, 11, 3, 4, 0, 16, 15, 15, 17, 8, 6, 8, 8, 5, 6, 7, 5, 9, 8, 8, 11, 0, 2, 0, 0, 3, 10, 0, 3, 4, 0, 5, 0, 4, 10, 10, 11, 10, 12, 21, 20, 15, 17, 12, 6, 13, 16, 5, 1, 19, 1, 2, 10, 11, 9, 10, 7, 0, 6, 0, 2, 17, 0, 0, 17, 7, 3, 2, 2, 1, 16, 13, 15, 5, 13, 2, 14, 12, 13, 8, 12, 16, 1, 2, 6, 7, 0, 8, 12, 21, 0, 6, 4, 7, 8, 8, 14, 11, 12, 0, 10, 2, 0, 6, 6, 11, 11, 16, 6, 16, 7, 10, 4, 18, 0, 3, 0, 1, 1, 16, 3, 16, 3, 9, 4, 7, 7, 4, 12, 3, 6, 6, 3, 3, 6, 1, 17, 18, 5, 6, 2, 7, 0, 8, 7, 5, 9, 14, 14, 8, 11, 0, 0, 1, 11, 18, 9, 10, 6, 14, 7, 4, 16, 13, 8, 16, 0, 5, 5, 6, 7, 10, 12, 10, 0, 4, 10, 6, 11, 8, 11, 9, 12, 4, 4, 9, 5, 9, 0, 9, 9, 4, 3, 1, 6, 18, 8, 19, 8, 8, 12, 7, 1, 12, 0, 0, 3, 6, 11, 8, 17, 14, 3, 3, 0, 0, 11, 11, 11, 20, 6, 0, 3, 5, 12, 0, 0, 5, 12, 13, 1, 0, 2, 2, 10, 10, 6, 12, 14, 1, 11, 15, 14, 3, 6, 6, 1, 1, 15, 15, 1, 3, 0, 3, 5, 0, 1, 7, 3, 3, 7, 7, 13, 5, 1, 1, 15, 2, 5, 15, 12, 12, 0, 2, 7, 9, 5, 5, 17, 18, 17, 17, 17, 0, 0, 14, 13, 20, 9, 10, 8, 10, 10, 15, 5, 13, 17, 12, 9, 9, 7, 4, 8, 7, 15, 8, 17, 17, 1, 7, 5, 4, 16, 16, 0, 6, 4, 0, 1, 6, 9, 2, 2, 3, 1, 9, 10, 0, 4, 1, 8, 0, 22, 15, 0, 7, 14, 14, 5, 5, 5, 5, 2, 2, 0, 4, 16, 0, 12, 21, 5, 5, 6, 5, 14, 5, 8, 6, 13, 10, 13, 0, 1, 4, 3, 13, 13, 13, 16, 16, 16, 16, 0, 1, 2, 15, 2, 2, 2, 2, 0, 12, 2, 10, 3, 7, 11, 8, 0, 0, 3, 18, 18, 3, 7, 3, 17, 5, 6, 16, 2, 2, 4, 13, 1, 12, 7, 5, 11, 11, 4, 2, 0, 0, 0, 0, 2, 13, 7, 8, 14, 0, 15, 9, 4, 10, 5, 18, 18, 20, 8, 8, 5, 5, 6, 0, 4, 4, 12, 0, 12, 12, 15, 15, 0, 0, 6, 12, 4, 22, 7, 0, 1, 16, 7, 10, 2, 9, 2, 2, 3, 13, 14, 2, 4, 1, 6, 21, 5, 6, 6, 3, 10, 15, 4, 0, 0, 0, 7, 0, 10, 2, 5, 0, 0, 2, 2, 0, 0, 2, 10, 7, 0, 3, 7, 6, 2, 6, 0, 0, 0, 17, 17, 14, 15, 15, 14, 8, 7, 8, 0, 8, 5, 6, 7, 8, 8, 10, 5, 12, 9, 14, 9, 18, 6, 6, 16, 16, 11, 6, 7, 6, 7, 10, 12, 14, 12, 13, 0, 1, 16, 17, 2, 0, 0, 2, 1, 8, 8, 5, 5, 4, 7, 15, 2, 1, 1, 1, 1, 11, 11, 6, 10, 9, 18, 21, 12, 6, 6, 4, 12, 14, 7, 13, 7, 12, 2, 0, 9, 10, 10, 15, 16, 2, 5, 0, 16, 12, 15, 10, 9, 11, 7, 15, 8, 4, 6, 6, 7, 8, 8, 3, 3, 2, 2, 3, 3, 3, 3, 11, 11, 8, 6, 18, 4, 1, 11, 12, 12, 0, 12, 20, 4, 2, 8, 7, 0, 11, 0, 7, 17, 10, 5, 11, 4, 0, 4, 4, 18, 0, 4, 4, 11, 6, 0, 9, 15, 7, 15, 12, 12, 12, 7, 7, 4, 4, 11, 16, 15, 15, 1, 21, 20, 1, 17, 16, 16, 16, 10, 18, 5, 2, 7, 6, 0, 7, 1, 18, 2, 7, 1, 0, 3, 15, 10, 3, 0, 0, 0, 4, 17, 20, 3, 3, 6, 6, 9, 18, 0, 1, 0, 10, 16, 16, 12, 16, 6, 6, 9, 9, 4, 8, 3, 3, 1, 5, 6, 10, 4, 2, 4, 4, 8, 8, 13, 13, 13, 2, 2, 2, 0, 2, 5, 3, 21, 10, 10, 8, 8, 8, 15, 13, 8, 13, 15, 4, 15, 15, 11, 6, 2, 2, 1, 7, 6, 11, 16, 0, 11, 9, 5, 2, 3, 15, 0, 0, 1, 0, 2, 2, 2, 4, 1, 1, 5, 4, 5, 5, 5, 0, 8, 6, 3, 18, 8, 2, 5, 4, 6, 1, 4, 6, 17, 6, 6, 5, 2, 2, 6, 3, 3, 3, 1, 2, 2, 14, 8, 0, 0, 6, 5, 7, 16, 17, 8, 13, 17, 17, 0, 2, 3, 17, 17, 18, 15, 13, 14, 18, 13, 14, 2, 9, 3, 2, 4, 5, 5, 6, 4, 4, 7, 9, 0, 3, 1, 22, 10, 0, 0, 2, 13, 21, 1, 7, 0, 1, 1, 2, 5, 2, 2, 11, 7, 9, 9, 4, 6, 21, 21, 5, 10, 0, 2, 0, 12, 13, 0, 1, 13, 21, 3, 10, 3, 2, 1, 0, 1, 18, 15, 10, 9, 11, 7, 2, 2, 4, 5, 7, 4, 0, 1, 0, 0, 1, 0, 5, 0, 14, 14, 18, 0, 4, 2, 1, 8, 15, 10, 17, 4, 0, 6, 9, 9, 11, 2, 0, 15, 18, 17, 11, 11, 9, 16, 16, 1, 2, 15, 11, 18, 14, 7, 8, 1, 14, 7, 12, 0, 0, 0, 0, 8, 8, 21, 0, 0, 6, 6, 0, 0, 16, 0, 0, 1, 1, 13, 0, 5, 10, 7, 10, 6, 2, 13, 6, 13, 20, 4, 6, 0, 13, 16, 0, 6, 5, 15, 7, 6, 6, 0, 0, 18, 15, 3, 3, 14, 14, 15, 17, 0, 0, 16, 0, 7, 8, 9, 0, 1, 4, 1, 2, 1, 0, 17, 14, 15, 21, 15, 15, 6, 3, 1, 4, 1, 2, 2, 2, 7, 3, 6, 1, 8, 0, 16, 16, 19, 16, 8, 15, 18, 18, 3, 5, 5, 6, 2, 6, 2, 8, 5, 8, 0, 12, 12, 7, 14, 6, 6, 13, 10, 10, 9, 3, 0, 12, 0, 0, 2, 2, 0, 0, 6, 6, 1, 1, 0, 10, 9, 9, 7, 15, 10, 4, 2, 0, 9, 2, 0, 15, 14, 1, 0, 3, 2, 4, 16, 16, 18, 0, 3, 12, 3, 3, 8, 15, 13, 6, 9, 0, 3, 3, 5, 4, 7, 0, 0, 0, 1, 2, 13, 13, 2, 9, 6, 8, 7, 12, 10, 6, 12, 15, 14, 8, 10, 10, 9, 12, 12, 12, 12, 12, 10, 15, 10, 1, 4, 5, 10, 12, 0, 10, 2, 20, 10, 17, 0, 0, 2, 2, 7, 1, 14, 13, 6, 2, 6, 19, 15, 5, 6, 6, 0, 0, 5, 5, 1, 13, 1, 17, 13, 18, 14, 1, 4, 0, 5, 5, 1, 1, 0, 4, 6, 18, 18, 15, 7, 7, 9, 13, 15, 15, 13, 13, 5, 18, 19, 19, 19, 14, 0, 1, 9, 15, 0, 10, 10, 8, 5, 5, 4, 4, 7, 6, 4, 0, 1, 1, 14, 3, 3, 2, 2, 7, 22, 16, 3, 10, 16, 0, 5, 8, 1, 6, 3, 13, 12, 5, 5, 6, 1, 19, 14, 6, 0, 0, 1, 8, 7, 12, 1, 1, 7, 10, 7, 3, 0, 0, 5, 5, 0, 0, 2, 1, 0, 17, 18, 17, 15, 15, 14, 10, 18, 12, 10, 10, 2, 6, 14, 14, 1, 21, 1, 16, 1, 0, 1, 1, 7, 14, 1, 0, 1, 1, 0, 14, 7, 11, 5, 6, 1, 1, 9, 4, 16, 0, 5, 3, 12, 11, 10, 9, 2, 6, 8, 1, 1, 14, 16, 16, 4, 19, 8, 1, 8, 8, 5, 6, 12, 12, 6, 6, 0, 1, 6, 6, 17, 22, 12, 12, 12, 14, 6, 7, 3, 1, 1, 2, 2, 12, 2, 6, 6, 0, 0, 6, 1, 7, 7, 20, 6, 2, 3, 4, 1, 0, 2, 2, 15, 17, 6, 0, 4, 6, 12, 14, 14, 18, 3, 3, 6, 5, 4, 16, 8, 6, 5, 1, 1, 10, 2, 0, 1, 6, 1, 4, 0, 16, 16, 0, 3, 7, 9, 14, 14, 21, 21, 4, 7, 4, 15, 13, 6, 16, 5, 8, 8, 8, 8, 8, 6, 8, 5, 5, 1, 10, 17, 16, 10, 4, 18, 18, 16, 15, 15, 1, 1, 5, 5, 0, 4, 0, 0, 5, 6, 2, 2, 0, 4, 0, 0, 7, 7, 8, 0, 10, 0, 1, 1, 6, 12, 9, 10, 18, 16, 14, 14, 10, 13, 13, 0, 8, 5, 0, 11, 5, 18, 8, 7, 0, 0, 2, 8, 9, 7, 2, 0, 14, 12, 12, 6, 0, 8, 6, 11, 3, 12, 16, 6, 10, 10, 12, 12, 15, 15, 20, 20, 17, 2, 1, 15, 2, 12, 7, 1, 8, 3, 6, 0, 0, 15, 7, 6, 21, 3, 7, 2, 10, 9, 5, 9, 11, 13, 0, 18, 4, 8, 3, 15, 18, 14, 15, 6, 6, 6, 14, 8, 6, 9, 9, 15, 20, 18, 18, 16, 16, 2, 2, 0, 20, 6, 9, 6, 6, 4, 6, 0, 1, 0, 0, 12, 12, 5, 6, 5, 16, 8, 8, 4, 4, 7, 19, 11, 1, 2, 13, 0, 11, 1, 10, 19, 10, 1, 1, 4, 4, 6, 9, 5, 2, 0, 0, 7, 2, 0, 6, 8, 18, 14, 15, 0, 0, 4, 0, 0, 2, 6, 1, 0, 0, 2, 0, 2, 11, 8, 8, 8, 11, 9, 4, 17, 21, 4, 15, 8, 12, 17, 16, 1, 1, 13, 1, 4, 8, 7, 7, 6, 6, 9, 1, 6, 5, 6, 4, 8, 10, 5, 4, 4, 7, 6, 5, 7, 7, 2, 1, 13, 13, 15, 15, 0, 6, 7, 9, 6, 7, 12, 14, 17, 12, 17, 3, 17, 1, 17, 5, 7, 4, 1, 5, 0, 11, 7, 7, 17, 6, 15, 15, 10, 10, 15, 1, 0, 0, 1, 21, 9, 4, 1, 9, 1, 0, 0, 6, 1, 12, 17, 1, 0, 6, 0, 7, 12, 9, 1, 11, 11, 10, 2, 16, 16, 13, 16, 16, 18, 13, 2, 8, 13, 20, 8, 7, 6, 20, 20, 1, 1, 3, 2, 9, 3, 0, 9, 4, 4, 13, 13, 15, 13, 0, 2, 1, 1, 6, 2, 11, 1, 0, 3, 1, 7, 0, 0, 9, 15, 7, 9, 17, 3, 1, 15, 0, 3, 1, 0, 6, 0, 0, 11, 7, 6, 14, 14, 0, 0, 1, 12, 8, 6, 5, 9, 8, 12, 19, 0, 4, 16, 7, 7, 6, 17, 17, 4, 0, 0, 0, 4, 12, 9, 5, 5, 7, 1, 0, 6, 8, 6, 12, 4, 1, 1, 10, 4, 13, 13, 15, 14, 14, 8, 10, 10, 7, 10, 1, 15, 6, 1, 6, 18, 0, 13, 6, 6, 6, 7, 8, 8, 8, 2, 10, 10, 7, 7, 9, 2, 2, 1, 2, 3, 8, 8, 18, 6, 6, 3, 6, 8, 2, 14, 2, 3, 6, 2, 17, 7, 11, 1, 0, 0, 7, 2, 1, 0, 0, 0, 15, 18, 8, 6, 2, 7, 6, 2, 9, 4, 8, 8, 0, 0, 0, 0, 2, 2, 6, 0, 1, 4, 5, 13, 14, 2, 1, 1, 4, 5, 1, 12, 12, 18, 13, 3, 9, 3, 2, 6, 6, 9, 9, 6, 6, 16, 20, 10, 6, 1, 13, 15, 12, 11, 6, 0, 0, 3, 3, 5, 5, 2, 2, 0, 0, 11, 11, 6, 16, 16, 6, 7, 6, 1, 9, 5, 11, 8, 8, 6, 5, 7, 0, 0, 6, 6, 6, 21, 19, 18, 18, 16, 16, 0, 0, 14, 14, 14, 14, 18, 18, 5, 3, 0, 0, 12, 3, 4, 4, 14, 14, 6, 11, 5, 4, 8, 8, 6, 14, 6, 6, 14, 5, 5, 0, 3, 3, 12, 10, 8, 14, 10, 10, 12, 8, 11, 11, 2, 2, 12, 10, 9, 8, 7, 0, 0, 5, 6, 0, 1, 0, 3, 14, 9, 2, 4, 4, 5, 7, 5, 5, 4, 14, 17, 16, 17, 20, 14, 6, 4, 3, 8, 6, 6, 5, 5, 5, 2, 1, 2, 0, 9, 0, 0, 0, 1, 9, 8, 9, 9, 0, 1, 1, 20, 0, 8, 8, 13, 13, 8, 8, 11, 11, 12, 1, 11, 10, 8, 8, 14, 18, 16, 20, 12, 12, 17, 6, 17, 18, 15, 13, 17, 17, 17, 17, 2, 13, 1};

localparam logic [2912:0][31:0] rectangle1_widths = {12, 12, 18, 9, 4, 12, 12, 4, 7, 12, 12, 19, 24, 6, 14, 14, 9, 6, 6, 4, 6, 24, 6, 10, 14, 24, 15, 5, 6, 3, 18, 13, 6, 6, 24, 14, 21, 4, 20, 6, 4, 22, 6, 6, 4, 19, 4, 4, 14, 18, 4, 6, 12, 12, 24, 18, 12, 4, 4, 24, 8, 3, 16, 12, 6, 9, 18, 16, 4, 18, 20, 14, 7, 9, 9, 8, 14, 12, 6, 6, 6, 6, 6, 18, 12, 24, 16, 6, 24, 4, 15, 4, 4, 6, 18, 4, 8, 10, 10, 18, 22, 18, 6, 4, 4, 20, 8, 6, 6, 12, 12, 6, 6, 9, 9, 6, 12, 20, 18, 18, 14, 10, 12, 18, 8, 18, 6, 12, 4, 19, 22, 11, 15, 12, 12, 5, 24, 12, 9, 6, 22, 17, 6, 6, 6, 6, 6, 8, 19, 6, 17, 3, 8, 9, 9, 10, 3, 24, 18, 6, 10, 9, 16, 9, 20, 9, 9, 10, 6, 12, 18, 22, 8, 6, 6, 11, 24, 22, 20, 2, 2, 2, 2, 3, 9, 9, 18, 8, 18, 12, 14, 6, 6, 9, 18, 5, 4, 18, 19, 4, 19, 6, 14, 20, 22, 7, 22, 22, 6, 9, 4, 12, 6, 18, 6, 16, 6, 24, 4, 4, 6, 6, 9, 14, 18, 15, 15, 16, 10, 15, 10, 6, 18, 18, 18, 14, 2, 2, 15, 21, 5, 24, 22, 15, 24, 18, 10, 10, 6, 20, 10, 16, 7, 6, 6, 12, 10, 6, 5, 24, 5, 6, 6, 6, 3, 13, 4, 9, 6, 6, 12, 6, 12, 8, 10, 6, 2, 6, 2, 2, 9, 9, 9, 9, 18, 24, 8, 4, 10, 3, 6, 6, 24, 13, 6, 16, 6, 6, 10, 6, 6, 6, 6, 6, 9, 6, 6, 5, 3, 18, 19, 6, 3, 3, 18, 6, 9, 20, 6, 22, 5, 18, 6, 24, 12, 12, 14, 8, 5, 3, 18, 20, 19, 6, 6, 6, 6, 6, 6, 15, 6, 6, 18, 12, 6, 6, 9, 13, 9, 6, 9, 3, 9, 10, 4, 4, 6, 18, 10, 22, 16, 18, 8, 6, 6, 6, 6, 6, 9, 9, 19, 19, 10, 10, 6, 6, 6, 9, 4, 14, 6, 18, 9, 21, 17, 11, 13, 9, 15, 6, 18, 24, 3, 24, 10, 18, 18, 16, 3, 18, 6, 6, 6, 18, 12, 6, 24, 5, 5, 6, 6, 19, 12, 4, 10, 10, 10, 9, 21, 9, 9, 4, 4, 9, 18, 6, 11, 6, 9, 6, 6, 9, 19, 6, 6, 4, 4, 18, 6, 6, 6, 18, 18, 11, 14, 15, 22, 24, 18, 12, 7, 22, 14, 24, 18, 22, 11, 6, 24, 10, 10, 24, 18, 16, 16, 18, 21, 6, 6, 9, 2, 6, 6, 6, 4, 24, 10, 6, 6, 9, 6, 10, 2, 15, 6, 6, 9, 14, 8, 7, 4, 6, 6, 21, 5, 4, 5, 11, 12, 24, 23, 18, 21, 6, 4, 8, 15, 10, 9, 6, 9, 9, 9, 9, 6, 18, 21, 6, 6, 6, 16, 10, 10, 10, 6, 12, 3, 6, 9, 8, 3, 4, 9, 24, 6, 6, 6, 12, 2, 12, 18, 18, 24, 4, 6, 6, 8, 16, 8, 8, 11, 24, 4, 4, 16, 6, 18, 6, 9, 8, 3, 18, 6, 6, 4, 4, 18, 12, 9, 9, 6, 6, 9, 3, 14, 3, 14, 14, 9, 9, 6, 6, 6, 6, 8, 9, 8, 10, 4, 6, 18, 8, 24, 3, 10, 10, 10, 24, 15, 12, 14, 4, 6, 6, 18, 14, 6, 6, 24, 6, 10, 6, 6, 11, 10, 6, 6, 4, 20, 10, 6, 10, 4, 10, 12, 8, 4, 9, 14, 19, 10, 16, 24, 18, 18, 18, 9, 23, 18, 12, 3, 10, 10, 6, 4, 6, 6, 9, 6, 3, 9, 3, 6, 18, 18, 8, 9, 9, 5, 14, 3, 15, 15, 6, 6, 6, 6, 6, 6, 8, 8, 10, 21, 12, 12, 12, 6, 20, 12, 8, 8, 20, 12, 16, 9, 12, 14, 9, 19, 6, 18, 4, 20, 22, 4, 4, 6, 6, 10, 12, 24, 4, 4, 17, 18, 14, 14, 3, 3, 14, 9, 18, 12, 8, 7, 22, 4, 7, 9, 22, 6, 8, 6, 6, 9, 18, 12, 4, 4, 6, 9, 8, 6, 6, 4, 19, 9, 12, 18, 4, 18, 4, 4, 4, 6, 4, 18, 20, 6, 8, 3, 14, 24, 18, 5, 5, 8, 8, 12, 6, 6, 12, 23, 19, 11, 8, 10, 9, 9, 9, 20, 9, 9, 8, 21, 10, 12, 23, 8, 18, 9, 9, 6, 6, 24, 18, 24, 18, 9, 9, 18, 6, 6, 5, 6, 6, 8, 21, 3, 11, 10, 12, 18, 22, 6, 6, 6, 6, 18, 3, 16, 6, 16, 18, 6, 8, 10, 10, 12, 8, 9, 24, 18, 9, 10, 4, 9, 6, 12, 20, 9, 9, 4, 8, 9, 12, 9, 6, 5, 21, 10, 6, 18, 8, 18, 9, 18, 12, 6, 4, 4, 24, 9, 9, 19, 22, 6, 20, 6, 16, 8, 6, 16, 16, 4, 8, 12, 6, 8, 6, 6, 21, 16, 7, 4, 6, 6, 4, 6, 12, 23, 6, 12, 10, 6, 9, 9, 18, 18, 12, 21, 12, 6, 19, 14, 18, 4, 11, 9, 4, 4, 18, 11, 20, 13, 22, 14, 10, 10, 6, 9, 8, 16, 14, 9, 18, 9, 24, 10, 18, 6, 11, 12, 4, 4, 6, 15, 6, 6, 6, 6, 16, 20, 4, 4, 18, 6, 9, 15, 19, 7, 9, 8, 18, 12, 9, 14, 22, 6, 10, 10, 16, 6, 8, 6, 8, 4, 8, 10, 14, 20, 4, 12, 12, 6, 8, 8, 9, 16, 6, 3, 5, 5, 10, 23, 21, 6, 12, 8, 24, 8, 8, 8, 5, 19, 24, 13, 24, 4, 6, 12, 12, 18, 9, 4, 4, 9, 9, 6, 6, 19, 18, 16, 9, 4, 15, 8, 6, 6, 12, 11, 21, 8, 6, 21, 19, 6, 6, 14, 9, 8, 22, 9, 18, 7, 16, 12, 4, 4, 4, 6, 6, 3, 6, 3, 12, 4, 3, 3, 10, 3, 6, 19, 18, 18, 6, 20, 20, 6, 24, 18, 6, 8, 8, 14, 4, 5, 8, 22, 6, 9, 19, 9, 18, 9, 24, 14, 9, 6, 13, 6, 21, 9, 9, 10, 24, 9, 6, 9, 6, 14, 14, 9, 6, 10, 4, 6, 6, 9, 9, 9, 4, 12, 9, 10, 10, 24, 9, 24, 11, 22, 6, 20, 14, 16, 19, 10, 4, 21, 6, 14, 6, 9, 4, 19, 20, 4, 8, 6, 6, 4, 4, 6, 6, 24, 6, 4, 4, 9, 6, 7, 14, 6, 4, 6, 6, 10, 14, 12, 12, 6, 20, 9, 6, 5, 16, 8, 6, 9, 9, 9, 9, 18, 18, 18, 19, 6, 15, 6, 6, 6, 22, 21, 18, 6, 18, 8, 18, 6, 6, 2, 2, 7, 9, 21, 7, 22, 24, 9, 12, 14, 14, 6, 6, 20, 9, 21, 14, 12, 9, 6, 6, 18, 6, 6, 6, 6, 6, 24, 18, 10, 12, 19, 4, 9, 15, 12, 6, 6, 16, 14, 20, 20, 6, 12, 12, 6, 6, 6, 6, 9, 15, 9, 9, 9, 9, 8, 4, 10, 4, 10, 18, 11, 12, 12, 9, 15, 12, 12, 12, 8, 8, 24, 8, 4, 4, 15, 24, 5, 18, 3, 4, 9, 20, 18, 10, 4, 6, 6, 6, 9, 18, 20, 4, 6, 18, 18, 6, 6, 6, 20, 20, 18, 6, 22, 6, 6, 24, 6, 6, 6, 6, 6, 9, 18, 9, 23, 18, 9, 8, 15, 8, 6, 8, 6, 4, 12, 8, 8, 6, 6, 12, 18, 8, 22, 12, 20, 20, 10, 18, 19, 6, 22, 7, 11, 10, 9, 6, 6, 6, 6, 6, 9, 18, 13, 8, 8, 8, 6, 6, 6, 5, 5, 6, 6, 12, 24, 2, 2, 2, 2, 6, 6, 18, 7, 12, 18, 20, 6, 18, 18, 6, 9, 18, 6, 12, 12, 6, 4, 9, 12, 6, 6, 9, 12, 20, 12, 3, 15, 6, 12, 8, 8, 9, 12, 6, 9, 8, 6, 24, 6, 5, 5, 6, 6, 6, 6, 18, 9, 10, 10, 6, 6, 10, 6, 18, 6, 9, 6, 4, 4, 12, 10, 22, 2, 24, 10, 8, 6, 5, 20, 12, 6, 10, 12, 6, 4, 6, 4, 4, 19, 2, 2, 2, 10, 4, 6, 16, 6, 6, 6, 12, 9, 9, 18, 22, 6, 6, 16, 9, 6, 6, 6, 24, 24, 6, 18, 18, 22, 9, 21, 12, 24, 4, 6, 6, 6, 6, 20, 12, 4, 12, 4, 3, 10, 12, 6, 4, 6, 6, 6, 4, 18, 22, 10, 10, 12, 12, 5, 21, 9, 12, 12, 8, 10, 10, 12, 10, 12, 4, 6, 6, 11, 6, 4, 4, 8, 16, 18, 16, 8, 9, 8, 8, 8, 8, 5, 7, 24, 8, 8, 24, 12, 12, 6, 8, 18, 18, 22, 12, 12, 12, 6, 9, 7, 9, 18, 4, 6, 6, 12, 14, 17, 12, 9, 24, 9, 18, 9, 9, 24, 20, 16, 4, 10, 6, 7, 7, 6, 19, 9, 9, 10, 18, 4, 4, 8, 12, 6, 12, 10, 21, 9, 6, 6, 12, 20, 10, 5, 4, 8, 24, 4, 18, 16, 6, 14, 8, 20, 9, 6, 4, 4, 8, 2, 9, 19, 9, 18, 6, 6, 4, 18, 14, 18, 9, 12, 7, 20, 9, 15, 6, 6, 9, 9, 12, 6, 8, 24, 6, 8, 24, 12, 9, 16, 4, 5, 9, 9, 6, 20, 17, 7, 23, 6, 4, 6, 18, 9, 2, 2, 18, 15, 18, 4, 10, 10, 6, 6, 6, 18, 6, 6, 11, 10, 10, 10, 6, 10, 16, 16, 22, 8, 6, 6, 6, 7, 8, 6, 3, 8, 19, 4, 18, 5, 4, 16, 18, 10, 12, 12, 22, 9, 12, 10, 8, 8, 18, 10, 21, 22, 6, 3, 12, 12, 22, 18, 22, 6, 6, 6, 18, 6, 12, 12, 18, 6, 6, 6, 18, 6, 6, 10, 5, 5, 9, 23, 8, 6, 9, 18, 11, 11, 24, 8, 14, 21, 24, 8, 21, 12, 4, 4, 6, 9, 19, 10, 18, 6, 17, 12, 6, 16, 5, 18, 6, 20, 15, 6, 6, 6, 9, 6, 6, 6, 6, 6, 6, 6, 9, 3, 14, 12, 4, 6, 4, 6, 14, 16, 6, 21, 6, 5, 16, 14, 4, 12, 12, 14, 18, 18, 24, 18, 9, 19, 24, 9, 9, 18, 18, 3, 8, 18, 3, 4, 10, 6, 10, 5, 12, 9, 8, 5, 14, 10, 4, 6, 18, 6, 6, 4, 6, 9, 14, 15, 8, 6, 6, 12, 12, 16, 18, 18, 24, 9, 24, 22, 9, 10, 6, 12, 12, 16, 10, 18, 9, 10, 18, 15, 15, 24, 6, 6, 6, 10, 18, 10, 10, 14, 9, 6, 6, 8, 4, 3, 16, 6, 6, 12, 12, 6, 6, 9, 9, 6, 6, 4, 12, 12, 12, 14, 20, 8, 13, 6, 6, 12, 15, 12, 18, 24, 3, 4, 4, 12, 17, 5, 5, 18, 12, 6, 6, 21, 6, 12, 16, 18, 15, 9, 15, 3, 3, 10, 16, 12, 9, 6, 6, 10, 18, 14, 14, 3, 5, 12, 20, 19, 9, 14, 14, 9, 18, 6, 18, 20, 20, 24, 20, 9, 9, 8, 8, 4, 20, 6, 21, 13, 12, 10, 5, 6, 18, 9, 21, 22, 18, 6, 6, 6, 6, 6, 4, 9, 9, 15, 3, 12, 20, 6, 18, 4, 4, 6, 6, 6, 6, 16, 6, 6, 18, 10, 10, 9, 6, 5, 8, 19, 12, 21, 16, 18, 10, 4, 18, 12, 6, 6, 6, 18, 12, 10, 10, 6, 6, 8, 12, 10, 10, 18, 4, 24, 6, 20, 19, 10, 21, 8, 10, 4, 6, 4, 4, 9, 16, 16, 24, 9, 14, 7, 8, 12, 4, 3, 9, 20, 24, 12, 8, 6, 10, 14, 10, 9, 24, 12, 22, 12, 9, 23, 19, 6, 18, 6, 4, 6, 6, 4, 8, 7, 18, 4, 4, 20, 6, 10, 4, 8, 8, 6, 6, 6, 6, 24, 10, 23, 19, 18, 9, 6, 6, 20, 6, 18, 9, 18, 18, 18, 10, 4, 4, 4, 12, 4, 10, 4, 3, 4, 6, 19, 9, 7, 14, 8, 8, 18, 9, 18, 6, 6, 4, 4, 4, 18, 6, 8, 18, 14, 15, 10, 4, 22, 6, 6, 4, 10, 8, 12, 12, 6, 6, 4, 19, 6, 8, 6, 6, 6, 24, 10, 10, 19, 19, 16, 24, 6, 6, 18, 18, 6, 6, 6, 4, 6, 10, 6, 6, 6, 6, 6, 15, 20, 4, 12, 6, 9, 6, 12, 18, 18, 18, 6, 12, 18, 4, 19, 15, 14, 22, 6, 18, 3, 20, 5, 12, 6, 8, 8, 12, 6, 3, 14, 12, 4, 15, 6, 10, 18, 15, 8, 24, 6, 8, 10, 18, 24, 6, 8, 18, 18, 18, 20, 14, 12, 21, 21, 18, 18, 4, 18, 4, 10, 11, 4, 9, 4, 8, 8, 12, 9, 12, 9, 12, 4, 14, 11, 6, 11, 9, 18, 12, 18, 18, 9, 9, 9, 6, 6, 6, 6, 6, 4, 6, 6, 18, 6, 15, 15, 4, 6, 8, 8, 24, 14, 8, 10, 8, 4, 6, 6, 18, 16, 16, 8, 16, 12, 9, 9, 16, 19, 9, 3, 24, 5, 19, 6, 24, 9, 10, 20, 7, 7, 2, 10, 12, 3, 12, 6, 9, 22, 22, 9, 4, 18, 24, 24, 18, 4, 10, 6, 6, 6, 6, 6, 6, 6, 10, 10, 9, 14, 10, 10, 3, 9, 5, 24, 12, 4, 9, 6, 6, 19, 4, 6, 18, 10, 18, 9, 24, 8, 4, 8, 10, 18, 19, 24, 8, 10, 6, 7, 12, 6, 15, 6, 7, 6, 6, 6, 4, 6, 6, 9, 18, 9, 9, 18, 18, 4, 4, 2, 16, 4, 10, 6, 7, 4, 6, 10, 18, 2, 2, 6, 6, 18, 9, 9, 10, 5, 5, 4, 4, 10, 14, 12, 24, 14, 6, 4, 14, 16, 21, 15, 6, 16, 16, 3, 3, 10, 6, 12, 5, 9, 11, 4, 9, 13, 4, 6, 10, 20, 9, 4, 4, 22, 9, 24, 16, 18, 6, 9, 9, 4, 7, 20, 19, 6, 6, 4, 9, 18, 2, 8, 18, 15, 12, 6, 20, 24, 9, 4, 4, 8, 6, 3, 12, 5, 5, 6, 6, 14, 3, 6, 4, 16, 7, 8, 6, 9, 3, 22, 18, 6, 9, 4, 4, 10, 3, 18, 18, 9, 9, 18, 6, 10, 18, 18, 9, 6, 18, 9, 10, 9, 3, 9, 11, 9, 11, 8, 20, 21, 12, 6, 8, 8, 8, 9, 8, 9, 9, 9, 9, 10, 6, 6, 10, 16, 19, 18, 9, 6, 6, 14, 8, 7, 12, 8, 22, 6, 6, 6, 17, 12, 18, 10, 10, 24, 6, 6, 19, 6, 10, 10, 9, 18, 18, 9, 9, 6, 4, 8, 18, 4, 12, 4, 18, 18, 6, 6, 4, 6, 12, 4, 6, 12, 8, 8, 9, 9, 18, 9, 18, 6, 9, 9, 14, 6, 12, 18, 6, 16, 3, 6, 4, 4, 5, 9, 18, 5, 17, 18, 24, 18, 6, 14, 3, 6, 6, 6, 21, 12, 9, 6, 8, 8, 8, 8, 12, 18, 20, 9, 8, 16, 10, 10, 15, 18, 10, 18, 10, 10, 18, 18, 18, 6, 8, 8, 8, 18, 9, 18, 6, 6, 18, 12, 6, 2, 10, 20, 12, 3, 3, 3, 18, 10, 14, 14, 9, 8, 4, 5, 9, 9, 12, 5, 3, 6, 7, 4, 14, 19, 6, 15, 10, 8, 12, 9, 14, 14, 13, 6, 17, 17, 8, 8, 24, 15, 18, 18, 3, 3, 6, 6, 11, 12, 12, 9, 12, 6, 9, 6, 9, 16, 10, 7, 11, 12, 8, 4, 3, 3, 18, 4, 3, 18, 3, 3, 5, 18, 20, 9, 19, 19, 9, 18, 14, 6, 9, 9, 6, 6, 6, 6, 12, 12, 4, 6, 3, 18, 16, 10, 9, 9, 10, 3, 12, 12, 8, 6, 12, 12, 6, 7, 18, 19, 12, 6, 6, 5, 5, 14, 3, 24, 20, 18, 6, 20, 6, 6, 6, 18, 15, 18, 3, 6, 6, 8, 8, 20, 13, 7, 7, 10, 10, 3, 18, 18, 9, 15, 12, 12, 6, 13, 22, 6, 6, 24, 10, 18, 10, 3, 12, 4, 4, 18, 9, 12, 9, 10, 10, 10, 10, 9, 9, 10, 10, 18, 18, 18, 7, 19, 16, 16, 12, 2, 2, 8, 8, 3, 12, 8, 12, 18, 18, 3, 18, 3, 3, 18, 18, 22, 21, 18, 18, 24, 16, 6, 8, 6, 6, 18, 10, 9, 9, 3, 3, 6, 6, 16, 9, 16, 18, 6, 6, 4, 6, 6, 18, 24, 9, 8, 13, 16, 14, 9, 16, 13, 13, 24, 10, 18, 18, 9, 22, 8, 8, 18, 5, 12, 18, 4, 6, 2, 2, 10, 18, 17, 12, 16, 5, 6, 6, 6, 13, 19, 6, 4, 6, 6, 6, 18, 4, 8, 8, 10, 10, 4, 4, 16, 16, 7, 3, 9, 17, 8, 8, 10, 22, 24, 12, 6, 6, 9, 22, 9, 18, 19, 18, 9, 9, 9, 9, 3, 24, 6};

localparam logic [2912:0][31:0] rectangle1_heights = {9, 7, 9, 6, 19, 16, 6, 10, 6, 6, 7, 12, 3, 15, 10, 9, 6, 10, 10, 9, 11, 13, 9, 6, 12, 3, 6, 14, 10, 12, 3, 6, 15, 15, 15, 12, 12, 10, 10, 13, 13, 19, 9, 11, 9, 3, 9, 9, 14, 2, 11, 9, 9, 6, 5, 6, 6, 13, 13, 23, 12, 14, 6, 6, 12, 6, 3, 12, 20, 2, 14, 12, 9, 6, 6, 10, 14, 5, 9, 9, 9, 9, 9, 4, 9, 6, 12, 6, 3, 9, 4, 9, 9, 12, 2, 10, 10, 6, 4, 2, 3, 3, 15, 10, 10, 6, 9, 9, 6, 6, 6, 9, 9, 6, 6, 10, 3, 2, 12, 24, 10, 12, 12, 3, 8, 6, 6, 18, 14, 2, 13, 4, 10, 6, 6, 12, 4, 4, 6, 6, 15, 9, 10, 8, 7, 22, 22, 16, 6, 12, 6, 14, 10, 11, 11, 18, 14, 8, 14, 6, 16, 6, 4, 6, 4, 6, 6, 6, 9, 6, 3, 3, 8, 6, 6, 6, 4, 12, 17, 24, 24, 22, 22, 18, 6, 4, 3, 18, 3, 4, 6, 6, 16, 16, 9, 8, 9, 3, 2, 9, 18, 9, 12, 2, 3, 9, 4, 4, 11, 6, 10, 12, 15, 3, 9, 6, 9, 14, 13, 13, 9, 9, 6, 6, 4, 4, 9, 4, 6, 10, 14, 9, 3, 3, 4, 6, 18, 18, 10, 4, 18, 6, 8, 9, 19, 3, 4, 4, 16, 4, 6, 9, 15, 13, 14, 10, 6, 14, 12, 5, 12, 12, 6, 6, 16, 6, 9, 6, 9, 9, 6, 9, 3, 21, 12, 9, 20, 9, 21, 23, 4, 4, 6, 6, 4, 19, 12, 10, 12, 19, 10, 12, 2, 4, 9, 4, 9, 9, 4, 9, 9, 9, 15, 15, 4, 7, 10, 8, 16, 3, 3, 9, 18, 18, 9, 14, 6, 16, 12, 16, 10, 3, 10, 4, 9, 5, 12, 10, 14, 16, 8, 2, 6, 9, 14, 12, 18, 18, 9, 6, 9, 9, 2, 6, 9, 9, 6, 6, 6, 15, 6, 14, 6, 4, 19, 19, 9, 3, 9, 4, 6, 22, 14, 20, 9, 9, 12, 12, 6, 6, 3, 3, 6, 12, 12, 12, 9, 12, 12, 8, 9, 3, 6, 23, 4, 18, 6, 6, 4, 9, 3, 4, 12, 3, 6, 3, 9, 9, 12, 4, 9, 10, 9, 21, 7, 9, 4, 12, 12, 9, 17, 9, 6, 19, 7, 12, 12, 6, 4, 6, 6, 14, 14, 6, 5, 11, 14, 9, 6, 9, 9, 4, 2, 9, 9, 9, 9, 7, 10, 9, 9, 3, 3, 12, 6, 4, 2, 24, 4, 9, 12, 6, 3, 16, 4, 2, 8, 6, 6, 10, 10, 4, 3, 6, 6, 3, 10, 24, 11, 6, 20, 24, 24, 14, 12, 14, 6, 9, 14, 15, 9, 14, 18, 6, 10, 9, 7, 3, 6, 12, 18, 9, 13, 3, 12, 10, 8, 9, 5, 5, 6, 3, 6, 12, 15, 10, 12, 6, 6, 16, 6, 6, 6, 6, 9, 3, 6, 6, 9, 9, 10, 16, 5, 5, 10, 6, 18, 9, 7, 10, 18, 9, 6, 3, 9, 10, 12, 12, 21, 8, 8, 3, 4, 9, 9, 22, 14, 15, 14, 14, 6, 9, 16, 16, 8, 9, 3, 9, 6, 10, 18, 3, 11, 11, 9, 9, 9, 4, 6, 6, 17, 17, 4, 18, 12, 12, 15, 15, 6, 6, 14, 9, 15, 15, 9, 21, 12, 12, 18, 9, 3, 10, 4, 20, 8, 8, 9, 3, 4, 6, 6, 10, 7, 6, 3, 18, 6, 6, 3, 7, 6, 6, 7, 12, 4, 9, 9, 15, 3, 6, 11, 9, 9, 4, 6, 10, 16, 4, 9, 8, 8, 18, 11, 5, 3, 3, 6, 10, 3, 3, 22, 6, 6, 12, 9, 9, 9, 6, 9, 19, 6, 19, 9, 3, 4, 10, 6, 8, 12, 6, 19, 20, 20, 6, 6, 14, 14, 7, 9, 10, 10, 6, 6, 6, 6, 6, 9, 6, 6, 10, 10, 13, 5, 6, 4, 5, 12, 6, 3, 9, 2, 18, 3, 3, 18, 23, 19, 9, 6, 12, 6, 10, 15, 6, 8, 6, 6, 18, 18, 4, 4, 9, 8, 5, 8, 4, 15, 8, 4, 4, 17, 18, 12, 9, 12, 2, 6, 11, 10, 17, 6, 9, 12, 12, 15, 3, 7, 9, 3, 12, 14, 9, 18, 18, 10, 11, 3, 3, 12, 8, 12, 14, 10, 2, 12, 12, 18, 18, 12, 9, 11, 12, 3, 3, 4, 5, 4, 9, 6, 6, 8, 18, 10, 5, 6, 14, 4, 4, 10, 3, 4, 4, 6, 6, 6, 3, 4, 3, 6, 6, 3, 10, 9, 8, 8, 11, 9, 6, 12, 12, 8, 3, 4, 22, 8, 9, 9, 14, 8, 14, 20, 10, 4, 4, 9, 5, 4, 4, 5, 10, 8, 3, 4, 6, 4, 12, 6, 9, 4, 3, 9, 4, 18, 12, 8, 5, 6, 9, 12, 6, 6, 15, 2, 6, 2, 6, 3, 5, 9, 9, 9, 4, 6, 6, 3, 12, 6, 3, 10, 6, 9, 14, 6, 8, 12, 10, 6, 9, 12, 9, 6, 3, 6, 6, 14, 9, 14, 16, 10, 5, 3, 12, 5, 4, 12, 6, 6, 13, 13, 6, 3, 6, 14, 2, 4, 4, 9, 4, 6, 23, 23, 3, 4, 3, 4, 15, 3, 4, 4, 9, 6, 10, 6, 6, 6, 2, 6, 3, 6, 3, 16, 6, 22, 10, 18, 9, 10, 9, 10, 10, 10, 9, 3, 13, 13, 7, 9, 6, 6, 2, 16, 6, 12, 3, 6, 4, 14, 6, 9, 10, 10, 6, 9, 14, 12, 12, 9, 16, 6, 14, 2, 16, 10, 4, 7, 16, 16, 6, 12, 8, 18, 14, 14, 6, 18, 3, 9, 6, 16, 4, 16, 16, 10, 8, 2, 9, 8, 3, 11, 9, 8, 6, 3, 6, 9, 9, 19, 19, 8, 8, 3, 4, 6, 6, 14, 12, 5, 9, 9, 8, 6, 3, 12, 12, 2, 3, 14, 14, 14, 6, 9, 4, 6, 3, 9, 4, 5, 9, 10, 10, 9, 9, 19, 9, 19, 4, 9, 19, 12, 5, 18, 12, 3, 3, 4, 9, 4, 4, 6, 8, 3, 6, 5, 5, 6, 15, 12, 14, 6, 6, 4, 3, 4, 3, 4, 3, 4, 6, 9, 4, 12, 3, 6, 7, 8, 3, 6, 9, 4, 6, 10, 10, 17, 20, 4, 9, 9, 16, 4, 4, 6, 10, 6, 8, 8, 8, 4, 6, 6, 4, 4, 18, 4, 14, 6, 3, 4, 15, 3, 6, 9, 9, 9, 21, 2, 3, 13, 8, 9, 9, 10, 10, 6, 6, 21, 13, 21, 20, 6, 9, 9, 3, 9, 10, 9, 9, 4, 14, 6, 12, 10, 8, 6, 9, 14, 6, 9, 10, 6, 6, 6, 6, 3, 3, 3, 2, 11, 6, 11, 11, 9, 4, 12, 3, 9, 3, 9, 3, 9, 9, 18, 18, 9, 6, 3, 9, 3, 16, 4, 8, 6, 6, 9, 9, 10, 8, 15, 8, 4, 6, 6, 6, 2, 11, 15, 13, 9, 9, 4, 4, 4, 3, 3, 20, 6, 4, 7, 9, 9, 6, 6, 4, 6, 9, 8, 8, 9, 16, 12, 12, 6, 22, 6, 6, 6, 6, 10, 16, 6, 10, 6, 2, 6, 10, 6, 4, 16, 13, 6, 9, 6, 6, 11, 10, 10, 21, 9, 6, 16, 3, 12, 9, 8, 2, 3, 6, 18, 9, 9, 9, 6, 2, 4, 12, 12, 22, 22, 11, 11, 9, 3, 2, 2, 9, 9, 9, 9, 6, 10, 9, 9, 9, 9, 6, 3, 6, 6, 3, 6, 10, 6, 10, 12, 10, 9, 18, 4, 10, 10, 14, 19, 6, 6, 10, 8, 6, 18, 12, 8, 3, 3, 9, 4, 12, 9, 8, 7, 9, 12, 6, 9, 23, 6, 3, 14, 12, 12, 7, 9, 12, 12, 15, 15, 9, 15, 8, 4, 19, 19, 20, 20, 12, 12, 14, 8, 12, 5, 3, 12, 3, 3, 9, 6, 4, 14, 6, 9, 6, 10, 6, 6, 9, 9, 6, 6, 3, 6, 24, 4, 12, 8, 14, 14, 10, 6, 9, 7, 10, 9, 12, 14, 8, 8, 6, 6, 9, 9, 6, 6, 8, 8, 12, 11, 4, 7, 3, 9, 7, 6, 11, 11, 18, 5, 3, 20, 4, 4, 10, 14, 8, 9, 8, 6, 4, 9, 8, 17, 6, 17, 17, 3, 18, 18, 18, 8, 9, 9, 8, 9, 9, 9, 6, 6, 6, 3, 6, 6, 6, 6, 4, 9, 9, 23, 3, 4, 23, 3, 3, 4, 6, 3, 6, 4, 15, 12, 9, 9, 9, 3, 6, 13, 4, 13, 18, 5, 8, 9, 9, 14, 14, 16, 10, 6, 4, 5, 5, 16, 16, 15, 2, 6, 4, 12, 12, 8, 8, 5, 8, 6, 18, 14, 14, 12, 16, 21, 21, 18, 8, 12, 12, 20, 6, 20, 20, 14, 14, 8, 9, 10, 11, 16, 6, 9, 12, 9, 10, 3, 2, 3, 9, 6, 6, 9, 6, 12, 6, 4, 16, 9, 9, 10, 6, 8, 21, 9, 3, 10, 3, 4, 6, 6, 6, 12, 15, 4, 8, 10, 10, 12, 8, 4, 4, 6, 2, 9, 9, 10, 13, 6, 3, 6, 5, 9, 9, 7, 6, 6, 4, 18, 9, 14, 6, 9, 3, 6, 9, 6, 10, 3, 6, 9, 11, 11, 10, 18, 6, 3, 6, 5, 9, 9, 15, 3, 6, 3, 6, 6, 8, 3, 6, 4, 6, 9, 6, 6, 6, 9, 10, 4, 6, 10, 6, 8, 6, 4, 10, 8, 12, 12, 9, 12, 16, 6, 2, 9, 9, 13, 2, 6, 24, 24, 10, 6, 3, 11, 4, 18, 16, 16, 6, 2, 6, 6, 6, 4, 7, 7, 6, 8, 3, 3, 14, 10, 12, 18, 9, 9, 10, 12, 12, 10, 2, 13, 3, 12, 15, 4, 3, 8, 6, 3, 4, 6, 5, 7, 10, 10, 6, 9, 6, 16, 22, 12, 18, 18, 4, 4, 6, 9, 9, 9, 3, 13, 4, 6, 3, 12, 9, 13, 2, 9, 9, 8, 8, 8, 6, 15, 12, 9, 4, 3, 6, 6, 6, 8, 6, 3, 3, 5, 3, 6, 10, 10, 12, 6, 2, 10, 12, 12, 9, 11, 13, 6, 12, 3, 6, 3, 10, 9, 9, 9, 6, 9, 9, 16, 16, 9, 9, 6, 6, 16, 12, 6, 20, 9, 9, 9, 4, 12, 9, 4, 9, 8, 16, 6, 15, 8, 4, 6, 10, 21, 21, 3, 6, 2, 2, 4, 4, 2, 3, 23, 6, 3, 23, 10, 12, 14, 9, 12, 10, 4, 10, 12, 24, 4, 10, 9, 3, 9, 9, 18, 11, 4, 8, 9, 10, 12, 12, 4, 10, 6, 9, 5, 22, 6, 8, 4, 6, 4, 9, 6, 6, 9, 6, 3, 6, 9, 3, 6, 6, 4, 12, 9, 12, 6, 9, 9, 8, 6, 7, 12, 12, 6, 14, 18, 12, 14, 14, 20, 20, 17, 17, 6, 6, 13, 13, 9, 7, 6, 6, 9, 3, 10, 9, 18, 9, 4, 12, 5, 3, 5, 18, 14, 9, 6, 4, 8, 8, 2, 5, 12, 12, 3, 12, 6, 9, 5, 6, 6, 11, 18, 18, 8, 8, 3, 13, 9, 9, 9, 2, 6, 6, 21, 12, 6, 3, 3, 6, 12, 18, 7, 4, 9, 4, 6, 6, 2, 8, 7, 7, 5, 5, 10, 2, 6, 3, 9, 5, 6, 8, 9, 6, 4, 3, 2, 3, 9, 9, 20, 20, 14, 9, 4, 4, 6, 18, 6, 4, 9, 14, 18, 18, 9, 9, 9, 6, 6, 11, 12, 3, 8, 6, 4, 12, 12, 8, 3, 6, 8, 8, 3, 14, 10, 3, 6, 9, 8, 8, 6, 6, 6, 6, 9, 9, 8, 6, 4, 4, 3, 10, 6, 9, 6, 8, 6, 14, 8, 4, 9, 10, 13, 13, 6, 6, 14, 4, 6, 4, 9, 10, 5, 13, 19, 6, 2, 4, 5, 14, 6, 24, 14, 8, 6, 3, 5, 4, 6, 6, 6, 12, 21, 3, 9, 12, 9, 9, 22, 12, 9, 4, 22, 22, 4, 7, 4, 15, 12, 12, 16, 16, 16, 16, 3, 4, 8, 3, 2, 6, 9, 9, 6, 14, 3, 7, 5, 5, 9, 10, 9, 9, 20, 3, 20, 8, 20, 19, 20, 9, 4, 6, 6, 8, 6, 6, 4, 6, 8, 9, 9, 18, 20, 20, 6, 9, 6, 8, 12, 7, 6, 10, 3, 10, 12, 18, 16, 12, 14, 6, 6, 6, 10, 3, 8, 22, 8, 8, 9, 4, 6, 6, 3, 3, 9, 5, 15, 9, 3, 2, 9, 9, 9, 10, 16, 10, 13, 13, 9, 11, 11, 6, 3, 9, 14, 9, 6, 9, 20, 3, 3, 3, 9, 15, 3, 18, 3, 4, 5, 14, 9, 3, 18, 3, 12, 5, 12, 10, 10, 6, 9, 20, 6, 13, 15, 4, 14, 6, 3, 8, 18, 3, 13, 10, 9, 3, 3, 11, 10, 3, 3, 10, 21, 3, 6, 4, 4, 3, 3, 18, 3, 18, 6, 9, 10, 6, 18, 10, 10, 5, 7, 5, 7, 5, 18, 12, 4, 10, 6, 6, 2, 13, 3, 3, 6, 6, 6, 16, 16, 10, 10, 24, 20, 9, 9, 5, 9, 8, 8, 9, 12, 18, 18, 6, 3, 15, 14, 10, 9, 8, 8, 12, 4, 15, 10, 6, 5, 4, 6, 12, 6, 6, 23, 6, 12, 18, 12, 8, 4, 6, 3, 20, 20, 18, 12, 8, 14, 16, 9, 4, 4, 6, 6, 9, 7, 6, 10, 21, 10, 8, 9, 12, 12, 12, 12, 9, 9, 4, 4, 6, 4, 4, 4, 19, 8, 12, 3, 4, 10, 6, 22, 22, 3, 15, 9, 3, 15, 3, 6, 14, 10, 9, 10, 10, 4, 2, 6, 16, 4, 9, 9, 6, 9, 8, 16, 12, 9, 9, 9, 18, 12, 12, 6, 4, 6, 6, 3, 3, 22, 22, 24, 4, 18, 14, 9, 9, 20, 9, 14, 6, 24, 24, 7, 7, 19, 6, 6, 8, 15, 15, 20, 20, 4, 4, 3, 3, 20, 9, 19, 3, 20, 9, 5, 6, 20, 20, 12, 12, 8, 6, 4, 15, 6, 10, 12, 4, 6, 18, 9, 6, 3, 6, 19, 19, 2, 6, 18, 8, 6, 10, 6, 6, 15, 10, 4, 3, 9, 9, 9, 9, 5, 20, 6, 2, 6, 6, 9, 4, 6, 4, 22, 22, 9, 9, 18, 6, 8, 8, 12, 12, 8, 14, 12, 18, 18, 20, 12, 14, 6, 18, 14, 2, 12, 7, 12, 12, 22, 20, 4, 4, 6, 6, 24, 12, 4, 6, 3, 8, 12, 3, 7, 6, 7, 19, 7, 9, 7, 6, 5, 19, 6, 14, 9, 5, 5, 5, 7, 10, 9, 9, 7, 7, 8, 12, 12, 12, 8, 3, 4, 6, 15, 6, 9, 20, 9, 5, 14, 4, 6, 7, 6, 18, 6, 4, 6, 12, 3, 6, 6, 3, 9, 6, 6, 6, 3, 3, 6, 6, 9, 12, 8, 3, 12, 3, 9, 3, 3, 20, 20, 18, 12, 6, 18, 9, 6, 20, 20, 6, 6, 3, 6, 3, 7, 6, 6, 6, 13, 6, 15, 7, 6, 12, 9, 24, 24, 12, 6, 6, 12, 6, 14, 2, 3, 9, 12, 12, 9, 10, 9, 7, 5, 8, 18, 10, 10, 10, 10, 5, 2, 6, 7, 16, 8, 4, 8, 4, 9, 8, 4, 12, 12, 7, 3, 3, 10, 24, 15, 24, 9, 6, 6, 9, 9, 4, 20, 23, 18, 6, 6, 5, 19, 18, 18, 3, 9, 7, 7, 6, 10, 10, 16, 6, 6, 9, 8, 12, 9, 6, 22, 3, 3, 24, 6, 14, 10, 5, 6, 14, 14, 4, 12, 6, 6, 9, 9, 10, 8, 8, 4, 18, 19, 16, 16, 6, 5, 5, 6, 5, 7, 6, 9, 6, 20, 12, 12, 6, 8, 10, 9, 22, 22, 4, 15, 12, 13, 24, 24, 8, 2, 3, 6, 10, 3, 4, 8, 4, 16, 16, 16, 14, 14, 22, 22, 20, 20, 9, 16, 12, 6, 8, 6, 6, 6, 8, 12, 9, 6, 5, 8, 6, 6, 6, 18, 3, 2, 6, 9, 9, 15, 15, 6, 14, 5, 3, 2, 10, 3, 11, 8, 9, 2, 6, 3, 18, 10, 10, 9, 9, 3, 4, 14, 14, 6, 6, 18, 3, 3, 10, 4, 6, 9, 12, 6, 13, 6, 6, 3, 6, 3, 6, 19, 16, 18, 18, 3, 4, 6, 4, 8, 8, 12, 12, 6, 6, 6, 6, 2, 3, 12, 9, 15, 4, 12, 15, 19, 19, 10, 10, 18, 6, 10, 10, 10, 10, 18, 3, 18, 18, 3, 3, 3, 10, 17, 17, 11, 6, 8, 7, 14, 14, 2, 6, 4, 6, 18, 18, 10, 9, 6, 6, 6, 3, 9, 6, 18, 9, 9, 9, 3, 4, 10, 9, 9, 9, 6, 6, 9, 9, 6, 9, 3, 3, 6, 4, 6, 15, 3, 10, 3, 6, 18, 6, 18, 18, 6, 12, 22, 6, 6, 18, 9, 9, 12, 4, 3, 8, 15, 14, 14, 14, 4, 20, 12, 12, 8, 8, 15, 15, 12, 12, 9, 21, 4, 9, 15, 15, 8, 6, 4, 3, 12, 12, 6, 10, 6, 2, 3, 3, 6, 6, 6, 6, 20, 8, 22};

localparam logic [2912:0][31:0] rectangle1_weights = {-128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128, -128};

localparam logic [2912:0][31:0] rectangle2_xs = {6, 10, 3, 8, 5, 6, 5, 11, 4, 6, 10, 1, 8, 9, 5, 5, 16, 9, 12, 4, 20, 8, 11, 7, 5, 8, 5, 9, 11, 6, 9, 5, 18, 4, 8, 5, 2, 10, 2, 2, 20, 11, 20, 2, 12, 0, 12, 10, 12, 1, 17, 0, 6, 10, 8, 4, 2, 19, 3, 8, 1, 14, 3, 6, 8, 15, 1, 4, 2, 3, 1, 5, 3, 14, 1, 15, 5, 10, 9, 11, 9, 12, 10, 9, 6, 8, 4, 11, 8, 11, 9, 11, 11, 9, 1, 10, 6, 7, 0, 6, 1, 6, 5, 20, 2, 12, 4, 14, 8, 17, 0, 14, 8, 8, 0, 12, 9, 2, 2, 3, 5, 14, 4, 4, 6, 3, 3, 10, 8, 3, 12, 8, 5, 16, 4, 19, 8, 6, 10, 9, 0, 4, 9, 18, 3, 18, 3, 16, 2, 9, 2, 14, 5, 18, 3, 8, 7, 8, 10, 14, 7, 13, 12, 13, 1, 13, 8, 8, 8, 7, 0, 1, 9, 12, 9, 7, 0, 13, 12, 14, 9, 14, 9, 18, 6, 13, 3, 13, 0, 6, 6, 10, 10, 4, 5, 9, 20, 2, 5, 2, 5, 2, 13, 0, 1, 2, 13, 0, 11, 10, 11, 6, 18, 3, 18, 1, 13, 0, 13, 9, 13, 10, 13, 2, 12, 5, 14, 4, 7, 5, 12, 9, 3, 0, 12, 4, 13, 10, 10, 8, 10, 0, 12, 4, 8, 11, 9, 10, 20, 1, 14, 3, 15, 11, 17, 3, 7, 4, 10, 8, 15, 3, 12, 6, 14, 1, 13, 10, 12, 9, 6, 9, 7, 8, 7, 0, 15, 0, 15, 8, 15, 0, 8, 0, 9, 8, 9, 12, 12, 6, 16, 2, 0, 4, 9, 0, 18, 0, 8, 10, 13, 9, 14, 8, 15, 8, 9, 7, 14, 2, 5, 11, 13, 10, 9, 8, 12, 1, 15, 1, 10, 3, 12, 8, 6, 10, 5, 4, 11, 7, 9, 2, 3, 10, 16, 9, 21, 0, 18, 3, 18, 0, 5, 6, 12, 10, 15, 3, 15, 5, 11, 8, 15, 9, 13, 9, 18, 1, 14, 1, 12, 1, 14, 0, 17, 5, 18, 3, 15, 0, 4, 2, 14, 6, 20, 1, 16, 7, 12, 4, 12, 8, 15, 7, 6, 1, 6, 0, 13, 9, 12, 8, 16, 0, 14, 7, 5, 4, 16, 6, 12, 11, 11, 12, 6, 10, 8, 14, 5, 11, 3, 3, 3, 20, 5, 13, 6, 12, 8, 9, 10, 13, 9, 14, 8, 20, 6, 18, 7, 18, 0, 9, 0, 17, 1, 14, 8, 9, 9, 14, 8, 6, 1, 10, 5, 5, 0, 8, 10, 6, 4, 12, 12, 12, 3, 2, 6, 14, 0, 19, 0, 12, 0, 13, 3, 6, 0, 15, 9, 12, 1, 15, 7, 19, 6, 8, 5, 14, 2, 18, 2, 17, 12, 14, 10, 14, 6, 6, 11, 12, 10, 16, 6, 9, 5, 10, 8, 6, 10, 8, 1, 9, 3, 2, 10, 8, 10, 0, 14, 9, 14, 1, 15, 0, 19, 2, 3, 9, 18, 0, 12, 2, 14, 5, 18, 5, 22, 8, 11, 7, 22, 12, 15, 0, 13, 9, 14, 6, 14, 6, 3, 3, 12, 12, 13, 8, 20, 3, 20, 0, 10, 8, 13, 9, 13, 0, 6, 3, 8, 2, 15, 3, 19, 3, 19, 3, 4, 6, 15, 0, 17, 5, 8, 6, 5, 10, 10, 0, 15, 0, 14, 11, 14, 8, 15, 3, 11, 6, 12, 0, 3, 3, 12, 1, 17, 2, 7, 8, 3, 10, 5, 11, 3, 18, 3, 9, 3, 13, 8, 13, 4, 13, 8, 7, 6, 16, 6, 11, 0, 13, 5, 10, 10, 14, 6, 12, 7, 8, 5, 3, 5, 5, 8, 3, 1, 5, 1, 1, 3, 6, 7, 14, 1, 13, 12, 13, 9, 15, 5, 15, 6, 15, 0, 5, 7, 17, 10, 15, 0, 14, 8, 13, 6, 13, 8, 17, 4, 12, 11, 11, 9, 8, 1, 9, 9, 18, 8, 2, 0, 18, 2, 2, 12, 13, 1, 11, 3, 12, 2, 18, 3, 22, 2, 1, 0, 19, 3, 20, 0, 13, 0, 10, 8, 4, 2, 14, 3, 17, 6, 10, 4, 2, 10, 5, 12, 0, 15, 5, 8, 1, 19, 8, 20, 9, 15, 2, 16, 2, 20, 3, 15, 0, 16, 2, 10, 1, 14, 3, 3, 10, 3, 2, 12, 10, 12, 11, 4, 0, 9, 8, 13, 5, 12, 1, 19, 0, 20, 0, 18, 9, 11, 0, 1, 1, 13, 4, 12, 4, 15, 1, 13, 5, 16, 5, 10, 7, 12, 0, 17, 0, 15, 0, 13, 8, 12, 2, 12, 1, 15, 0, 6, 10, 12, 8, 12, 8, 13, 1, 15, 6, 18, 11, 12, 0, 11, 11, 12, 8, 9, 10, 4, 11, 5, 8, 15, 12, 12, 7, 11, 3, 14, 8, 9, 1, 11, 9, 12, 1, 6, 1, 8, 2, 11, 7, 14, 9, 14, 7, 4, 9, 7, 11, 2, 8, 3, 11, 0, 10, 2, 20, 2, 12, 0, 14, 0, 12, 8, 4, 10, 14, 2, 14, 2, 5, 9, 12, 6, 12, 0, 18, 5, 10, 2, 13, 6, 11, 7, 18, 11, 10, 0, 15, 4, 13, 7, 14, 7, 12, 6, 16, 0, 16, 5, 5, 5, 9, 9, 13, 5, 19, 3, 5, 0, 2, 5, 1, 10, 8, 11, 12, 4, 12, 3, 5, 4, 6, 10, 0, 0, 3, 2, 7, 5, 10, 9, 18, 9, 12, 11, 13, 9, 4, 2, 13, 9, 9, 1, 8, 3, 5, 8, 9, 0, 6, 4, 13, 5, 12, 11, 14, 5, 12, 0, 20, 9, 12, 10, 14, 7, 12, 2, 18, 1, 6, 12, 14, 6, 11, 1, 9, 7, 17, 2, 7, 1, 8, 11, 3, 20, 8, 20, 0, 8, 5, 4, 8, 6, 0, 20, 10, 12, 0, 6, 0, 20, 2, 18, 3, 13, 8, 5, 9, 6, 9, 10, 1, 11, 7, 14, 5, 13, 0, 12, 1, 2, 2, 20, 1, 14, 0, 15, 1, 9, 0, 16, 12, 7, 11, 12, 10, 15, 3, 16, 3, 16, 12, 10, 7, 11, 11, 12, 11, 3, 2, 12, 5, 14, 0, 10, 8, 5, 11, 11, 9, 5, 10, 10, 7, 12, 0, 12, 2, 12, 1, 12, 0, 5, 6, 14, 5, 9, 8, 11, 6, 17, 8, 8, 4, 12, 9, 16, 1, 11, 3, 7, 12, 12, 3, 12, 3, 13, 5, 11, 9, 17, 2, 12, 0, 12, 5, 12, 9, 2, 5, 4, 2, 7, 0, 2, 6, 6, 11, 15, 8, 3, 2, 19, 1, 14, 4, 14, 8, 14, 4, 8, 3, 20, 2, 8, 9, 16, 12, 11, 12, 12, 10, 14, 5, 18, 6, 13, 1, 15, 9, 10, 3, 16, 9, 15, 0, 13, 2, 5, 1, 5, 1, 16, 9, 16, 6, 18, 1, 9, 0, 14, 3, 16, 3, 11, 11, 15, 8, 17, 3, 3, 0, 2, 0, 13, 5, 12, 5, 18, 0, 13, 5, 9, 12, 6, 9, 13, 8, 6, 2, 20, 2, 14, 8, 8, 12, 9, 11, 4, 10, 8, 7, 12, 0, 18, 0, 16, 1, 12, 9, 12, 8, 12, 4, 15, 3, 15, 4, 15, 0, 15, 0, 14, 3, 7, 10, 8, 12, 7, 0, 16, 7, 10, 11, 12, 3, 16, 0, 0, 0, 10, 10, 4, 8, 9, 9, 6, 11, 8, 4, 8, 7, 1, 15, 7, 13, 9, 3, 0, 10, 6, 15, 0, 20, 2, 13, 0, 2, 1, 18, 0, 17, 0, 0, 2, 12, 9, 17, 5, 15, 0, 15, 0, 5, 0, 13, 8, 13, 8, 13, 10, 12, 11, 13, 7, 14, 12, 12, 1, 20, 0, 14, 0, 13, 0, 6, 0, 14, 1, 13, 4, 17, 5, 16, 3, 14, 10, 11, 0, 4, 5, 19, 0, 8, 3, 17, 4, 16, 3, 18, 1, 17, 0, 15, 8, 22, 1, 20, 2, 3, 6, 7, 11, 4, 9, 4, 3, 18, 2, 13, 7, 13, 10, 12, 0, 11, 2, 13, 5, 9, 5, 3, 6, 12, 8, 9, 1, 19, 1, 9, 6, 12, 10, 14, 4, 8, 6, 19, 0, 17, 1, 18, 0, 3, 2, 14, 5, 10, 11, 7, 12, 5, 10, 11, 9, 14, 8, 12, 7, 2, 1, 8, 7, 6, 17, 4, 2, 6, 9, 7, 10, 8, 18, 3, 18, 4, 5, 11, 15, 7, 12, 12, 12, 2, 14, 10, 14, 3, 14, 1, 3, 1, 18, 0, 5, 6, 14, 4, 17, 8, 8, 5, 3, 0, 12, 0, 9, 2, 0, 10, 10, 8, 13, 11, 2, 1, 13, 12, 10, 7, 14, 10, 11, 10, 20, 1, 17, 9, 12, 12, 14, 5, 16, 4, 10, 1, 15, 12, 12, 8, 19, 0, 14, 6, 13, 9, 13, 8, 7, 4, 17, 3, 14, 2, 3, 4, 19, 10, 19, 1, 15, 5, 10, 4, 0, 8, 14, 0, 6, 1, 18, 4, 6, 1, 1, 2, 18, 0, 12, 7, 9, 7, 12, 7, 12, 10, 15, 3, 4, 6, 8, 12, 11, 2, 8, 0, 0, 2, 12, 10, 7, 9, 17, 0, 19, 1, 12, 3, 12, 12, 12, 10, 14, 10, 13, 7, 7, 9, 0, 11, 3, 15, 2, 13, 4, 20, 8, 12, 2, 3, 3, 13, 5, 17, 2, 12, 10, 12, 10, 12, 12, 12, 0, 9, 7, 14, 8, 13, 1, 9, 2, 15, 0, 9, 2, 15, 4, 17, 0, 15, 0, 15, 3, 20, 8, 13, 0, 0, 5, 11, 4, 10, 8, 11, 4, 14, 2, 4, 8, 1, 9, 13, 10, 4, 6, 14, 9, 9, 9, 9, 11, 9, 12, 14, 8, 18, 3, 18, 0, 13, 10, 11, 8, 16, 5, 7, 9, 13, 3, 20, 7, 15, 0, 19, 1, 12, 1, 3, 8, 5, 9, 11, 4, 6, 5, 17, 11, 1, 10, 10, 11, 11, 9, 15, 0, 2, 0, 9, 9, 18, 0, 12, 3, 2, 5, 12, 10, 5, 9, 7, 9, 4, 0, 11, 11, 6, 11, 12, 5, 14, 5, 14, 0, 16, 4, 8, 0, 13, 0, 12, 6, 10, 1, 0, 6, 9, 1, 10, 7, 9, 10, 3, 7, 3, 10, 3, 10, 4, 5, 8, 9, 3, 2, 9, 11, 11, 16, 7, 16, 6, 19, 3, 14, 0, 9, 6, 14, 4, 7, 9, 14, 12, 14, 5, 4, 11, 3, 4, 16, 4, 13, 10, 15, 12, 12, 3, 12, 8, 6, 0, 4, 0, 15, 0, 6, 3, 13, 6, 6, 10, 10, 7, 17, 2, 11, 1, 15, 1, 10, 11, 7, 10, 15, 3, 15, 7, 12, 9, 15, 5, 8, 7, 12, 9, 7, 10, 13, 9, 9, 0, 14, 0, 12, 1, 7, 11, 16, 2, 8, 0, 5, 2, 14, 3, 9, 4, 12, 9, 13, 0, 14, 2, 11, 7, 13, 7, 17, 4, 13, 10, 18, 12, 17, 5, 16, 4, 18, 4, 15, 0, 20, 2, 16, 9, 12, 0, 5, 0, 12, 5, 10, 8, 6, 3, 16, 6, 8, 6, 10, 11, 14, 0, 16, 3, 6, 4, 17, 2, 2, 4, 18, 8, 6, 6, 14, 8, 15, 6, 14, 4, 7, 8, 13, 9, 8, 0, 17, 0, 21, 0, 12, 1, 5, 1, 6, 5, 14, 1, 11, 0, 13, 1, 0, 1, 14, 7, 12, 8, 13, 11, 9, 7, 6, 10, 10, 6, 15, 8, 11, 8, 1, 0, 15, 7, 20, 2, 14, 2, 12, 1, 7, 8, 12, 2, 14, 3, 17, 5, 13, 9, 13, 12, 12, 11, 20, 1, 7, 6, 9, 1, 19, 4, 3, 1, 9, 4, 6, 4, 15, 9, 12, 6, 15, 3, 14, 1, 14, 0, 15, 3, 9, 1, 13, 1, 6, 8, 0, 0, 14, 1, 14, 8, 10, 11, 10, 9, 14, 8, 11, 3, 13, 0, 12, 11, 10, 8, 11, 10, 12, 10, 4, 0, 11, 1, 11, 6, 14, 7, 12, 12, 11, 1, 9, 0, 1, 1, 9, 9, 11, 11, 18, 4, 15, 1, 14, 3, 15, 7, 14, 12, 7, 0, 19, 1, 16, 6, 17, 5, 0, 7, 1, 1, 6, 1, 15, 3, 4, 0, 6, 7, 12, 6, 9, 4, 20, 2, 13, 12, 13, 1, 13, 2, 13, 2, 3, 7, 17, 5, 16, 0, 15, 0, 9, 4, 12, 10, 13, 9, 14, 8, 10, 0, 13, 9, 14, 0, 1, 10, 16, 10, 12, 8, 13, 2, 11, 7, 13, 0, 12, 8, 12, 6, 14, 0, 14, 0, 4, 1, 4, 8, 3, 11, 0, 6, 2, 18, 0, 11, 9, 7, 3, 18, 7, 18, 3, 9, 2, 10, 5, 11, 10, 12, 4, 6, 9, 9, 11, 10, 2, 21, 0, 5, 12, 1, 10, 6, 9, 2, 5, 12, 9, 18, 2, 16, 1, 12, 4, 10, 5, 14, 7, 7, 2, 5, 7, 0, 2, 20, 5, 5, 0, 13, 0, 4, 2, 12, 12, 6, 0, 10, 7, 11, 7, 21, 3, 21, 7, 9, 0, 15, 1, 13, 7, 13, 10, 13, 10, 13, 10, 5, 0, 11, 2, 15, 1, 10, 0, 6, 0, 13, 2, 13, 8, 13, 9, 12, 3, 16, 6, 10, 7, 12, 7, 10, 3, 16, 4, 0, 11, 10, 12, 17, 5, 16, 5, 3, 4, 4, 3, 16, 6, 14, 7, 4, 0, 10, 6, 0, 0, 3, 9, 12, 6, 8, 2, 12, 5, 14, 10, 12, 7, 17, 9, 13, 0, 12, 9, 10, 9, 0, 8, 9, 9, 15, 10, 15, 6, 19, 2, 12, 10, 14, 5, 11, 3, 10, 5, 20, 7, 4, 8, 6, 19, 3, 20, 2, 5, 10, 11, 0, 7, 1, 11, 0, 17, 12, 17, 7, 13, 0, 8, 6, 7, 0, 13, 3, 12, 2, 9, 6, 14, 5, 12, 6, 17, 4, 14, 0, 13, 2, 6, 0, 21, 1, 15, 11, 13, 7, 14, 3, 22, 7, 12, 11, 15, 8, 13, 8, 9, 8, 12, 3, 19, 0, 22, 0, 7, 11, 10, 0, 14, 2, 13, 8, 15, 7, 11, 11, 15, 1, 16, 5, 12, 4, 6, 9, 15, 6, 12, 7, 6, 10, 12, 3, 4, 2, 13, 9, 1, 0, 0, 3, 3, 5, 16, 5, 10, 6, 12, 2, 12, 10, 13, 6, 9, 2, 14, 3, 10, 2, 17, 2, 0, 7, 17, 5, 11, 8, 11, 5, 15, 4, 15, 6, 12, 9, 12, 4, 4, 5, 14, 9, 12, 10, 12, 2, 12, 9, 12, 8, 7, 1, 13, 2, 15, 0, 15, 6, 8, 1, 6, 10, 12, 3, 18, 1, 18, 11, 18, 6, 18, 6, 16, 12, 9, 6, 11, 6, 16, 4, 18, 8, 18, 3, 15, 6, 18, 0, 13, 7, 4, 0, 15, 3, 9, 8, 5, 3, 5, 10, 4, 2, 8, 18, 3, 4, 6, 13, 4, 12, 8, 13, 8, 3, 0, 14, 0, 14, 0, 6, 0, 14, 8, 15, 8, 10, 7, 7, 12, 11, 7, 21, 0, 15, 0, 18, 7, 16, 0, 18, 2, 14, 1, 9, 5, 5, 11, 12, 9, 12, 10, 12, 9, 13, 3, 12, 9, 13, 9, 11, 7, 5, 8, 4, 0, 0, 0, 11, 3, 12, 10, 12, 7, 9, 10, 11, 9, 19, 1, 15, 5, 6, 10, 12, 10, 14, 3, 7, 7, 14, 7, 18, 9, 13, 6, 10, 0, 3, 4, 16, 8, 16, 7, 15, 3, 18, 0, 13, 2, 17, 1, 8, 0, 15, 1, 20, 3, 9, 9, 7, 10, 11, 4, 10, 3, 15, 0, 6, 9, 12, 10, 16, 10, 6, 0, 17, 5, 14, 1, 7, 10, 14, 3, 9, 3, 6, 1, 16, 0, 12, 8, 10, 0, 21, 2, 20, 2, 8, 8, 11, 9, 7, 12, 11, 8, 11, 4, 12, 0, 12, 4, 12, 11, 15, 8, 13, 10, 12, 9, 17, 6, 10, 2, 2, 7, 3, 2, 15, 8, 10, 7, 18, 3, 20, 2, 17, 5, 16, 4, 11, 12, 12, 3, 13, 0, 8, 9, 19, 9, 6, 10, 5, 12, 3, 15, 4, 11, 9, 5, 4, 11, 10, 16, 3, 13, 8, 8, 10, 5, 2, 2, 11, 9, 9, 5, 2, 6, 6, 20, 2, 10, 10, 3, 5, 17, 0, 9, 10, 11, 0, 6, 4, 9, 5, 6, 7, 11, 12, 18, 0, 0, 0, 6, 0, 20, 4, 21, 1, 3, 0, 18, 7, 17, 2, 19, 0, 15, 0, 14, 0, 5, 0, 12, 5, 4, 3, 4, 10, 16, 7, 17, 3, 12, 5, 14, 6, 15, 0, 12, 0, 12, 9, 6, 0, 2, 7, 12, 6, 8, 4, 12, 10, 18, 3, 6, 5, 12, 0, 12, 11, 11, 1, 14, 1, 7, 0, 12, 12, 12, 10, 9, 1, 0, 6, 12, 5, 4, 4, 8, 1, 10, 1, 12, 1, 5, 0, 9, 1, 8, 8, 5, 9, 6, 2, 12, 10, 14, 8, 9, 12, 5, 4, 14, 9, 14, 8, 11, 5, 5, 9, 11, 2, 18, 3, 12, 5, 20, 0, 18, 1, 15, 5, 6, 2, 14, 10, 13, 3, 13, 3, 16, 0, 0, 12, 21, 0, 15, 1, 15, 0, 3, 0, 15, 0, 12, 3, 17, 0, 12};

localparam logic [2912:0][31:0] rectangle2_ys = {7, 4, 12, 20, 5, 13, 11, 19, 3, 8, 4, 12, 2, 14, 11, 3, 11, 5, 8, 5, 0, 6, 6, 20, 13, 3, 11, 13, 5, 12, 21, 8, 1, 1, 8, 6, 16, 1, 13, 1, 2, 5, 4, 3, 1, 7, 1, 1, 5, 11, 13, 7, 7, 5, 1, 12, 17, 3, 3, 1, 11, 14, 12, 8, 13, 17, 18, 10, 1, 1, 5, 12, 17, 17, 17, 6, 5, 0, 3, 6, 0, 6, 6, 8, 3, 0, 11, 6, 20, 6, 13, 6, 6, 18, 23, 12, 12, 8, 16, 19, 2, 17, 4, 4, 4, 16, 12, 0, 10, 8, 8, 0, 0, 16, 18, 8, 19, 11, 9, 0, 6, 5, 5, 15, 17, 19, 0, 6, 1, 3, 8, 11, 12, 16, 16, 5, 2, 10, 5, 20, 12, 4, 5, 1, 1, 0, 0, 7, 12, 13, 17, 14, 6, 8, 8, 15, 14, 14, 10, 15, 0, 0, 3, 0, 1, 0, 0, 20, 3, 5, 11, 11, 11, 11, 11, 12, 13, 4, 0, 0, 0, 1, 1, 6, 16, 16, 19, 4, 18, 2, 11, 5, 13, 4, 3, 19, 0, 1, 23, 0, 12, 1, 5, 2, 3, 11, 12, 12, 7, 1, 7, 10, 6, 16, 8, 5, 0, 4, 0, 0, 6, 7, 19, 18, 18, 20, 15, 6, 8, 14, 9, 6, 7, 11, 16, 6, 0, 0, 7, 20, 14, 2, 1, 3, 0, 21, 7, 7, 8, 15, 17, 3, 11, 1, 2, 14, 8, 2, 8, 17, 11, 1, 16, 16, 14, 14, 1, 0, 2, 2, 20, 6, 7, 10, 8, 4, 2, 6, 3, 0, 10, 10, 16, 16, 10, 0, 7, 6, 9, 0, 0, 0, 12, 11, 11, 14, 15, 15, 7, 7, 0, 0, 3, 3, 4, 10, 19, 17, 13, 18, 19, 0, 4, 4, 3, 1, 19, 3, 5, 2, 19, 22, 14, 2, 7, 6, 12, 14, 13, 14, 7, 4, 14, 6, 6, 9, 6, 6, 5, 20, 5, 5, 11, 2, 0, 0, 14, 8, 14, 5, 8, 13, 14, 12, 1, 1, 12, 22, 16, 13, 6, 0, 7, 4, 0, 0, 12, 12, 14, 14, 15, 14, 17, 0, 1, 1, 17, 9, 7, 4, 6, 10, 17, 1, 11, 6, 17, 17, 7, 15, 8, 14, 16, 4, 19, 13, 3, 6, 11, 7, 6, 8, 15, 1, 8, 5, 2, 11, 11, 6, 1, 4, 18, 4, 16, 7, 7, 2, 20, 14, 2, 0, 0, 17, 8, 3, 12, 7, 8, 7, 7, 6, 23, 17, 17, 11, 11, 9, 17, 0, 0, 18, 18, 12, 6, 6, 1, 0, 15, 11, 16, 2, 20, 0, 13, 11, 7, 8, 9, 0, 0, 1, 18, 15, 15, 17, 18, 0, 4, 5, 14, 0, 0, 7, 7, 5, 15, 0, 7, 2, 2, 2, 6, 5, 6, 0, 3, 7, 7, 13, 6, 17, 0, 2, 8, 8, 8, 3, 6, 0, 12, 21, 8, 5, 7, 12, 7, 19, 20, 14, 20, 20, 11, 11, 3, 18, 17, 20, 6, 6, 0, 0, 0, 0, 3, 11, 0, 0, 8, 12, 0, 6, 2, 3, 7, 6, 1, 10, 3, 5, 4, 1, 13, 5, 1, 2, 10, 9, 10, 10, 17, 7, 1, 1, 5, 12, 17, 15, 16, 13, 11, 6, 5, 5, 1, 1, 15, 11, 4, 4, 0, 0, 19, 11, 8, 8, 12, 12, 2, 2, 6, 7, 6, 6, 3, 0, 13, 7, 6, 3, 15, 14, 12, 2, 16, 16, 3, 0, 10, 5, 16, 19, 6, 0, 2, 12, 0, 11, 20, 11, 14, 11, 11, 8, 17, 0, 0, 7, 1, 20, 7, 17, 2, 3, 6, 8, 12, 10, 5, 20, 0, 2, 11, 3, 17, 18, 15, 14, 8, 8, 2, 19, 20, 3, 6, 0, 0, 10, 11, 5, 8, 5, 6, 22, 10, 4, 8, 9, 10, 6, 5, 4, 4, 10, 10, 2, 2, 4, 4, 4, 4, 20, 20, 2, 2, 5, 11, 9, 5, 14, 14, 11, 9, 6, 21, 5, 5, 4, 7, 13, 8, 2, 19, 10, 2, 0, 3, 2, 7, 0, 3, 19, 14, 14, 5, 6, 6, 5, 5, 12, 12, 3, 3, 1, 11, 14, 11, 11, 20, 4, 3, 11, 0, 0, 11, 23, 10, 1, 0, 3, 17, 16, 12, 12, 7, 6, 8, 11, 7, 6, 9, 0, 5, 5, 5, 4, 17, 17, 13, 17, 16, 9, 0, 12, 9, 9, 6, 6, 5, 6, 13, 5, 3, 16, 19, 13, 10, 9, 16, 14, 10, 0, 11, 2, 4, 0, 19, 8, 10, 17, 18, 18, 11, 11, 3, 5, 0, 17, 17, 17, 18, 8, 6, 12, 12, 5, 9, 9, 11, 13, 8, 8, 11, 11, 6, 0, 0, 3, 10, 7, 13, 4, 2, 5, 0, 4, 10, 10, 11, 10, 12, 21, 20, 17, 19, 18, 6, 16, 18, 6, 4, 21, 7, 2, 10, 11, 9, 10, 11, 0, 8, 0, 3, 20, 1, 0, 18, 7, 3, 2, 2, 1, 18, 15, 16, 5, 13, 3, 14, 12, 16, 8, 12, 20, 7, 2, 6, 7, 0, 11, 12, 21, 3, 9, 11, 7, 8, 16, 14, 11, 13, 0, 10, 4, 0, 6, 6, 11, 11, 16, 7, 16, 14, 11, 6, 18, 0, 5, 0, 1, 1, 17, 5, 17, 5, 9, 4, 7, 7, 4, 12, 3, 6, 9, 5, 4, 6, 2, 19, 19, 5, 8, 13, 12, 6, 11, 7, 5, 9, 14, 14, 11, 12, 0, 0, 1, 14, 20, 11, 11, 14, 16, 11, 5, 16, 15, 8, 16, 0, 5, 5, 6, 10, 10, 18, 10, 0, 4, 12, 6, 12, 16, 11, 11, 12, 4, 4, 9, 5, 9, 0, 16, 16, 7, 9, 1, 6, 18, 8, 19, 8, 8, 17, 11, 2, 12, 4, 1, 3, 6, 11, 8, 18, 16, 3, 3, 0, 0, 11, 11, 12, 20, 8, 0, 10, 11, 12, 0, 0, 5, 14, 14, 1, 0, 3, 3, 10, 10, 6, 14, 17, 1, 13, 16, 17, 3, 6, 6, 1, 1, 18, 18, 1, 3, 0, 3, 5, 0, 7, 7, 3, 3, 8, 8, 13, 5, 1, 1, 15, 2, 6, 15, 12, 12, 2, 7, 11, 9, 5, 8, 19, 19, 19, 18, 19, 1, 2, 16, 16, 22, 13, 10, 8, 10, 10, 15, 7, 16, 19, 15, 9, 9, 7, 4, 8, 7, 15, 8, 19, 19, 1, 12, 5, 4, 16, 16, 0, 8, 4, 2, 1, 15, 11, 9, 5, 4, 3, 14, 11, 0, 7, 1, 11, 7, 23, 16, 0, 11, 17, 17, 5, 5, 8, 8, 2, 2, 0, 4, 18, 0, 15, 21, 5, 5, 6, 5, 16, 5, 8, 6, 13, 10, 15, 3, 8, 6, 6, 13, 15, 15, 18, 18, 17, 17, 1, 2, 2, 15, 2, 2, 5, 2, 0, 13, 2, 11, 6, 8, 11, 8, 0, 0, 6, 20, 19, 6, 8, 3, 19, 5, 6, 16, 5, 5, 4, 13, 1, 12, 7, 5, 11, 11, 5, 2, 0, 0, 0, 0, 2, 13, 7, 8, 15, 10, 17, 9, 4, 13, 8, 18, 18, 20, 8, 8, 5, 5, 6, 0, 8, 8, 14, 11, 14, 14, 17, 17, 0, 0, 8, 17, 6, 22, 9, 0, 1, 18, 7, 10, 2, 12, 5, 5, 3, 13, 19, 9, 7, 1, 14, 21, 11, 6, 6, 4, 10, 17, 4, 0, 0, 0, 7, 1, 10, 8, 5, 0, 0, 2, 2, 0, 1, 3, 11, 10, 3, 6, 10, 8, 2, 6, 0, 0, 0, 19, 18, 16, 17, 16, 16, 8, 7, 8, 0, 8, 5, 6, 7, 8, 8, 10, 5, 12, 9, 14, 9, 18, 6, 6, 16, 17, 12, 9, 7, 10, 10, 10, 12, 17, 16, 16, 0, 1, 18, 18, 9, 0, 0, 2, 1, 8, 8, 10, 10, 7, 12, 15, 2, 1, 1, 1, 1, 11, 11, 13, 14, 13, 18, 22, 12, 7, 7, 7, 14, 14, 7, 13, 7, 12, 7, 0, 12, 13, 13, 17, 19, 3, 5, 0, 16, 18, 15, 10, 9, 16, 9, 15, 8, 4, 9, 6, 7, 12, 12, 6, 6, 5, 5, 5, 5, 3, 3, 11, 11, 8, 6, 19, 4, 1, 11, 12, 12, 0, 12, 21, 4, 2, 10, 7, 0, 15, 3, 7, 20, 12, 5, 11, 4, 0, 4, 4, 19, 9, 13, 13, 11, 6, 0, 9, 18, 7, 18, 14, 14, 14, 8, 9, 7, 7, 14, 18, 18, 18, 1, 21, 20, 1, 18, 17, 16, 18, 10, 18, 7, 7, 13, 6, 0, 7, 2, 18, 2, 7, 1, 0, 3, 15, 10, 3, 0, 0, 0, 4, 17, 20, 3, 3, 6, 6, 14, 19, 2, 1, 0, 10, 16, 16, 12, 16, 6, 6, 9, 9, 10, 8, 10, 10, 1, 5, 10, 14, 4, 2, 4, 4, 8, 8, 17, 16, 18, 2, 2, 2, 3, 2, 8, 3, 22, 11, 11, 11, 8, 8, 15, 15, 14, 13, 15, 4, 15, 15, 11, 8, 6, 9, 4, 7, 11, 12, 18, 2, 13, 12, 5, 7, 5, 19, 5, 5, 1, 4, 4, 4, 4, 4, 1, 1, 5, 4, 5, 5, 7, 0, 11, 6, 3, 18, 8, 4, 11, 4, 13, 1, 4, 7, 19, 9, 6, 5, 3, 2, 6, 3, 3, 3, 1, 2, 3, 16, 8, 0, 0, 11, 6, 9, 17, 19, 8, 17, 18, 19, 2, 5, 6, 19, 19, 18, 18, 13, 14, 18, 13, 17, 2, 9, 5, 7, 8, 9, 9, 9, 8, 12, 10, 10, 0, 3, 1, 23, 10, 0, 0, 2, 13, 21, 1, 7, 0, 1, 1, 5, 6, 5, 5, 13, 7, 9, 9, 4, 6, 21, 21, 5, 10, 0, 2, 0, 15, 13, 0, 7, 13, 22, 3, 11, 7, 7, 3, 1, 1, 18, 15, 10, 9, 11, 7, 2, 2, 4, 8, 9, 4, 11, 7, 0, 0, 1, 2, 7, 3, 14, 14, 19, 0, 4, 2, 2, 12, 15, 10, 18, 4, 0, 6, 13, 13, 13, 7, 6, 18, 20, 18, 13, 13, 9, 20, 18, 2, 2, 15, 11, 18, 19, 12, 12, 1, 15, 7, 12, 0, 3, 0, 0, 11, 14, 21, 0, 1, 6, 6, 0, 0, 18, 0, 0, 1, 1, 16, 3, 5, 10, 15, 10, 8, 2, 16, 6, 16, 22, 10, 6, 2, 16, 20, 0, 6, 10, 15, 7, 6, 6, 0, 0, 19, 17, 4, 4, 16, 16, 16, 18, 0, 3, 17, 0, 12, 12, 9, 3, 7, 4, 3, 2, 5, 0, 19, 19, 15, 22, 15, 15, 6, 3, 3, 8, 4, 2, 2, 2, 7, 3, 6, 1, 8, 0, 18, 20, 19, 18, 8, 15, 18, 18, 6, 7, 6, 9, 5, 7, 4, 10, 5, 8, 0, 12, 14, 10, 17, 6, 6, 13, 10, 10, 9, 3, 0, 12, 0, 0, 2, 2, 0, 0, 8, 8, 1, 1, 0, 10, 11, 11, 10, 16, 10, 7, 8, 0, 11, 6, 0, 15, 14, 1, 0, 3, 2, 6, 20, 20, 19, 0, 3, 12, 4, 3, 8, 15, 13, 6, 9, 0, 9, 9, 5, 4, 7, 0, 0, 0, 4, 3, 13, 13, 2, 13, 8, 9, 8, 14, 14, 12, 12, 17, 17, 8, 10, 10, 9, 12, 12, 12, 12, 12, 10, 15, 10, 1, 7, 5, 12, 16, 0, 10, 4, 20, 11, 18, 0, 0, 2, 2, 7, 1, 16, 15, 8, 8, 6, 19, 18, 5, 6, 6, 0, 0, 5, 5, 1, 13, 1, 18, 17, 20, 16, 1, 8, 0, 6, 5, 1, 5, 1, 11, 11, 18, 18, 15, 11, 11, 9, 15, 17, 17, 16, 16, 5, 18, 21, 21, 20, 19, 2, 4, 9, 19, 2, 10, 10, 8, 5, 5, 4, 4, 7, 6, 4, 0, 1, 1, 17, 3, 3, 2, 2, 7, 22, 16, 3, 10, 19, 0, 5, 8, 1, 6, 3, 13, 14, 7, 7, 10, 8, 19, 14, 6, 0, 0, 1, 14, 10, 12, 1, 1, 7, 10, 7, 8, 0, 0, 5, 5, 0, 0, 3, 3, 4, 18, 19, 19, 18, 18, 17, 10, 19, 12, 10, 10, 2, 6, 14, 14, 1, 21, 1, 16, 1, 0, 1, 1, 9, 16, 4, 4, 4, 4, 0, 16, 7, 11, 5, 6, 1, 1, 9, 4, 16, 0, 5, 3, 14, 16, 11, 9, 2, 6, 8, 1, 1, 16, 19, 19, 4, 20, 12, 12, 12, 12, 8, 8, 14, 14, 7, 7, 3, 1, 11, 6, 18, 23, 15, 15, 15, 19, 14, 12, 3, 1, 1, 2, 2, 14, 3, 6, 6, 0, 0, 6, 1, 7, 7, 20, 6, 2, 4, 4, 2, 2, 2, 2, 15, 18, 12, 1, 8, 6, 12, 14, 14, 18, 6, 3, 6, 5, 9, 16, 8, 8, 6, 5, 10, 11, 2, 0, 4, 7, 2, 4, 0, 17, 17, 0, 3, 7, 9, 14, 14, 21, 21, 4, 8, 4, 17, 16, 11, 18, 5, 8, 8, 8, 8, 8, 6, 8, 11, 11, 3, 10, 19, 18, 11, 4, 19, 19, 18, 17, 17, 1, 1, 5, 5, 0, 4, 0, 0, 5, 6, 2, 2, 0, 4, 0, 0, 9, 7, 8, 0, 10, 0, 1, 1, 10, 14, 14, 10, 18, 16, 16, 16, 14, 15, 15, 0, 10, 9, 9, 11, 5, 20, 10, 8, 10, 10, 11, 8, 9, 14, 2, 0, 16, 12, 12, 6, 0, 8, 8, 11, 3, 12, 16, 6, 10, 10, 12, 12, 15, 15, 20, 20, 19, 4, 3, 15, 2, 12, 11, 1, 10, 3, 6, 0, 0, 16, 12, 6, 22, 8, 8, 2, 17, 9, 5, 9, 11, 13, 1, 18, 12, 10, 6, 18, 18, 17, 19, 14, 10, 9, 17, 8, 6, 9, 9, 17, 20, 20, 20, 17, 17, 2, 2, 0, 20, 6, 9, 9, 9, 4, 9, 0, 1, 0, 0, 12, 12, 5, 6, 5, 16, 13, 13, 4, 4, 7, 19, 11, 2, 2, 13, 0, 11, 1, 10, 19, 10, 1, 1, 10, 10, 6, 12, 7, 7, 2, 5, 13, 4, 2, 6, 8, 20, 15, 17, 0, 0, 5, 2, 9, 6, 8, 1, 0, 0, 7, 5, 2, 12, 8, 8, 8, 11, 9, 14, 20, 22, 4, 17, 11, 12, 19, 18, 1, 1, 16, 1, 10, 8, 11, 11, 6, 6, 9, 8, 10, 5, 12, 14, 14, 10, 5, 4, 4, 8, 10, 5, 13, 13, 13, 1, 13, 13, 17, 17, 0, 10, 9, 9, 7, 7, 12, 15, 17, 14, 17, 3, 17, 4, 17, 8, 7, 4, 1, 5, 0, 11, 7, 7, 17, 6, 15, 15, 10, 10, 15, 1, 0, 0, 1, 22, 9, 6, 6, 9, 4, 0, 3, 6, 1, 14, 20, 1, 0, 12, 0, 7, 14, 9, 1, 11, 11, 11, 5, 18, 18, 15, 17, 17, 20, 15, 2, 8, 17, 20, 8, 7, 6, 20, 20, 1, 1, 3, 6, 9, 3, 0, 9, 4, 4, 15, 15, 15, 15, 1, 2, 1, 1, 6, 2, 11, 1, 0, 6, 7, 7, 0, 0, 13, 17, 9, 13, 19, 3, 2, 16, 0, 9, 7, 0, 6, 0, 0, 11, 7, 6, 14, 14, 0, 0, 1, 12, 8, 6, 5, 9, 8, 12, 19, 0, 4, 16, 7, 7, 6, 18, 18, 4, 0, 0, 0, 4, 14, 9, 8, 8, 7, 1, 0, 15, 10, 6, 12, 4, 1, 1, 10, 4, 13, 13, 15, 14, 19, 16, 12, 12, 10, 14, 7, 15, 9, 1, 6, 19, 0, 13, 6, 6, 6, 7, 8, 8, 10, 2, 13, 13, 10, 10, 9, 2, 2, 1, 2, 3, 8, 8, 20, 6, 6, 3, 6, 8, 2, 17, 2, 3, 6, 6, 19, 7, 11, 1, 0, 0, 7, 7, 7, 0, 0, 0, 19, 19, 9, 8, 7, 8, 8, 2, 9, 4, 8, 8, 0, 0, 0, 0, 2, 2, 6, 0, 7, 4, 5, 15, 16, 2, 1, 7, 7, 5, 1, 16, 14, 18, 16, 12, 9, 4, 2, 6, 6, 14, 14, 6, 13, 16, 20, 11, 6, 2, 13, 19, 15, 12, 8, 1, 0, 3, 3, 5, 5, 3, 4, 7, 7, 11, 11, 12, 17, 17, 11, 9, 6, 4, 9, 7, 11, 11, 11, 7, 7, 8, 2, 0, 6, 6, 6, 22, 21, 18, 20, 16, 16, 0, 0, 16, 16, 16, 16, 19, 19, 5, 6, 5, 2, 12, 3, 4, 4, 14, 14, 12, 11, 5, 4, 8, 8, 12, 15, 12, 12, 15, 6, 6, 0, 3, 3, 12, 13, 12, 14, 10, 10, 13, 10, 13, 13, 2, 2, 12, 13, 9, 10, 9, 1, 0, 5, 6, 0, 4, 3, 4, 16, 9, 5, 7, 7, 7, 9, 8, 8, 4, 17, 18, 17, 19, 20, 17, 11, 5, 8, 8, 6, 6, 5, 14, 14, 2, 1, 13, 2, 9, 9, 0, 0, 1, 11, 9, 13, 14, 0, 1, 1, 20, 0, 8, 8, 13, 13, 13, 13, 15, 15, 15, 8, 13, 13, 13, 13, 14, 18, 16, 20, 12, 12, 19, 6, 19, 19, 16, 14, 19, 19, 19, 19, 2, 17, 1};

localparam logic [2912:0][31:0] rectangle2_widths = {12, 4, 18, 9, 2, 12, 12, 4, 7, 12, 4, 19, 8, 6, 14, 14, 3, 2, 2, 2, 2, 8, 2, 10, 14, 8, 15, 5, 2, 3, 6, 13, 3, 3, 8, 7, 21, 2, 10, 2, 2, 11, 2, 2, 2, 19, 2, 2, 7, 18, 2, 6, 12, 4, 8, 18, 6, 2, 2, 8, 8, 3, 8, 12, 6, 9, 18, 16, 2, 18, 10, 14, 7, 9, 9, 4, 7, 4, 6, 2, 2, 2, 2, 6, 12, 8, 16, 3, 8, 2, 5, 2, 2, 6, 18, 4, 8, 10, 10, 18, 22, 18, 3, 2, 2, 10, 4, 2, 3, 6, 6, 2, 2, 9, 9, 2, 6, 20, 9, 9, 7, 5, 6, 18, 8, 18, 3, 4, 2, 19, 11, 11, 5, 4, 4, 5, 8, 12, 3, 6, 22, 17, 2, 3, 3, 3, 3, 4, 19, 6, 17, 3, 4, 3, 3, 10, 3, 8, 9, 6, 5, 3, 8, 3, 10, 3, 3, 10, 2, 12, 18, 22, 4, 3, 3, 11, 12, 11, 10, 1, 1, 1, 1, 1, 9, 9, 18, 4, 18, 6, 14, 3, 6, 3, 18, 5, 2, 18, 19, 2, 19, 2, 7, 20, 22, 7, 11, 11, 2, 3, 4, 12, 6, 18, 6, 8, 2, 12, 2, 2, 2, 2, 9, 7, 9, 5, 5, 16, 10, 5, 5, 2, 18, 18, 9, 7, 1, 1, 5, 7, 5, 12, 11, 15, 8, 9, 5, 5, 3, 10, 10, 16, 7, 2, 3, 6, 10, 3, 5, 8, 5, 3, 6, 6, 3, 13, 2, 3, 3, 3, 12, 2, 6, 8, 10, 6, 1, 6, 1, 1, 9, 9, 9, 9, 6, 8, 8, 2, 5, 1, 2, 3, 24, 13, 6, 16, 6, 6, 5, 2, 2, 2, 2, 2, 9, 3, 6, 5, 3, 18, 19, 2, 1, 1, 6, 2, 9, 10, 3, 11, 5, 18, 2, 8, 12, 4, 14, 4, 5, 3, 6, 20, 19, 2, 3, 2, 3, 3, 6, 15, 6, 6, 18, 12, 2, 2, 9, 13, 9, 3, 3, 3, 9, 5, 2, 2, 6, 18, 10, 11, 8, 9, 4, 3, 2, 2, 3, 3, 9, 9, 19, 19, 10, 5, 3, 3, 6, 9, 4, 14, 2, 6, 9, 7, 17, 11, 13, 9, 5, 6, 6, 8, 3, 24, 10, 6, 18, 16, 3, 6, 2, 2, 2, 9, 6, 2, 8, 5, 5, 2, 3, 19, 6, 2, 5, 5, 5, 3, 7, 9, 3, 2, 2, 9, 6, 2, 11, 6, 9, 6, 6, 9, 19, 6, 6, 2, 2, 6, 6, 2, 2, 18, 18, 11, 7, 15, 22, 8, 9, 12, 7, 11, 7, 12, 9, 22, 11, 6, 24, 5, 5, 12, 18, 8, 8, 18, 21, 2, 2, 3, 2, 2, 2, 3, 2, 8, 10, 2, 3, 3, 2, 5, 1, 5, 2, 2, 3, 7, 4, 7, 2, 6, 2, 7, 5, 4, 5, 11, 4, 8, 23, 6, 21, 2, 4, 8, 5, 10, 9, 6, 9, 9, 9, 9, 2, 18, 21, 6, 6, 6, 8, 5, 5, 5, 3, 6, 1, 2, 3, 4, 1, 2, 9, 24, 2, 2, 2, 12, 1, 12, 18, 18, 12, 2, 2, 2, 4, 16, 4, 4, 11, 8, 2, 2, 8, 6, 18, 6, 9, 4, 3, 18, 2, 2, 2, 2, 9, 12, 9, 9, 2, 2, 9, 3, 14, 3, 14, 14, 9, 9, 2, 2, 2, 2, 4, 3, 8, 5, 2, 6, 18, 4, 12, 1, 5, 5, 10, 8, 15, 4, 14, 4, 3, 3, 18, 14, 3, 3, 8, 3, 10, 3, 3, 11, 10, 2, 2, 4, 20, 10, 3, 10, 2, 5, 6, 4, 4, 9, 14, 19, 5, 8, 8, 9, 18, 18, 9, 23, 18, 6, 1, 10, 10, 2, 2, 2, 2, 3, 3, 1, 9, 1, 6, 18, 6, 4, 3, 3, 5, 7, 1, 5, 5, 3, 3, 3, 3, 3, 2, 4, 4, 10, 21, 6, 6, 6, 6, 20, 6, 4, 4, 10, 6, 8, 9, 4, 7, 3, 19, 6, 18, 2, 20, 22, 2, 2, 3, 2, 10, 6, 12, 4, 4, 17, 9, 7, 7, 1, 1, 14, 9, 18, 4, 4, 7, 22, 4, 7, 9, 22, 2, 8, 3, 2, 9, 18, 6, 2, 2, 2, 9, 8, 6, 6, 4, 19, 3, 12, 18, 4, 9, 2, 2, 2, 2, 2, 18, 20, 6, 8, 3, 7, 12, 18, 5, 5, 4, 4, 6, 2, 2, 6, 23, 19, 11, 4, 5, 9, 9, 9, 10, 3, 3, 4, 7, 5, 12, 23, 4, 18, 9, 9, 3, 3, 12, 18, 12, 18, 9, 9, 18, 2, 2, 5, 6, 2, 8, 21, 3, 11, 5, 6, 6, 22, 6, 2, 2, 3, 6, 3, 16, 2, 16, 6, 2, 4, 5, 5, 4, 4, 3, 8, 6, 9, 10, 4, 3, 6, 12, 20, 9, 9, 4, 4, 3, 4, 3, 2, 5, 7, 10, 2, 18, 8, 18, 3, 18, 4, 2, 2, 2, 12, 9, 9, 19, 11, 3, 20, 2, 8, 8, 3, 8, 16, 4, 4, 6, 2, 4, 6, 3, 7, 16, 7, 4, 2, 3, 4, 2, 4, 23, 2, 4, 10, 2, 3, 3, 6, 6, 4, 21, 4, 6, 19, 14, 6, 2, 11, 3, 2, 2, 18, 11, 20, 13, 11, 7, 5, 5, 2, 3, 4, 8, 14, 9, 18, 3, 24, 10, 18, 3, 11, 12, 4, 4, 6, 5, 2, 2, 2, 2, 16, 20, 2, 2, 6, 6, 9, 15, 19, 7, 9, 8, 18, 4, 9, 7, 11, 2, 5, 5, 8, 6, 4, 6, 4, 2, 4, 10, 7, 20, 4, 6, 12, 3, 4, 4, 3, 8, 3, 1, 5, 5, 10, 23, 7, 2, 6, 4, 8, 4, 4, 8, 5, 19, 8, 13, 24, 2, 2, 6, 6, 18, 9, 2, 2, 3, 3, 3, 3, 19, 6, 16, 3, 4, 15, 4, 2, 2, 6, 11, 21, 4, 3, 21, 19, 3, 3, 7, 9, 8, 11, 9, 18, 7, 8, 6, 2, 2, 2, 6, 6, 1, 2, 1, 6, 2, 1, 3, 5, 1, 2, 19, 18, 9, 2, 10, 10, 3, 8, 18, 3, 4, 4, 14, 4, 5, 4, 11, 6, 9, 19, 9, 18, 9, 24, 14, 9, 6, 13, 6, 7, 3, 3, 5, 8, 9, 6, 9, 6, 7, 7, 3, 3, 5, 2, 2, 3, 9, 9, 3, 4, 4, 3, 5, 5, 12, 9, 12, 11, 11, 6, 20, 14, 16, 19, 10, 4, 21, 3, 14, 2, 9, 4, 19, 20, 2, 8, 6, 6, 2, 2, 6, 6, 8, 2, 2, 2, 9, 2, 7, 7, 3, 2, 2, 3, 10, 7, 6, 6, 2, 10, 9, 6, 5, 16, 8, 2, 9, 9, 9, 9, 18, 18, 18, 19, 2, 5, 2, 2, 6, 11, 7, 18, 2, 18, 8, 18, 2, 2, 1, 1, 7, 9, 21, 7, 22, 12, 9, 6, 7, 7, 6, 6, 10, 3, 7, 7, 6, 3, 3, 3, 18, 2, 2, 2, 2, 2, 8, 9, 5, 6, 19, 4, 9, 5, 4, 6, 6, 8, 7, 10, 10, 2, 4, 4, 2, 2, 6, 6, 9, 15, 9, 9, 9, 9, 4, 2, 10, 4, 10, 9, 11, 6, 6, 9, 5, 6, 6, 12, 8, 8, 12, 4, 4, 4, 15, 8, 5, 6, 3, 2, 3, 20, 6, 10, 2, 2, 2, 2, 3, 18, 10, 4, 3, 9, 9, 2, 2, 2, 20, 20, 18, 6, 22, 6, 6, 24, 2, 2, 2, 2, 2, 9, 18, 9, 23, 18, 9, 4, 5, 4, 3, 4, 2, 2, 6, 4, 4, 3, 3, 6, 9, 4, 11, 6, 10, 10, 5, 18, 19, 6, 11, 7, 11, 5, 3, 6, 6, 6, 2, 2, 9, 18, 13, 4, 4, 4, 2, 3, 3, 5, 5, 6, 6, 6, 12, 1, 1, 1, 1, 2, 2, 18, 7, 12, 9, 20, 3, 18, 18, 6, 9, 9, 3, 6, 4, 3, 4, 3, 12, 6, 6, 9, 12, 20, 4, 1, 5, 6, 6, 4, 4, 9, 12, 2, 3, 4, 6, 8, 3, 5, 5, 6, 6, 6, 6, 18, 9, 5, 5, 3, 3, 5, 3, 18, 2, 3, 3, 2, 2, 4, 5, 22, 1, 8, 10, 4, 3, 5, 20, 6, 6, 10, 4, 3, 2, 3, 2, 2, 19, 2, 2, 2, 5, 2, 2, 8, 6, 2, 6, 12, 9, 9, 18, 22, 6, 6, 16, 9, 6, 6, 2, 8, 8, 2, 18, 18, 11, 9, 7, 6, 24, 4, 6, 2, 2, 2, 20, 6, 2, 6, 2, 1, 5, 4, 2, 2, 3, 3, 3, 2, 9, 11, 5, 5, 4, 4, 5, 21, 9, 6, 6, 4, 5, 5, 4, 5, 6, 2, 3, 3, 11, 3, 4, 4, 4, 8, 18, 16, 4, 3, 4, 4, 4, 4, 5, 7, 24, 4, 4, 12, 12, 6, 6, 4, 18, 18, 22, 12, 6, 6, 2, 9, 7, 3, 6, 2, 2, 2, 6, 14, 17, 12, 9, 12, 9, 18, 9, 9, 24, 20, 8, 4, 10, 6, 7, 7, 3, 19, 9, 9, 10, 9, 2, 2, 4, 4, 3, 6, 10, 7, 9, 2, 3, 6, 10, 10, 5, 2, 8, 12, 2, 18, 16, 6, 7, 4, 20, 3, 2, 2, 2, 4, 1, 3, 19, 9, 6, 2, 2, 4, 18, 14, 18, 9, 6, 7, 20, 9, 15, 6, 6, 9, 9, 6, 6, 4, 8, 3, 4, 24, 6, 3, 16, 4, 5, 9, 9, 6, 20, 17, 7, 23, 2, 2, 2, 18, 3, 1, 1, 6, 5, 6, 2, 5, 5, 2, 2, 6, 18, 6, 6, 11, 5, 5, 5, 3, 5, 8, 8, 11, 4, 3, 2, 2, 7, 4, 3, 3, 4, 19, 2, 18, 5, 4, 16, 18, 5, 6, 6, 11, 3, 4, 5, 4, 4, 9, 10, 21, 11, 6, 3, 6, 6, 11, 18, 22, 6, 2, 2, 18, 3, 6, 4, 18, 6, 2, 2, 18, 2, 2, 5, 5, 5, 9, 23, 8, 6, 9, 18, 11, 11, 12, 8, 14, 21, 12, 4, 7, 6, 4, 4, 6, 3, 19, 5, 9, 2, 17, 4, 3, 16, 5, 6, 3, 20, 5, 2, 2, 2, 9, 2, 2, 2, 2, 6, 6, 3, 3, 3, 7, 12, 2, 6, 2, 6, 14, 16, 2, 21, 6, 5, 8, 7, 4, 6, 6, 7, 9, 6, 8, 18, 9, 19, 24, 9, 9, 18, 18, 1, 8, 18, 1, 4, 10, 3, 10, 5, 6, 9, 4, 5, 7, 10, 4, 2, 18, 2, 2, 2, 2, 9, 14, 15, 4, 3, 3, 6, 4, 8, 6, 6, 12, 9, 24, 11, 9, 5, 2, 6, 6, 16, 10, 18, 9, 10, 18, 15, 15, 12, 2, 2, 3, 10, 18, 10, 5, 7, 3, 3, 3, 4, 2, 1, 8, 2, 2, 4, 4, 2, 2, 9, 9, 2, 2, 2, 4, 12, 12, 14, 20, 4, 13, 6, 2, 12, 15, 4, 6, 8, 1, 2, 2, 6, 17, 5, 5, 18, 4, 3, 2, 21, 3, 6, 8, 9, 5, 3, 5, 3, 3, 5, 8, 6, 3, 2, 2, 10, 18, 7, 7, 1, 5, 12, 20, 19, 9, 14, 14, 3, 18, 6, 9, 10, 10, 12, 10, 3, 3, 4, 4, 2, 10, 3, 7, 13, 4, 10, 5, 2, 6, 9, 7, 22, 18, 2, 2, 2, 2, 3, 2, 9, 9, 15, 3, 6, 10, 6, 9, 2, 2, 2, 2, 2, 3, 8, 2, 3, 18, 10, 10, 9, 3, 5, 4, 19, 6, 7, 16, 18, 10, 4, 6, 4, 3, 6, 6, 9, 12, 10, 10, 6, 6, 4, 6, 10, 10, 18, 4, 24, 6, 10, 19, 10, 7, 4, 5, 2, 2, 2, 2, 3, 8, 8, 12, 3, 7, 7, 4, 4, 2, 1, 3, 10, 12, 4, 4, 6, 5, 7, 5, 3, 12, 4, 11, 12, 9, 23, 19, 6, 6, 2, 2, 2, 2, 2, 8, 7, 9, 2, 2, 10, 3, 5, 4, 4, 4, 2, 2, 2, 2, 24, 10, 23, 19, 18, 9, 6, 6, 20, 3, 18, 3, 6, 6, 6, 5, 2, 2, 2, 6, 2, 5, 2, 1, 2, 2, 19, 9, 7, 14, 8, 8, 9, 9, 6, 2, 2, 2, 2, 2, 9, 2, 4, 9, 7, 5, 10, 4, 22, 2, 3, 2, 5, 4, 6, 12, 6, 6, 2, 19, 6, 8, 6, 6, 6, 24, 10, 10, 19, 19, 16, 8, 6, 2, 18, 18, 6, 6, 6, 4, 6, 10, 2, 3, 2, 3, 3, 15, 20, 2, 6, 2, 3, 2, 6, 9, 9, 6, 2, 4, 18, 2, 19, 15, 7, 11, 2, 18, 3, 20, 5, 4, 3, 4, 4, 6, 6, 1, 7, 4, 4, 5, 3, 10, 18, 15, 8, 24, 2, 4, 10, 18, 24, 2, 4, 18, 18, 9, 10, 7, 6, 7, 7, 6, 6, 2, 18, 2, 10, 11, 4, 9, 2, 4, 4, 4, 3, 4, 3, 4, 4, 14, 11, 2, 11, 9, 18, 4, 18, 18, 9, 9, 9, 3, 3, 2, 2, 2, 2, 2, 2, 6, 2, 5, 5, 2, 3, 4, 4, 24, 7, 4, 5, 4, 2, 3, 3, 18, 16, 16, 4, 8, 4, 9, 9, 16, 19, 9, 1, 24, 5, 19, 3, 12, 9, 10, 20, 7, 7, 2, 5, 6, 3, 6, 2, 9, 11, 11, 3, 2, 6, 24, 8, 6, 2, 5, 2, 3, 3, 3, 3, 2, 2, 5, 5, 9, 14, 10, 5, 1, 3, 5, 8, 12, 2, 3, 2, 2, 19, 4, 2, 18, 10, 18, 3, 24, 4, 2, 4, 5, 9, 19, 8, 8, 10, 6, 7, 6, 6, 15, 6, 7, 6, 6, 2, 2, 3, 3, 9, 9, 9, 9, 18, 18, 2, 2, 1, 8, 2, 5, 6, 7, 2, 6, 5, 9, 1, 1, 3, 3, 6, 3, 3, 5, 5, 5, 2, 2, 5, 7, 6, 24, 7, 2, 2, 7, 8, 7, 5, 3, 8, 8, 3, 3, 5, 6, 12, 5, 9, 11, 4, 9, 13, 2, 2, 10, 20, 9, 2, 2, 22, 9, 24, 16, 18, 2, 3, 3, 4, 7, 10, 19, 2, 2, 2, 3, 6, 2, 8, 18, 5, 12, 6, 10, 24, 9, 2, 2, 8, 2, 3, 6, 5, 5, 3, 3, 7, 3, 6, 2, 16, 7, 8, 3, 3, 1, 11, 18, 6, 3, 4, 4, 10, 1, 9, 9, 9, 9, 9, 6, 10, 9, 18, 3, 2, 18, 3, 10, 3, 1, 3, 11, 3, 11, 4, 10, 7, 6, 2, 4, 4, 4, 3, 4, 3, 3, 3, 3, 5, 3, 3, 5, 8, 19, 9, 9, 6, 3, 14, 4, 7, 4, 4, 22, 6, 3, 3, 17, 6, 9, 10, 5, 8, 3, 3, 19, 6, 10, 10, 9, 18, 18, 9, 9, 2, 2, 8, 6, 2, 6, 2, 6, 6, 3, 3, 2, 6, 6, 2, 2, 6, 4, 4, 9, 9, 6, 9, 18, 3, 3, 3, 7, 2, 6, 6, 3, 16, 3, 2, 2, 2, 5, 9, 18, 5, 17, 9, 24, 18, 2, 14, 3, 2, 2, 2, 7, 4, 3, 3, 4, 4, 4, 4, 6, 9, 10, 3, 4, 8, 5, 5, 5, 6, 5, 6, 5, 5, 6, 18, 18, 2, 4, 4, 4, 6, 9, 9, 6, 6, 9, 6, 3, 2, 10, 10, 4, 1, 1, 1, 6, 5, 7, 7, 3, 4, 4, 5, 9, 9, 12, 5, 3, 2, 7, 2, 7, 19, 3, 5, 5, 4, 6, 3, 7, 7, 13, 3, 17, 17, 8, 8, 12, 5, 6, 9, 1, 1, 2, 2, 11, 4, 4, 3, 6, 3, 3, 6, 3, 8, 5, 7, 11, 6, 4, 2, 1, 1, 9, 4, 3, 9, 1, 1, 5, 18, 20, 9, 19, 19, 9, 6, 7, 3, 3, 3, 2, 2, 2, 2, 4, 4, 2, 3, 3, 9, 8, 10, 9, 3, 5, 3, 12, 4, 4, 6, 12, 6, 6, 7, 6, 19, 6, 2, 2, 5, 5, 7, 3, 8, 10, 18, 2, 20, 2, 6, 6, 18, 15, 18, 1, 2, 2, 4, 4, 20, 13, 7, 7, 5, 5, 3, 18, 18, 9, 15, 6, 12, 3, 13, 11, 6, 6, 24, 10, 18, 10, 1, 6, 2, 2, 18, 9, 6, 9, 5, 5, 5, 5, 9, 9, 10, 10, 18, 18, 9, 7, 19, 16, 8, 6, 1, 1, 4, 4, 3, 6, 4, 6, 9, 9, 3, 18, 3, 3, 18, 18, 22, 7, 6, 6, 8, 16, 6, 4, 3, 3, 18, 10, 9, 9, 1, 1, 2, 6, 8, 9, 16, 18, 2, 3, 2, 2, 6, 18, 24, 9, 4, 13, 16, 14, 9, 16, 13, 13, 12, 10, 18, 18, 9, 11, 8, 8, 18, 5, 6, 9, 2, 3, 2, 2, 5, 9, 17, 12, 8, 5, 2, 2, 2, 13, 19, 6, 4, 3, 3, 3, 9, 2, 4, 4, 5, 5, 4, 4, 16, 16, 7, 3, 9, 17, 8, 8, 5, 11, 12, 6, 3, 3, 9, 11, 9, 18, 19, 18, 9, 9, 9, 9, 1, 24, 3};

localparam logic [2912:0][31:0] rectangle2_heights = {3, 7, 3, 2, 19, 8, 3, 5, 3, 2, 7, 4, 3, 5, 5, 3, 6, 10, 10, 9, 11, 13, 9, 2, 6, 3, 3, 7, 10, 6, 3, 2, 15, 15, 15, 6, 4, 10, 10, 13, 13, 19, 9, 11, 9, 1, 9, 9, 7, 1, 11, 3, 3, 6, 5, 2, 3, 13, 13, 23, 4, 7, 3, 2, 6, 2, 1, 6, 20, 1, 7, 4, 3, 2, 2, 5, 7, 5, 3, 9, 9, 9, 9, 4, 3, 6, 4, 6, 3, 9, 4, 9, 9, 6, 1, 5, 5, 2, 2, 1, 1, 1, 15, 10, 10, 3, 9, 9, 6, 3, 3, 9, 9, 2, 2, 10, 3, 1, 6, 24, 5, 6, 6, 1, 4, 3, 6, 18, 14, 1, 13, 2, 10, 6, 6, 4, 4, 2, 6, 3, 5, 3, 10, 8, 7, 22, 22, 16, 2, 4, 2, 7, 5, 11, 11, 9, 7, 8, 14, 3, 8, 6, 4, 6, 2, 6, 6, 2, 9, 2, 1, 1, 8, 6, 6, 2, 2, 6, 17, 24, 24, 22, 22, 18, 2, 2, 1, 9, 1, 4, 3, 6, 8, 16, 3, 4, 9, 1, 1, 9, 6, 9, 6, 1, 1, 3, 2, 2, 11, 6, 5, 6, 5, 1, 3, 3, 9, 7, 13, 13, 9, 9, 2, 3, 2, 4, 9, 2, 2, 10, 7, 9, 1, 1, 2, 3, 18, 18, 10, 4, 9, 3, 4, 3, 19, 3, 4, 4, 8, 2, 2, 3, 5, 13, 14, 5, 2, 14, 4, 5, 4, 6, 3, 3, 8, 2, 9, 6, 9, 9, 2, 9, 3, 7, 4, 3, 20, 3, 21, 23, 2, 2, 2, 2, 4, 19, 6, 10, 6, 19, 10, 6, 1, 2, 3, 2, 3, 3, 4, 9, 9, 9, 15, 15, 2, 7, 5, 4, 8, 1, 1, 9, 18, 18, 9, 14, 3, 8, 6, 8, 5, 1, 10, 4, 3, 5, 4, 5, 7, 8, 8, 1, 2, 9, 14, 12, 9, 9, 3, 2, 3, 3, 1, 2, 9, 9, 2, 2, 2, 15, 6, 7, 2, 4, 19, 19, 3, 1, 3, 2, 3, 11, 7, 10, 9, 9, 6, 6, 2, 2, 1, 1, 2, 6, 6, 6, 3, 6, 6, 4, 9, 3, 2, 23, 2, 6, 2, 2, 4, 3, 3, 4, 6, 1, 2, 3, 3, 3, 6, 4, 9, 10, 9, 21, 7, 9, 4, 4, 4, 9, 17, 3, 3, 19, 7, 6, 6, 6, 4, 2, 6, 14, 14, 2, 5, 11, 7, 3, 2, 3, 3, 2, 1, 3, 3, 9, 9, 7, 5, 9, 9, 1, 1, 6, 3, 2, 1, 24, 4, 3, 4, 3, 3, 8, 2, 1, 4, 3, 2, 5, 5, 2, 1, 3, 3, 1, 5, 24, 11, 6, 10, 24, 24, 7, 12, 14, 2, 9, 7, 15, 9, 7, 18, 6, 10, 9, 7, 3, 6, 6, 9, 3, 13, 3, 4, 5, 4, 3, 5, 5, 2, 3, 2, 12, 5, 5, 12, 2, 2, 8, 2, 2, 2, 2, 9, 1, 2, 3, 3, 3, 5, 8, 5, 5, 10, 3, 18, 9, 7, 5, 18, 9, 2, 1, 9, 10, 12, 6, 21, 4, 4, 1, 2, 9, 9, 22, 7, 5, 7, 7, 3, 9, 16, 16, 4, 3, 1, 3, 2, 5, 6, 1, 11, 11, 9, 9, 9, 2, 2, 2, 17, 17, 2, 6, 6, 6, 5, 5, 2, 2, 14, 9, 15, 15, 9, 21, 4, 6, 9, 3, 1, 5, 2, 20, 4, 4, 3, 3, 2, 6, 3, 5, 7, 6, 1, 6, 6, 6, 3, 7, 2, 6, 7, 4, 2, 9, 9, 5, 1, 2, 11, 3, 9, 4, 3, 5, 8, 2, 3, 4, 8, 18, 11, 5, 1, 1, 2, 5, 1, 3, 22, 2, 2, 12, 9, 9, 9, 6, 9, 19, 2, 19, 3, 1, 4, 5, 6, 8, 4, 3, 19, 20, 20, 6, 6, 7, 7, 7, 9, 10, 10, 2, 2, 6, 6, 3, 3, 2, 3, 5, 5, 13, 5, 3, 2, 5, 6, 6, 1, 3, 1, 9, 1, 1, 9, 23, 19, 9, 2, 6, 3, 5, 5, 3, 4, 3, 3, 18, 18, 2, 2, 3, 8, 5, 4, 2, 5, 4, 2, 2, 17, 9, 6, 9, 6, 1, 3, 11, 10, 17, 2, 3, 4, 4, 5, 1, 7, 3, 1, 6, 14, 9, 18, 18, 10, 11, 1, 1, 4, 4, 6, 7, 5, 1, 4, 4, 9, 9, 6, 9, 11, 6, 1, 1, 2, 5, 4, 3, 2, 2, 4, 18, 10, 5, 6, 7, 2, 2, 5, 1, 2, 2, 6, 6, 3, 1, 2, 1, 2, 2, 1, 10, 9, 4, 4, 11, 3, 2, 6, 4, 4, 3, 4, 11, 4, 9, 9, 7, 8, 7, 10, 10, 2, 4, 9, 5, 4, 4, 5, 5, 8, 3, 4, 2, 2, 6, 6, 3, 2, 1, 3, 2, 6, 6, 8, 5, 6, 9, 4, 6, 2, 15, 1, 3, 1, 6, 1, 5, 9, 9, 9, 2, 2, 2, 1, 6, 6, 1, 10, 3, 3, 7, 3, 4, 6, 5, 3, 9, 6, 3, 6, 3, 3, 3, 7, 9, 7, 8, 10, 5, 1, 12, 5, 2, 12, 6, 6, 13, 13, 6, 1, 6, 7, 1, 2, 4, 9, 2, 6, 23, 23, 1, 2, 1, 2, 15, 3, 4, 4, 9, 6, 5, 3, 3, 2, 1, 6, 1, 2, 1, 8, 2, 11, 5, 6, 3, 10, 9, 10, 10, 10, 3, 1, 13, 13, 7, 3, 2, 2, 1, 8, 2, 4, 1, 6, 2, 7, 3, 9, 5, 5, 3, 3, 7, 6, 6, 9, 8, 2, 7, 1, 8, 5, 2, 7, 8, 8, 6, 6, 8, 18, 7, 7, 3, 6, 3, 9, 3, 8, 4, 8, 8, 5, 4, 1, 9, 4, 1, 11, 9, 4, 3, 1, 2, 9, 9, 19, 19, 8, 8, 1, 4, 2, 6, 7, 6, 5, 9, 9, 4, 2, 1, 6, 6, 1, 1, 7, 7, 7, 2, 3, 2, 2, 1, 3, 4, 5, 9, 10, 10, 3, 3, 19, 9, 19, 4, 9, 19, 6, 5, 18, 12, 1, 1, 2, 9, 2, 2, 6, 8, 1, 6, 5, 5, 2, 5, 4, 7, 3, 3, 2, 1, 2, 1, 2, 1, 2, 2, 3, 2, 4, 3, 6, 7, 4, 3, 2, 3, 2, 3, 5, 5, 17, 10, 4, 9, 9, 8, 2, 2, 6, 5, 6, 8, 4, 4, 2, 2, 3, 2, 2, 9, 2, 7, 3, 1, 2, 5, 1, 6, 3, 9, 3, 7, 1, 1, 13, 4, 3, 3, 10, 10, 3, 3, 21, 13, 21, 20, 2, 9, 3, 3, 9, 10, 9, 9, 2, 7, 3, 6, 10, 4, 2, 3, 7, 2, 3, 10, 2, 2, 2, 2, 1, 1, 1, 1, 11, 6, 11, 11, 3, 2, 12, 1, 9, 1, 3, 1, 9, 9, 18, 18, 3, 2, 1, 3, 1, 8, 2, 4, 3, 3, 3, 3, 5, 8, 15, 8, 4, 6, 6, 6, 1, 11, 15, 13, 9, 9, 4, 4, 4, 3, 1, 10, 2, 4, 7, 3, 3, 3, 3, 2, 3, 9, 8, 8, 9, 16, 4, 4, 2, 11, 2, 2, 2, 2, 5, 16, 2, 5, 2, 2, 2, 5, 3, 2, 16, 13, 3, 3, 3, 3, 11, 5, 5, 7, 3, 6, 8, 3, 6, 9, 8, 1, 3, 2, 9, 9, 9, 9, 6, 1, 2, 6, 6, 11, 11, 11, 11, 9, 1, 1, 1, 3, 3, 3, 3, 2, 10, 9, 9, 9, 9, 2, 1, 2, 2, 1, 2, 5, 6, 5, 12, 5, 9, 9, 4, 5, 5, 7, 19, 3, 3, 5, 4, 3, 9, 6, 4, 1, 1, 3, 2, 4, 3, 4, 7, 3, 4, 3, 9, 23, 2, 1, 7, 6, 6, 7, 9, 6, 6, 5, 5, 3, 5, 4, 2, 19, 19, 20, 20, 12, 12, 7, 4, 4, 5, 1, 6, 1, 1, 3, 2, 2, 7, 3, 9, 6, 5, 6, 3, 3, 3, 2, 3, 1, 6, 24, 4, 6, 4, 7, 7, 5, 2, 9, 7, 5, 3, 12, 14, 4, 4, 3, 3, 3, 3, 2, 2, 4, 4, 12, 11, 4, 7, 1, 9, 7, 6, 11, 11, 18, 5, 1, 20, 4, 2, 5, 7, 4, 3, 4, 3, 2, 9, 8, 17, 6, 17, 17, 1, 9, 9, 9, 4, 9, 9, 4, 3, 9, 3, 2, 2, 2, 1, 2, 3, 3, 3, 2, 3, 3, 23, 3, 4, 23, 1, 1, 2, 2, 3, 3, 2, 5, 6, 9, 9, 9, 1, 3, 13, 4, 13, 18, 5, 8, 9, 9, 7, 7, 8, 10, 3, 4, 5, 5, 16, 16, 5, 1, 2, 4, 6, 6, 4, 4, 5, 4, 3, 9, 7, 7, 6, 8, 7, 7, 9, 4, 4, 4, 10, 6, 10, 10, 7, 7, 4, 3, 5, 11, 8, 3, 3, 6, 3, 5, 1, 1, 1, 3, 3, 3, 9, 2, 6, 6, 4, 16, 9, 9, 5, 2, 4, 7, 3, 3, 5, 1, 2, 2, 2, 3, 6, 5, 2, 4, 5, 5, 6, 4, 2, 2, 2, 2, 9, 9, 5, 13, 6, 3, 2, 5, 3, 9, 7, 3, 3, 2, 6, 9, 7, 3, 9, 1, 2, 3, 3, 5, 1, 6, 9, 11, 11, 5, 18, 6, 1, 2, 5, 9, 9, 5, 1, 2, 1, 2, 3, 4, 1, 2, 2, 3, 3, 2, 2, 3, 3, 5, 4, 6, 5, 3, 4, 6, 2, 5, 4, 4, 4, 3, 4, 8, 3, 1, 9, 9, 13, 1, 6, 24, 24, 10, 6, 3, 11, 4, 18, 16, 16, 3, 1, 3, 3, 2, 4, 7, 7, 6, 4, 3, 3, 7, 5, 6, 18, 9, 3, 5, 6, 6, 5, 1, 13, 1, 4, 5, 2, 1, 4, 3, 3, 4, 6, 5, 7, 10, 10, 3, 3, 2, 8, 11, 6, 9, 9, 2, 2, 2, 3, 9, 9, 1, 13, 4, 6, 1, 4, 9, 13, 1, 9, 9, 4, 4, 4, 2, 5, 6, 3, 2, 1, 2, 2, 3, 4, 2, 1, 3, 5, 3, 3, 5, 5, 4, 6, 1, 5, 12, 12, 3, 11, 13, 3, 6, 3, 6, 1, 10, 9, 9, 9, 2, 9, 9, 16, 16, 3, 3, 6, 6, 8, 6, 2, 20, 3, 9, 3, 2, 6, 9, 2, 3, 4, 8, 3, 5, 4, 4, 3, 5, 21, 21, 1, 2, 1, 1, 2, 2, 1, 1, 23, 3, 1, 23, 5, 4, 7, 3, 6, 5, 2, 5, 4, 24, 2, 5, 9, 1, 9, 9, 9, 11, 2, 4, 3, 5, 12, 12, 4, 10, 3, 9, 5, 11, 2, 4, 2, 2, 4, 9, 3, 3, 3, 2, 1, 3, 3, 1, 2, 2, 2, 12, 9, 6, 2, 3, 3, 4, 3, 7, 6, 6, 6, 14, 18, 12, 14, 14, 20, 20, 17, 17, 2, 2, 13, 13, 9, 7, 2, 2, 3, 1, 5, 3, 6, 9, 2, 4, 5, 3, 5, 18, 14, 9, 3, 2, 4, 4, 1, 5, 6, 12, 1, 6, 3, 9, 5, 6, 6, 11, 6, 6, 4, 4, 3, 13, 9, 9, 3, 1, 3, 3, 21, 4, 2, 1, 1, 2, 4, 6, 7, 2, 3, 2, 3, 3, 2, 4, 7, 7, 5, 5, 10, 2, 6, 3, 3, 5, 2, 4, 9, 6, 2, 3, 1, 1, 9, 9, 20, 20, 7, 9, 2, 2, 2, 6, 3, 2, 3, 7, 9, 9, 9, 9, 9, 6, 3, 11, 6, 1, 4, 2, 2, 6, 4, 8, 1, 3, 8, 4, 1, 7, 5, 3, 6, 9, 4, 4, 3, 2, 2, 2, 3, 3, 8, 3, 2, 2, 1, 5, 2, 3, 3, 4, 2, 14, 8, 4, 9, 10, 13, 13, 6, 3, 7, 2, 6, 4, 3, 5, 5, 13, 19, 6, 2, 2, 5, 7, 3, 12, 7, 4, 6, 3, 5, 2, 2, 2, 2, 4, 7, 3, 9, 12, 9, 9, 11, 6, 3, 2, 11, 11, 2, 7, 4, 5, 6, 6, 16, 16, 16, 16, 1, 2, 4, 1, 1, 2, 3, 3, 3, 7, 1, 7, 5, 5, 9, 5, 9, 9, 10, 3, 10, 4, 10, 19, 10, 9, 2, 2, 3, 4, 3, 3, 2, 2, 8, 9, 9, 9, 10, 10, 3, 9, 6, 4, 6, 7, 2, 5, 1, 10, 6, 9, 8, 6, 7, 2, 3, 3, 10, 1, 4, 11, 4, 4, 3, 2, 2, 2, 1, 1, 3, 5, 5, 9, 1, 1, 3, 3, 3, 5, 8, 5, 13, 13, 9, 11, 11, 2, 1, 9, 7, 9, 6, 9, 10, 3, 3, 3, 9, 15, 1, 9, 1, 2, 5, 14, 9, 1, 6, 1, 4, 5, 6, 5, 5, 3, 3, 20, 3, 13, 5, 4, 7, 2, 1, 4, 9, 1, 13, 5, 3, 1, 1, 11, 5, 1, 1, 5, 21, 3, 3, 4, 4, 3, 3, 9, 1, 9, 2, 3, 5, 2, 9, 5, 5, 5, 7, 5, 7, 5, 6, 6, 2, 10, 2, 2, 1, 13, 1, 1, 2, 2, 2, 16, 16, 10, 10, 24, 10, 9, 9, 5, 9, 8, 8, 9, 6, 18, 18, 2, 3, 15, 14, 5, 9, 8, 8, 4, 2, 5, 5, 3, 5, 2, 2, 4, 2, 2, 23, 2, 4, 9, 6, 4, 2, 2, 1, 10, 10, 9, 12, 4, 7, 8, 9, 2, 2, 3, 6, 9, 7, 2, 10, 21, 10, 4, 9, 6, 6, 6, 6, 9, 9, 4, 4, 2, 2, 2, 4, 19, 8, 4, 3, 2, 10, 6, 22, 22, 1, 5, 9, 1, 5, 1, 6, 7, 5, 9, 5, 5, 2, 1, 6, 8, 2, 3, 3, 3, 3, 4, 8, 4, 3, 3, 9, 9, 6, 6, 2, 2, 2, 2, 1, 1, 11, 11, 24, 4, 9, 7, 3, 3, 10, 3, 7, 6, 24, 24, 7, 7, 19, 6, 6, 4, 5, 5, 10, 10, 4, 4, 3, 1, 10, 9, 19, 3, 10, 9, 5, 6, 10, 10, 6, 6, 4, 3, 2, 5, 2, 5, 6, 2, 2, 9, 9, 2, 1, 2, 19, 19, 1, 2, 9, 4, 2, 10, 6, 6, 5, 5, 2, 1, 9, 9, 9, 9, 5, 10, 3, 1, 6, 2, 3, 2, 2, 2, 11, 11, 3, 9, 6, 3, 4, 4, 6, 6, 4, 7, 4, 9, 6, 10, 6, 7, 6, 18, 7, 1, 4, 7, 6, 6, 11, 20, 2, 2, 2, 2, 12, 4, 2, 3, 1, 8, 12, 1, 7, 2, 7, 19, 7, 3, 7, 3, 5, 19, 6, 7, 9, 5, 5, 5, 7, 5, 9, 9, 7, 7, 4, 6, 6, 6, 8, 1, 2, 2, 5, 6, 3, 10, 3, 5, 14, 2, 3, 7, 6, 6, 3, 2, 2, 6, 3, 6, 6, 1, 3, 2, 2, 2, 1, 1, 2, 2, 9, 12, 4, 3, 12, 3, 9, 3, 3, 10, 10, 9, 4, 3, 9, 9, 3, 10, 10, 2, 2, 3, 2, 1, 7, 6, 6, 3, 13, 3, 15, 7, 3, 6, 9, 24, 24, 4, 2, 2, 4, 2, 7, 1, 1, 9, 6, 6, 9, 10, 9, 7, 5, 8, 9, 5, 5, 5, 5, 5, 2, 3, 7, 8, 4, 4, 4, 4, 9, 4, 4, 6, 6, 7, 1, 1, 10, 24, 15, 24, 9, 2, 3, 3, 3, 2, 10, 23, 9, 2, 3, 5, 19, 18, 18, 3, 9, 7, 7, 6, 5, 5, 8, 2, 2, 3, 4, 6, 9, 3, 22, 3, 1, 24, 6, 7, 5, 5, 6, 7, 7, 2, 6, 3, 3, 3, 3, 5, 8, 8, 2, 18, 19, 16, 16, 2, 5, 5, 6, 5, 7, 6, 3, 6, 10, 6, 4, 2, 4, 5, 9, 22, 22, 2, 5, 6, 13, 24, 24, 4, 1, 1, 2, 5, 1, 2, 8, 4, 16, 16, 16, 14, 14, 22, 22, 20, 20, 9, 16, 6, 3, 4, 2, 2, 6, 4, 6, 3, 6, 5, 4, 2, 3, 3, 9, 3, 1, 3, 9, 9, 5, 5, 3, 7, 5, 3, 1, 10, 1, 11, 4, 3, 1, 2, 1, 18, 10, 10, 9, 9, 1, 2, 7, 7, 6, 6, 6, 1, 1, 5, 2, 3, 3, 6, 2, 13, 3, 3, 1, 2, 1, 2, 19, 8, 9, 9, 1, 2, 3, 2, 4, 4, 6, 6, 2, 2, 2, 2, 1, 1, 6, 3, 5, 2, 12, 15, 19, 19, 5, 5, 6, 3, 5, 5, 5, 5, 6, 1, 6, 6, 1, 1, 1, 10, 17, 17, 11, 3, 4, 7, 7, 7, 1, 2, 2, 2, 18, 18, 10, 3, 3, 2, 2, 1, 9, 6, 9, 9, 3, 3, 1, 2, 5, 3, 3, 3, 2, 2, 3, 3, 3, 3, 1, 1, 2, 2, 3, 5, 1, 5, 3, 3, 9, 6, 9, 9, 6, 12, 11, 2, 3, 9, 9, 9, 12, 2, 1, 4, 5, 7, 7, 7, 2, 10, 6, 6, 4, 4, 5, 5, 4, 4, 3, 7, 2, 3, 5, 5, 4, 3, 4, 3, 6, 6, 2, 5, 2, 1, 1, 1, 2, 2, 2, 2, 20, 4, 11};

localparam logic [2912:0][31:0] rectangle2_weights = {384, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 256, 384, 384, 384, 384, 256, 384, 256, 256, 384, 256, 384, 384, 256, 256, 384, 256, 384, 256, 256, 384, 256, 256, 384, 384, 256, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 384, 256, 256, 256, 384, 384, 256, 256, 384, 256, 384, 384, 256, 256, 256, 256, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 256, 384, 256, 256, 256, 256, 256, 256, 384, 256, 256, 384, 384, 256, 256, 256, 256, 256, 384, 256, 256, 256, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 256, 256, 384, 256, 256, 256, 256, 384, 384, 384, 384, 384, 256, 384, 256, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 256, 256, 384, 384, 256, 256, 384, 256, 256, 256, 384, 256, 384, 256, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 384, 256, 256, 256, 256, 256, 256, 256, 384, 384, 256, 384, 256, 384, 256, 256, 256, 256, 384, 384, 256, 256, 384, 256, 256, 384, 384, 256, 256, 384, 384, 256, 256, 384, 384, 256, 256, 384, 384, 384, 256, 384, 256, 256, 256, 384, 384, 384, 256, 256, 384, 384, 256, 384, 384, 256, 384, 384, 384, 256, 256, 256, 256, 384, 384, 256, 256, 256, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 256, 256, 384, 256, 384, 384, 384, 256, 256, 256, 256, 384, 256, 384, 256, 256, 384, 384, 256, 384, 384, 384, 256, 384, 256, 256, 256, 256, 384, 384, 384, 384, 256, 256, 256, 384, 384, 256, 256, 256, 384, 256, 384, 384, 256, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 384, 384, 256, 256, 256, 384, 256, 384, 384, 256, 384, 256, 256, 384, 384, 384, 384, 256, 384, 384, 384, 384, 384, 384, 256, 384, 256, 384, 256, 256, 256, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 256, 256, 384, 384, 384, 384, 384, 256, 256, 256, 384, 256, 256, 256, 384, 384, 384, 384, 256, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 384, 256, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 256, 256, 384, 384, 384, 256, 384, 384, 384, 384, 256, 256, 384, 384, 256, 256, 384, 256, 384, 384, 384, 384, 256, 256, 256, 256, 384, 256, 384, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 256, 256, 384, 256, 256, 384, 256, 384, 384, 384, 256, 384, 384, 256, 256, 384, 384, 384, 256, 384, 384, 256, 256, 384, 384, 384, 384, 256, 256, 256, 256, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 384, 256, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 256, 256, 256, 256, 256, 256, 384, 384, 384, 256, 384, 256, 384, 384, 384, 384, 384, 256, 256, 256, 256, 384, 256, 256, 384, 384, 256, 384, 256, 256, 256, 384, 256, 256, 256, 384, 384, 384, 384, 256, 384, 384, 384, 384, 256, 256, 256, 256, 384, 384, 384, 384, 256, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 256, 256, 384, 384, 256, 256, 384, 256, 256, 384, 384, 256, 384, 256, 256, 256, 256, 384, 384, 256, 256, 384, 256, 384, 256, 256, 384, 256, 384, 384, 384, 384, 384, 256, 384, 256, 256, 256, 256, 256, 256, 384, 256, 256, 256, 384, 256, 384, 384, 384, 256, 384, 256, 384, 384, 384, 384, 256, 384, 384, 384, 256, 384, 384, 384, 384, 384, 384, 256, 384, 384, 384, 256, 384, 384, 384, 256, 256, 256, 256, 256, 384, 256, 256, 384, 384, 256, 256, 256, 384, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 384, 384, 384, 256, 256, 384, 384, 256, 256, 256, 384, 384, 256, 256, 256, 384, 256, 256, 256, 256, 384, 384, 256, 256, 384, 384, 256, 256, 256, 384, 256, 256, 256, 384, 256, 256, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 384, 256, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 256, 256, 256, 384, 384, 256, 384, 384, 256, 256, 256, 384, 384, 384, 256, 384, 384, 256, 384, 256, 256, 256, 256, 384, 256, 256, 256, 256, 256, 384, 256, 384, 384, 384, 384, 384, 384, 256, 256, 384, 384, 384, 256, 384, 256, 256, 384, 256, 256, 384, 384, 256, 384, 256, 256, 384, 256, 384, 384, 256, 256, 256, 384, 256, 384, 384, 384, 384, 256, 256, 384, 384, 256, 384, 384, 256, 384, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 384, 384, 384, 384, 256, 256, 256, 384, 384, 384, 256, 256, 384, 384, 256, 384, 256, 256, 256, 256, 256, 256, 384, 256, 384, 256, 384, 256, 256, 256, 384, 256, 256, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 384, 256, 256, 384, 256, 256, 384, 256, 384, 256, 256, 256, 256, 256, 384, 384, 256, 256, 256, 384, 256, 384, 384, 384, 384, 256, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 256, 256, 256, 384, 256, 256, 256, 384, 256, 256, 256, 256, 256, 384, 256, 256, 256, 256, 256, 256, 256, 256, 384, 256, 256, 384, 256, 256, 256, 384, 384, 384, 256, 256, 384, 256, 256, 256, 256, 256, 384, 256, 384, 256, 384, 256, 256, 384, 384, 256, 256, 384, 384, 256, 256, 384, 384, 384, 384, 256, 256, 256, 384, 384, 256, 384, 384, 256, 256, 256, 384, 256, 256, 256, 384, 384, 256, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 384, 256, 256, 384, 256, 256, 384, 384, 384, 384, 256, 384, 256, 256, 256, 384, 384, 256, 256, 256, 384, 384, 384, 256, 256, 256, 256, 384, 256, 384, 256, 384, 256, 384, 384, 256, 384, 384, 384, 384, 256, 384, 384, 384, 256, 256, 256, 256, 384, 256, 256, 256, 384, 256, 256, 256, 384, 256, 384, 384, 256, 256, 256, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 384, 384, 256, 384, 384, 384, 384, 256, 384, 256, 256, 384, 384, 256, 256, 256, 256, 384, 384, 256, 256, 384, 384, 384, 256, 256, 256, 384, 256, 256, 256, 256, 256, 384, 256, 384, 384, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 256, 384, 384, 256, 256, 384, 256, 256, 256, 384, 384, 384, 384, 384, 384, 256, 256, 256, 384, 256, 384, 384, 384, 384, 384, 256, 256, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 256, 256, 384, 256, 384, 256, 384, 256, 256, 256, 384, 256, 256, 384, 256, 256, 256, 256, 256, 384, 384, 384, 256, 384, 256, 256, 384, 256, 384, 384, 256, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 256, 256, 256, 384, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 384, 384, 384, 256, 384, 384, 256, 384, 384, 384, 256, 384, 384, 384, 384, 256, 256, 256, 256, 384, 256, 256, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 384, 384, 256, 256, 384, 256, 384, 256, 384, 384, 384, 384, 256, 256, 256, 384, 256, 256, 384, 256, 384, 384, 384, 256, 384, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 256, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 384, 384, 384, 256, 256, 256, 384, 256, 384, 256, 384, 256, 256, 256, 256, 384, 256, 256, 256, 384, 256, 256, 256, 256, 256, 384, 256, 256, 256, 256, 256, 384, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 256, 256, 384, 256, 384, 384, 384, 384, 256, 256, 256, 256, 384, 256, 384, 384, 256, 256, 256, 256, 256, 256, 256, 256, 256, 384, 384, 384, 256, 384, 256, 256, 256, 256, 256, 384, 256, 256, 256, 256, 256, 256, 256, 384, 384, 256, 256, 384, 384, 256, 384, 256, 256, 256, 256, 256, 384, 256, 256, 256, 256, 384, 256, 384, 256, 384, 256, 384, 384, 256, 256, 384, 384, 256, 384, 384, 256, 384, 384, 256, 384, 256, 384, 384, 256, 256, 384, 256, 384, 384, 256, 256, 384, 256, 256, 256, 256, 256, 256, 256, 256, 384, 256, 256, 256, 256, 384, 256, 256, 384, 384, 384, 384, 256, 256, 256, 256, 384, 256, 256, 256, 256, 384, 384, 384, 256, 256, 384, 384, 384, 256, 256, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 384, 384, 256, 256, 384, 384, 384, 256, 384, 256, 384, 256, 256, 256, 256, 384, 256, 256, 256, 384, 384, 384, 384, 256, 256, 256, 384, 256, 384, 256, 384, 256, 256, 384, 384, 384, 256, 256, 256, 384, 384, 256, 256, 256, 256, 384, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 384, 384, 384, 256, 256, 256, 256, 256, 256, 384, 384, 384, 256, 384, 256, 256, 256, 256, 384, 384, 256, 256, 256, 256, 384, 384, 256, 256, 256, 256, 256, 256, 256, 384, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 384, 256, 384, 384, 256, 256, 256, 384, 384, 256, 384, 256, 384, 384, 384, 256, 256, 384, 384, 256, 256, 384, 256, 256, 256, 384, 384, 256, 256, 256, 384, 384, 384, 256, 256, 256, 384, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 256, 256, 384, 256, 384, 256, 384, 256, 256, 384, 256, 384, 256, 256, 256, 384, 256, 256, 256, 256, 384, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 256, 384, 384, 256, 384, 256, 384, 256, 256, 256, 256, 384, 256, 256, 256, 384, 384, 384, 384, 256, 384, 256, 256, 384, 256, 256, 256, 256, 384, 256, 384, 384, 256, 384, 256, 256, 384, 256, 384, 256, 256, 384, 384, 384, 256, 384, 384, 384, 384, 256, 384, 384, 256, 384, 384, 384, 256, 256, 384, 256, 256, 256, 256, 384, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 384, 256, 384, 384, 384, 256, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 384, 384, 256, 256, 256, 256, 384, 384, 384, 384, 384, 256, 256, 256, 384, 384, 384, 384, 256, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 256, 256, 256, 256, 256, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 256, 384, 384, 256, 384, 256, 384, 384, 384, 384, 384, 256, 256, 256, 256, 384, 384, 256, 256, 384, 256, 256, 256, 384, 384, 384, 256, 256, 384, 256, 384, 256, 384, 256, 256, 384, 256, 384, 256, 384, 256, 384, 256, 256, 384, 384, 256, 256, 256, 256, 384, 384, 384, 384, 384, 256, 256, 256, 256, 384, 256, 384, 384, 256, 256, 384, 384, 256, 256, 256, 384, 256, 256, 384, 256, 256, 256, 384, 256, 384, 256, 384, 256, 384, 384, 256, 256, 384, 256, 256, 256, 256, 256, 384, 256, 384, 256, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 256, 256, 384, 256, 256, 256, 256, 256, 256, 384, 256, 256, 384, 384, 384, 384, 384, 256, 256, 384, 256, 384, 384, 384, 256, 256, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 256, 256, 384, 256, 384, 256, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 256, 256, 256, 256, 384, 256, 256, 256, 384, 384, 256, 384, 384, 256, 256, 256, 256, 256, 384, 256, 256, 256, 384, 256, 256, 256, 256, 384, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 384, 256, 256, 256, 384, 256, 384, 256, 256, 384, 384, 256, 256, 384, 384, 384, 256, 256, 256, 384, 384, 384, 384, 256, 384, 256, 256, 256, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 384, 384, 256, 384, 384, 384, 256, 384, 384, 256, 256, 384, 384, 256, 384, 384, 384, 384, 256, 384, 384, 256, 256, 256, 256, 384, 384, 384, 384, 256, 384, 256, 384, 384, 256, 384, 256, 256, 256, 384, 384, 384, 384, 384, 384, 256, 256, 384, 384, 384, 256, 384, 384, 384, 384, 384, 384, 256, 256, 384, 384, 384, 256, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 384, 256, 256, 384, 256, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 384, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 256, 256, 384, 256, 384, 384, 384, 384, 256, 256, 384, 256, 256, 256, 256, 384, 384, 256, 256, 384, 256, 256, 256, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 256, 384, 384, 256, 384, 256, 256, 384, 384, 384, 384, 256, 256, 256, 384, 256, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 384, 384, 256, 384, 256, 256, 256, 256, 256, 256, 384, 384, 384, 256, 384, 384, 256, 256, 256, 256, 256, 384, 256, 384, 256, 256, 256, 384, 384, 256, 256, 256, 256, 256, 256, 256, 256, 384, 384, 256, 256, 256, 384, 256, 384, 384, 384, 384, 256, 256, 256, 384, 256, 256, 384, 384, 384, 384, 384, 256, 256, 384, 384, 384, 256, 384, 384, 256, 256, 256, 384, 384, 384, 256, 384, 256, 256, 256, 384, 384, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 384, 256, 256, 256, 384, 384, 256, 256, 384, 384, 256, 256, 256, 384, 256, 256, 384, 384, 256, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 384, 256, 384, 256, 256, 256, 384, 256, 384, 384, 384, 384, 256, 256, 256, 256, 256, 384, 256, 384, 384, 256, 384, 256, 384, 384, 256, 256, 256, 256, 256, 384, 256, 256, 384, 256, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 384, 256, 256, 256, 384, 384, 256, 256, 256, 384, 256, 256, 384, 256, 256, 256, 384, 384, 384, 384, 384, 256, 384, 384, 256, 384, 256, 384, 256, 256, 256, 384, 256, 256, 384, 384, 384, 384, 384, 256, 256, 384, 384, 256, 256, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 256, 256, 384, 256, 256, 256, 256, 384, 384, 256, 384, 256, 256, 384, 384, 384, 384, 256, 256, 256, 384, 384, 256, 384, 384, 256, 256, 256, 256, 384, 256, 384, 384, 384, 384, 384, 256, 256, 256, 384, 256, 256, 256, 384, 384, 384, 256, 256, 384, 256, 256, 256, 384, 256, 384, 256, 256, 256, 384, 256, 256, 256, 256, 256, 256, 384, 384, 256, 384, 384, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 384, 384, 384, 256, 256, 384, 384, 256, 256, 256, 384, 384, 256, 384, 256, 256, 384, 384, 256, 256, 384, 384, 256, 384, 256, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 384, 384, 384, 256, 256, 384, 384, 256, 256, 384, 256, 256, 256, 384, 256, 256, 384, 384, 384, 384, 256, 256, 384, 256, 256, 384, 384, 384, 256, 384, 256, 384, 384, 384, 384, 384, 256, 256, 384, 256, 256, 256, 256, 256, 384, 384, 384, 256, 256, 256, 384, 256, 384, 256, 256, 256, 384, 384, 384, 384, 384, 256, 256, 256, 384, 256, 256, 256, 256, 256, 256, 256, 384, 384, 384, 384, 256, 384, 256, 384, 384, 256, 256, 256, 256, 256, 256, 256, 384, 256, 256, 256, 256, 256, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 256, 256, 256, 256, 256, 256, 384, 256, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 256, 256, 384, 384, 384, 384, 384, 384, 384, 256, 384, 384, 384, 384, 256, 256, 384, 384, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 384, 256, 256, 384, 384, 384, 256, 384, 256, 384, 256, 256, 256, 256, 256, 256, 256, 256, 256, 384, 384, 384, 384, 384, 384, 256, 384, 384, 384, 256, 256, 256, 256, 256, 256, 384, 256, 384, 256, 384, 384, 384, 384, 384, 384, 384, 256, 256};

localparam logic [2912:0][31:0] rectangle3_xs = {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 11, 6, 0, 0, 0, 0, 0, 0, 0, 11, 0, 12, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 2, 11, 0, 0, 0, 0, 0, 0, 0, 9, 0, 12, 0, 0, 0, 0, 0, 9, 3, 0, 0, 0, 0, 0, 7, 0, 0, 0, 3, 11, 0, 0, 0, 0, 0, 12, 1, 0, 0, 0, 0, 0, 17, 11, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 12, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 18, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 4, 10, 10, 3, 0, 0, 15, 6, 0, 0, 0, 0, 0, 11, 17, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 8, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 1, 0, 0, 12, 0, 0, 0, 0, 14, 5, 0, 0, 5, 11, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 5, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 11, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 16, 4, 0, 0, 0, 0, 5, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 10, 0, 0, 7, 0, 0, 12, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 7, 0, 0, 0, 0, 0, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 6, 14, 6, 0, 0, 5, 0, 0, 10, 0, 0, 0, 0, 20, 0, 0, 2, 0, 0, 0, 0, 7, 12, 0, 0, 0, 11, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 16, 4, 12, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 12, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 6, 0, 11, 10, 0, 0, 8, 12, 0, 4, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 11, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 1, 0, 9, 10, 4, 0, 16, 0, 8, 0, 10, 0, 5, 0, 0, 7, 0, 0, 10, 10, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 16, 0, 16, 4, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 8, 4, 0, 0, 17, 4, 7, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 4, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 9, 8, 0, 6, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 12, 12, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 11, 5, 12, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 6, 10, 0, 0, 0, 6, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 10, 0, 9, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 9, 0, 9, 0, 10, 0, 9, 11, 11, 0, 6, 10, 16, 11, 8, 10, 3, 5, 0, 0, 0, 12, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 4, 0, 0, 14, 7, 0, 0, 0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 4, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 15, 5, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 14, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 17, 4, 14, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 14, 5, 0, 11, 7, 11, 10, 11, 0, 7, 0, 0, 10, 10, 0, 0, 15, 0, 15, 5, 11, 9, 0, 0, 0, 0, 10, 12, 0, 7, 0, 8, 0, 0, 0, 0, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 9, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 13, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 16, 0, 0, 4, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 2, 7, 17, 0, 0, 0, 15, 4, 0, 5, 0, 0, 0, 0, 0, 0, 0, 10, 11, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 11, 0, 0, 12, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 6, 0, 9, 0, 5, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 7, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 11, 0, 0, 0, 0, 5, 0, 0, 12, 0, 0, 1, 0, 0, 0, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 12, 6, 0, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 14, 0, 0, 7, 12, 0, 0, 0, 0, 0, 0, 0, 9, 12, 0, 0, 0, 0, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 3, 11, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 6, 12, 0, 12, 15, 7, 0, 0, 0, 0, 4, 0, 17, 0, 0, 0, 0, 4, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 5, 12, 0, 0, 0, 12, 0, 0, 0, 0, 0, 12, 0, 5, 0, 11, 7, 12, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 12, 13, 9, 4, 0, 0, 0, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 9, 0, 0, 11, 0, 11, 6, 11, 0, 11, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 12, 11, 11, 5, 0, 0, 9, 6, 0, 0, 0, 0, 0, 13, 12, 7, 12, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 14, 6, 10, 0, 0, 11, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 4, 0, 0, 3, 0, 0, 6, 0, 0, 0, 0, 19, 0, 19, 0, 0, 0, 0, 3, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 11, 0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 10, 0, 12, 9, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 13, 12, 4, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 8, 14, 7, 0, 9, 0, 0, 0, 0, 19, 3, 0, 0, 11, 12, 0, 0, 20, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 20, 2, 0, 0, 0, 0, 7, 0, 0, 0, 7, 0, 0, 0, 7, 9, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 15, 7, 0, 0, 0, 11, 0, 0, 12, 9, 5, 0, 0, 6, 0, 0, 0, 12, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 4, 11, 0, 0, 6, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 13, 3, 10, 12, 0, 0, 6, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 12, 4, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 3, 13, 0, 12, 9, 0, 6, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 15, 5, 11, 9, 0, 0, 2, 0, 10, 11, 0, 12, 0, 0, 13, 0, 8, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 4, 8, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 0, 0, 7, 10, 0, 6, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 10, 8, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 5, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 10, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 19, 3, 0, 0, 12, 0, 12, 7, 14, 5, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 13, 7, 0, 11, 10, 12, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 11, 10, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 6, 3, 7, 16, 4, 13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 0, 0, 18, 3, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9};

localparam logic [2912:0][31:0] rectangle3_ys = {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 15, 0, 11, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 14, 14, 0, 0, 0, 0, 0, 0, 0, 8, 0, 11, 0, 0, 0, 0, 0, 21, 20, 0, 0, 0, 0, 0, 16, 0, 0, 0, 18, 9, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 16, 17, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 10, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 15, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 9, 11, 14, 14, 0, 0, 18, 18, 0, 0, 0, 0, 0, 6, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 13, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 5, 0, 8, 15, 0, 0, 0, 0, 5, 5, 3, 0, 18, 18, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 14, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 14, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 17, 0, 17, 17, 0, 0, 0, 0, 9, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 15, 0, 0, 19, 14, 0, 20, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 9, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 8, 19, 19, 0, 0, 9, 0, 0, 11, 0, 0, 0, 0, 11, 0, 0, 11, 0, 0, 0, 0, 6, 6, 0, 0, 0, 9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 5, 0, 0, 0, 15, 15, 11, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 7, 0, 0, 15, 0, 0, 0, 0, 0, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 11, 0, 0, 0, 15, 0, 15, 15, 0, 0, 7, 9, 0, 6, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 19, 0, 10, 10, 9, 0, 17, 0, 16, 0, 12, 0, 13, 0, 0, 16, 0, 0, 12, 12, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 21, 16, 0, 16, 16, 0, 0, 0, 0, 0, 0, 0, 0, 15, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 7, 6, 0, 0, 17, 17, 13, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 14, 14, 0, 14, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 20, 20, 2, 0, 7, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 11, 12, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 9, 9, 19, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 21, 22, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 5, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 12, 0, 11, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 13, 0, 13, 0, 15, 0, 13, 13, 17, 0, 15, 12, 19, 13, 21, 15, 12, 20, 0, 0, 0, 9, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 14, 14, 0, 0, 0, 0, 19, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 16, 14, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 17, 16, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 8, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 16, 20, 20, 0, 20, 9, 15, 16, 16, 0, 16, 0, 0, 10, 9, 0, 0, 14, 0, 14, 14, 15, 15, 0, 0, 0, 0, 10, 5, 0, 8, 0, 8, 0, 0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 21, 11, 0, 0, 0, 0, 4, 0, 0, 0, 0, 9, 10, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 18, 0, 0, 18, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 12, 15, 6, 0, 0, 0, 18, 6, 0, 18, 0, 0, 0, 0, 0, 0, 0, 5, 21, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 12, 0, 0, 9, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 0, 19, 0, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 9, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 7, 0, 0, 0, 0, 9, 0, 0, 11, 0, 0, 21, 0, 0, 0, 21, 21, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 18, 0, 0, 0, 10, 9, 0, 16, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 9, 0, 0, 9, 11, 0, 0, 0, 0, 0, 0, 0, 9, 8, 0, 0, 0, 0, 0, 0, 16, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 13, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 9, 21, 0, 12, 15, 15, 0, 0, 0, 0, 4, 0, 7, 0, 0, 0, 0, 7, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 11, 2, 0, 0, 0, 8, 0, 0, 0, 0, 0, 18, 0, 17, 0, 12, 12, 12, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 14, 12, 12, 9, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 11, 0, 0, 11, 0, 11, 20, 11, 0, 11, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 15, 11, 11, 12, 0, 0, 4, 11, 0, 0, 0, 0, 0, 8, 15, 16, 7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 19, 19, 21, 0, 0, 9, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 5, 0, 0, 5, 0, 0, 12, 0, 0, 0, 0, 13, 0, 13, 0, 0, 0, 0, 14, 13, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 15, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 9, 0, 0, 0, 0, 0, 0, 0, 13, 0, 10, 0, 0, 14, 15, 0, 0, 0, 0, 0, 0, 0, 20, 0, 16, 16, 18, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 14, 16, 15, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 15, 15, 15, 0, 22, 0, 0, 0, 0, 13, 13, 0, 0, 15, 16, 0, 0, 14, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 14, 14, 0, 0, 0, 0, 12, 0, 0, 0, 11, 0, 0, 0, 11, 11, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 12, 12, 0, 0, 0, 11, 0, 0, 12, 12, 13, 0, 0, 14, 0, 0, 0, 17, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 15, 15, 0, 0, 12, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 19, 7, 6, 6, 0, 0, 11, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 12, 0, 12, 12, 0, 12, 14, 14, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 19, 19, 5, 5, 0, 0, 11, 0, 13, 13, 0, 16, 0, 0, 8, 0, 13, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 9, 11, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 11, 0, 0, 15, 15, 0, 8, 0, 0, 0, 0, 14, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 12, 0, 0, 11, 16, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 9, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 5, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 15, 15, 0, 0, 21, 0, 20, 20, 6, 6, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 19, 19, 0, 14, 10, 9, 13, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 17, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 9, 15, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 8, 22, 10, 14, 14, 17, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 21, 0, 0, 18, 18, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12};

localparam logic [2912:0][31:0] rectangle3_widths = {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 9, 0, 7, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 8, 0, 12, 0, 0, 0, 0, 0, 7, 9, 0, 0, 0, 0, 0, 5, 0, 0, 0, 9, 7, 0, 0, 0, 0, 0, 12, 11, 0, 0, 0, 0, 0, 3, 10, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 3, 11, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 9, 4, 3, 0, 0, 3, 3, 0, 0, 0, 0, 0, 5, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 11, 0, 12, 9, 0, 0, 0, 0, 5, 5, 12, 0, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 0, 6, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 4, 0, 4, 4, 0, 0, 0, 0, 8, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 4, 12, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 7, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 6, 4, 4, 0, 0, 8, 0, 0, 7, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, 0, 0, 6, 12, 0, 0, 0, 9, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 0, 0, 0, 4, 4, 6, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 5, 0, 0, 4, 0, 0, 0, 0, 0, 12, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 11, 0, 0, 0, 8, 0, 3, 8, 0, 0, 4, 6, 0, 4, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 11, 0, 5, 5, 8, 0, 4, 0, 4, 0, 4, 0, 7, 0, 0, 6, 0, 0, 4, 4, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 4, 3, 0, 0, 3, 3, 7, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 7, 7, 0, 3, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 5, 5, 12, 0, 12, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 6, 6, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 6, 7, 7, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 6, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 10, 0, 3, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 4, 0, 4, 0, 2, 0, 4, 4, 3, 0, 6, 9, 4, 11, 6, 10, 10, 5, 0, 0, 0, 11, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 3, 3, 0, 0, 0, 0, 6, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 9, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 4, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 5, 5, 0, 5, 6, 2, 3, 3, 0, 3, 0, 0, 4, 8, 0, 0, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 4, 12, 0, 6, 0, 4, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 0, 0, 0, 0, 12, 0, 0, 0, 0, 7, 4, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 4, 0, 0, 4, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 11, 4, 3, 0, 0, 0, 4, 3, 0, 4, 0, 0, 0, 0, 0, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 11, 0, 0, 6, 6, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 0, 6, 0, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 6, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 4, 0, 0, 0, 0, 8, 0, 0, 12, 0, 0, 11, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 3, 0, 0, 0, 5, 7, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 10, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 6, 10, 0, 9, 2, 2, 0, 0, 0, 0, 8, 0, 3, 0, 0, 0, 0, 3, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 12, 0, 0, 0, 4, 0, 0, 0, 0, 0, 12, 0, 4, 0, 5, 7, 5, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 9, 2, 2, 10, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 5, 0, 0, 2, 0, 2, 5, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 2, 2, 2, 9, 0, 0, 9, 7, 0, 0, 0, 0, 0, 3, 2, 5, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 4, 6, 0, 0, 7, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 4, 0, 0, 9, 0, 0, 6, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, 0, 2, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 0, 0, 0, 0, 0, 0, 0, 6, 0, 6, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 5, 0, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 4, 5, 9, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 0, 9, 0, 0, 0, 0, 2, 2, 0, 0, 2, 5, 0, 0, 2, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 2, 2, 0, 0, 0, 0, 7, 0, 0, 0, 8, 0, 0, 0, 8, 8, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 2, 2, 0, 0, 0, 6, 0, 0, 3, 3, 7, 0, 0, 2, 0, 0, 0, 3, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 5, 3, 3, 5, 0, 0, 9, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 6, 9, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 0, 6, 2, 0, 6, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 4, 4, 4, 0, 0, 10, 0, 4, 8, 0, 5, 0, 0, 5, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 9, 6, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 0, 0, 7, 7, 0, 3, 0, 0, 0, 0, 12, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 6, 4, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 6, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 2, 2, 0, 0, 6, 0, 5, 5, 5, 5, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 6, 4, 6, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 9, 2, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 9, 2, 4, 4, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 0, 0, 3, 3, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3};

localparam logic [2912:0][31:0] rectangle3_heights = {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 6, 0, 5, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 7, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 7, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 8, 2, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 6, 8, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 11, 7, 10, 0, 0, 6, 6, 0, 0, 0, 0, 0, 6, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 0, 8, 2, 0, 0, 0, 0, 5, 5, 2, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 7, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 0, 3, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 7, 0, 7, 7, 0, 0, 0, 0, 4, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 9, 0, 0, 5, 2, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 3, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 3, 5, 5, 0, 0, 3, 0, 0, 6, 0, 0, 0, 0, 9, 0, 0, 9, 0, 0, 0, 0, 6, 3, 0, 0, 0, 4, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 9, 9, 6, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 7, 0, 0, 5, 0, 0, 0, 0, 0, 3, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 6, 0, 0, 0, 3, 0, 7, 3, 0, 0, 5, 3, 0, 6, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 0, 5, 5, 3, 0, 7, 0, 6, 0, 8, 0, 7, 0, 0, 5, 0, 0, 8, 8, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 0, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 6, 6, 0, 0, 7, 7, 7, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 5, 5, 0, 10, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 4, 4, 2, 0, 3, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 6, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 4, 3, 3, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 5, 3, 0, 0, 0, 3, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 2, 0, 6, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 5, 0, 5, 0, 9, 0, 5, 5, 7, 0, 3, 3, 5, 4, 3, 9, 6, 4, 0, 0, 0, 2, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 6, 6, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 2, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 7, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 8, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 4, 4, 0, 4, 3, 9, 7, 7, 0, 8, 0, 0, 9, 4, 0, 0, 10, 0, 10, 10, 7, 7, 0, 0, 0, 0, 8, 3, 0, 6, 0, 5, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 5, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 0, 0, 5, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 7, 5, 6, 0, 0, 0, 5, 6, 0, 5, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 8, 0, 0, 9, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 3, 0, 4, 0, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 5, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 5, 0, 0, 0, 0, 3, 0, 0, 11, 0, 0, 2, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 6, 0, 0, 0, 4, 3, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 6, 0, 0, 6, 3, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 3, 2, 0, 7, 9, 9, 0, 0, 0, 0, 3, 0, 6, 0, 0, 0, 0, 6, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 2, 0, 0, 0, 5, 0, 0, 0, 0, 0, 2, 0, 7, 0, 12, 7, 4, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 2, 11, 11, 2, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 5, 0, 0, 10, 0, 10, 4, 10, 0, 10, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 9, 10, 10, 3, 0, 0, 4, 6, 0, 0, 0, 0, 0, 6, 9, 8, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 5, 3, 0, 0, 3, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 5, 0, 0, 5, 0, 0, 3, 0, 0, 0, 0, 9, 0, 9, 0, 0, 0, 0, 9, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 0, 0, 0, 4, 0, 8, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 4, 0, 6, 6, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 5, 5, 2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 9, 6, 6, 0, 2, 0, 0, 0, 0, 11, 11, 0, 0, 9, 7, 0, 0, 10, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 10, 10, 0, 0, 0, 0, 10, 0, 0, 0, 10, 0, 0, 0, 10, 10, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 11, 11, 0, 0, 0, 3, 0, 0, 6, 6, 4, 0, 0, 9, 0, 0, 0, 7, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 12, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 4, 6, 6, 6, 0, 0, 2, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 9, 0, 3, 9, 0, 3, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 5, 5, 5, 0, 0, 3, 0, 8, 4, 0, 4, 0, 0, 4, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 2, 10, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 7, 7, 0, 6, 0, 0, 0, 0, 5, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 6, 0, 0, 4, 5, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 9, 0, 0, 3, 0, 4, 4, 6, 6, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 3, 5, 5, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 2, 10, 6, 6, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 6, 6, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11};

localparam logic [2912:0][31:0] rectangle3_weights = {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 256, 256, 0, 0, 256, 256, 0, 0, 0, 0, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 0, 256, 256, 0, 0, 0, 0, 256, 256, 256, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 256, 0, 256, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 256, 256, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 256, 256, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 256, 256, 0, 0, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 256, 256, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 256, 0, 0, 0, 256, 0, 256, 256, 0, 0, 256, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 256, 256, 256, 0, 256, 0, 256, 0, 256, 0, 256, 0, 0, 256, 0, 0, 256, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 256, 0, 0, 256, 256, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 256, 0, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 256, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 0, 256, 0, 256, 0, 256, 256, 256, 0, 256, 256, 256, 256, 256, 256, 256, 256, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 256, 256, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 256, 0, 256, 256, 256, 256, 256, 0, 256, 0, 0, 256, 256, 0, 0, 256, 0, 256, 256, 256, 256, 0, 0, 0, 0, 256, 256, 0, 256, 0, 256, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 0, 0, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 256, 256, 0, 0, 0, 256, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 256, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 256, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 256, 256, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 256, 0, 256, 256, 256, 0, 0, 0, 0, 256, 0, 256, 0, 0, 0, 0, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 256, 0, 256, 256, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 256, 256, 256, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 0, 256, 0, 256, 256, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 256, 256, 256, 0, 0, 256, 256, 0, 0, 0, 0, 0, 256, 256, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 256, 0, 0, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 256, 0, 256, 0, 0, 0, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 256, 0, 0, 0, 0, 256, 256, 0, 0, 256, 256, 0, 0, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 256, 0, 0, 0, 0, 256, 0, 0, 0, 256, 0, 0, 0, 256, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 256, 0, 0, 0, 256, 0, 0, 256, 256, 256, 0, 0, 256, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 256, 256, 256, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 256, 256, 0, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 256, 256, 0, 0, 256, 0, 256, 256, 0, 256, 0, 0, 256, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 256, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 256, 256, 0, 256, 0, 0, 0, 0, 256, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 256, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 0, 0, 256, 0, 256, 256, 256, 256, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 256, 256, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 256, 256, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 256, 256, 256, 256, 256, 256, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 256, 0, 0, 256, 256, 0, 256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256};

localparam logic [2912:0][31:0] feature_threshold = {-4, 2, 3, 1, 2, 13, 0, -2, 1, -3, 3, 3, 12, 5, -2, 1, 2, -1, -1, 2, -3, -18, 2, 1, 12, 9, 4, 2, 2, 0, 4, -1, 6, 6, -9, -6, 11, 0, 15, -7, -5, 48, 2, 2, 5, -1, 0, 4, -10, 0, 3, -6, -8, 2, 19, 1, 1, 2, 3, -36, 1, -5, 2, -1, 4, -5, -1, -8, -5, 0, -17, 3, -4, 3, 3, -1, 6, 7, 0, 2, -3, -1, -2, -9, 5, 24, 10, 0, 11, 1, 1, -3, 1, 4, 0, 4, -1, -1, -3, 0, -2, -1, 10, 4, 3, -4, -4, 3, 1, -5, -2, -3, -3, 2, -2, -4, 2, 0, 11, 33, -5, -2, 0, -1, 0, -6, -3, -10, 3, 0, 15, 0, 9, -6, -6, 4, 12, 2, 2, 0, 4, 0, -2, 3, 4, -6, -9, 8, 1, 5, 0, -4, -2, 5, 3, 7, -2, -23, 23, -1, 8, -4, -6, 5, -3, -8, -4, 1, 0, 3, -1, 2, -6, 3, 0, 2, -4, 9, 30, -2, 1, 2, -1, 1, 1, 2, 0, -14, 1, 4, 4, 1, 3, 2, 3, -2, -5, -1, 0, -4, 8, 1, 1, 0, 1, 1, 4, 3, 1, 4, 0, -5, -5, 0, -7, -1, 4, -14, -1, -1, -1, -2, -3, 2, -3, -5, -8, 3, 0, 6, 7, -1, -2, 3, -3, 2, -1, -1, 16, 6, 7, -5, -9, 17, -27, -8, 8, -3, -4, -2, 2, 6, 2, 2, 6, 2, -2, 5, -7, -9, 2, -1, -5, 0, -3, 0, 0, 5, 8, 0, 0, -1, -3, -13, -1, 5, -2, -6, 3, -1, 5, 0, 1, 1, -7, -29, -2, -2, -5, -1, -2, 4, 3, 1, -3, -1, -5, -3, 0, -3, -4, -2, -8, -2, -3, -4, -3, 0, -4, 2, 1, -1, 0, -1, -6, -8, -4, -19, -2, 19, 7, 0, -6, 17, -12, 2, 4, 2, 2, -4, 18, -1, 2, 3, 6, -1, 5, -4, -5, 0, 4, 4, 1, 0, 5, 3, -2, -1, 3, 8, 5, 3, -4, 1, 3, -2, 6, 0, -11, 2, 5, -26, -2, 5, 0, -2, -6, -4, -6, -4, -1, -1, 1, 7, 4, -2, -4, -10, 0, 12, 5, 7, -3, 42, 1, 21, -1, -2, 10, 2, -10, -9, -1, 4, -4, -10, 0, 4, 1, 13, -1, 1, 3, 36, -6, -2, 18, 4, 2, 3, 7, 2, 1, 4, -6, 2, 1, -6, 11, -1, 5, -1, -1, 1, 12, -4, -8, -5, -1, 6, -5, -3, 0, -4, 2, 0, 0, -12, -10, 2, -3, -2, 1, 13, -5, 3, 0, -37, 12, 15, -9, -4, -6, 23, -2, 1, 1, -3, -9, -8, 3, -2, -1, -5, -5, -2, -3, -11, -1, -5, 6, -18, -8, 1, 0, 35, -3, 5, 1, 4, -5, -12, -1, 2, -4, -3, 6, -3, -3, 8, 2, -2, -3, -3, 5, -1, -4, 5, 3, 26, 2, 5, -4, -5, -8, -2, 9, -3, -3, 0, 5, 4, 1, -1, -4, -1, -7, 1, 4, -4, 6, -1, 8, -6, 2, 4, -3, 4, 7, -4, 3, -3, 4, -1, -1, 0, -5, -4, 1, -12, 3, 0, 4, 2, 0, -6, -6, -14, -16, -6, -6, -16, -3, -2, -6, 7, -1, 2, 1, 1, 1, 1, -4, -5, -4, 0, 24, 1, 3, -3, 1, 7, 0, 2, 2, 4, 1, 18, 2, -2, -1, -2, -13, -1, 6, -15, 1, 3, -2, 7, -1, 1, -2, -3, 2, -2, 4, 12, 3, 2, 0, -1, 3, -5, -1, -3, -3, 2, 12, -4, -2, 0, 2, -2, -1, -3, -2, -5, -1, -2, -6, -8, 0, 3, 3, 3, -4, 0, 7, -12, 2, 29, -23, -9, 2, 1, -2, 2, 2, -5, 2, -3, -3, -1, 2, -4, -4, -2, 5, -2, 0, 2, 4, 0, 11, -8, 6, 5, 5, 8, -3, -21, 9, 1, 0, 10, -7, 1, -2, 12, 1, 1, 4, -7, -9, -1, 9, -9, -3, 3, -6, 24, -6, 3, 1, 3, -12, -2, 2, 4, 1, -7, -2, 3, 6, 2, 21, 2, -2, 10, 5, 4, 2, 6, 4, 5, -2, 2, 1, 4, 0, 6, 4, 4, 1, -1, 2, 1, 0, -2, 4, 1, 1, 3, -3, 0, 1, 3, -7, -8, -4, -5, 16, -1, -8, 1, -2, 2, 1, -1, 27, -3, 8, -1, 6, -3, -1, 0, 6, 0, -4, 11, -17, -1, -2, -3, -7, -11, -7, -1, 7, -9, -3, 1, 3, -3, -3, -7, 1, -3, -11, 17, 2, 1, -6, 7, -1, -7, 6, 1, 3, -2, -5, 0, 3, 1, 4, -1, 7, -3, -2, 2, 4, 4, 0, -6, 10, 3, 0, -11, -2, -1, 12, 70, 5, 3, 7, -2, -16, 0, 15, 5, 1, -3, -4, -1, -7, -2, -1, -6, 8, -2, 6, 0, 6, 4, 4, -1, 2, 0, -7, -2, -7, 7, -3, 0, -5, -3, 4, 15, -3, 2, 0, 0, 0, 5, -2, 0, -5, -4, 3, 4, -2, 2, 0, 13, 0, 1, -5, -3, 2, -1, 3, -3, 0, -5, 4, 6, 5, 6, -2, 10, 13, -2, -2, -2, -3, 1, -3, 1, -2, 3, 11, 3, -5, -10, -2, 15, 20, -6, -1, 12, 2, 0, 4, -4, 0, -8, 0, 3, -7, 1, 2, -1, 5, -51, -3, -2, -2, 3, 2, -3, 8, 14, -4, 0, -1, -1, 3, 1, -6, 0, 15, 2, 7, -1, 16, -1, 2, -6, -4, -3, -2, -2, 0, -6, 5, 1, -2, 1, 6, 1, 0, 1, -6, -3, 4, 6, 0, -3, 2, 2, 8, -5, -11, 6, 3, -1, 3, -11, 3, -2, 4, 0, 7, -14, -1, 10, -12, 6, -2, 11, 10, -4, 2, 7, 3, 1, -5, 20, -9, -4, -8, 1, -1, -17, 7, -1, 4, 5, -4, -2, -1, 1, -6, 3, 4, -9, 4, 0, 0, 4, -2, 5, 0, -5, -3, 1, -3, 3, -5, -1, 7, 3, 0, 2, 14, 5, -1, 3, -4, 3, 1, 1, 3, 10, 1, 0, 0, 4, -4, 3, -3, 1, 2, 4, 1, -1, -1, -3, -5, -2, 1, -1, 3, -3, -9, -3, -6, -14, 2, -1, -1, -5, 1, -4, 7, -5, -3, -1, 2, 1, -3, 1, 5, 2, -3, 1, 1, -1, -1, 13, 7, 2, -4, -7, -1, 4, 0, 1, 10, 7, -3, 1, -4, 5, 2, -6, -3, 2, 13, -2, 5, 3, -4, 1, -6, -5, 6, 7, 2, -12, 1, 5, 6, -2, -5, -5, 3, 1, -17, 1, 1, -8, 0, 0, 3, 1, 3, -5, 3, 2, -3, -2, 58, 2, -3, -6, -2, -3, 3, -3, 0, 2, -3, 0, 0, -4, -1, 4, -4, 2, -4, 1, 8, -8, -12, -5, 3, -3, -5, -2, 1, -1, -1, 0, -4, -2, -1, -4, 2, -2, -11, 1, -4, 0, -14, 2, 1, -3, -2, -1, 9, -2, 0, -7, -1, 27, 2, 5, 3, -4, 8, 3, -10, 2, -9, 17, -6, -4, 0, -3, 0, 2, 3, -6, -3, 3, 24, -10, -6, -2, 0, -13, -3, 8, -3, 4, 5, -3, 3, -3, -3, 0, 14, 6, 6, 0, 9, 5, -3, 54, 1, -2, -2, -2, 0, 12, -2, -3, -3, -2, 4, 7, 1, -2, 29, 14, 0, 11, 3, -2, 42, 1, 6, -5, -10, 28, 2, 7, 1, 1, -3, 0, 7, -1, -5, -3, -2, -3, 7, 0, 1, -7, -2, -4, -38, -5, -7, 4, -1, -1, 0, 7, -16, 12, 5, 0, 1, 3, -2, -1, -1, 3, -2, 2, -6, 1, 1, 2, 12, 6, 1, -5, 3, 1, 8, 1, 2, -6, 7, 3, 5, -3, -11, 1, 10, -12, -4, 1, -1, 3, -2, 3, -2, 4, -1, 3, -4, 0, 4, 1, 4, 1, 6, -4, 3, 3, 1, -7, 4, -4, 2, -6, 11, 3, 2, -2, 0, 2, -1, -2, -13, -12, -5, 0, 14, 0, 4, 1, -2, -2, 3, 6, -3, 5, 3, -3, 10, -2, -3, -9, -1, 3, -5, 3, 6, 5, 10, 4, 1, -8, -9, -15, 0, -6, 7, -4, 3, -18, 7, 3, -2, -3, -3, 2, 7, 2, -3, 0, -1, 12, -8, 2, -3, -1, -1, -4, -3, -5, 1, 21, 12, 5, 2, 18, 2, -1, -1, 0, 4, -2, 0, 0, 0, 1, 2, -7, 12, 3, 0, -4, -3, 3, -4, -3, -2, -8, -6, -3, -1, 1, -3, -2, -2, 4, 5, -3, -8, -1, 0, -3, -2, -3, 20, 9, -1, -2, -4, 3, 12, 4, 0, -5, -3, -2, 4, -4, -1, -3, -2, -5, 4, 1, 2, 6, 0, 3, -2, 5, -10, -2, 4, -15, 15, 1, -9, 23, 1, -2, 2, 3, 8, -4, -3, 2, 4, -1, -2, -2, 9, 1, -5, 1, 22, 15, -3, -7, 29, 1, -15, 5, 3, -5, -17, -5, -4, 2, -5, -9, -3, 5, 13, -10, -3, -1, 0, 0, 2, -3, -1, 0, -6, 1, 4, -1, -3, -4, 6, 6, 3, 1, 12, 22, -6, 14, -2, 4, 3, 3, 11, 11, -7, -8, -3, 7, 0, 13, -1, 6, -1, 2, 3, -4, 0, 0, 1, 8, -4, 6, -4, 16, 1, 4, 3, 1, -2, 0, 5, -6, 4, -5, -5, 2, -3, -3, 2, -6, -1, 6, -2, 0, 0, -4, -1, -4, 1, 1, 12, -4, -2, 2, 2, -10, -2, 3, 0, -6, -1, -1, 1, 3, 3, -7, 3, 3, -2, -6, -9, 1, -4, -2, -6, 7, 5, 0, -4, 13, -5, -6, -15, -15, 9, 1, 3, 0, 4, -1, 3, 2, -1, -5, -12, -3, -3, -1, 9, 4, -6, -3, -2, -6, -3, -4, -1, -6, 2, 0, 3, -10, 6, -16, 2, 2, 5, 2, 2, 1, 5, -1, 4, -3, 3, 0, -5, 1, 6, 0, -1, -1, 0, -11, 6, 0, -2, 6, -4, -4, 1, 0, 14, 9, 0, 25, 20, -6, 7, 6, -5, -5, -5, 2, 0, 4, -1, 1, 12, 2, 1, -2, -1, 4, -2, -2, -5, 4, 8, 1, -5, 0, 1, 11, -4, -3, 5, 0, -1, 17, -2, -10, -2, -7, 0, 3, -3, -1, -5, 28, -2, 9, 7, 5, 8, 1, 8, -5, -1, 14, 2, 4, -3, -1, -1, -2, 2, 1, 2, 4, 3, 1, -7, 9, -3, -2, -5, 3, -1, 3, -9, 6, 1, 2, -1, -14, 6, -3, 2, 6, -4, 5, 24, -1, 1, -1, -1, 1, -3, 0, 0, 1, -3, 10, 2, -3, 4, 2, 11, -5, 0, -7, 3, -3, 1, 44, 1, 4, 0, 0, 7, -1, -2, -1, -1, -6, 2, 0, 0, 1, -1, 7, 2, 22, 7, -41, -3, 10, 3, 1, 4, -6, -7, 2, -6, -8, 1, 4, 8, 1, 0, 4, 4, 6, -3, -7, -3, 14, -5, 2, 3, 6, 5, 5, 2, -2, 0, -18, -1, -3, -18, -11, 0, -1, -2, -7, 2, 2, 0, -11, 4, -1, -3, 1, -4, -25, -14, -2, 0, 8, -7, -5, 11, -1, 1, 1, -2, 0, -9, -1, 0, -5, -4, -10, 5, -4, 6, 33, 0, -11, -1, -17, 5, 13, -2, -8, 3, 3, 2, 3, -5, -1, 2, -4, -2, 3, -13, -2, -2, -2, -16, 2, 4, 1, 1, 5, -10, -9, 8, 3, -10, -2, 1, -3, 0, -2, 1, 7, -14, 3, 0, 0, -3, 11, -1, 10, 1, -1, 4, -3, -7, -5, -1, 2, -5, -3, -3, -6, -3, 2, -4, 9, 0, -1, -2, -2, -1, 2, -6, -3, -3, 1, 3, 2, -1, -3, -8, -6, 1, -7, 41, 10, -2, 6, 1, -4, -4, 0, -2, -1, -7, 0, 2, 2, 2, -2, 0, -2, -2, 2, -1, -1, 1, 3, 4, -2, 3, 53, -5, -1, 2, -1, 2, -1, -2, -6, 6, -5, 0, -6, -1, -6, 13, -2, 1, -2, 9, -2, -1, -7, 0, -6, -15, -2, -1, 7, 9, -2, -2, -5, -2, -1, -16, 6, 4, 1, -8, 0, -9, 13, 2, -1, -1, -8, 5, -5, 6, 6, 8, -8, 4, 0, -1, 6, 2, 6, 25, 2, 0, 3, -2, -1, -2, 6, 3, -2, -22, -15, -10, -2, -8, 1, 5, -5, -1, -3, 0, 2, 2, -8, 7, 3, -2, -13, 15, -2, -4, 2, -15, 0, 4, 3, -4, 5, -9, -5, 6, 8, 2, -4, -2, 9, 0, 2, 0, -1, 6, -4, 13, 0, 5, 0, 3, -1, 0, -2, -4, 0, -7, -8, 4, 4, -3, 2, 6, 24, 4, 2, -1, -1, 2, 3, -3, -2, 1, 0, -6, 7, 1, -7, 7, -2, 1, -3, -8, 0, 5, -2, -5, 13, 11, 5, 8, 19, 0, -4, 1, 6, -9, -40, 4, 1, -4, -1, 4, -4, 3, 2, -5, 1, -9, -1, -2, -2, -1, -7, 4, -1, -1, 10, -1, 4, 5, 2, -6, -2, -2, -5, 4, -1, 2, 9, 68, -2, 0, 6, -6, -12, 5, -2, -2, -7, -1, -9, -3, 2, -6, 6, 2, -12, 9, 7, -2, 3, 2, -7, -2, 1, 4, -3, 1, 11, -1, 1, -1, 1, 0, 5, -1, 4, -1, 11, 1, -2, -3, 14, -1, -7, 13, 3, -2, -41, 26, -9, 5, -9, 8, 5, 1, -6, -9, -5, 0, 2, 1, -4, 12, 0, 2, -18, -12, -1, 2, 9, -5, 66, -4, -5, 1, -2, 1, -18, 23, 1, 14, -4, -3, 0, -4, 2, 2, -2, -2, -4, -13, 5, -37, 20, 0, -3, 5, 7, 1, -7, 3, 3, 5, -13, 11, 2, 4, -8, 9, -4, -2, 3, 13, 3, 4, 5, -6, -5, 0, 5, 3, 0, -1, 2, 5, -9, -8, 4, 5, -4, -4, 0, -9, -10, 1, -5, -8, 2, -7, -6, 2, -3, -5, -5, -2, 0, -1, 5, 0, -3, 3, -2, 1, -1, 7, 7, -2, 12, -2, 4, 4, 2, -6, -1, -8, -9, 2, -1, 1, 0, 26, -2, -2, -3, -3, -3, 6, -6, 3, -6, -2, 2, 0, -6, -2, -2, -29, -16, 1, 1, 37, -30, 8, 1, -4, -2, -6, -10, 4, -12, -2, -1, 0, -1, -5, 4, -1, 0, 5, -3, 0, -2, 85, 14, 2, -3, -10, -7, -3, -6, -2, 3, 4, 3, -3, 8, 19, 7, 1, 0, -4, 3, 0, -2, -11, -2, -2, 2, -2, 2, -1, -3, -4, 1, -1, 2, 5, -7, -7, 0, 38, -11, -7, 5, -1, 0, -9, 1, -1, 2, 3, -2, -9, -2, 3, 2, -3, 1, 29, -5, -2, 5, 1, 12, -5, 1, 10, 4, -4, -1, 1, 14, -15, -5, -4, -16, 30, -4, 5, 9, 1, 7, -6, -5, -13, -16, -15, 4, 1, 7, 0, -4, -20, 1, 6, 3, 9, 1, -7, 14, 3, 4, 5, -1, 0, 3, -4, 10, -2, -2, -3, 3, 19, 0, 1, -1, -5, 3, -4, -2, -2, 1, -2, 2, -4, 0, 0, 6, -1, -6, 3, -3, 6, 8, -5, 0, 3, -2, -1, -2, -1, -16, -11, 8, -4, -10, -2, -1, -2, 0, 4, 4, 4, -2, -11, 1, 7, -1, -2, 7, -3, -9, -2, 4, 7, 5, -16, 0, 1, 6, -10, 1, -2, 4, -4, -9, -2, 6, 4, -4, 5, -3, 8, 4, 5, -3, -3, -1, -7, -3, 1, 4, -3, -1, 3, 4, 2, 14, -2, 1, -1, -11, 0, 47, 28, -2, -6, 2, -4, -1, 17, 4, 6, 0, -3, -4, 2, 0, 0, -4, -4, 20, 11, 0, 1, 5, 10, 0, -1, 15, -1, -4, 3, 6, -3, 3, 1, -30, -3, -1, 1, -5, -2, -16, 9, 11, 2, 10, 2, -11, 9, -10, 12, -5, -1, 0, 2, -3, 7, 0, -2, 4, 0, 11, -5, 10, 5, 3, -9, 6, 10, 8, 4, 2, 3, 4, -2, -1, -4, -1, 41, -2, -1, -4, -1, 1, 1, 25, 1, -9, -4, 1, 12, -8, -22, 1, -5, 16, 11, 11, 7, 1, 2, 7, -3, 6, 3, 1, -4, 4, 0, -12, 2, 3, 0, -1, 2, 0, -10, 6, 0, 2, 5, -2, 7, 1, 6, 3, 20, -1, 0, -3, -1, -4, -3, 0, -1, -2, -1, -1, -5, 1, -1, 1, -1, 6, 2, 21, 0, 0, -3, -2, 2, 7, -5, -4, -5, -4, -11, 54, 8, -2, -1, -7, -2, 6, 0, -11, -3, 6, 0, 1, -2, 1, 3, -3, 8, -10, 1, -3, -5, 1, -2, 1, -9, 1, 14, 5, -14, -15, 2, -1, -4, 2, -5, 3, -3, -2, -15, -11, -3, -1, 1, -4, 1, 2, -2, 36, -30, -14, 16, -8, 2, 0, 4, -6, 1, 3, -3, 4, 2, 1, 5, -2, 7, 1, -3, -1, 4, 3, -1, 4, 1, -11, -2, 0, -2, -10, -30, -13, 0, 3, -14, 2, 9, 2, 1, 1, 1, 0, 0, -4, 2, -8, -3, 4, 2, 0, -5, 2, 10, -30, 18, 1, -7, -7, -3, 3, -2, 0, 1, -1, 1, 3, -1, 1, -4, 6, -5, 5, -9, 5, -5, -3, -20, 1, 3, 10, 0, -2, -4, 6, 0, 6, 14, -5, 4, -7, 2, 9, -2, -1, 0, 2, -5, 3, 7, -2, 0, 10, -3};

localparam logic [2912:0][31:0] feature_above = {-284, 170, 136, 151, 161, -240, 56, 57, 109, -201, 151, 90, 221, -279, 58, 69, 119, -85, -38, 174, -25, -68, 146, 99, -194, 188, 128, -204, 106, 54, 135, -172, 186, 155, -59, 20, -200, 30, 164, -39, -7, 197, 120, 123, -379, -56, 51, -339, 36, 30, 138, 13, -137, 98, 177, 66, 75, 150, 122, -18, 35, 30, -172, -115, -209, 23, -49, 32, -38, 81, 7, 50, 13, -161, -305, -35, -146, -162, 35, 91, 5, -6, -45, 27, 139, 180, 95, 48, 162, 59, -123, 6, 69, -191, -67, -205, 20, -92, 9, 87, 10, -28, 168, 156, 109, 38, -42, -107, -86, 18, 10, 25, 9, 100, 16, 2, 68, 50, -271, 126, 12, -19, -74, -22, -82, 32, -35, 30, -162, 39, 68, 31, 66, -2, -33, -76, 134, 71, 82, 68, 46, 46, -64, 109, 146, -23, -40, 134, 25, -170, -90, 29, -66, 79, 61, -88, 15, -7, 106, -23, -198, 31, -41, -106, 7, 17, 5, 63, -73, 82, 8, -128, 5, -133, -69, 57, 0, -83, 103, 27, -135, -110, 8, 81, 72, -193, 48, 16, 87, 122, 63, 64, -160, 76, 39, 29, -13, 24, -60, -34, 53, 76, -59, 18, -125, 23, -170, -268, 66, -164, -59, 6, 44, 55, 21, -60, -214, 5, 30, 13, -24, -49, 25, 65, 30, -41, -2, 133, -107, 58, -192, -49, -14, -215, 31, 60, 23, 9, -198, 48, -159, 7, 29, 157, -6, -28, -243, 1, -11, 8, -98, 105, 38, 74, 115, 65, -90, 91, 34, -49, 33, -75, 22, -112, 30, -72, 49, -178, -137, 25, 56, -57, 29, -1, -67, -193, 24, 0, -284, 8, -152, 16, 91, -135, 25, -32, -27, -36, 31, 7, 25, 135, -220, 8, 4, -62, 21, 5, 41, -34, 19, 5, 20, -54, 24, 0, 40, -83, 20, 196, 83, 5, -13, -44, -2, -4, 21, 0, -23, -164, -194, 42, 19, 142, -79, 51, 37, 58, -87, 8, -221, 16, -104, 86, 108, -61, 121, -40, 23, 32, -55, -205, 48, 32, -185, -174, 35, -104, -96, 104, 110, -127, 20, -90, -52, 9, -92, 34, 19, -138, 156, 2, -20, 90, 43, 10, 6, -31, 16, -3, -15, -34, -83, -159, 130, -46, 26, -3, -38, 139, 156, -136, 22, 66, 32, -296, -42, 9, -221, 130, 19, -37, -43, -300, 20, -4, 30, 118, 40, -347, -4, 29, -134, 98, 36, -33, 140, 68, 52, 95, 94, 49, 47, 102, -42, -124, -136, 17, 77, -27, -188, 26, 13, -51, -206, -17, 1, 33, -92, -211, 3, -13, -69, 26, -129, -35, -68, 27, -5, -91, 2, -8, 102, -88, -28, 160, 19, -2, 138, 146, -1, 31, -26, -156, 7, 37, -86, 2, 3, 4, 76, 34, -43, 20, -3, -6, -57, 18, -49, 8, 102, 15, -1, 52, -49, 98, -29, -186, 33, 62, -28, 19, -26, 35, -24, 20, -210, 31, -1, -58, 56, 32, 3, 0, 195, -28, 3, 82, 74, 168, 37, 68, -57, -35, 26, 9, -67, 6, 24, -88, -108, -175, 33, 8, -2, -42, 26, 29, -137, 5, -92, -68, 125, -30, 59, -341, 3, -278, 96, 1, 127, -32, -78, 4, -17, -67, 19, 0, -79, -27, 61, 14, -192, 104, -9, 6, -1, -24, 12, -35, 20, -30, 25, 3, -2, -222, -7, -99, 86, 40, 33, 53, 2, -27, 5, 22, 105, 3, -44, 0, 32, -183, 43, 17, -40, 91, 25, -114, -35, 3, -22, -26, 15, -58, 50, -26, 26, -131, -12, -247, -9, 24, 28, -24, 48, -34, 74, 129, 72, 40, -143, 42, 67, -4, 15, 27, -36, -90, 94, 20, -44, -17, -123, -60, -67, 28, 8, 28, 6, 22, -28, 23, 7, 67, 72, -90, 6, 33, 74, 25, 27, 99, -32, -5, 141, 92, 6, -48, 143, 25, -149, 21, -2, -11, 76, 17, -4, 2, 68, 21, -96, -84, -157, 55, -153, 18, 69, 72, -102, 190, -4, 4, 38, -49, -68, 269, -5, 46, -23, -166, 18, 50, -92, 8, -21, -21, 94, 26, -38, 52, -22, 89, 0, 69, -96, 43, -5, 2, 93, -63, 99, 9, -24, -205, 152, 50, -206, 69, -41, -132, -101, -107, -80, 201, 49, 67, -36, -39, -112, -26, 10, 73, 57, 87, 25, -91, 15, 26, 47, 16, 74, -67, 61, -199, 24, -57, -27, 67, 4, -29, 19, 2, -126, 3, 25, 49, -19, -36, 77, -48, 132, -29, -152, 6, 137, -22, -9, 51, -156, -91, 23, -198, 21, -2, 30, 7, -2, -27, 24, -51, -329, -2, 21, 42, -62, -29, 24, -27, -77, -3, 8, -197, 48, 18, -2, -157, 0, -2, -159, 66, -91, 0, 19, -60, -53, 56, -122, -39, -253, -1, -4, 50, 75, -121, 27, -4, 149, -143, 27, -20, 23, 6, -96, -214, 98, -113, -315, -38, 21, -48, 76, 71, 52, -30, 20, -44, 12, 4, -7, -3, 117, -37, 68, -57, -328, -142, 73, 16, 112, 27, 7, -1, 22, -178, 0, -53, 2, -25, 66, 90, -86, 46, 24, 34, 34, -138, -36, 31, -32, 1, 91, -184, 6, -57, 44, -172, -66, -93, -3, 25, -112, -31, -160, -11, -62, 23, 80, 118, 99, -139, -30, 79, 129, 6, 1, 2, -37, -21, -1, -38, -4, -91, -194, -50, -3, 19, -53, 53, 71, 2, -38, -59, -66, 27, 184, -5, 17, 14, 29, 48, -25, 75, -86, -10, 149, 6, -28, 26, 5, 46, 25, 31, 163, -276, -21, 27, -25, 28, -128, 63, -22, -96, 70, -65, -123, 22, -168, 2, 31, 20, -2, 8, -6, 20, 7, 1, -171, 48, -19, 33, -134, 51, 4, 48, -27, 23, -83, -127, 4, 0, 60, 73, -244, -1, -7, -157, -139, -47, 30, 20, -243, 3, 78, 24, 275, 17, -66, 158, -4, 206, -1, 122, 248, -89, 39, 73, 74, 55, -26, 141, 7, -43, 29, 8, 24, -33, 91, 10, 116, 93, 27, -2, -15, -98, 5, 76, 42, -33, -72, -67, 38, 32, -60, -145, -34, -2, 20, -90, 30, 58, 18, -33, -227, 69, 43, -149, -319, 123, -33, -129, 25, -128, 53, 50, -46, 119, 43, 12, 31, -161, 22, -112, 17, 28, -65, 59, 71, 2, -22, 1, 14, -24, 105, -44, -178, 0, 15, -3, 15, -27, 68, -40, -7, -2, 54, 5, 81, 1, -8, 11, -51, 66, 18, 80, -349, -138, 4, 56, -31, -39, 33, -251, 95, 34, 22, -33, -37, -226, -3, 132, -160, -220, 26, 26, 26, 214, -45, -23, 16, -148, -599, -19, 44, 39, 3, 28, 20, -1, -88, 156, -53, -2, 25, -54, 100, -4, 8, -24, -101, 75, -38, 53, 22, 3, -53, 46, 110, 13, -89, 5, -89, -124, 0, -42, 93, 39, -13, -28, -20, -3, -49, -35, 34, 71, 4, 8, -27, 8, 36, -113, 20, 54, 20, 16, 105, -22, 19, -4, -89, -3, 19, 5, 103, -32, 25, 17, 24, -45, 27, -2, -58, 2, 4, 35, 22, 9, 15, 142, 59, -24, 18, 1, -141, 0, 45, -4, -19, -317, -56, 90, 79, -3, -138, -91, 4, 22, 2, 144, 22, -23, -31, 0, 33, 33, 75, -28, 20, -145, 159, -24, 16, 1, -15, -7, -5, -138, 0, -108, -102, -27, 55, 0, 29, -49, -102, 52, 102, 15, 160, 99, 20, -236, -20, 0, 22, 1, 32, -235, -49, 3, -2, -36, -180, 102, -11, -28, -165, 70, -21, 68, -22, 5, -132, 41, -209, -26, -86, 116, -164, 97, 29, 40, -49, 35, -155, -40, -26, 26, 5, 20, 151, 42, 53, 23, -57, -14, -5, -6, -26, -145, 2, 29, 5, -143, -19, -507, -126, -96, 39, 67, -1, 30, 10, -86, -27, -134, 0, 79, -109, -65, -163, 348, 20, 18, 44, 62, -257, -14, -149, 18, 79, -96, 128, -4, -24, 37, 76, 23, -27, 77, -3, 73, -35, 32, -26, -97, -33, -37, 4, -34, -147, 38, -170, 90, -58, -8, 56, 90, 31, 15, -140, 10, 15, 21, -109, 54, -83, 20, -44, 101, -29, -1, -8, 26, -29, 32, 93, 37, -143, 85, -34, 24, -141, -375, -35, -80, -47, 25, -249, 24, -20, 14, 3, 126, -6, -151, -120, -192, 200, -87, 14, 4, -22, 17, -67, 17, 62, 1, 69, -3, 64, -28, 2, 9, -1, -37, -286, 52, -26, 35, 11, -140, -19, -54, -26, 4, -28, 18, -2, 16, -81, -60, 250, -271, 63, 98, 51, -81, -74, -88, 35, 31, 35, 15, 31, -85, 54, -24, -117, 50, 57, 0, 22, -103, 23, -27, 28, -24, 19, -30, 28, -77, 20, 2, -12, -179, -63, -2, 0, -38, 26, 6, 19, -34, 133, -151, -7, -31, 22, -137, -171, 58, -48, 2, 30, -41, -131, -22, 31, -27, 22, -4, 129, -77, 48, -92, 41, -99, -8, 74, 16, -7, -81, -23, -272, 11, 2, -141, -49, -22, -49, 45, -117, -3, 0, 44, 45, 5, -7, -41, 1280, 43, 23, 21, -197, -128, 2, -26, 139, 25, 9, -108, 47, -35, 14, -30, 22, -107, -22, -19, 2, -97, 98, -1, 28, -46, 33, 4, -86, -19, 27, 6, 17, 51, -91, -37, 0, -1, -151, -238, 50, -142, 126, -89, 9, -320, 19, -274, 100, -92, -175, 93, 25, -5, 0, -233, 27, -181, -15, 33, 22, -78, 39, -29, 27, 9, 67, -63, 10, 64, -75, 77, 28, 78, 65, 53, 12, 30, 23, 5, -105, 29, -25, 103, 3, -10, 54, 20, 1, -116, -33, 34, 13, 29, -34, 18, -93, 66, -139, 19, 4, 32, 60, 17, -31, -79, 4, 22, -35, 31, 18, -31, -121, 12, -110, 49, 4, 6, -31, 32, -30, -26, -5, 77, 115, -35, 3, 82, -30, 4, 4, 21, -254, 49, -118, 29, 69, -16, 41, -78, -4, 4, -6, 1, -19, 22, 61, -45, -5, 20, -26, 11, -1, 18, 1, 19, -58, 36, 86, 12, 43, 18, -87, 69, 101, -61, -78, 53, 95, -17, 79, 19, -140, 29, 7, -27, 79, 32, 5, 0, -43, 1, 62, -22, 1, 41, -22, -1, 61, -34, -131, 73, -54, 369, 267, 18, 69, -200, -19, 17, -7, 74, 3, 48, -29, -52, -217, -59, 20, 4, -24, -61, -34, 7, -17, -87, -94, 39, -4, 42, 56, -609, -8, -4, -98, -11, -3, -285, -31, 16, -25, 18, 4, -18, -6, -9, -5, 105, -24, 78, 56, 70, 59, -126, 91, -28, 32, -138, 66, -159, 26, -45, 26, 3, 70, 34, -131, -112, 103, 29, 18, -245, -42, 0, 21, 107, -9, -148, 19, 65, 37, -114, -6, -3, 124, -22, 35, -228, -3, -90, 42, -39, 74, 6, 24, -88, 20, -77, 48, 66, 18, 151, 117, -7, -128, -1, -216, -20, -24, -2, -33, -40, 54, 119, 52, -127, 33, 15, -132, 4, 0, -44, 19, 4, 24, 10, 29, 8, 28, -56, 49, 51, -34, -9, 20, 99, -77, -79, -91, -9, 11, 35, -8, -8, 65, 39, -64, 50, 26, -68, -80, 182, 20, -21, 19, 54, 19, 34, 55, 89, -43, -173, -8, -5, 30, -27, 27, -1, 6, -30, 35, 10, -3, -5, 64, 34, 41, -18, -4, -2, 6, 41, 22, -19, 16, -3, 21, 144, 5, -26, 69, 0, 54, 16, 28, -53, 14, -38, 32, -30, 20, -7, -298, -1, -86, -162, 2, -3, -4, -18, 48, -434, 2, -23, -40, 42, -23, -145, 9, -2, -24, -2, 2, -53, 15, -25, -3, -3, 8, 0, 63, 65, -21, -145, 11, -19, 110, 43, 15, -31, -38, 0, -18, -36, -36, 78, -53, 38, 18, -88, 16, -131, 27, 62, 40, -38, -128, 3, -4, -34, -48, 53, 17, 0, -27, -1, -7, -94, 21, -119, 32, 9, 21, -3, -20, 94, 23, -2, -5, 54, -126, 27, 38, -31, 18, -26, 51, -7, 159, 77, 20, -58, 29, -31, 5, 18, 11, -4, 7, -43, -52, -105, -42, 6, 28, -28, 23, -112, 3, 7, 44, -84, 75, -41, -30, -206, 19, 2, 71, -48, -55, 6, 6, -23, -38, -6, 24, -23, -8, -8, -181, -7, 57, -24, 104, 0, 7, -26, 29, -33, 17, 2, 18, -72, -38, 2, 0, -5, -32, -23, 19, 44, -129, 11, 8, 11, 15, 243, 33, 6, -5, -9, 110, -20, -327, -91, 211, -22, -10, 13, 34, -109, -72, 124, -141, 105, 37, -100, 26, 8, -23, 142, 89, -32, 15, -7, 6, -44, 15, -56, -93, -23, 5, -27, 36, 70, -14, -21, -101, 85, 21, -20, -575, 2, 17, -94, 18, 10, 54, 83, 18, -300, 11, -7, 94, 89, -26, -23, 24, 420, 30, 38, -17, -37, -87, -2, 139, 25, -73, 18, -71, -29, 25, -44, 12, 0, 3, -6, -66, -153, 5, 63, 51, 88, 33, 40, -35, -35, -113, -70, 3, 27, -87, 30, -27, 86, -103, 2, 60, -8, -130, 1, 0, 32, -120, 1, -46, -209, -217, 66, 122, -148, -42, 0, -99, 95, -24, 4, -164, 85, -3, 30, 110, 4, -124, 66, -23, 41, -8, 3, -37, 30, -33, 8, 210, -57, -30, 103, -42, -182, 75, 50, -20, 1, -4, 21, 70, -2, 97, -95, 197, 26, 7, 38, -36, 11, 32, 2, -32, 11, -52, 22, -5, -103, -22, -252, -132, 16, 95, -57, -22, -16, -43, 19, -4, 42, -107, 23, 9, -48, -27, 58, 10, -36, -71, -27, 9, 97, -41, -146, 24, 21, -3, 68, -36, 8, 65, -186, 3, 15, -131, 24, -106, 18, 61, -78, 15, 8, -18, 8, -69, 50, -69, 5, 293, -77, 48, 6, -9, -6, -102, -81, -5, -202, -6, -4, 22, 21, 72, 15, 119, -21, 130, 4, -1, -15, -9, -86, -95, -3, -27, 18, -9, -290, -19, 53, -53, 8, 59, -169, 25, 10, 59, -64, -197, 15, -188, -14, 73, 12, 111, 7, -36, 38, 78, 50, 75, 82, -19, -37, 67, -114, 57, 23, -38, 205, -68, -54, 17, 126, -72, -1, 17, 12, -5, -4, 29, -4, 16, 33, 20, 0, -71, -22, 5, -2, -2, 18, 30, -166, -24, -25, -42, -1, 76, -30, 94, 140, 22, 129, -7, -120, 70, 52, 4, -45, 22, -26, -63, -2, -21, -53, 91, -39, 3, -21, 26, 1, 112, -22, -78, -25, 21, -98, -15, -5, 24, 1, 16, -25, 31, -50, -3840, -8, -90, 8, 0, -18, 0, -2, -54, -26, 23, 4, 39, -34, 9, -110, -6, -58, -60, -6, 37, -1, -451, 188, -167, -1, 11, -22, 32, -31, 26, -136, 64, 53, 17, 75, -403, 89, 39, -41, 7, 118, 26, 3, 17, -25, 20, -71, -6, -121, -1, -3, 14, 1, -11, 145, 98, -8, 12, 11, -141, -26, 18, -158, 2, -41, 29, 65, 9, 20, -23, 7, -9, -25, -110, -145, 20, -79, 89, -19, 22, 79, 54, 160, 18, 76, -101, -182, 4, -29, 41, 83, 14, 3, 4, -33, 116, 1, -123, 175, 28, -113, 8, -19, 16, -8, 14, 47, 35, 138, 26, 3, 7, 27, -200, 67, -168, -65, 8, 394, 50, 58, 55, -85, 36, 57, -32, 44, 4, -8, -31, -62, 92, -44, -105, 24, -4, -69, -5, 20, -28, 78, -2, -35, -5, -7, -70, 62, -42, 16, 69, 6, 53, 88, -29, -28, -93, 24, -59, 31, 4, 10, -24, -3840, -6, 20, -32, 24, -25, 29, -85, 83, 45, 27, -23, 39, 128, -8, -39, -120, -3, 11, -40, -108, -171, -78, -5, 42, 38, -192, -6, -19, -5, 77, -5, 7, -34, 46, 66, 0, 79, 23, -247, 79, 57, 31, -19, -23, -24, 29, -66, 45, -28, -37, 34, -64, -99, -41, -29, 66, 6, 1, 9, -243, -183, 23, -21, -36, -2, -1, 325, 37, 84, 35, -32, 7, 60, 33, 9, 22, -23, 306, 80, -8, 14, -117, 191, 25, 0, 134, 35, 7, -124, -45, -7, 36, 27, 15, -29, -13, 10, 21, -22, 16, -142, -617, -82, 314, -65, 14, -181, 5, 43, 6, 0, 46, 56, -6, -118, 26, -30, 34, 6, -362, -20, -255, 167, -6, -26, -122, -271, -206, 90, -51, 57, -202, -5, -2, 3, -8, -108, 21, 1, 17, -21, 71, -138, 150, 49, 14, -24, 24, 122, 5, -8, 54, -27, -272, -190, 41, 24, 36, 34, -78, 3, 62, -119, 44, -8, 82, -51, -59, 28, 54, -81, -39, 52, -100, 21, -102, 33, -91, 95, -31, -17, 18, 115, -110, 109, -38, 25, -33, 28, -6, 24, 40, 21, -80, 25, -2, -4, 27, 24, 7, 25, 122, 32, -210, -12, -46, 26, -24, 105, -59, 18, -26, 7, -28, 18, 229, -242, -7, -13, -6, -12, -183, 41, -4, -2, 140, 40, -88, -1, 16, 50, -26, 116, -25, -66, -4, 16, -81, 8, 40, 22, 45, -95, 53, 0, -21, -67, 0, 8, 19, 17, -175, -1, -40, 11, -23, 18, -30, -3, -3, 59, 51, 4, 56, 9, -27, 46, -20, 36, -47, 53, -22, -84, -59, 9, -129, 54, 34, -133, -3, 200, 19, 0, -5, -112, 76, -7, -174, 33, -18, 22, 37, 26, -20, 10, 10, -47, -118, 10, 92, -112, -76, 62, 43, 40, 23, -38, -18, 71, -8, 25, 38, 86, 0, 15, -65, -28, -19, 51, 15, 11, -24, 20, -137, 7, -8, 85, 8, -32, 51, -12, -59, 19, 202, 10, 60, 15, -107, 10, -23, 16, 35, -55, 75, -5, -3, 18, -53, 27, 81, -66, -23, 88, -20, -31, -113, 23, -21, 44, 111, 15, -115, -139, -4, 28, 215, 0};

localparam logic [2912:0][31:0] feature_below = {267, -239, -193, -112, -100, 71, -216, -189, -110, 159, -207, -249, -71, 34, -342, -139, -45, 119, 148, -54, 187, 143, -45, -78, 50, -130, -211, 59, -84, -179, -65, 47, -39, -52, 135, -208, 36, -130, -21, 194, 226, -40, -13, -52, 22, 114, -48, 8, -224, -120, -7, -234, 148, -200, -74, -187, -107, -40, -56, 191, -123, -313, 22, 62, 23, -251, 127, -330, 184, -63, -298, -108, -185, 23, 9, 50, 19, 32, -97, -47, -297, 54, 142, -426, -156, -62, -138, -154, -56, -24, 39, 160, -76, 36, 62, 34, -168, 58, -222, -25, -206, 95, -34, -8, -45, -134, 106, 26, 26, -166, -168, -135, -176, -5, -128, 185, -48, -74, 2, -10, -147, 48, 34, 97, 29, -162, 111, -178, 8, -69, -45, -75, -43, 89, 110, 25, -114, -161, -110, -96, -162, -126, 82, -31, -44, 141, 201, -35, -140, 39, 33, -158, 52, -12, -53, 32, -120, 159, -42, 45, 7, -131, 132, 28, -204, -132, -189, -31, 37, -30, -155, 31, -175, 27, 42, -36, -296, 37, -35, -196, 10, 18, -141, 2, -44, 26, -52, -285, -37, -114, -143, -129, 33, -73, -71, -165, 223, -135, 73, 167, -59, -53, 46, -114, 38, -102, 20, 4, -50, 11, 71, -237, -62, -58, -108, 45, 24, -160, -104, -119, 72, 103, -109, -52, -196, 81, 75, -33, 37, -51, 27, 56, 120, 1, -130, -48, -103, -135, 26, -49, 27, -131, -132, -27, 113, 134, 18, -213, 102, -123, 25, -133, -158, -97, -50, -92, 71, -57, -140, 107, -33, 40, -134, 21, -88, 32, -65, 5, 18, -115, -58, 43, -101, -292, 50, 4, -139, -241, 19, -130, 20, -99, -15, 9, -225, 123, 60, 91, -141, -140, -34, -28, 24, -119, 251, 27, -150, -144, -22, 106, -148, -134, -140, 54, -118, -204, -85, 25, -81, -24, -14, -138, 44, 61, 125, -278, -82, -189, 54, 3, 20, -52, -255, -80, 130, -131, -146, -73, 39, -220, 30, -156, 42, -41, -14, 51, 0, 96, -106, -76, 20, 4, -67, -68, 26, 6, -117, 12, 27, -35, -13, 8, -119, 17, 25, -146, 22, -61, -277, 6, -4, -169, 47, -33, -10, -101, 218, 99, -191, -273, 73, 87, 32, 2, -1, 58, -122, -258, 51, -32, -7, 6, -63, -38, -77, -4, 48, -128, 18, -27, -169, 63, 54, -4, -101, -288, -33, -29, -37, -4, 76, -61, 29, -33, -77, 91, -72, -91, -143, -52, -49, -90, -70, -13, 108, 34, 20, -255, -41, 76, 3, -56, -114, 27, 2, 129, -188, -104, 15, 17, -151, 81, 24, -119, 5, 47, 25, -215, -394, 27, -147, 107, -36, 23, 123, 1, -68, 105, -25, -3, -174, -83, 108, 25, -93, -46, 7, 60, -145, 126, -36, -82, 48, -167, -262, 99, 22, -192, 37, 177, -29, -203, -153, -20, 33, -11, 96, 16, -47, -10, 100, -115, 106, 2, 145, -74, -3, -70, -157, 19, -36, -31, -110, 89, -21, 56, -125, -116, -101, -39, -115, -54, 59, 117, -188, -134, 37, -165, -110, 21, 20, 3, -21, -125, 126, 61, -123, -67, 22, -145, 33, 25, -7, 136, -24, -4, 128, -4, 0, -196, 4, 98, 21, -125, 59, 33, -103, -168, 26, 125, -24, -87, 24, -30, 32, -133, 66, 207, 382, 77, -79, 85, -144, -138, 104, -3, 87, 7, -17, -48, -75, -39, 76, 124, 117, -77, 6, -120, 23, -165, -6, -2, -34, -66, 53, -32, -29, 8, 24, -121, 47, 123, -393, 29, 0, 122, -13, 1, 83, -5, 89, -52, -83, 125, -13, 78, -130, -53, -75, -119, 15, -74, -49, 151, -110, -96, 118, 34, -36, -79, 74, 42, 11, 44, 30, -95, -116, -44, -120, -68, 118, -91, -111, -29, -39, 34, -151, -70, -35, -117, -56, 3, 101, 103, -26, -6, -116, 45, -25, -179, 0, -63, -156, 48, -38, -184, -289, 48, -38, -128, 6, 19, -2, -18, -2, -222, -31, 1, 5, 10, -217, 81, -43, 29, 25, 12, -223, -31, 151, 18, -70, -28, 8, 88, 223, 39, -27, -102, 48, -2, 155, -3, -136, -4, 5, -10, -246, 62, -25, 25, -25, 232, 100, 20, -21, -13, -5, -7, 36, 16, 3, 24, 9, 6, -35, 7, 49, 20, 3, 21, -79, -109, -104, -47, -152, 42, -65, -134, -65, -127, -12, 30, -13, 0, -84, 36, 20, -37, 175, 156, -105, -156, 15, -150, -137, -46, 63, 75, -10, 35, -1, 105, 17, -116, 1, 228, 73, -41, 25, 9, -50, -3, -246, -164, -52, -93, 74, 117, -66, 31, 21, -175, -219, -40, 19, 95, -52, 104, 42, -161, 177, -5, -24, -57, 87, -2, 43, -136, 19, -31, 17, -134, -194, 18, 37, -35, 24, 42, 15, -142, 103, -34, 2, 2, -39, -206, 10, -1, -31, 245, -32, -89, 23, -4, 8, 1, 19, 50, -199, 28, -6, -33, -23, 70, -89, 38, 118, -102, 42, -176, 8, 46, -20, 17, 14, -1, 0, -60, -1, -44, 192, -127, -74, -4, 51, 23, 70, 87, -115, -72, 46, -71, -137, -92, -60, 27, 86, -122, 104, 158, -39, 27, -116, 29, -51, 24, 20, 28, -189, -22, 5, 43, 1, 58, 20, -167, -31, 4, -29, 26, 88, -1, -26, 61, -142, 130, 53, 27, -148, 45, -197, 26, -3, 22, -153, -140, 36, -6, -34, 77, 49, 17, 15, -44, -22, 78, -62, -515, -50, -11, 147, -3, 5, 72, -22, 162, 86, -53, -117, 0, -48, -54, -21, 19, 176, -43, 98, -89, -2, -13, 137, 24, -28, 33, -1, -37, -5, 42, -45, -184, -151, 283, -239, -98, -81, 109, -4, -25, 264, -15, -2, -5, -85, -7, 78, -73, 7, 22, -86, 38, -36, -14, -7, 58, -260, 22, -3, 39, -40, -230, -7, 27, -26, -122, -18, -140, 13, 8, -172, 6, -131, 11, -19, 84, -116, -64, -54, -61, 65, -30, 52, 58, -109, -119, -164, 75, -7, -111, -10, -32, -144, -186, 69, 9, 146, -32, -5, 75, 20, 22, -19, -51, 36, 0, 53, -183, -32, 6, -120, -35, -132, 81, 21, -32, -37, -1, 14, -25, 40, -1, -59, -2, -10, -34, 23, -24, -19, -67, -49, -1, -74, 3, -83, -43, 19, -32, -14, -125, 49, -133, -705, 122, 1, 29, 21, -111, -361, -166, -104, 84, 1, 39, 33, -184, -22, -83, -7, -118, 69, -70, 20, -31, -65, -28, 15, -2, 156, -32, 29, 32, -42, -7, 0, -39, -31, 60, 49, -6, 27, -22, 15, -6, -52, -42, -93, -20, 25, 105, -55, -4, 14, 279, -6, -42, 147, -50, -215, -125, 27, -21, 30, -119, -94, 18, 1, -152, 311, 92, 20, -104, 119, -72, -101, -181, 49, -52, -31, -112, 20, -147, 20, 5, 56, 56, -12, -49, 114, 110, 77, -203, 22, 65, -55, -40, 135, -92, 32, -88, -76, 6, -79, -39, -176, -72, 1, 200, -202, -199, 22, -167, -177, -91, -5, 74, -63, -63, -77, 30, -10, -154, 30, -104, 79, -38, -78, -68, -165, -22, -14, 131, -100, -113, 15, -104, -9, -165, 61, -8, 22, -26, -9, -163, 16, 2, 79, -46, 67, -22, -152, 107, 45, -113, -18, -37, -4, 89, -83, -4, -1, 109, -266, -110, 49, -221, 70, -5, 75, -2, 19, 66, -3, -110, -58, 17, 17, -32, 3, -50, 11, -23, -79, -6, 23, -108, -24, -102, -30, -7, 34, -86, 86, 39, 19, -24, 24, 58, 17, -27, 41, -26, 20, -80, 21, -32, 20, 73, 73, -49, 28, -37, -83, -37, 58, -66, 2, 50, 152, -87, -109, -141, -25, -52, -38, -167, 30, 37, -310, 113, 103, 19, -104, -91, -93, 22, 354, 15, -1, 30, -40, -6, -149, -35, -69, 23, 80, 31, -120, -10, 5, 22, -4, 12, -51, -29, -35, -14, -6, 19, -3, -103, -27, 26, -23, 64, 150, -8, -30, -105, 78, -5, -147, -1, 48, -13, 86, 20, 49, 19, -87, 33, -4, -45, -5, -3, 14, 60, -36, -3, -42, -157, -2, 84, -67, -100, 0, -7, 2, -80, 23, 6, 58, 43, -299, -85, 59, -34, -24, -3, -4, 1, 54, -3, -4, 14, 37, 15, 19, -69, -8, -58, 155, -295, -92, 9, -157, 17, -4, 17, -19, 25, -48, 104, 107, -121, 6, -249, -27, 77, -28, 81, -30, 23, -89, 44, -112, 30, -8, -25, 124, -8, -58, 15, 232, 30, 63, 78, 51, -109, -101, -86, 5, 18, -18, 18, -26, -60, -121, 42, 35, 30, -74, -78, -72, -103, -104, 18, -21, 185, 17, -43, -15, -127, -62, 5, -139, 122, -133, 115, -130, 79, -11, 8, -120, -108, 78, -4, 17, -145, 97, 38, 3, -109, -8, 46, 0, -4, 76, 76, -150, -2, 21, -29, 35, -97, -29, 25, 21, 164, -69, 81, -64, -152, 3, 4, -27, 0, -28, -1, 57, -26, -98, -181, 25, 108, 16, -60, 66, -4, 31, 125, 26, -33, 22, -110, 72, -33, 1, -77, 54, 29, 12, -34, -93, -45, 15, -1, 26, 74, 2, -42, 176, 0, -2, 48, -352, 61, -74, -1, 45, 182, 31, -1, -2, -116, -27, 25, -12, -71, 24, 248, -34, -70, -328, -32, 21, 28, 40, -122, 16, -8, 5, -6, 5, 4, 132, -9, -76, -8, 7, -1, 19, -23, -76, -138, 100, -8, -2, -7, 44, -34, -17, 4, 3, 58, -25, -69, -2, 9, 87, -26, 91, -47, -110, -35, -44, -41, -88, -27, -63, 172, 6, -91, 129, -2, -105, 69, -43, -153, -114, 21, 80, -36, -82, -98, 58, -98, 6, -6, -3, -123, -90, -36, -32, -89, 59, 23, -81, -132, 44, -37, -57, 23, -1, 212, -1, 0, -79, 90, 50, -3, 60, 41, -157, 6, -21, 43, -109, 7, 67, 80, -79, -108, -8, -23, -4, -31, -30, 50, -34, 22, -139, 92, -152, 81, 169, -43, -33, 18, -149, -51, 63, 240, -114, -149, -86, -61, 15, -10, -26, 118, -34, -69, 2, -2, -23, 27, 3, -2, -24, 52, -26, -217, -4, -26, -58, 30, -23, -35, -59, 53, 19, 96, -24, 45, -82, 2, 135, 38, -28, 31, -4, -1, 10, 10, -18, -238, -24, 18, 206, -104, -178, 4, -71, 3, 57, 23, -8, 26, -41, 111, 82, 22, 31, 69, 306, 20, 0, -15, -135, -26, -27, 14, -220, 83, -1, 25, -111, 18, 43, -320, 65, -375, -77, 43, -142, 57, -133, 4, 68, -69, -64, -42, -41, 14, -18, 121, -70, 2, -40, -1, -98, 31, -12, -101, -13, -52, 26, 0, -1, -47, -183, -5, 34, -107, -63, -24, 30, -5, -228, -28, -23, -1, 39, -122, 4, 125, -3, -7, 84, 3, -1, 44, -1, -67, -75, 3, -47, 5, -19, -28, -139, -20, 6, -198, 21, -99, 14, 142, 35, -103, 18, 25, -6, -21, -16, -4, -8, -47, 15, -67, 83, 22, -25, -65, -9, -52, -27, -64, -26, 23, 2, -27, 32, -244, -91, -22, 24, 1, 22, -289, 308, -35, 40, -186, -2, -30, 18, -28, -15, 3, 23, -19, -67, 113, -62, -27, -9, -32, 1, -23, 17, -6, 22, -145, -29, 58, -19, -87, 83, 57, -11, -60, 37, -155, -6, -34, -17, 249, 20, -91, 118, -29, -93, 160, -185, -100, -109, -19, 70, 47, -4, -79, -8, -44, -39, 10, -125, 24, -8, 42, -38, -155, 17, -85, 21, -7, 26, -101, 37, 221, 2, -10, 41, 98, 24, -30, 22, -6, 103, -105, 19, -93, 73, 5, -254, 64, 51, -98, 111, -72, 5, -25, 24, -6, 181, 169, 6, -27, -160, 33, 29, -110, 40, 32, 34, -69, 92, -75, -95, 23, -138, 3, -58, -35, -63, 53, 21, -141, 83, 54, 45, -37, -169, -112, 33, -127, 81, 3, -72, 0, -12, -84, -60, -136, 65, -39, -143, -111, 84, -29, 23, -42, -15, 49, -114, 69, -7, -195, 10, -25, -82, 11, -55, 51, 68, -50, 112, -149, 140, 18, 17, -2, 23, -68, -14, 50, -33, -3, 101, -61, -22, 0, 2, 26, 24, -8, -42, -80, -4, 25, 26, -73, 96, 109, 21, -170, -8, 98, 29, -204, 15, -168, 0, 84, 9, -86, 43, 58, -6, 34, -106, -86, -9, 4, 17, -76, 52, -139, 37, 84, -251, -29, 20, -50, 220, -49, -396, -18, -8, -72, 32, -335, 8, 120, 18, -2, 8, 91, 19, -48, -30, -4, 24, -20, 19, -21, -9, -3, -23, -58, 34, -20, 9, 35, -394, -187, 113, 18, -132, 10, 15, 86, 27, 57, 5, -25, 17, 108, 22, -23, -18, 134, 14, -101, -78, -2, -262, -54, 3, -22, -28, -9, 165, -149, 9, -23, 28, 79, -59, -16, -39, -29, 32, 37, 25, -97, 11, -34, 17, -52, 21, 40, -34, 20, 147, -91, 53, -171, 18, -6, 82, -28, -103, -41, -82, -59, 59, 47, 3, 22, -123, -91, 9, -96, 87, -16, 9, 122, -36, 49, 0, 109, -118, -70, -1, 92, 25, 15, -7, -14, -23, 21, 26, 120, 0, 0, 93, 128, -6, 2, -121, -56, -23, 74, -3, -18, 125, -11, -265, 56, 37, -73, 44, 72, -19, 31, 55, 3, 23, 19, -25, 0, 162, 83, -132, -61, -27, 66, -27, 23, -19, -36, -57, 5, 51, 282, -36, 44, 37, 82, 10, -57, -126, 29, 107, 15, -5, -173, -23, 16, 103, 21, 20, -236, -103, -18, -3, -94, -58, 27, 51, -3, -64, 23, 6, 22, -59, 7, 19, 18, -37, -39, -126, 6, 30, 60, -27, 21, -72, -456, -5, -72, -4, -68, -28, 18, -44, 123, 223, 178, 7, -12, 5, 122, -17, 29, -28, 165, -506, 48, -3, 22, -120, 17, -146, 63, -40, -49, -24, -76, -20, 41, -20, 97, -113, 31, -240, 17, -3, 60, 51, -200, -246, 17, 131, -12, 14, 77, -24, 15, -36, 93, -25, 20, -7, -206, -8, 21, -23, 595, -22, 117, 28, -115, -48, -49, -23, -29, 91, 61, -24, 5, -30, -59, 43, -21, 29, 19, -190, -25, 17, -139, -76, -63, 76, -151, -78, -146, -211, -40, -89, -92, 29, 132, 58, -109, 74, -48, -34, -4, 26, 86, 22, -107, -4, 54, 9, -20, -91, -21, 50, 2, 6, -35, 108, 20, -119, 66, 18, -115, 25, 12, -8, 31, 78, 116, -40, -85, 8, 102, 24, 75, -33, -2, 26, -137, -74, -85, -62, 74, -7, 16, 14, -222, 17, -60, 89, 216, 102, -130, 18, 65, -20, -70, -22, 32, 119, -4, 45, 9, 18, -132, -25, -99, 17, -20, 19, -91, 142, 119, -25, 54, -66, -6, 7, -30, -113, -26, 17, -22, 7, 20, 91, -20, -44, -71, -462, 66, -11, 4, 30, -5, 59, -98, -479, -82, 25, -21, 3, -217, 152, -52, 20, 63, -31, -6, 56, 24, -56, -26, 40, -40, 18, -65, 61, 58, 17, -5, -44, 1, 10, 149, -41, -23, 0, -19, -51, -23, 19, -8, 44, 40, -5, -23, -129, -69, 62, 34, 5, -77, 20, -19, 2, -2, 46, 153, -79, -234, -3840, -31, -4, -20, -8, -83, 139, -33, 18, -27, 19, 4, 162, -16, -88, -61, -60, 33, -62, -31, 97, -45, -101, 60, 86, 32, -28, 36, 7, -128, -153, 19, -182, -36, 61, -8, -110, 21, -150, 34, 5, -5, 37, -180, -27, 43, -32, 5, 68, 32, 1, -64, 11, -67, -81, 165, 107, 14, -173, -173, 52, -34, 75, -21, 2, -2, -31, -69, 96, -21, -22, 30, 32, 17, -107, 302, 24, 19, -6, 23, -126, -21, -31, 18, -133, 25, -116, -4, -128, 94, 36, 1, -26, 83, -24, -37, -9, -2, -27, -46, 139, 27, 66, -56, 4, 2, 44, 42, -32, 18, -2, 24, 45, -5, -55, 85, -63, 17, -7, -74, 125, 23, -104, 36, -17, -9, -23, -20, 37, 57, -25, -1, -54, -109, 107, 13, -24, 32, -45, 21, -19, -27, -91, 4, -35, 46, -6, 17, -138, 3, -33, -227, 38, 25, -55, -65, 100, -81, -6, 15, -2, 11, 5, -243, -8, 114, -28, 74, -69, -10, -26, 53, -4, -15, 42, -3, -56, 15, 117, 14, -18, 26, 42, 20, -10, 15, -21, 29, -25, 15, -115, 46, -59, 30, -4, -65, -69, -114, 103, 2, -6, 9, -25, -696, 57, -2, -19, 59, -211, -5, 44, 16, -8, 2, -35, -23, -41, 16, -64, 6, -5, 0, -196, 5, 13, 80, -119, -52, 12, 48, -30, 5, -64, 4, -64, 5, -8, 62, 17, -57, 4, 2, 2, 37, -52, 42, -68, -185, -101, -34, -70, 3, -64, -101, 102, -42, -35, -68, -72, -22, -12, -7, 30, 23, -55, 74, 4, 9, -161, 68, 149, 50, -94, -18, 15, -181, 57, -178, 66, -7, -10, -111, 67, -21, -22, -1, 81, -43, -4, 83, 7, 84, 25, -119, -87, 2, 129, -30, -93, -28, 21, -31, 65, 116, 18, -85, 103, -43, -71, -8, 44, 36, 150, 105, -24, 42, 25, -120, 3, -27, 95, -25, 89, 50, -9, 122, -7, 10, 7, 92, 18, 5, 69, -6, 4, -33, 20, -94, 11, -45, 36, -108, 19, -24, 57, -7, -40, 210, -100, -30, -46, 100, 151, -60, 28, -5, 54, -21, 20, -1, -4, -29, -8, -38, 28, 156, 2, -191, -49, -27, 0, -80, -54, 3, 17, 151, 4, -41, 108, 47, -67, -8, 101, -150, 5, -46, 27, -24, 33, 4, -127, -17, 43, -23, -126, -4, 149, 82, -30, -28, 21, -22, 33, -98, -35, 10, -5, -23, 24, 90, 9, 96, 25, -6, -57, 83, -7, -20, -78, -6, 14, -102, -24, -17, 62};

