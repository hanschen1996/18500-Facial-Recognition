/** @file vj_weights.vh
 *  @brief Viola-Jones weights data structure
 */

// assume we use haarcascade_frontalface_default.xml
`define NUM_STAGE 25
`define NUM_FEATURE 2913
`define WINDOW_SIZE 24
`define LAPTOP_WIDTH 160
`define LAPTOP_HEIGHT 120
`define PYRAMID_LEVELS 9

`define PYRAMID_WIDTHS {32'd37,32'd44,32'd53,32'd64,32'd77,32'd92,32'd111,32'd133,32'd160}
`define PYRAMID_HEIGHTS {32'd27,32'd33,32'd40,32'd48,32'd57,32'd69,32'd83,32'd99,32'd120}

`define PYRAMID_X_MAPPINGS {{32'd687,32'd683,32'd678,32'd674,32'd670,32'd665,32'd661,32'd657,32'd652,32'd648,32'd644,32'd640,32'd635,32'd631,32'd627,32'd622,32'd618,32'd614,32'd609,32'd605,32'd601,32'd596,32'd592,32'd588,32'd583,32'd579,32'd575,32'd570,32'd566,32'd562,32'd557,32'd553,32'd549,32'd544,32'd540,32'd536,32'd531,32'd527,32'd523,32'd518,32'd514,32'd510,32'd505,32'd501,32'd497,32'd492,32'd488,32'd484,32'd480,32'd475,32'd471,32'd467,32'd462,32'd458,32'd454,32'd449,32'd445,32'd441,32'd436,32'd432,32'd428,32'd423,32'd419,32'd415,32'd410,32'd406,32'd402,32'd397,32'd393,32'd389,32'd384,32'd380,32'd376,32'd371,32'd367,32'd363,32'd358,32'd354,32'd350,32'd345,32'd341,32'd337,32'd332,32'd328,32'd324,32'd320,32'd315,32'd311,32'd307,32'd302,32'd298,32'd294,32'd289,32'd285,32'd281,32'd276,32'd272,32'd268,32'd263,32'd259,32'd255,32'd250,32'd246,32'd242,32'd237,32'd233,32'd229,32'd224,32'd220,32'd216,32'd211,32'd207,32'd203,32'd198,32'd194,32'd190,32'd185,32'd181,32'd177,32'd172,32'd168,32'd164,32'd160,32'd155,32'd151,32'd147,32'd142,32'd138,32'd134,32'd129,32'd125,32'd121,32'd116,32'd112,32'd108,32'd103,32'd99,32'd95,32'd90,32'd86,32'd82,32'd77,32'd73,32'd69,32'd64,32'd60,32'd56,32'd51,32'd47,32'd43,32'd38,32'd34,32'd30,32'd25,32'd21,32'd17,32'd12,32'd8,32'd4,32'd0},{32'd578,32'd574,32'd570,32'd567,32'd563,32'd560,32'd556,32'd552,32'd549,32'd545,32'd541,32'd538,32'd534,32'd530,32'd527,32'd523,32'd520,32'd516,32'd512,32'd509,32'd505,32'd501,32'd498,32'd494,32'd490,32'd487,32'd483,32'd480,32'd476,32'd472,32'd469,32'd465,32'd461,32'd458,32'd454,32'd450,32'd447,32'd443,32'd440,32'd436,32'd432,32'd429,32'd425,32'd421,32'd418,32'd414,32'd410,32'd407,32'd403,32'd400,32'd396,32'd392,32'd389,32'd385,32'd381,32'd378,32'd374,32'd370,32'd367,32'd363,32'd360,32'd356,32'd352,32'd349,32'd345,32'd341,32'd338,32'd334,32'd330,32'd327,32'd323,32'd320,32'd316,32'd312,32'd309,32'd305,32'd301,32'd298,32'd294,32'd290,32'd287,32'd283,32'd280,32'd276,32'd272,32'd269,32'd265,32'd261,32'd258,32'd254,32'd250,32'd247,32'd243,32'd240,32'd236,32'd232,32'd229,32'd225,32'd221,32'd218,32'd214,32'd210,32'd207,32'd203,32'd200,32'd196,32'd192,32'd189,32'd185,32'd181,32'd178,32'd174,32'd170,32'd167,32'd163,32'd160,32'd156,32'd152,32'd149,32'd145,32'd141,32'd138,32'd134,32'd130,32'd127,32'd123,32'd120,32'd116,32'd112,32'd109,32'd105,32'd101,32'd98,32'd94,32'd90,32'd87,32'd83,32'd80,32'd76,32'd72,32'd69,32'd65,32'd61,32'd58,32'd54,32'd50,32'd47,32'd43,32'd40,32'd36,32'd32,32'd29,32'd25,32'd21,32'd18,32'd14,32'd10,32'd7,32'd3,32'd0},{32'd480,32'd476,32'd473,32'd470,32'd467,32'd464,32'd461,32'd458,32'd455,32'd452,32'd449,32'd446,32'd443,32'd440,32'd437,32'd434,32'd431,32'd428,32'd425,32'd422,32'd419,32'd416,32'd413,32'd410,32'd407,32'd404,32'd401,32'd398,32'd395,32'd392,32'd389,32'd386,32'd383,32'd380,32'd377,32'd374,32'd371,32'd368,32'd365,32'd362,32'd359,32'd356,32'd353,32'd350,32'd347,32'd344,32'd341,32'd338,32'd335,32'd332,32'd329,32'd326,32'd323,32'd320,32'd316,32'd313,32'd310,32'd307,32'd304,32'd301,32'd298,32'd295,32'd292,32'd289,32'd286,32'd283,32'd280,32'd277,32'd274,32'd271,32'd268,32'd265,32'd262,32'd259,32'd256,32'd253,32'd250,32'd247,32'd244,32'd241,32'd238,32'd235,32'd232,32'd229,32'd226,32'd223,32'd220,32'd217,32'd214,32'd211,32'd208,32'd205,32'd202,32'd199,32'd196,32'd193,32'd190,32'd187,32'd184,32'd181,32'd178,32'd175,32'd172,32'd169,32'd166,32'd163,32'd160,32'd156,32'd153,32'd150,32'd147,32'd144,32'd141,32'd138,32'd135,32'd132,32'd129,32'd126,32'd123,32'd120,32'd117,32'd114,32'd111,32'd108,32'd105,32'd102,32'd99,32'd96,32'd93,32'd90,32'd87,32'd84,32'd81,32'd78,32'd75,32'd72,32'd69,32'd66,32'd63,32'd60,32'd57,32'd54,32'd51,32'd48,32'd45,32'd42,32'd39,32'd36,32'd33,32'd30,32'd27,32'd24,32'd21,32'd18,32'd15,32'd12,32'd9,32'd6,32'd3,32'd0},{32'd397,32'd395,32'd392,32'd390,32'd387,32'd385,32'd382,32'd380,32'd377,32'd375,32'd372,32'd370,32'd367,32'd365,32'd362,32'd360,32'd357,32'd355,32'd352,32'd350,32'd347,32'd345,32'd342,32'd340,32'd337,32'd335,32'd332,32'd330,32'd327,32'd325,32'd322,32'd320,32'd317,32'd315,32'd312,32'd310,32'd307,32'd305,32'd302,32'd300,32'd297,32'd295,32'd292,32'd290,32'd287,32'd285,32'd282,32'd280,32'd277,32'd275,32'd272,32'd270,32'd267,32'd265,32'd262,32'd260,32'd257,32'd255,32'd252,32'd250,32'd247,32'd245,32'd242,32'd240,32'd237,32'd235,32'd232,32'd230,32'd227,32'd225,32'd222,32'd220,32'd217,32'd215,32'd212,32'd210,32'd207,32'd205,32'd202,32'd200,32'd197,32'd195,32'd192,32'd190,32'd187,32'd185,32'd182,32'd180,32'd177,32'd175,32'd172,32'd170,32'd167,32'd165,32'd162,32'd160,32'd157,32'd155,32'd152,32'd150,32'd147,32'd145,32'd142,32'd140,32'd137,32'd135,32'd132,32'd130,32'd127,32'd125,32'd122,32'd120,32'd117,32'd115,32'd112,32'd110,32'd107,32'd105,32'd102,32'd100,32'd97,32'd95,32'd92,32'd90,32'd87,32'd85,32'd82,32'd80,32'd77,32'd75,32'd72,32'd70,32'd67,32'd65,32'd62,32'd60,32'd57,32'd55,32'd52,32'd50,32'd47,32'd45,32'd42,32'd40,32'd37,32'd35,32'd32,32'd30,32'd27,32'd25,32'd22,32'd20,32'd17,32'd15,32'd12,32'd10,32'd7,32'd5,32'd2,32'd0},{32'd330,32'd328,32'd326,32'd324,32'd322,32'd320,32'd317,32'd315,32'd313,32'd311,32'd309,32'd307,32'd305,32'd303,32'd301,32'd299,32'd297,32'd295,32'd292,32'd290,32'd288,32'd286,32'd284,32'd282,32'd280,32'd278,32'd276,32'd274,32'd272,32'd270,32'd268,32'd265,32'd263,32'd261,32'd259,32'd257,32'd255,32'd253,32'd251,32'd249,32'd247,32'd245,32'd243,32'd241,32'd238,32'd236,32'd234,32'd232,32'd230,32'd228,32'd226,32'd224,32'd222,32'd220,32'd218,32'd216,32'd214,32'd211,32'd209,32'd207,32'd205,32'd203,32'd201,32'd199,32'd197,32'd195,32'd193,32'd191,32'd189,32'd187,32'd184,32'd182,32'd180,32'd178,32'd176,32'd174,32'd172,32'd170,32'd168,32'd166,32'd164,32'd162,32'd160,32'd157,32'd155,32'd153,32'd151,32'd149,32'd147,32'd145,32'd143,32'd141,32'd139,32'd137,32'd135,32'd132,32'd130,32'd128,32'd126,32'd124,32'd122,32'd120,32'd118,32'd116,32'd114,32'd112,32'd110,32'd108,32'd105,32'd103,32'd101,32'd99,32'd97,32'd95,32'd93,32'd91,32'd89,32'd87,32'd85,32'd83,32'd81,32'd78,32'd76,32'd74,32'd72,32'd70,32'd68,32'd66,32'd64,32'd62,32'd60,32'd58,32'd56,32'd54,32'd51,32'd49,32'd47,32'd45,32'd43,32'd41,32'd39,32'd37,32'd35,32'd33,32'd31,32'd29,32'd27,32'd24,32'd22,32'd20,32'd18,32'd16,32'd14,32'd12,32'd10,32'd8,32'd6,32'd4,32'd2,32'd0},{32'd276,32'd274,32'd273,32'd271,32'd269,32'd267,32'd266,32'd264,32'd262,32'd260,32'd259,32'd257,32'd255,32'd253,32'd252,32'd250,32'd248,32'd246,32'd245,32'd243,32'd241,32'd240,32'd238,32'd236,32'd234,32'd233,32'd231,32'd229,32'd227,32'd226,32'd224,32'd222,32'd220,32'd219,32'd217,32'd215,32'd213,32'd212,32'd210,32'd208,32'd206,32'd205,32'd203,32'd201,32'd200,32'd198,32'd196,32'd194,32'd193,32'd191,32'd189,32'd187,32'd186,32'd184,32'd182,32'd180,32'd179,32'd177,32'd175,32'd173,32'd172,32'd170,32'd168,32'd166,32'd165,32'd163,32'd161,32'd160,32'd158,32'd156,32'd154,32'd153,32'd151,32'd149,32'd147,32'd146,32'd144,32'd142,32'd140,32'd139,32'd137,32'd135,32'd133,32'd132,32'd130,32'd128,32'd126,32'd125,32'd123,32'd121,32'd120,32'd118,32'd116,32'd114,32'd113,32'd111,32'd109,32'd107,32'd106,32'd104,32'd102,32'd100,32'd99,32'd97,32'd95,32'd93,32'd92,32'd90,32'd88,32'd86,32'd85,32'd83,32'd81,32'd80,32'd78,32'd76,32'd74,32'd73,32'd71,32'd69,32'd67,32'd66,32'd64,32'd62,32'd60,32'd59,32'd57,32'd55,32'd53,32'd52,32'd50,32'd48,32'd46,32'd45,32'd43,32'd41,32'd40,32'd38,32'd36,32'd34,32'd33,32'd31,32'd29,32'd27,32'd26,32'd24,32'd22,32'd20,32'd19,32'd17,32'd15,32'd13,32'd12,32'd10,32'd8,32'd6,32'd5,32'd3,32'd1,32'd0},{32'd229,32'd227,32'd226,32'd224,32'd223,32'd221,32'd220,32'd219,32'd217,32'd216,32'd214,32'd213,32'd211,32'd210,32'd209,32'd207,32'd206,32'd204,32'd203,32'd201,32'd200,32'd198,32'd197,32'd196,32'd194,32'd193,32'd191,32'd190,32'd188,32'd187,32'd185,32'd184,32'd183,32'd181,32'd180,32'd178,32'd177,32'd175,32'd174,32'd172,32'd171,32'd170,32'd168,32'd167,32'd165,32'd164,32'd162,32'd161,32'd160,32'd158,32'd157,32'd155,32'd154,32'd152,32'd151,32'd149,32'd148,32'd147,32'd145,32'd144,32'd142,32'd141,32'd139,32'd138,32'd136,32'd135,32'd134,32'd132,32'd131,32'd129,32'd128,32'd126,32'd125,32'd123,32'd122,32'd121,32'd119,32'd118,32'd116,32'd115,32'd113,32'd112,32'd110,32'd109,32'd108,32'd106,32'd105,32'd103,32'd102,32'd100,32'd99,32'd98,32'd96,32'd95,32'd93,32'd92,32'd90,32'd89,32'd87,32'd86,32'd85,32'd83,32'd82,32'd80,32'd79,32'd77,32'd76,32'd74,32'd73,32'd72,32'd70,32'd69,32'd67,32'd66,32'd64,32'd63,32'd61,32'd60,32'd59,32'd57,32'd56,32'd54,32'd53,32'd51,32'd50,32'd49,32'd47,32'd46,32'd44,32'd43,32'd41,32'd40,32'd38,32'd37,32'd36,32'd34,32'd33,32'd31,32'd30,32'd28,32'd27,32'd25,32'd24,32'd23,32'd21,32'd20,32'd18,32'd17,32'd15,32'd14,32'd12,32'd11,32'd10,32'd8,32'd7,32'd5,32'd4,32'd2,32'd1,32'd0},{32'd191,32'd190,32'd188,32'd187,32'd186,32'd185,32'd184,32'd182,32'd181,32'd180,32'd179,32'd178,32'd176,32'd175,32'd174,32'd173,32'd172,32'd170,32'd169,32'd168,32'd167,32'd166,32'd164,32'd163,32'd162,32'd161,32'd160,32'd158,32'd157,32'd156,32'd155,32'd153,32'd152,32'd151,32'd150,32'd149,32'd147,32'd146,32'd145,32'd144,32'd143,32'd141,32'd140,32'd139,32'd138,32'd137,32'd135,32'd134,32'd133,32'd132,32'd131,32'd129,32'd128,32'd127,32'd126,32'd125,32'd123,32'd122,32'd121,32'd120,32'd119,32'd117,32'd116,32'd115,32'd114,32'd113,32'd111,32'd110,32'd109,32'd108,32'd107,32'd105,32'd104,32'd103,32'd102,32'd101,32'd99,32'd98,32'd97,32'd96,32'd95,32'd93,32'd92,32'd91,32'd90,32'd89,32'd87,32'd86,32'd85,32'd84,32'd83,32'd81,32'd80,32'd79,32'd78,32'd76,32'd75,32'd74,32'd73,32'd72,32'd70,32'd69,32'd68,32'd67,32'd66,32'd64,32'd63,32'd62,32'd61,32'd60,32'd58,32'd57,32'd56,32'd55,32'd54,32'd52,32'd51,32'd50,32'd49,32'd48,32'd46,32'd45,32'd44,32'd43,32'd42,32'd40,32'd39,32'd38,32'd37,32'd36,32'd34,32'd33,32'd32,32'd31,32'd30,32'd28,32'd27,32'd26,32'd25,32'd24,32'd22,32'd21,32'd20,32'd19,32'd18,32'd16,32'd15,32'd14,32'd13,32'd12,32'd10,32'd9,32'd8,32'd7,32'd6,32'd4,32'd3,32'd2,32'd1,32'd0}}
`define PYRAMID_Y_MAPPINGS {{32'd528,32'd524,32'd520,32'd515,32'd511,32'd506,32'd502,32'd497,32'd493,32'd488,32'd484,32'd480,32'd475,32'd471,32'd466,32'd462,32'd457,32'd453,32'd448,32'd444,32'd440,32'd435,32'd431,32'd426,32'd422,32'd417,32'd413,32'd408,32'd404,32'd400,32'd395,32'd391,32'd386,32'd382,32'd377,32'd373,32'd368,32'd364,32'd360,32'd355,32'd351,32'd346,32'd342,32'd337,32'd333,32'd328,32'd324,32'd320,32'd315,32'd311,32'd306,32'd302,32'd297,32'd293,32'd288,32'd284,32'd280,32'd275,32'd271,32'd266,32'd262,32'd257,32'd253,32'd248,32'd244,32'd240,32'd235,32'd231,32'd226,32'd222,32'd217,32'd213,32'd208,32'd204,32'd200,32'd195,32'd191,32'd186,32'd182,32'd177,32'd173,32'd168,32'd164,32'd160,32'd155,32'd151,32'd146,32'd142,32'd137,32'd133,32'd128,32'd124,32'd120,32'd115,32'd111,32'd106,32'd102,32'd97,32'd93,32'd88,32'd84,32'd80,32'd75,32'd71,32'd66,32'd62,32'd57,32'd53,32'd48,32'd44,32'd40,32'd35,32'd31,32'd26,32'd22,32'd17,32'd13,32'd8,32'd4,32'd0},{32'd432,32'd429,32'd425,32'd421,32'd418,32'd414,32'd410,32'd407,32'd403,32'd400,32'd396,32'd392,32'd389,32'd385,32'd381,32'd378,32'd374,32'd370,32'd367,32'd363,32'd360,32'd356,32'd352,32'd349,32'd345,32'd341,32'd338,32'd334,32'd330,32'd327,32'd323,32'd320,32'd316,32'd312,32'd309,32'd305,32'd301,32'd298,32'd294,32'd290,32'd287,32'd283,32'd280,32'd276,32'd272,32'd269,32'd265,32'd261,32'd258,32'd254,32'd250,32'd247,32'd243,32'd240,32'd236,32'd232,32'd229,32'd225,32'd221,32'd218,32'd214,32'd210,32'd207,32'd203,32'd200,32'd196,32'd192,32'd189,32'd185,32'd181,32'd178,32'd174,32'd170,32'd167,32'd163,32'd160,32'd156,32'd152,32'd149,32'd145,32'd141,32'd138,32'd134,32'd130,32'd127,32'd123,32'd120,32'd116,32'd112,32'd109,32'd105,32'd101,32'd98,32'd94,32'd90,32'd87,32'd83,32'd80,32'd76,32'd72,32'd69,32'd65,32'd61,32'd58,32'd54,32'd50,32'd47,32'd43,32'd40,32'd36,32'd32,32'd29,32'd25,32'd21,32'd18,32'd14,32'd10,32'd7,32'd3,32'd0},{32'd357,32'd354,32'd351,32'd348,32'd345,32'd342,32'd339,32'd336,32'd333,32'd330,32'd327,32'd324,32'd321,32'd318,32'd315,32'd312,32'd309,32'd306,32'd303,32'd300,32'd297,32'd294,32'd291,32'd288,32'd285,32'd282,32'd279,32'd276,32'd273,32'd270,32'd267,32'd264,32'd261,32'd258,32'd255,32'd252,32'd249,32'd246,32'd243,32'd240,32'd237,32'd234,32'd231,32'd228,32'd225,32'd222,32'd219,32'd216,32'd213,32'd210,32'd207,32'd204,32'd201,32'd198,32'd195,32'd192,32'd189,32'd186,32'd183,32'd180,32'd177,32'd174,32'd171,32'd168,32'd165,32'd162,32'd159,32'd156,32'd153,32'd150,32'd147,32'd144,32'd141,32'd138,32'd135,32'd132,32'd129,32'd126,32'd123,32'd120,32'd117,32'd114,32'd111,32'd108,32'd105,32'd102,32'd99,32'd96,32'd93,32'd90,32'd87,32'd84,32'd81,32'd78,32'd75,32'd72,32'd69,32'd66,32'd63,32'd60,32'd57,32'd54,32'd51,32'd48,32'd45,32'd42,32'd39,32'd36,32'd33,32'd30,32'd27,32'd24,32'd21,32'd18,32'd15,32'd12,32'd9,32'd6,32'd3,32'd0},{32'd297,32'd295,32'd292,32'd290,32'd287,32'd285,32'd282,32'd280,32'd277,32'd275,32'd272,32'd270,32'd267,32'd265,32'd262,32'd260,32'd257,32'd255,32'd252,32'd250,32'd247,32'd245,32'd242,32'd240,32'd237,32'd235,32'd232,32'd230,32'd227,32'd225,32'd222,32'd220,32'd217,32'd215,32'd212,32'd210,32'd207,32'd205,32'd202,32'd200,32'd197,32'd195,32'd192,32'd190,32'd187,32'd185,32'd182,32'd180,32'd177,32'd175,32'd172,32'd170,32'd167,32'd165,32'd162,32'd160,32'd157,32'd155,32'd152,32'd150,32'd147,32'd145,32'd142,32'd140,32'd137,32'd135,32'd132,32'd130,32'd127,32'd125,32'd122,32'd120,32'd117,32'd115,32'd112,32'd110,32'd107,32'd105,32'd102,32'd100,32'd97,32'd95,32'd92,32'd90,32'd87,32'd85,32'd82,32'd80,32'd77,32'd75,32'd72,32'd70,32'd67,32'd65,32'd62,32'd60,32'd57,32'd55,32'd52,32'd50,32'd47,32'd45,32'd42,32'd40,32'd37,32'd35,32'd32,32'd30,32'd27,32'd25,32'd22,32'd20,32'd17,32'd15,32'd12,32'd10,32'd7,32'd5,32'd2,32'd0},{32'd250,32'd248,32'd246,32'd244,32'd242,32'd240,32'd237,32'd235,32'd233,32'd231,32'd229,32'd227,32'd225,32'd223,32'd221,32'd218,32'd216,32'd214,32'd212,32'd210,32'd208,32'd206,32'd204,32'd202,32'd200,32'd197,32'd195,32'd193,32'd191,32'd189,32'd187,32'd185,32'd183,32'd181,32'd178,32'd176,32'd174,32'd172,32'd170,32'd168,32'd166,32'd164,32'd162,32'd160,32'd157,32'd155,32'd153,32'd151,32'd149,32'd147,32'd145,32'd143,32'd141,32'd138,32'd136,32'd134,32'd132,32'd130,32'd128,32'd126,32'd124,32'd122,32'd120,32'd117,32'd115,32'd113,32'd111,32'd109,32'd107,32'd105,32'd103,32'd101,32'd98,32'd96,32'd94,32'd92,32'd90,32'd88,32'd86,32'd84,32'd82,32'd80,32'd77,32'd75,32'd73,32'd71,32'd69,32'd67,32'd65,32'd63,32'd61,32'd58,32'd56,32'd54,32'd52,32'd50,32'd48,32'd46,32'd44,32'd42,32'd40,32'd37,32'd35,32'd33,32'd31,32'd29,32'd27,32'd25,32'd23,32'd21,32'd18,32'd16,32'd14,32'd12,32'd10,32'd8,32'd6,32'd4,32'd2,32'd0},{32'd206,32'd205,32'd203,32'd201,32'd200,32'd198,32'd196,32'd194,32'd193,32'd191,32'd189,32'd187,32'd186,32'd184,32'd182,32'd180,32'd179,32'd177,32'd175,32'd173,32'd172,32'd170,32'd168,32'd166,32'd165,32'd163,32'd161,32'd160,32'd158,32'd156,32'd154,32'd153,32'd151,32'd149,32'd147,32'd146,32'd144,32'd142,32'd140,32'd139,32'd137,32'd135,32'd133,32'd132,32'd130,32'd128,32'd126,32'd125,32'd123,32'd121,32'd120,32'd118,32'd116,32'd114,32'd113,32'd111,32'd109,32'd107,32'd106,32'd104,32'd102,32'd100,32'd99,32'd97,32'd95,32'd93,32'd92,32'd90,32'd88,32'd86,32'd85,32'd83,32'd81,32'd80,32'd78,32'd76,32'd74,32'd73,32'd71,32'd69,32'd67,32'd66,32'd64,32'd62,32'd60,32'd59,32'd57,32'd55,32'd53,32'd52,32'd50,32'd48,32'd46,32'd45,32'd43,32'd41,32'd40,32'd38,32'd36,32'd34,32'd33,32'd31,32'd29,32'd27,32'd26,32'd24,32'd22,32'd20,32'd19,32'd17,32'd15,32'd13,32'd12,32'd10,32'd8,32'd6,32'd5,32'd3,32'd1,32'd0},{32'd172,32'd170,32'd169,32'd167,32'd166,32'd164,32'd163,32'd161,32'd160,32'd159,32'd157,32'd156,32'd154,32'd153,32'd151,32'd150,32'd148,32'd147,32'd146,32'd144,32'd143,32'd141,32'd140,32'd138,32'd137,32'd135,32'd134,32'd133,32'd131,32'd130,32'd128,32'd127,32'd125,32'd124,32'd122,32'd121,32'd120,32'd118,32'd117,32'd115,32'd114,32'd112,32'd111,32'd109,32'd108,32'd106,32'd105,32'd104,32'd102,32'd101,32'd99,32'd98,32'd96,32'd95,32'd93,32'd92,32'd91,32'd89,32'd88,32'd86,32'd85,32'd83,32'd82,32'd80,32'd79,32'd78,32'd76,32'd75,32'd73,32'd72,32'd70,32'd69,32'd67,32'd66,32'd65,32'd63,32'd62,32'd60,32'd59,32'd57,32'd56,32'd54,32'd53,32'd52,32'd50,32'd49,32'd47,32'd46,32'd44,32'd43,32'd41,32'd40,32'd39,32'd37,32'd36,32'd34,32'd33,32'd31,32'd30,32'd28,32'd27,32'd26,32'd24,32'd23,32'd21,32'd20,32'd18,32'd17,32'd15,32'd14,32'd13,32'd11,32'd10,32'd8,32'd7,32'd5,32'd4,32'd2,32'd1,32'd0},{32'd144,32'd143,32'd141,32'd140,32'd139,32'd138,32'd136,32'd135,32'd134,32'd133,32'd132,32'd130,32'd129,32'd128,32'd127,32'd126,32'd124,32'd123,32'd122,32'd121,32'd120,32'd118,32'd117,32'd116,32'd115,32'd113,32'd112,32'd111,32'd110,32'd109,32'd107,32'd106,32'd105,32'd104,32'd103,32'd101,32'd100,32'd99,32'd98,32'd96,32'd95,32'd94,32'd93,32'd92,32'd90,32'd89,32'd88,32'd87,32'd86,32'd84,32'd83,32'd82,32'd81,32'd80,32'd78,32'd77,32'd76,32'd75,32'd73,32'd72,32'd71,32'd70,32'd69,32'd67,32'd66,32'd65,32'd64,32'd63,32'd61,32'd60,32'd59,32'd58,32'd56,32'd55,32'd54,32'd53,32'd52,32'd50,32'd49,32'd48,32'd47,32'd46,32'd44,32'd43,32'd42,32'd41,32'd40,32'd38,32'd37,32'd36,32'd35,32'd33,32'd32,32'd31,32'd30,32'd29,32'd27,32'd26,32'd25,32'd24,32'd23,32'd21,32'd20,32'd19,32'd18,32'd16,32'd15,32'd14,32'd13,32'd12,32'd10,32'd9,32'd8,32'd7,32'd6,32'd4,32'd3,32'd2,32'd1,32'd0}}

`define STAGE_NUM_FEATURE {32'd2913,32'd2713,32'd2502,32'd2303,32'd2122,32'd1925,32'd1729,32'd1560,32'd1405,32'd1246,32'd1109,32'd973,32'd838,32'd711,32'd596,32'd497,32'd406,32'd323,32'd251,32'd189,32'd136,32'd84,32'd52,32'd25,32'd9,32'd0}
// thresholds are negative values
`define STAGE_THRESHOLD {32'd4294967143,32'd4294967123,32'd4294967129,32'd4294967126,32'd4294967128,32'd4294967132,32'd4294967130,32'd4294967122,32'd4294967112,32'd4294967116,32'd4294967121,32'd4294967106,32'd4294967113,32'd4294967106,32'd4294967098,32'd4294967109,32'd4294967099,32'd4294967097,32'd4294967090,32'd4294967085,32'd4294967071,32'd4294967068,32'd4294967058,32'd4294967041,32'd4294967038}

`define RECTANGLE1_XS {32'd9,32'd0,32'd16,32'd3,32'd12,32'd0,32'd15,32'd0,32'd3,32'd0,32'd15,32'd1,32'd15,32'd0,32'd18,32'd6,32'd0,32'd0,32'd11,32'd3,32'd13,32'd3,32'd13,32'd10,32'd14,32'd2,32'd6,32'd5,32'd15,32'd1,32'd13,32'd0,32'd16,32'd5,32'd3,32'd3,32'd15,32'd2,32'd11,32'd9,32'd5,32'd5,32'd9,32'd6,32'd12,32'd9,32'd6,32'd4,32'd5,32'd3,32'd9,32'd8,32'd14,32'd7,32'd10,32'd2,32'd6,32'd9,32'd5,32'd8,32'd8,32'd1,32'd9,32'd0,32'd5,32'd1,32'd0,32'd1,32'd10,32'd1,32'd8,32'd4,32'd4,32'd5,32'd8,32'd6,32'd0,32'd1,32'd9,32'd8,32'd10,32'd9,32'd10,32'd0,32'd7,32'd1,32'd6,32'd1,32'd9,32'd10,32'd11,32'd0,32'd12,32'd5,32'd6,32'd3,32'd15,32'd6,32'd12,32'd4,32'd0,32'd0,32'd6,32'd0,32'd2,32'd0,32'd6,32'd9,32'd12,32'd0,32'd12,32'd0,32'd6,32'd6,32'd10,32'd5,32'd12,32'd3,32'd13,32'd6,32'd16,32'd4,32'd4,32'd3,32'd4,32'd5,32'd3,32'd0,32'd5,32'd0,32'd14,32'd0,32'd15,32'd0,32'd14,32'd2,32'd12,32'd7,32'd12,32'd0,32'd3,32'd1,32'd19,32'd4,32'd19,32'd0,32'd6,32'd0,32'd0,32'd0,32'd18,32'd1,32'd11,32'd7,32'd6,32'd5,32'd9,32'd4,32'd6,32'd0,32'd11,32'd5,32'd9,32'd0,32'd17,32'd5,32'd3,32'd6,32'd10,32'd0,32'd18,32'd5,32'd6,32'd2,32'd5,32'd9,32'd9,32'd9,32'd2,32'd0,32'd5,32'd0,32'd0,32'd8,32'd6,32'd3,32'd16,32'd8,32'd9,32'd4,32'd5,32'd3,32'd11,32'd4,32'd9,32'd3,32'd12,32'd1,32'd6,32'd6,32'd9,32'd14,32'd6,32'd8,32'd0,32'd5,32'd3,32'd12,32'd9,32'd11,32'd0,32'd12,32'd3,32'd15,32'd0,32'd18,32'd0,32'd15,32'd4,32'd10,32'd2,32'd15,32'd2,32'd3,32'd7,32'd2,32'd2,32'd10,32'd5,32'd16,32'd0,32'd12,32'd10,32'd4,32'd7,32'd14,32'd9,32'd8,32'd4,32'd12,32'd0,32'd7,32'd4,32'd8,32'd8,32'd8,32'd9,32'd7,32'd6,32'd7,32'd4,32'd8,32'd0,32'd18,32'd1,32'd20,32'd0,32'd4,32'd3,32'd0,32'd0,32'd16,32'd1,32'd6,32'd3,32'd9,32'd3,32'd7,32'd7,32'd7,32'd1,32'd9,32'd0,32'd17,32'd0,32'd6,32'd8,32'd16,32'd8,32'd12,32'd9,32'd6,32'd0,32'd15,32'd3,32'd10,32'd4,32'd8,32'd3,32'd7,32'd4,32'd3,32'd2,32'd19,32'd0,32'd11,32'd0,32'd8,32'd1,32'd17,32'd2,32'd4,32'd0,32'd18,32'd3,32'd15,32'd1,32'd16,32'd4,32'd16,32'd2,32'd3,32'd0,32'd4,32'd6,32'd8,32'd3,32'd13,32'd1,32'd9,32'd7,32'd7,32'd3,32'd10,32'd7,32'd2,32'd1,32'd6,32'd5,32'd11,32'd1,32'd15,32'd9,32'd8,32'd6,32'd2,32'd5,32'd10,32'd8,32'd12,32'd3,32'd9,32'd0,32'd0,32'd0,32'd4,32'd8,32'd5,32'd7,32'd11,32'd7,32'd13,32'd7,32'd12,32'd3,32'd13,32'd3,32'd6,32'd8,32'd5,32'd6,32'd9,32'd8,32'd5,32'd5,32'd3,32'd1,32'd14,32'd2,32'd14,32'd0,32'd14,32'd7,32'd12,32'd0,32'd13,32'd0,32'd18,32'd1,32'd5,32'd10,32'd7,32'd5,32'd4,32'd8,32'd15,32'd6,32'd14,32'd0,32'd6,32'd0,32'd14,32'd0,32'd14,32'd0,32'd3,32'd5,32'd13,32'd0,32'd7,32'd4,32'd4,32'd6,32'd4,32'd0,32'd18,32'd8,32'd2,32'd0,32'd6,32'd5,32'd3,32'd5,32'd5,32'd9,32'd3,32'd6,32'd0,32'd4,32'd7,32'd10,32'd0,32'd13,32'd3,32'd12,32'd0,32'd15,32'd8,32'd15,32'd0,32'd16,32'd2,32'd9,32'd6,32'd2,32'd2,32'd16,32'd6,32'd15,32'd6,32'd15,32'd10,32'd15,32'd1,32'd15,32'd3,32'd10,32'd7,32'd6,32'd1,32'd8,32'd6,32'd6,32'd0,32'd15,32'd2,32'd4,32'd0,32'd7,32'd8,32'd12,32'd6,32'd12,32'd2,32'd1,32'd9,32'd9,32'd9,32'd14,32'd5,32'd4,32'd4,32'd12,32'd9,32'd5,32'd6,32'd12,32'd4,32'd15,32'd5,32'd11,32'd6,32'd11,32'd5,32'd15,32'd7,32'd0,32'd2,32'd17,32'd2,32'd5,32'd3,32'd14,32'd2,32'd3,32'd3,32'd13,32'd8,32'd10,32'd2,32'd2,32'd6,32'd10,32'd2,32'd13,32'd3,32'd3,32'd3,32'd0,32'd0,32'd1,32'd7,32'd13,32'd2,32'd4,32'd3,32'd10,32'd10,32'd6,32'd7,32'd12,32'd6,32'd15,32'd9,32'd6,32'd4,32'd7,32'd5,32'd16,32'd1,32'd7,32'd8,32'd6,32'd0,32'd7,32'd1,32'd13,32'd0,32'd7,32'd0,32'd10,32'd4,32'd7,32'd0,32'd20,32'd0,32'd19,32'd3,32'd9,32'd5,32'd3,32'd5,32'd13,32'd7,32'd15,32'd2,32'd7,32'd7,32'd20,32'd3,32'd14,32'd7,32'd11,32'd3,32'd15,32'd1,32'd19,32'd0,32'd6,32'd2,32'd13,32'd0,32'd14,32'd4,32'd14,32'd6,32'd10,32'd5,32'd14,32'd6,32'd9,32'd2,32'd12,32'd3,32'd13,32'd0,32'd7,32'd6,32'd0,32'd0,32'd4,32'd7,32'd13,32'd10,32'd13,32'd0,32'd8,32'd1,32'd7,32'd0,32'd9,32'd10,32'd5,32'd0,32'd18,32'd0,32'd19,32'd6,32'd0,32'd4,32'd4,32'd19,32'd0,32'd10,32'd3,32'd11,32'd0,32'd14,32'd8,32'd10,32'd2,32'd16,32'd6,32'd12,32'd8,32'd10,32'd7,32'd3,32'd0,32'd0,32'd3,32'd10,32'd6,32'd1,32'd0,32'd13,32'd7,32'd11,32'd7,32'd6,32'd5,32'd14,32'd5,32'd12,32'd2,32'd8,32'd6,32'd0,32'd9,32'd3,32'd0,32'd0,32'd5,32'd10,32'd0,32'd4,32'd7,32'd14,32'd2,32'd8,32'd3,32'd4,32'd4,32'd3,32'd2,32'd16,32'd3,32'd13,32'd7,32'd10,32'd4,32'd0,32'd0,32'd16,32'd3,32'd10,32'd2,32'd7,32'd5,32'd4,32'd4,32'd14,32'd3,32'd10,32'd7,32'd11,32'd5,32'd13,32'd2,32'd13,32'd0,32'd6,32'd0,32'd6,32'd1,32'd15,32'd2,32'd9,32'd0,32'd5,32'd10,32'd9,32'd7,32'd9,32'd7,32'd9,32'd7,32'd9,32'd1,32'd15,32'd0,32'd9,32'd7,32'd19,32'd3,32'd19,32'd1,32'd5,32'd0,32'd3,32'd0,32'd6,32'd2,32'd3,32'd2,32'd4,32'd0,32'd11,32'd0,32'd5,32'd5,32'd16,32'd0,32'd0,32'd7,32'd5,32'd2,32'd7,32'd7,32'd9,32'd5,32'd6,32'd4,32'd11,32'd1,32'd10,32'd2,32'd14,32'd9,32'd8,32'd5,32'd2,32'd9,32'd6,32'd8,32'd1,32'd5,32'd5,32'd0,32'd19,32'd2,32'd6,32'd9,32'd3,32'd0,32'd6,32'd4,32'd10,32'd7,32'd9,32'd5,32'd10,32'd2,32'd9,32'd0,32'd18,32'd5,32'd18,32'd1,32'd7,32'd9,32'd11,32'd0,32'd18,32'd2,32'd6,32'd0,32'd9,32'd3,32'd0,32'd4,32'd1,32'd4,32'd0,32'd14,32'd0,32'd14,32'd6,32'd12,32'd8,32'd12,32'd0,32'd13,32'd7,32'd11,32'd2,32'd7,32'd8,32'd7,32'd10,32'd13,32'd8,32'd1,32'd0,32'd14,32'd4,32'd6,32'd0,32'd10,32'd6,32'd5,32'd9,32'd11,32'd10,32'd10,32'd2,32'd3,32'd0,32'd6,32'd0,32'd16,32'd5,32'd17,32'd7,32'd3,32'd0,32'd11,32'd1,32'd11,32'd1,32'd11,32'd6,32'd11,32'd0,32'd20,32'd4,32'd3,32'd0,32'd6,32'd4,32'd6,32'd0,32'd4,32'd3,32'd15,32'd1,32'd6,32'd1,32'd1,32'd7,32'd0,32'd3,32'd15,32'd4,32'd14,32'd1,32'd15,32'd0,32'd7,32'd9,32'd4,32'd7,32'd13,32'd3,32'd14,32'd1,32'd13,32'd2,32'd16,32'd9,32'd9,32'd3,32'd9,32'd1,32'd1,32'd0,32'd9,32'd1,32'd7,32'd0,32'd9,32'd7,32'd7,32'd6,32'd11,32'd1,32'd7,32'd0,32'd4,32'd7,32'd11,32'd8,32'd7,32'd8,32'd10,32'd4,32'd9,32'd0,32'd5,32'd3,32'd8,32'd6,32'd14,32'd7,32'd10,32'd6,32'd10,32'd1,32'd14,32'd1,32'd4,32'd0,32'd0,32'd8,32'd6,32'd1,32'd13,32'd1,32'd9,32'd3,32'd15,32'd0,32'd14,32'd1,32'd5,32'd3,32'd15,32'd3,32'd8,32'd3,32'd15,32'd4,32'd6,32'd4,32'd2,32'd1,32'd3,32'd0,32'd19,32'd1,32'd9,32'd6,32'd7,32'd1,32'd17,32'd9,32'd4,32'd9,32'd11,32'd7,32'd11,32'd5,32'd15,32'd3,32'd14,32'd2,32'd6,32'd8,32'd7,32'd1,32'd12,32'd0,32'd11,32'd0,32'd18,32'd5,32'd13,32'd0,32'd1,32'd1,32'd11,32'd2,32'd13,32'd6,32'd10,32'd6,32'd6,32'd0,32'd9,32'd1,32'd13,32'd4,32'd12,32'd4,32'd11,32'd1,32'd0,32'd1,32'd3,32'd0,32'd11,32'd1,32'd11,32'd5,32'd6,32'd1,32'd5,32'd1,32'd12,32'd0,32'd20,32'd0,32'd10,32'd0,32'd8,32'd7,32'd11,32'd5,32'd7,32'd4,32'd9,32'd6,32'd15,32'd3,32'd11,32'd1,32'd6,32'd0,32'd12,32'd4,32'd2,32'd0,32'd14,32'd0,32'd6,32'd3,32'd16,32'd0,32'd8,32'd9,32'd10,32'd5,32'd0,32'd0,32'd12,32'd3,32'd6,32'd6,32'd10,32'd5,32'd8,32'd0,32'd5,32'd0,32'd12,32'd5,32'd16,32'd0,32'd18,32'd0,32'd15,32'd2,32'd16,32'd0,32'd12,32'd3,32'd15,32'd4,32'd17,32'd8,32'd13,32'd4,32'd14,32'd4,32'd6,32'd7,32'd11,32'd2,32'd14,32'd0,32'd11,32'd7,32'd0,32'd4,32'd9,32'd3,32'd14,32'd2,32'd5,32'd0,32'd8,32'd2,32'd10,32'd9,32'd7,32'd1,32'd1,32'd0,32'd14,32'd0,32'd3,32'd3,32'd5,32'd6,32'd7,32'd6,32'd12,32'd7,32'd8,32'd5,32'd15,32'd7,32'd10,32'd5,32'd13,32'd3,32'd13,32'd10,32'd7,32'd4,32'd10,32'd1,32'd15,32'd1,32'd11,32'd2,32'd14,32'd7,32'd10,32'd9,32'd6,32'd6,32'd12,32'd3,32'd6,32'd0,32'd15,32'd0,32'd4,32'd0,32'd6,32'd0,32'd6,32'd3,32'd5,32'd6,32'd9,32'd10,32'd6,32'd4,32'd16,32'd4,32'd3,32'd9,32'd4,32'd5,32'd14,32'd10,32'd14,32'd7,32'd7,32'd4,32'd14,32'd3,32'd9,32'd0,32'd14,32'd1,32'd17,32'd4,32'd14,32'd7,32'd14,32'd9,32'd9,32'd4,32'd2,32'd0,32'd3,32'd8,32'd5,32'd1,32'd6,32'd3,32'd8,32'd3,32'd7,32'd3,32'd7,32'd9,32'd7,32'd10,32'd1,32'd2,32'd2,32'd0,32'd1,32'd10,32'd6,32'd0,32'd0,32'd13,32'd0,32'd8,32'd4,32'd16,32'd0,32'd14,32'd5,32'd14,32'd5,32'd10,32'd9,32'd6,32'd9,32'd9,32'd0,32'd4,32'd5,32'd7,32'd6,32'd5,32'd8,32'd10,32'd5,32'd2,32'd3,32'd1,32'd0,32'd12,32'd9,32'd9,32'd0,32'd2,32'd0,32'd6,32'd5,32'd11,32'd6,32'd6,32'd7,32'd1,32'd5,32'd11,32'd5,32'd6,32'd4,32'd11,32'd9,32'd5,32'd6,32'd3,32'd1,32'd12,32'd1,32'd15,32'd0,32'd13,32'd5,32'd17,32'd3,32'd2,32'd1,32'd7,32'd5,32'd16,32'd3,32'd11,32'd5,32'd13,32'd0,32'd18,32'd3,32'd18,32'd6,32'd12,32'd7,32'd9,32'd9,32'd3,32'd4,32'd3,32'd8,32'd14,32'd3,32'd4,32'd8,32'd13,32'd7,32'd1,32'd8,32'd4,32'd2,32'd14,32'd4,32'd11,32'd8,32'd10,32'd4,32'd8,32'd5,32'd0,32'd0,32'd13,32'd0,32'd16,32'd3,32'd9,32'd0,32'd15,32'd0,32'd17,32'd4,32'd15,32'd2,32'd9,32'd0,32'd15,32'd2,32'd9,32'd1,32'd13,32'd6,32'd12,32'd1,32'd9,32'd0,32'd9,32'd11,32'd8,32'd8,32'd12,32'd8,32'd9,32'd2,32'd13,32'd5,32'd13,32'd3,32'd3,32'd0,32'd0,32'd8,32'd20,32'd4,32'd13,32'd2,32'd9,32'd0,32'd9,32'd0,32'd2,32'd7,32'd1,32'd13,32'd6,32'd10,32'd8,32'd12,32'd3,32'd12,32'd3,32'd12,32'd1,32'd16,32'd0,32'd17,32'd9,32'd7,32'd10,32'd4,32'd2,32'd0,32'd0,32'd8,32'd2,32'd11,32'd0,32'd8,32'd6,32'd4,32'd3,32'd9,32'd8,32'd10,32'd5,32'd6,32'd4,32'd9,32'd7,32'd10,32'd0,32'd12,32'd2,32'd1,32'd1,32'd6,32'd4,32'd18,32'd1,32'd6,32'd0,32'd10,32'd4,32'd0,32'd4,32'd10,32'd5,32'd11,32'd1,32'd15,32'd7,32'd15,32'd4,32'd3,32'd2,32'd10,32'd3,32'd17,32'd4,32'd7,32'd8,32'd10,32'd9,32'd7,32'd6,32'd10,32'd0,32'd14,32'd8,32'd6,32'd6,32'd15,32'd1,32'd10,32'd0,32'd12,32'd0,32'd14,32'd1,32'd3,32'd7,32'd14,32'd1,32'd17,32'd8,32'd9,32'd6,32'd14,32'd6,32'd10,32'd6,32'd13,32'd1,32'd2,32'd9,32'd11,32'd6,32'd10,32'd10,32'd0,32'd2,32'd2,32'd0,32'd1,32'd0,32'd3,32'd3,32'd0,32'd0,32'd15,32'd4,32'd14,32'd6,32'd5,32'd0,32'd18,32'd1,32'd3,32'd1,32'd14,32'd3,32'd14,32'd8,32'd14,32'd2,32'd10,32'd10,32'd7,32'd7,32'd15,32'd11,32'd5,32'd2,32'd18,32'd0,32'd18,32'd5,32'd6,32'd7,32'd9,32'd6,32'd2,32'd4,32'd14,32'd6,32'd7,32'd0,32'd0,32'd2,32'd2,32'd8,32'd6,32'd14,32'd6,32'd8,32'd8,32'd5,32'd9,32'd7,32'd8,32'd10,32'd5,32'd9,32'd2,32'd3,32'd0,32'd18,32'd1,32'd17,32'd0,32'd19,32'd3,32'd0,32'd4,32'd10,32'd7,32'd10,32'd6,32'd9,32'd1,32'd15,32'd1,32'd9,32'd3,32'd11,32'd2,32'd3,32'd5,32'd9,32'd5,32'd13,32'd2,32'd8,32'd0,32'd12,32'd6,32'd7,32'd7,32'd4,32'd2,32'd18,32'd3,32'd4,32'd9,32'd4,32'd2,32'd7,32'd6,32'd3,32'd0,32'd18,32'd0,32'd22,32'd7,32'd15,32'd0,32'd11,32'd1,32'd18,32'd3,32'd16,32'd4,32'd14,32'd1,32'd8,32'd0,32'd15,32'd5,32'd4,32'd0,32'd9,32'd8,32'd14,32'd3,32'd16,32'd2,32'd12,32'd4,32'd13,32'd1,32'd14,32'd0,32'd6,32'd0,32'd3,32'd0,32'd8,32'd0,32'd16,32'd1,32'd6,32'd9,32'd11,32'd7,32'd9,32'd5,32'd10,32'd8,32'd9,32'd5,32'd9,32'd3,32'd9,32'd0,32'd5,32'd0,32'd15,32'd0,32'd15,32'd3,32'd15,32'd7,32'd10,32'd0,32'd0,32'd0,32'd17,32'd0,32'd18,32'd1,32'd2,32'd0,32'd11,32'd0,32'd18,32'd0,32'd6,32'd6,32'd10,32'd0,32'd3,32'd6,32'd11,32'd5,32'd13,32'd1,32'd7,32'd2,32'd4,32'd5,32'd11,32'd6,32'd3,32'd9,32'd0,32'd4,32'd10,32'd10,32'd0,32'd0,32'd0,32'd16,32'd3,32'd6,32'd5,32'd5,32'd7,32'd10,32'd0,32'd7,32'd3,32'd8,32'd10,32'd7,32'd1,32'd10,32'd0,32'd15,32'd0,32'd15,32'd4,32'd15,32'd3,32'd15,32'd2,32'd10,32'd4,32'd8,32'd7,32'd2,32'd1,32'd9,32'd0,32'd18,32'd0,32'd8,32'd2,32'd8,32'd10,32'd4,32'd5,32'd9,32'd3,32'd0,32'd6,32'd12,32'd0,32'd18,32'd0,32'd6,32'd5,32'd13,32'd6,32'd6,32'd5,32'd2,32'd2,32'd3,32'd0,32'd18,32'd5,32'd5,32'd5,32'd13,32'd0,32'd2,32'd0,32'd3,32'd3,32'd17,32'd7,32'd15,32'd9,32'd9,32'd3,32'd16,32'd3,32'd12,32'd0,32'd2,32'd1,32'd18,32'd4,32'd14,32'd4,32'd14,32'd1,32'd5,32'd1,32'd5,32'd2,32'd13,32'd0,32'd15,32'd7,32'd16,32'd3,32'd10,32'd9,32'd15,32'd1,32'd11,32'd6,32'd12,32'd5,32'd14,32'd7,32'd10,32'd10,32'd11,32'd5,32'd16,32'd7,32'd8,32'd0,32'd20,32'd1,32'd0,32'd4,32'd14,32'd6,32'd14,32'd4,32'd14,32'd1,32'd19,32'd2,32'd3,32'd8,32'd15,32'd9,32'd6,32'd3,32'd2,32'd0,32'd7,32'd2,32'd4,32'd5,32'd2,32'd9,32'd1,32'd5,32'd0,32'd0,32'd0,32'd2,32'd12,32'd6,32'd7,32'd5,32'd10,32'd3,32'd12,32'd3,32'd10,32'd10,32'd7,32'd3,32'd8,32'd1,32'd9,32'd9,32'd12,32'd4,32'd8,32'd0,32'd12,32'd3,32'd8,32'd1,32'd9,32'd5,32'd14,32'd6,32'd5,32'd0,32'd12,32'd1,32'd12,32'd2,32'd12,32'd0,32'd1,32'd7,32'd10,32'd10,32'd5,32'd5,32'd11,32'd8,32'd5,32'd0,32'd10,32'd0,32'd4,32'd3,32'd3,32'd2,32'd3,32'd9,32'd11,32'd6,32'd11,32'd6,32'd10,32'd6,32'd15,32'd1,32'd15,32'd3,32'd15,32'd8,32'd12,32'd9,32'd7,32'd4,32'd16,32'd0,32'd9,32'd1,32'd15,32'd0,32'd7,32'd1,32'd17,32'd2,32'd2,32'd1,32'd8,32'd0,32'd13,32'd5,32'd12,32'd5,32'd11,32'd1,32'd10,32'd6,32'd6,32'd3,32'd5,32'd5,32'd13,32'd0,32'd15,32'd0,32'd20,32'd0,32'd6,32'd0,32'd6,32'd8,32'd20,32'd0,32'd6,32'd0,32'd4,32'd5,32'd8,32'd0,32'd16,32'd0,32'd16,32'd3,32'd9,32'd1,32'd1,32'd7,32'd2,32'd17,32'd6,32'd9,32'd1,32'd8,32'd6,32'd10,32'd9,32'd6,32'd1,32'd18,32'd2,32'd5,32'd7,32'd10,32'd8,32'd8,32'd9,32'd16,32'd0,32'd4,32'd5,32'd9,32'd9,32'd1,32'd5,32'd13,32'd0,32'd6,32'd0,32'd9,32'd8,32'd5,32'd3,32'd8,32'd1,32'd3,32'd7,32'd13,32'd2,32'd4,32'd7,32'd11,32'd9,32'd10,32'd4,32'd18,32'd9,32'd10,32'd5,32'd7,32'd2,32'd3,32'd0,32'd0,32'd7,32'd6,32'd4,32'd5,32'd3,32'd8,32'd1,32'd10,32'd6,32'd8,32'd3,32'd1,32'd5,32'd2,32'd0,32'd5,32'd1,32'd19,32'd2,32'd13,32'd7,32'd3,32'd5,32'd5,32'd5,32'd12,32'd0,32'd12,32'd0,32'd6,32'd4,32'd11,32'd5,32'd13,32'd0,32'd13,32'd0,32'd6,32'd9,32'd18,32'd7,32'd9,32'd6,32'd13,32'd2,32'd3,32'd2,32'd18,32'd0,32'd10,32'd6,32'd8,32'd9,32'd5,32'd2,32'd11,32'd2,32'd6,32'd8,32'd4,32'd5,32'd1,32'd0,32'd14,32'd0,32'd0,32'd0,32'd20,32'd0,32'd6,32'd0,32'd8,32'd3,32'd8,32'd2,32'd9,32'd7,32'd2,32'd4,32'd5,32'd11,32'd5,32'd11,32'd7,32'd11,32'd2,32'd8,32'd1,32'd6,32'd1,32'd9,32'd9,32'd11,32'd1,32'd3,32'd0,32'd11,32'd3,32'd7,32'd2,32'd12,32'd8,32'd13,32'd2,32'd5,32'd9,32'd4,32'd10,32'd3,32'd8,32'd10,32'd9,32'd11,32'd0,32'd6,32'd5,32'd13,32'd6,32'd15,32'd1,32'd13,32'd6,32'd12,32'd8,32'd10,32'd8,32'd6,32'd0,32'd15,32'd1,32'd0,32'd2,32'd0,32'd5,32'd13,32'd0,32'd15,32'd0,32'd13,32'd0,32'd12,32'd7,32'd3,32'd1,32'd13,32'd2,32'd3,32'd1,32'd15,32'd4,32'd12,32'd0,32'd13,32'd1,32'd1,32'd0,32'd9,32'd7,32'd12,32'd0,32'd16,32'd0,32'd19,32'd1,32'd0,32'd5,32'd13,32'd8,32'd9,32'd0,32'd4,32'd9,32'd10,32'd8,32'd12,32'd0,32'd3,32'd10,32'd3,32'd3,32'd11,32'd1,32'd10,32'd2,32'd16,32'd0,32'd15,32'd1,32'd20,32'd0,32'd10,32'd2,32'd15,32'd7,32'd17,32'd8,32'd17,32'd1,32'd8,32'd5,32'd15,32'd0,32'd12,32'd1,32'd6,32'd2,32'd4,32'd10,32'd5,32'd16,32'd3,32'd7,32'd2,32'd4,32'd8,32'd10,32'd0,32'd7,32'd0,32'd18,32'd0,32'd19,32'd0,32'd1,32'd2,32'd20,32'd3,32'd18,32'd2,32'd9,32'd3,32'd7,32'd1,32'd5,32'd6,32'd2,32'd2,32'd14,32'd0,32'd2,32'd8,32'd12,32'd3,32'd9,32'd1,32'd8,32'd5,32'd11,32'd9,32'd12,32'd4,32'd14,32'd5,32'd13,32'd1,32'd8,32'd7,32'd7,32'd0,32'd12,32'd7,32'd13,32'd1,32'd5,32'd0,32'd14,32'd6,32'd14,32'd2,32'd12,32'd7,32'd11,32'd10,32'd11,32'd1,32'd14,32'd6,32'd6,32'd3,32'd1,32'd1,32'd5,32'd1,32'd3,32'd0,32'd5,32'd0,32'd3,32'd5,32'd8,32'd7,32'd8,32'd6,32'd14,32'd8,32'd10,32'd2,32'd13,32'd0,32'd11,32'd4,32'd14,32'd6,32'd7,32'd5,32'd13,32'd4,32'd13,32'd0,32'd13,32'd0,32'd9,32'd3,32'd18,32'd0,32'd11,32'd5,32'd6,32'd3,32'd0,32'd7,32'd2,32'd12,32'd0,32'd0,32'd3,32'd3,32'd0,32'd10,32'd6,32'd11,32'd0,32'd15,32'd6,32'd12,32'd9,32'd12,32'd0,32'd15,32'd0,32'd10,32'd10,32'd5,32'd6,32'd8,32'd3,32'd15,32'd0,32'd15,32'd6,32'd4,32'd1,32'd19,32'd1,32'd17,32'd3,32'd15,32'd2,32'd8,32'd3,32'd6,32'd0,32'd5,32'd7,32'd13,32'd0,32'd10,32'd0,32'd16,32'd3,32'd16,32'd6,32'd11,32'd10,32'd0,32'd3,32'd3,32'd6,32'd14,32'd6,32'd12,32'd7,32'd11,32'd0,32'd15,32'd10,32'd21,32'd7,32'd8,32'd6,32'd21,32'd5,32'd18,32'd0,32'd14,32'd2,32'd4,32'd0,32'd18,32'd9,32'd3,32'd2,32'd17,32'd0,32'd15,32'd1,32'd14,32'd9,32'd14,32'd0,32'd5,32'd8,32'd10,32'd0,32'd3,32'd3,32'd1,32'd0,32'd6,32'd6,32'd8,32'd10,32'd5,32'd2,32'd4,32'd16,32'd10,32'd12,32'd7,32'd6,32'd3,32'd12,32'd8,32'd9,32'd11,32'd12,32'd0,32'd15,32'd2,32'd12,32'd5,32'd0,32'd4,32'd16,32'd5,32'd13,32'd1,32'd9,32'd7,32'd13,32'd0,32'd6,32'd3,32'd5,32'd0,32'd0,32'd0,32'd14,32'd0,32'd14,32'd6,32'd2,32'd3,32'd0,32'd5,32'd1,32'd4,32'd6,32'd1,32'd0,32'd0,32'd5,32'd5,32'd10,32'd1,32'd6,32'd6,32'd12,32'd9,32'd3,32'd6,32'd14,32'd1,32'd17,32'd0,32'd9,32'd0,32'd18,32'd7,32'd18,32'd6,32'd18,32'd2,32'd14,32'd7,32'd13,32'd7,32'd9,32'd1,32'd9,32'd6,32'd8,32'd0,32'd20,32'd3,32'd3,32'd0,32'd9,32'd5,32'd14,32'd0,32'd8,32'd6,32'd3,32'd9,32'd9,32'd10,32'd0,32'd16,32'd4,32'd5,32'd1,32'd14,32'd0,32'd16,32'd0,32'd6,32'd9,32'd8,32'd0,32'd6,32'd1,32'd6,32'd0,32'd15,32'd2,32'd10,32'd4,32'd12,32'd7,32'd16,32'd1,32'd17,32'd6,32'd14,32'd2,32'd4,32'd0,32'd15,32'd3,32'd15,32'd3,32'd15,32'd0,32'd10,32'd1,32'd4,32'd1,32'd14,32'd1,32'd18,32'd7,32'd13,32'd4,32'd15,32'd8,32'd8,32'd2,32'd15,32'd3,32'd15,32'd8,32'd10,32'd6,32'd5,32'd0,32'd18,32'd3,32'd18,32'd0,32'd18,32'd7,32'd16,32'd8,32'd3,32'd2,32'd3,32'd7,32'd11,32'd4,32'd5,32'd6,32'd6,32'd0,32'd10,32'd3,32'd10,32'd1,32'd12,32'd1,32'd12,32'd6,32'd3,32'd9,32'd12,32'd9,32'd5,32'd2,32'd14,32'd7,32'd9,32'd5,32'd15,32'd6,32'd12,32'd7,32'd11,32'd8,32'd8,32'd0,32'd18,32'd0,32'd9,32'd4,32'd0,32'd2,32'd14,32'd5,32'd7,32'd10,32'd9,32'd0,32'd3,32'd0,32'd8,32'd0,32'd15,32'd7,32'd15,32'd0,32'd15,32'd0,32'd7,32'd8,32'd7,32'd7,32'd6,32'd6,32'd12,32'd7,32'd13,32'd1,32'd14,32'd6,32'd12,32'd3,32'd15,32'd0,32'd10,32'd1,32'd7,32'd3,32'd17,32'd9,32'd15,32'd3,32'd14,32'd1,32'd17,32'd5,32'd9,32'd2,32'd0,32'd4,32'd1,32'd0,32'd10,32'd1,32'd5,32'd9,32'd13,32'd4,32'd3,32'd0,32'd3,32'd7,32'd7,32'd0,32'd7,32'd4,32'd9,32'd0,32'd3,32'd2,32'd13,32'd8,32'd11,32'd7,32'd13,32'd0,32'd11,32'd1,32'd18,32'd3,32'd18,32'd6,32'd11,32'd7,32'd9,32'd0,32'd2,32'd2,32'd1,32'd0,32'd6,32'd0,32'd5,32'd0,32'd5,32'd2,32'd20,32'd9,32'd5,32'd1,32'd10,32'd7,32'd6,32'd0,32'd0,32'd9,32'd3,32'd13,32'd6,32'd17,32'd8,32'd14,32'd8,32'd14,32'd2,32'd2,32'd0,32'd7,32'd6,32'd12,32'd5,32'd1,32'd0,32'd7,32'd6,32'd8,32'd5,32'd10,32'd1,32'd10,32'd4,32'd10,32'd7,32'd14,32'd1,32'd0,32'd7,32'd8,32'd0,32'd15,32'd5,32'd14,32'd2,32'd9,32'd2,32'd16,32'd0,32'd18,32'd0,32'd18,32'd7,32'd4,32'd0,32'd9,32'd7,32'd6,32'd0,32'd19,32'd0,32'd12,32'd0,32'd8,32'd1,32'd3,32'd6,32'd6,32'd0,32'd3,32'd6,32'd4,32'd4,32'd9,32'd5,32'd3,32'd2,32'd2,32'd3,32'd10,32'd0,32'd8,32'd6,32'd12,32'd0,32'd11,32'd5,32'd12,32'd0,32'd2,32'd0,32'd20,32'd2,32'd6,32'd1,32'd6,32'd0,32'd7,32'd6,32'd10,32'd1,32'd9,32'd9,32'd11,32'd4,32'd11,32'd0,32'd11,32'd4,32'd0,32'd6,32'd3,32'd8,32'd10,32'd7,32'd9,32'd9,32'd6,32'd5,32'd11,32'd1,32'd14,32'd3,32'd5,32'd1,32'd3,32'd0,32'd4,32'd1,32'd15,32'd8,32'd6,32'd3,32'd14,32'd1,32'd0,32'd1,32'd19,32'd2,32'd4,32'd0,32'd6,32'd6,32'd0,32'd17,32'd1,32'd5,32'd8,32'd12,32'd0,32'd12,32'd0,32'd18,32'd0,32'd20,32'd0,32'd2,32'd8,32'd2,32'd5,32'd0,32'd1,32'd18,32'd5,32'd3,32'd6,32'd9,32'd9,32'd5,32'd0,32'd5,32'd7,32'd9,32'd0,32'd18,32'd2,32'd10,32'd7,32'd13,32'd5,32'd5,32'd9,32'd0,32'd1,32'd6,32'd6,32'd4,32'd11,32'd5,32'd6,32'd3,32'd8,32'd3,32'd6,32'd6}
`define RECTANGLE1_YS {32'd1,32'd13,32'd2,32'd17,32'd17,32'd17,32'd17,32'd13,32'd15,32'd18,32'd17,32'd6,32'd17,32'd12,32'd12,32'd20,32'd16,32'd18,32'd14,32'd8,32'd8,32'd10,32'd11,32'd1,32'd12,32'd11,32'd11,32'd8,32'd8,32'd13,32'd13,32'd8,32'd8,32'd0,32'd20,32'd1,32'd1,32'd0,32'd9,32'd9,32'd8,32'd9,32'd1,32'd0,32'd0,32'd0,32'd9,32'd0,32'd2,32'd1,32'd2,32'd5,32'd5,32'd5,32'd6,32'd6,32'd8,32'd3,32'd4,32'd6,32'd14,32'd20,32'd17,32'd16,32'd17,32'd14,32'd4,32'd5,32'd5,32'd7,32'd5,32'd4,32'd4,32'd2,32'd9,32'd14,32'd3,32'd0,32'd1,32'd0,32'd6,32'd5,32'd0,32'd0,32'd7,32'd8,32'd9,32'd10,32'd12,32'd2,32'd2,32'd11,32'd11,32'd8,32'd12,32'd10,32'd10,32'd14,32'd8,32'd10,32'd12,32'd3,32'd3,32'd0,32'd5,32'd5,32'd14,32'd6,32'd6,32'd14,32'd6,32'd8,32'd8,32'd4,32'd5,32'd11,32'd6,32'd14,32'd14,32'd4,32'd4,32'd3,32'd12,32'd0,32'd0,32'd3,32'd5,32'd18,32'd18,32'd14,32'd14,32'd14,32'd14,32'd0,32'd0,32'd16,32'd16,32'd18,32'd18,32'd19,32'd21,32'd6,32'd6,32'd6,32'd0,32'd0,32'd7,32'd5,32'd6,32'd8,32'd8,32'd11,32'd5,32'd9,32'd1,32'd6,32'd7,32'd6,32'd16,32'd16,32'd6,32'd11,32'd11,32'd0,32'd0,32'd2,32'd2,32'd5,32'd5,32'd3,32'd3,32'd0,32'd0,32'd6,32'd11,32'd12,32'd15,32'd13,32'd1,32'd6,32'd10,32'd20,32'd16,32'd6,32'd6,32'd9,32'd9,32'd6,32'd6,32'd2,32'd3,32'd9,32'd3,32'd13,32'd18,32'd12,32'd12,32'd1,32'd5,32'd4,32'd1,32'd1,32'd2,32'd14,32'd13,32'd5,32'd4,32'd1,32'd0,32'd6,32'd2,32'd2,32'd0,32'd0,32'd0,32'd0,32'd8,32'd8,32'd4,32'd9,32'd2,32'd6,32'd7,32'd2,32'd6,32'd8,32'd18,32'd15,32'd0,32'd0,32'd0,32'd1,32'd2,32'd7,32'd0,32'd0,32'd1,32'd11,32'd7,32'd17,32'd2,32'd6,32'd3,32'd2,32'd14,32'd2,32'd8,32'd6,32'd3,32'd6,32'd6,32'd18,32'd8,32'd8,32'd3,32'd2,32'd1,32'd2,32'd2,32'd9,32'd7,32'd7,32'd10,32'd10,32'd2,32'd8,32'd8,32'd8,32'd7,32'd6,32'd6,32'd6,32'd13,32'd0,32'd18,32'd6,32'd1,32'd6,32'd15,32'd1,32'd10,32'd7,32'd10,32'd10,32'd8,32'd14,32'd14,32'd15,32'd13,32'd13,32'd4,32'd10,32'd1,32'd1,32'd4,32'd12,32'd6,32'd8,32'd6,32'd0,32'd1,32'd7,32'd5,32'd5,32'd9,32'd12,32'd4,32'd0,32'd0,32'd0,32'd4,32'd17,32'd17,32'd6,32'd7,32'd7,32'd16,32'd4,32'd0,32'd19,32'd12,32'd8,32'd9,32'd5,32'd6,32'd8,32'd12,32'd1,32'd0,32'd0,32'd14,32'd14,32'd6,32'd7,32'd11,32'd0,32'd0,32'd6,32'd0,32'd1,32'd3,32'd0,32'd15,32'd1,32'd3,32'd17,32'd9,32'd7,32'd15,32'd9,32'd0,32'd0,32'd7,32'd1,32'd3,32'd0,32'd1,32'd11,32'd2,32'd6,32'd1,32'd1,32'd2,32'd0,32'd13,32'd15,32'd13,32'd13,32'd4,32'd4,32'd9,32'd0,32'd3,32'd9,32'd2,32'd3,32'd1,32'd1,32'd20,32'd20,32'd6,32'd7,32'd8,32'd20,32'd13,32'd8,32'd2,32'd13,32'd18,32'd16,32'd16,32'd13,32'd16,32'd16,32'd2,32'd10,32'd11,32'd11,32'd1,32'd9,32'd12,32'd7,32'd0,32'd6,32'd0,32'd1,32'd17,32'd12,32'd1,32'd6,32'd0,32'd0,32'd1,32'd9,32'd1,32'd4,32'd9,32'd21,32'd1,32'd0,32'd0,32'd1,32'd15,32'd10,32'd10,32'd15,32'd15,32'd6,32'd17,32'd7,32'd7,32'd11,32'd0,32'd5,32'd1,32'd4,32'd7,32'd5,32'd17,32'd1,32'd17,32'd3,32'd17,32'd12,32'd17,32'd14,32'd12,32'd7,32'd6,32'd9,32'd7,32'd6,32'd0,32'd15,32'd15,32'd13,32'd13,32'd1,32'd2,32'd7,32'd7,32'd5,32'd6,32'd7,32'd4,32'd4,32'd5,32'd10,32'd8,32'd4,32'd6,32'd5,32'd6,32'd1,32'd9,32'd6,32'd6,32'd7,32'd7,32'd8,32'd4,32'd1,32'd13,32'd1,32'd1,32'd16,32'd17,32'd12,32'd8,32'd15,32'd4,32'd21,32'd17,32'd4,32'd9,32'd11,32'd8,32'd8,32'd8,32'd11,32'd2,32'd0,32'd2,32'd0,32'd0,32'd1,32'd6,32'd2,32'd0,32'd0,32'd4,32'd0,32'd0,32'd15,32'd14,32'd18,32'd8,32'd6,32'd0,32'd2,32'd7,32'd0,32'd0,32'd2,32'd5,32'd9,32'd6,32'd4,32'd4,32'd1,32'd1,32'd10,32'd19,32'd10,32'd1,32'd11,32'd0,32'd13,32'd2,32'd1,32'd11,32'd19,32'd7,32'd4,32'd4,32'd8,32'd8,32'd16,32'd5,32'd6,32'd5,32'd12,32'd12,32'd0,32'd0,32'd1,32'd0,32'd6,32'd4,32'd6,32'd6,32'd9,32'd6,32'd20,32'd0,32'd2,32'd2,32'd16,32'd16,32'd18,32'd18,32'd20,32'd15,32'd9,32'd9,32'd6,32'd8,32'd14,32'd6,32'd6,32'd6,32'd15,32'd14,32'd18,32'd15,32'd3,32'd8,32'd4,32'd18,32'd0,32'd13,32'd11,32'd9,32'd5,32'd9,32'd10,32'd2,32'd7,32'd3,32'd21,32'd6,32'd7,32'd15,32'd0,32'd0,32'd6,32'd3,32'd8,32'd1,32'd7,32'd12,32'd2,32'd15,32'd1,32'd2,32'd17,32'd20,32'd20,32'd15,32'd15,32'd12,32'd12,32'd10,32'd10,32'd6,32'd16,32'd12,32'd3,32'd11,32'd6,32'd8,32'd0,32'd6,32'd12,32'd12,32'd14,32'd0,32'd2,32'd7,32'd9,32'd8,32'd2,32'd0,32'd0,32'd7,32'd8,32'd18,32'd5,32'd11,32'd0,32'd5,32'd8,32'd0,32'd13,32'd13,32'd10,32'd14,32'd14,32'd16,32'd18,32'd10,32'd9,32'd12,32'd6,32'd1,32'd1,32'd0,32'd10,32'd0,32'd8,32'd7,32'd7,32'd0,32'd0,32'd4,32'd0,32'd2,32'd2,32'd6,32'd5,32'd0,32'd0,32'd4,32'd0,32'd5,32'd5,32'd1,32'd1,32'd15,32'd15,32'd16,32'd18,32'd18,32'd4,32'd10,32'd16,32'd17,32'd10,32'd1,32'd5,32'd5,32'd8,32'd6,32'd8,32'd8,32'd8,32'd8,32'd8,32'd5,32'd16,32'd6,32'd13,32'd15,32'd4,32'd7,32'd4,32'd21,32'd21,32'd14,32'd14,32'd9,32'd7,32'd3,32'd0,32'd16,32'd16,32'd0,32'd4,32'd1,32'd6,32'd1,32'd0,32'd2,32'd10,32'd1,32'd1,32'd5,32'd6,32'd8,32'd16,32'd4,32'd5,32'd6,32'd3,32'd3,32'd18,32'd14,32'd14,32'd12,32'd6,32'd4,32'd0,32'd6,32'd17,32'd15,32'd2,32'd2,32'd0,32'd1,32'd4,32'd3,32'd2,32'd6,32'd20,32'd7,32'd7,32'd1,32'd6,32'd0,32'd0,32'd6,32'd6,32'd2,32'd12,32'd2,32'd2,32'd1,32'd1,32'd3,32'd7,32'd6,32'd14,32'd12,32'd12,32'd12,32'd22,32'd17,32'd6,32'd6,32'd1,32'd0,32'd6,32'd6,32'd12,32'd12,32'd6,32'd5,32'd8,32'd8,32'd1,32'd8,32'd19,32'd4,32'd16,32'd16,32'd14,32'd1,32'd1,32'd8,32'd6,32'd2,32'd9,32'd10,32'd11,32'd12,32'd3,32'd5,32'd0,32'd16,32'd4,32'd9,32'd1,32'd1,32'd6,32'd5,32'd11,32'd7,32'd14,32'd0,32'd1,32'd1,32'd0,32'd1,32'd14,32'd7,32'd1,32'd1,32'd0,32'd1,32'd16,32'd1,32'd21,32'd1,32'd14,32'd14,32'd6,32'd2,32'd10,32'd10,32'd12,32'd18,32'd10,32'd14,32'd15,32'd15,32'd17,32'd18,32'd17,32'd0,32'd1,32'd2,32'd0,32'd0,32'd5,32'd5,32'd0,32'd0,32'd3,32'd7,32'd10,32'd7,32'd1,32'd1,32'd12,32'd7,32'd8,32'd1,32'd0,32'd0,32'd6,32'd14,32'd19,32'd1,32'd6,32'd5,32'd5,32'd12,32'd13,32'd3,32'd6,32'd1,32'd8,32'd5,32'd0,32'd16,32'd10,32'd3,32'd16,32'd22,32'd7,32'd2,32'd2,32'd3,32'd3,32'd14,32'd1,32'd1,32'd0,32'd4,32'd6,32'd7,32'd4,32'd4,32'd5,32'd5,32'd8,32'd10,32'd10,32'd0,32'd15,32'd9,32'd1,32'd0,32'd14,32'd19,32'd19,32'd19,32'd18,32'd5,32'd13,32'd13,32'd15,32'd15,32'd13,32'd9,32'd7,32'd7,32'd15,32'd18,32'd18,32'd6,32'd4,32'd0,32'd1,32'd1,32'd5,32'd5,32'd0,32'd4,32'd1,32'd14,32'd18,32'd13,32'd17,32'd1,32'd13,32'd1,32'd5,32'd5,32'd0,32'd0,32'd6,32'd6,32'd5,32'd15,32'd19,32'd6,32'd2,32'd6,32'd13,32'd14,32'd1,32'd7,32'd2,32'd2,32'd0,32'd0,32'd17,32'd10,32'd20,32'd2,32'd10,32'd0,32'd12,32'd10,32'd5,32'd4,32'd1,32'd10,32'd15,32'd10,32'd12,32'd12,32'd12,32'd12,32'd12,32'd9,32'd10,32'd10,32'd8,32'd14,32'd15,32'd12,32'd6,32'd10,32'd12,32'd7,32'd8,32'd6,32'd9,32'd2,32'd13,32'd13,32'd2,32'd1,32'd0,32'd0,32'd0,32'd7,32'd4,32'd5,32'd3,32'd3,32'd0,32'd9,32'd6,32'd13,32'd15,32'd8,32'd3,32'd3,32'd12,32'd3,32'd0,32'd18,32'd16,32'd16,32'd4,32'd2,32'd3,32'd0,32'd1,32'd14,32'd15,32'd0,32'd2,32'd9,32'd0,32'd2,32'd4,32'd10,32'd15,32'd7,32'd9,32'd9,32'd10,32'd0,32'd1,32'd1,32'd6,32'd6,32'd0,32'd0,32'd2,32'd2,32'd0,32'd0,32'd12,32'd0,32'd3,32'd9,32'd10,32'd10,32'd13,32'd6,32'd6,32'd14,32'd7,32'd12,32'd12,32'd0,32'd8,32'd5,32'd8,32'd2,32'd6,32'd2,32'd6,32'd5,32'd5,32'd3,32'd18,32'd18,32'd15,32'd8,32'd16,32'd19,32'd16,32'd16,32'd0,32'd8,32'd1,32'd6,32'd3,32'd7,32'd2,32'd2,32'd2,32'd1,32'd4,32'd1,32'd3,32'd6,32'd15,32'd15,32'd21,32'd15,32'd14,32'd17,32'd0,32'd1,32'd2,32'd1,32'd4,32'd1,32'd0,32'd9,32'd8,32'd7,32'd0,32'd16,32'd0,32'd0,32'd17,32'd15,32'd14,32'd14,32'd3,32'd3,32'd15,32'd18,32'd0,32'd0,32'd6,32'd6,32'd7,32'd15,32'd5,32'd6,32'd0,32'd16,32'd13,32'd0,32'd6,32'd4,32'd20,32'd13,32'd6,32'd13,32'd2,32'd6,32'd10,32'd7,32'd10,32'd5,32'd0,32'd13,32'd1,32'd1,32'd0,32'd0,32'd16,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd21,32'd8,32'd8,32'd0,32'd0,32'd0,32'd0,32'd12,32'd7,32'd14,32'd1,32'd8,32'd7,32'd14,32'd18,32'd11,32'd15,32'd2,32'd1,32'd16,32'd16,32'd9,32'd11,32'd11,32'd17,32'd18,32'd15,32'd0,32'd2,32'd11,32'd9,32'd9,32'd6,32'd0,32'd4,32'd17,32'd10,32'd15,32'd8,32'd1,32'd2,32'd4,32'd0,32'd18,32'd14,32'd14,32'd0,32'd5,32'd0,32'd1,32'd0,32'd0,32'd1,32'd0,32'd4,32'd7,32'd5,32'd4,32'd2,32'd2,32'd7,32'd11,32'd9,32'd10,32'd15,32'd18,32'd1,32'd0,32'd1,32'd2,32'd3,32'd10,32'd3,32'd21,32'd13,32'd1,32'd0,32'd13,32'd12,32'd0,32'd2,32'd0,32'd10,32'd5,32'd21,32'd21,32'd6,32'd4,32'd9,32'd9,32'd7,32'd11,32'd2,32'd2,32'd5,32'd2,32'd1,32'd1,32'd0,32'd7,32'd1,32'd21,32'd13,32'd2,32'd0,32'd0,32'd10,32'd22,32'd1,32'd3,32'd0,32'd9,32'd7,32'd4,32'd4,32'd6,32'd5,32'd5,32'd4,32'd2,32'd3,32'd9,32'd2,32'd14,32'd13,32'd18,32'd14,32'd13,32'd15,32'd18,32'd17,32'd17,32'd3,32'd2,32'd0,32'd17,32'd17,32'd13,32'd8,32'd17,32'd16,32'd7,32'd5,32'd6,32'd0,32'd0,32'd8,32'd14,32'd2,32'd2,32'd1,32'd3,32'd3,32'd3,32'd6,32'd2,32'd2,32'd5,32'd6,32'd6,32'd17,32'd6,32'd4,32'd1,32'd6,32'd4,32'd5,32'd2,32'd8,32'd18,32'd3,32'd6,32'd8,32'd0,32'd5,32'd5,32'd5,32'd4,32'd5,32'd1,32'd1,32'd4,32'd2,32'd2,32'd2,32'd0,32'd1,32'd0,32'd0,32'd15,32'd3,32'd2,32'd5,32'd9,32'd11,32'd0,32'd16,32'd11,32'd6,32'd7,32'd1,32'd2,32'd2,32'd6,32'd11,32'd15,32'd15,32'd4,32'd15,32'd13,32'd8,32'd13,32'd15,32'd8,32'd8,32'd8,32'd10,32'd10,32'd21,32'd3,32'd5,32'd2,32'd0,32'd2,32'd2,32'd2,32'd13,32'd13,32'd13,32'd8,32'd8,32'd4,32'd4,32'd2,32'd4,32'd10,32'd6,32'd5,32'd1,32'd3,32'd3,32'd8,32'd4,32'd9,32'd9,32'd6,32'd6,32'd16,32'd12,32'd16,32'd16,32'd10,32'd0,32'd1,32'd0,32'd18,32'd9,32'd6,32'd6,32'd3,32'd3,32'd20,32'd17,32'd4,32'd0,32'd0,32'd0,32'd3,32'd10,32'd15,32'd3,32'd0,32'd1,32'd7,32'd2,32'd18,32'd1,32'd7,32'd0,32'd6,32'd7,32'd2,32'd5,32'd18,32'd10,32'd16,32'd16,32'd16,32'd17,32'd1,32'd20,32'd21,32'd1,32'd15,32'd15,32'd16,32'd11,32'd4,32'd4,32'd7,32'd7,32'd12,32'd12,32'd12,32'd15,32'd7,32'd15,32'd9,32'd0,32'd6,32'd11,32'd4,32'd4,32'd0,32'd18,32'd4,32'd4,32'd0,32'd4,32'd11,32'd5,32'd10,32'd17,32'd7,32'd0,32'd11,32'd0,32'd7,32'd8,32'd2,32'd4,32'd20,32'd12,32'd0,32'd12,32'd12,32'd11,32'd1,32'd4,32'd18,32'd6,32'd8,32'd11,32'd11,32'd3,32'd3,32'd3,32'd3,32'd2,32'd2,32'd3,32'd3,32'd8,32'd8,32'd7,32'd6,32'd6,32'd4,32'd8,32'd15,32'd7,32'd11,32'd9,32'd10,32'd15,32'd12,32'd16,32'd0,32'd5,32'd2,32'd16,32'd15,32'd10,32'd10,32'd9,32'd0,32'd2,32'd12,32'd7,32'd13,32'd7,32'd14,32'd12,32'd4,32'd6,32'd6,32'd12,32'd21,32'd18,32'd9,32'd10,32'd6,32'd11,32'd11,32'd1,32'd1,32'd1,32'd1,32'd2,32'd15,32'd7,32'd4,32'd5,32'd5,32'd8,32'd8,32'd1,32'd2,32'd0,32'd0,32'd2,32'd17,32'd16,32'd1,32'd0,32'd13,32'd12,32'd14,32'd12,32'd10,32'd7,32'd6,32'd7,32'd6,32'd11,32'd16,32'd16,32'd6,32'd6,32'd18,32'd9,32'd14,32'd9,32'd12,32'd5,32'd10,32'd8,32'd8,32'd7,32'd6,32'd5,32'd8,32'd0,32'd8,32'd7,32'd8,32'd14,32'd15,32'd15,32'd14,32'd17,32'd17,32'd0,32'd0,32'd0,32'd6,32'd2,32'd6,32'd7,32'd3,32'd0,32'd7,32'd10,32'd2,32'd0,32'd0,32'd2,32'd2,32'd0,32'd0,32'd5,32'd2,32'd10,32'd0,32'd7,32'd0,32'd0,32'd0,32'd4,32'd15,32'd10,32'd3,32'd6,32'd6,32'd5,32'd21,32'd6,32'd1,32'd4,32'd2,32'd14,32'd13,32'd3,32'd2,32'd2,32'd9,32'd2,32'd10,32'd7,32'd16,32'd1,32'd0,32'd7,32'd22,32'd4,32'd12,32'd6,32'd0,32'd0,32'd15,32'd15,32'd12,32'd12,32'd0,32'd12,32'd4,32'd4,32'd0,32'd6,32'd5,32'd5,32'd8,32'd8,32'd20,32'd18,32'd18,32'd5,32'd10,32'd4,32'd9,32'd15,32'd0,32'd14,32'd8,32'd7,32'd13,32'd2,32'd0,32'd0,32'd0,32'd0,32'd2,32'd4,32'd11,32'd11,32'd5,32'd7,32'd12,32'd1,32'd13,32'd4,32'd2,32'd2,32'd16,32'd6,32'd5,32'd17,32'd3,32'd7,32'd3,32'd18,32'd18,32'd3,32'd0,32'd0,32'd8,32'd11,32'd7,32'd3,32'd10,32'd2,32'd12,32'd0,32'd2,32'd2,32'd2,32'd2,32'd15,32'd2,32'd1,32'd0,32'd16,32'd16,32'd16,32'd16,32'd13,32'd13,32'd13,32'd3,32'd4,32'd1,32'd0,32'd13,32'd10,32'd13,32'd6,32'd8,32'd5,32'd14,32'd5,32'd6,32'd5,32'd5,32'd21,32'd12,32'd0,32'd16,32'd4,32'd0,32'd2,32'd2,32'd5,32'd5,32'd5,32'd5,32'd14,32'd14,32'd7,32'd0,32'd15,32'd22,32'd0,32'd8,32'd1,32'd4,32'd0,32'd10,32'd9,32'd1,32'd3,32'd2,32'd2,32'd9,32'd6,32'd1,32'd0,32'd4,32'd6,32'd0,32'd16,32'd16,32'd4,32'd5,32'd7,32'd1,32'd17,32'd17,32'd8,32'd15,32'd7,32'd8,32'd4,32'd7,32'd9,32'd9,32'd12,32'd17,32'd13,32'd5,32'd15,32'd10,32'd10,32'd8,32'd10,32'd9,32'd20,32'd13,32'd14,32'd0,32'd0,32'd17,32'd17,32'd17,32'd18,32'd17,32'd5,32'd5,32'd9,32'd7,32'd2,32'd0,32'd12,32'd12,32'd15,32'd5,32'd2,32'd15,32'd1,32'd1,32'd5,32'd13,32'd7,32'd7,32'd3,32'd3,32'd7,32'd1,32'd0,32'd5,32'd3,32'd0,32'd3,32'd1,32'd15,32'd15,32'd1,32'd1,32'd6,32'd6,32'd3,32'd14,32'd15,32'd11,32'd1,32'd14,32'd12,32'd6,32'd10,32'd10,32'd2,32'd2,32'd0,32'd1,32'd13,32'd12,32'd5,32'd0,32'd0,32'd12,32'd5,32'd3,32'd0,32'd6,32'd20,32'd11,32'd11,32'd11,32'd0,32'd0,32'd3,32'd3,32'd14,32'd17,32'd8,32'd11,32'd6,32'd3,32'd0,32'd0,32'd12,32'd1,32'd7,32'd12,32'd8,32'd8,32'd19,32'd8,32'd18,32'd6,32'd1,32'd3,32'd4,32'd9,32'd9,32'd0,32'd9,32'd5,32'd9,32'd4,32'd4,32'd12,32'd9,32'd11,32'd8,32'd11,32'd6,32'd10,32'd4,32'd0,32'd10,32'd12,32'd10,32'd7,32'd6,32'd5,32'd5,32'd0,32'd16,32'd8,32'd13,32'd16,32'd4,32'd7,32'd14,32'd6,32'd10,32'd9,32'd18,32'd11,32'd1,32'd0,32'd0,32'd11,32'd8,32'd14,32'd14,32'd9,32'd5,32'd7,32'd8,32'd0,32'd7,32'd2,32'd6,32'd5,32'd18,32'd17,32'd1,32'd6,32'd3,32'd3,32'd6,32'd6,32'd3,32'd12,32'd4,32'd7,32'd7,32'd4,32'd9,32'd3,32'd16,32'd3,32'd16,32'd1,32'd1,32'd0,32'd3,32'd0,32'd18,32'd4,32'd10,32'd7,32'd16,32'd6,32'd16,32'd11,32'd11,32'd6,32'd6,32'd0,32'd2,32'd10,32'd0,32'd12,32'd11,32'd14,32'd8,32'd8,32'd7,32'd4,32'd6,32'd0,32'd21,32'd12,32'd8,32'd0,32'd7,32'd6,32'd2,32'd1,32'd16,32'd12,32'd8,32'd13,32'd12,32'd14,32'd2,32'd13,32'd5,32'd15,32'd13,32'd16,32'd1,32'd2,32'd2,32'd3,32'd7,32'd17,32'd0,32'd0,32'd17,32'd2,32'd0,32'd6,32'd0,32'd7,32'd10,32'd9,32'd11,32'd10,32'd2,32'd1,32'd19,32'd1,32'd5,32'd16,32'd13,32'd6,32'd12,32'd17,32'd15,32'd20,32'd21,32'd12,32'd10,32'd11,32'd10,32'd10,32'd4,32'd0,32'd5,32'd0,32'd4,32'd3,32'd0,32'd10,32'd3,32'd0,32'd0,32'd2,32'd0,32'd11,32'd8,32'd8,32'd9,32'd5,32'd7,32'd6,32'd5,32'd8,32'd8,32'd6,32'd8,32'd17,32'd15,32'd15,32'd16,32'd0,32'd4,32'd3,32'd11,32'd11,32'd16,32'd16,32'd16,32'd10,32'd6,32'd17,32'd0,32'd4,32'd2,32'd11,32'd0,32'd10,32'd12,32'd14,32'd6,32'd10,32'd13,32'd17,32'd15,32'd2,32'd5,32'd13,32'd6,32'd5,32'd6,32'd6,32'd5,32'd5,32'd11,32'd0,32'd9,32'd10,32'd13,32'd9,32'd16,32'd16,32'd4,32'd5,32'd5,32'd5,32'd0,32'd9,32'd0,32'd6,32'd8,32'd8,32'd5,32'd2,32'd8,32'd8,32'd13,32'd15,32'd3,32'd0,32'd1,32'd10,32'd22,32'd5,32'd0,32'd0,32'd2,32'd3,32'd2,32'd18,32'd7,32'd6,32'd12,32'd7,32'd1,32'd3,32'd0,32'd10,32'd10,32'd5,32'd5,32'd6,32'd6,32'd5,32'd11,32'd9,32'd14,32'd3,32'd0,32'd5,32'd2,32'd3,32'd0,32'd2,32'd9,32'd18,32'd2,32'd7,32'd10,32'd6,32'd4,32'd5,32'd5,32'd19,32'd6,32'd9,32'd11,32'd14,32'd14,32'd5,32'd7,32'd8,32'd5,32'd2,32'd2,32'd18,32'd18,32'd4,32'd4,32'd4,32'd4,32'd2,32'd2,32'd10,32'd10,32'd4,32'd4,32'd5,32'd6,32'd6,32'd9,32'd8,32'd4,32'd10,32'd21,32'd3,32'd5,32'd6,32'd5,32'd11,32'd10,32'd0,32'd0,32'd6,32'd3,32'd18,32'd17,32'd2,32'd8,32'd7,32'd9,32'd13,32'd17,32'd16,32'd3,32'd11,32'd2,32'd0,32'd16,32'd2,32'd8,32'd4,32'd8,32'd6,32'd3,32'd2,32'd14,32'd7,32'd18,32'd0,32'd2,32'd0,32'd0,32'd15,32'd4,32'd11,32'd11,32'd12,32'd11,32'd20,32'd11,32'd0,32'd6,32'd1,32'd0,32'd6,32'd14,32'd13,32'd5,32'd8,32'd0,32'd0,32'd16,32'd16,32'd2,32'd12,32'd14,32'd14,32'd0,32'd6,32'd7,32'd9,32'd0,32'd3,32'd6,32'd6,32'd7,32'd6,32'd0,32'd0,32'd7,32'd7,32'd2,32'd2,32'd5,32'd17,32'd0,32'd0,32'd2,32'd2,32'd9,32'd15,32'd1,32'd1,32'd5,32'd5,32'd5,32'd5,32'd13,32'd14,32'd12,32'd16,32'd9,32'd5,32'd1,32'd1,32'd7,32'd14,32'd10,32'd10,32'd4,32'd10,32'd2,32'd1,32'd5,32'd13,32'd0,32'd0,32'd1,32'd3,32'd4,32'd1,32'd6,32'd7,32'd2,32'd0,32'd6,32'd0,32'd12,32'd8,32'd0,32'd0,32'd11,32'd3,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd17,32'd15,32'd17,32'd3,32'd9,32'd9,32'd18,32'd18,32'd6,32'd18,32'd17,32'd7,32'd7,32'd2,32'd5,32'd6,32'd21,32'd10,32'd0,32'd6,32'd0,32'd4,32'd3,32'd4,32'd2,32'd0,32'd14,32'd6,32'd7,32'd7,32'd7,32'd3,32'd0,32'd6,32'd5,32'd6,32'd2,32'd2,32'd2,32'd7,32'd0,32'd13,32'd5,32'd7,32'd7,32'd0,32'd0,32'd4,32'd5,32'd4,32'd0,32'd13,32'd16,32'd15,32'd15,32'd17,32'd1,32'd0,32'd0,32'd7,32'd5,32'd3,32'd10,32'd13,32'd0,32'd20,32'd2,32'd12,32'd8,32'd15,32'd0,32'd0,32'd4,32'd6,32'd6,32'd17,32'd17,32'd0,32'd0,32'd12,32'd9,32'd11,32'd11,32'd14,32'd14,32'd22,32'd4,32'd4,32'd4,32'd6,32'd4,32'd5,32'd3,32'd8,32'd15,32'd0,32'd0,32'd2,32'd12,32'd20,32'd2,32'd7,32'd7,32'd16,32'd4,32'd18,32'd1,32'd1,32'd6,32'd7,32'd7,32'd2,32'd5,32'd8,32'd1,32'd15,32'd8,32'd6,32'd7,32'd5,32'd3,32'd0,32'd13,32'd17,32'd3,32'd10,32'd14,32'd8,32'd12,32'd7,32'd15,32'd15,32'd0,32'd9,32'd1,32'd15,32'd10,32'd6,32'd0,32'd1,32'd3,32'd14,32'd1,32'd1,32'd0,32'd15,32'd13,32'd14,32'd12,32'd12,32'd12,32'd12,32'd0,32'd0,32'd4,32'd7,32'd0,32'd6,32'd13,32'd13,32'd21,32'd9,32'd1,32'd1,32'd12,32'd12,32'd6,32'd8,32'd5,32'd12,32'd6,32'd12,32'd0,32'd0,32'd0,32'd10,32'd2,32'd2,32'd18,32'd2,32'd6,32'd6,32'd9,32'd6,32'd6,32'd12,32'd3,32'd7,32'd6,32'd6,32'd14,32'd8,32'd6,32'd4,32'd2,32'd14,32'd21,32'd14,32'd2,32'd5,32'd3,32'd16,32'd1,32'd3,32'd4,32'd4,32'd0,32'd18,32'd17,32'd5,32'd13,32'd14,32'd10,32'd2,32'd3,32'd3,32'd0,32'd0,32'd7,32'd7,32'd12,32'd12,32'd12,32'd8,32'd9,32'd11,32'd0,32'd0,32'd0,32'd9,32'd6,32'd1,32'd0,32'd10,32'd14,32'd14,32'd8,32'd8,32'd0,32'd3,32'd3,32'd2,32'd1,32'd4,32'd3,32'd7,32'd6,32'd18,32'd2,32'd2,32'd0,32'd1,32'd12,32'd6,32'd13,32'd13,32'd1,32'd7,32'd17,32'd4,32'd2,32'd6,32'd14,32'd2,32'd1,32'd6,32'd0,32'd15,32'd15,32'd8,32'd7,32'd7,32'd21,32'd0,32'd0,32'd1,32'd2,32'd5,32'd20,32'd7,32'd0,32'd0,32'd6,32'd16,32'd10,32'd6,32'd6,32'd9,32'd14,32'd6,32'd4,32'd15,32'd20,32'd18,32'd18,32'd17,32'd7,32'd6,32'd0,32'd0,32'd4,32'd0,32'd5,32'd5,32'd15,32'd1,32'd4,32'd2,32'd1,32'd7,32'd12,32'd12,32'd8,32'd2,32'd1,32'd5,32'd1,32'd6,32'd0,32'd22,32'd0,32'd0,32'd15,32'd0,32'd4,32'd5,32'd5,32'd8,32'd2,32'd17,32'd4,32'd18,32'd14,32'd14,32'd6,32'd1,32'd1,32'd0,32'd0,32'd0,32'd4,32'd13,32'd10,32'd11,32'd11,32'd11,32'd10,32'd10,32'd3,32'd3,32'd18,32'd0,32'd0,32'd1,32'd0,32'd3,32'd0,32'd0,32'd12,32'd10,32'd14,32'd7,32'd6,32'd8,32'd8,32'd6,32'd7,32'd15,32'd9,32'd10,32'd7,32'd0,32'd0,32'd1,32'd1,32'd5,32'd1,32'd7,32'd17,32'd5,32'd8,32'd2,32'd1,32'd16,32'd16,32'd12,32'd9,32'd8,32'd2,32'd1,32'd6,32'd0,32'd16,32'd13,32'd14,32'd5,32'd5,32'd6,32'd0,32'd9,32'd10,32'd19,32'd8,32'd16,32'd14,32'd0,32'd0,32'd8,32'd8,32'd10,32'd0,32'd12,32'd16,32'd4,32'd4,32'd4,32'd16,32'd1,32'd18,32'd14,32'd6,32'd7,32'd7,32'd22,32'd12,32'd6,32'd6,32'd13,32'd6,32'd20,32'd6,32'd7,32'd0,32'd0,32'd8,32'd6,32'd6,32'd0,32'd6,32'd0,32'd0,32'd5,32'd6,32'd15,32'd15,32'd14,32'd8,32'd5,32'd0,32'd1,32'd4,32'd17,32'd15,32'd7,32'd6,32'd12,32'd7,32'd7,32'd1,32'd3,32'd3,32'd17,32'd10,32'd1,32'd5,32'd4,32'd4,32'd13,32'd10,32'd5,32'd1,32'd1,32'd6,32'd1,32'd3,32'd4,32'd5,32'd2,32'd1,32'd13,32'd1,32'd12,32'd6,32'd8,32'd1,32'd1,32'd6,32'd21,32'd6,32'd5,32'd6,32'd8,32'd3,32'd7,32'd18,32'd6,32'd6,32'd0,32'd5,32'd8,32'd5,32'd11,32'd0,32'd6,32'd9,32'd2,32'd8,32'd4,32'd6,32'd0,32'd14,32'd8,32'd5,32'd5,32'd18,32'd9,32'd4,32'd4}
`define RECTANGLE1_WIDTHS {32'd6,32'd24,32'd3,32'd9,32'd9,32'd9,32'd9,32'd18,32'd19,32'd18,32'd9,32'd22,32'd9,32'd6,32'd6,32'd12,32'd24,32'd22,32'd10,32'd8,32'd8,32'd17,32'd9,32'd3,32'd7,32'd16,32'd16,32'd4,32'd4,32'd10,32'd10,32'd8,32'd8,32'd4,32'd18,32'd6,32'd6,32'd6,32'd4,32'd6,32'd19,32'd13,32'd6,32'd6,32'd6,32'd5,32'd16,32'd12,32'd17,32'd18,32'd10,32'd2,32'd2,32'd6,32'd4,32'd18,32'd12,32'd5,32'd18,32'd8,32'd8,32'd22,32'd9,32'd18,32'd18,32'd10,32'd24,32'd13,32'd13,32'd16,32'd9,32'd14,32'd16,32'd13,32'd8,32'd9,32'd24,32'd18,32'd6,32'd6,32'd4,32'd6,32'd6,32'd18,32'd16,32'd9,32'd16,32'd6,32'd6,32'd3,32'd3,32'd9,32'd9,32'd10,32'd18,32'd6,32'd6,32'd8,32'd6,32'd16,32'd24,32'd18,32'd18,32'd21,32'd22,32'd18,32'd18,32'd3,32'd3,32'd18,32'd3,32'd18,32'd18,32'd12,32'd8,32'd12,32'd3,32'd8,32'd8,32'd2,32'd2,32'd12,32'd16,32'd16,32'd19,32'd7,32'd18,32'd18,32'd18,32'd10,32'd10,32'd9,32'd9,32'd10,32'd10,32'd10,32'd10,32'd9,32'd12,32'd9,32'd18,32'd4,32'd4,32'd12,32'd3,32'd10,32'd18,32'd10,32'd24,32'd6,32'd6,32'd22,32'd13,32'd6,32'd12,32'd12,32'd15,32'd9,32'd18,32'd18,32'd3,32'd10,32'd10,32'd7,32'd7,32'd13,32'd20,32'd8,32'd8,32'd6,32'd6,32'd3,32'd18,32'd15,32'd18,32'd6,32'd6,32'd6,32'd20,32'd6,32'd18,32'd20,32'd24,32'd3,32'd14,32'd5,32'd5,32'd6,32'd6,32'd12,32'd19,32'd18,32'd7,32'd6,32'd12,32'd12,32'd6,32'd8,32'd12,32'd12,32'd3,32'd10,32'd9,32'd9,32'd10,32'd16,32'd18,32'd3,32'd6,32'd4,32'd12,32'd12,32'd6,32'd6,32'd6,32'd6,32'd9,32'd9,32'd6,32'd14,32'd18,32'd9,32'd19,32'd19,32'd9,32'd20,32'd18,32'd5,32'd3,32'd3,32'd18,32'd3,32'd4,32'd18,32'd3,32'd3,32'd4,32'd8,32'd12,32'd11,32'd7,32'd10,32'd16,32'd9,32'd6,32'd9,32'd6,32'd12,32'd9,32'd12,32'd12,32'd11,32'd6,32'd6,32'd3,32'd3,32'd18,32'd18,32'd15,32'd24,32'd8,32'd8,32'd17,32'd17,32'd6,32'd13,32'd14,32'd14,32'd9,32'd12,32'd8,32'd10,32'd15,32'd6,32'd19,32'd14,32'd4,32'd7,32'd6,32'd3,32'd5,32'd12,32'd9,32'd9,32'd5,32'd4,32'd8,32'd9,32'd14,32'd14,32'd10,32'd18,32'd3,32'd3,32'd3,32'd12,32'd20,32'd10,32'd2,32'd6,32'd12,32'd18,32'd6,32'd6,32'd18,32'd9,32'd18,32'd8,32'd8,32'd8,32'd6,32'd18,32'd18,32'd18,32'd10,32'd10,32'd18,32'd10,32'd18,32'd15,32'd10,32'd10,32'd16,32'd8,32'd9,32'd20,32'd18,32'd12,32'd8,32'd8,32'd8,32'd8,32'd6,32'd9,32'd12,32'd21,32'd6,32'd6,32'd6,32'd3,32'd14,32'd6,32'd18,32'd24,32'd18,32'd17,32'd5,32'd18,32'd9,32'd5,32'd4,32'd4,32'd6,32'd3,32'd16,32'd6,32'd18,32'd12,32'd6,32'd14,32'd9,32'd9,32'd6,32'd18,32'd9,32'd18,32'd9,32'd9,32'd8,32'd8,32'd12,32'd6,32'd4,32'd12,32'd6,32'd4,32'd6,32'd6,32'd18,32'd18,32'd4,32'd12,32'd4,32'd18,32'd8,32'd4,32'd6,32'd9,32'd9,32'd18,32'd18,32'd9,32'd10,32'd10,32'd6,32'd19,32'd6,32'd6,32'd24,32'd10,32'd10,32'd18,32'd12,32'd17,32'd6,32'd6,32'd6,32'd22,32'd8,32'd12,32'd7,32'd8,32'd14,32'd6,32'd6,32'd9,32'd18,32'd19,32'd16,32'd10,32'd6,32'd6,32'd10,32'd9,32'd9,32'd9,32'd9,32'd8,32'd9,32'd8,32'd8,32'd8,32'd6,32'd12,32'd21,32'd20,32'd8,32'd11,32'd9,32'd11,32'd9,32'd3,32'd9,32'd10,32'd9,32'd18,32'd6,32'd9,32'd18,32'd18,32'd10,32'd6,32'd18,32'd9,32'd9,32'd18,32'd18,32'd3,32'd10,32'd4,32'd4,32'd9,32'd6,32'd18,32'd22,32'd3,32'd9,32'd6,32'd8,32'd7,32'd16,32'd4,32'd6,32'd3,32'd14,32'd6,32'd6,32'd5,32'd5,32'd12,32'd3,32'd6,32'd8,32'd4,32'd4,32'd9,32'd24,32'd20,32'd6,32'd12,32'd15,32'd18,32'd8,32'd2,32'd18,32'd9,32'd4,32'd6,32'd6,32'd19,32'd20,32'd7,32'd4,32'd9,32'd9,32'd6,32'd18,32'd16,32'd24,32'd9,32'd22,32'd4,32'd4,32'd9,32'd20,32'd10,32'd6,32'd4,32'd13,32'd9,32'd4,32'd11,32'd9,32'd5,32'd12,32'd6,32'd10,32'd3,32'd3,32'd16,32'd16,32'd6,32'd15,32'd21,32'd16,32'd14,32'd4,32'd6,32'd14,32'd24,32'd12,32'd14,32'd10,32'd4,32'd4,32'd5,32'd5,32'd10,32'd9,32'd9,32'd18,32'd6,32'd6,32'd2,32'd2,32'd18,32'd10,32'd6,32'd4,32'd7,32'd6,32'd10,32'd4,32'd16,32'd2,32'd4,32'd4,32'd18,32'd18,32'd9,32'd9,32'd18,32'd9,32'd6,32'd6,32'd4,32'd6,32'd6,32'd6,32'd7,32'd6,32'd15,32'd6,32'd12,32'd7,32'd6,32'd10,32'd8,32'd24,32'd19,32'd18,32'd10,32'd8,32'd4,32'd8,32'd24,32'd9,32'd18,32'd10,32'd18,32'd6,32'd4,32'd19,32'd6,32'd6,32'd9,32'd4,32'd12,32'd24,32'd5,32'd9,32'd3,32'd10,32'd10,32'd14,32'd9,32'd10,32'd10,32'd6,32'd6,32'd6,32'd6,32'd6,32'd6,32'd6,32'd10,32'd4,32'd18,32'd24,32'd24,32'd18,32'd4,32'd9,32'd22,32'd22,32'd9,32'd6,32'd12,32'd3,32'd12,32'd10,32'd2,32'd7,32'd7,32'd20,32'd10,32'd9,32'd24,32'd6,32'd19,32'd5,32'd24,32'd3,32'd9,32'd19,32'd16,32'd9,32'd9,32'd12,32'd16,32'd8,32'd16,32'd16,32'd18,32'd6,32'd6,32'd4,32'd8,32'd10,32'd8,32'd14,32'd24,32'd8,32'd8,32'd6,32'd4,32'd15,32'd15,32'd6,32'd18,32'd6,32'd6,32'd4,32'd6,32'd6,32'd6,32'd6,32'd6,32'd9,32'd9,32'd9,32'd18,32'd18,32'd12,32'd18,32'd9,32'd11,32'd6,32'd11,32'd14,32'd4,32'd12,32'd9,32'd12,32'd9,32'd12,32'd8,32'd8,32'd4,32'd9,32'd4,32'd11,32'd10,32'd4,32'd18,32'd4,32'd18,32'd18,32'd21,32'd21,32'd12,32'd14,32'd20,32'd18,32'd18,32'd18,32'd8,32'd6,32'd24,32'd18,32'd10,32'd8,32'd6,32'd24,32'd8,32'd15,32'd18,32'd10,32'd6,32'd15,32'd4,32'd12,32'd14,32'd3,32'd6,32'd12,32'd8,32'd8,32'd6,32'd12,32'd5,32'd20,32'd3,32'd18,32'd6,32'd22,32'd14,32'd15,32'd19,32'd4,32'd18,32'd12,32'd6,32'd18,32'd18,32'd18,32'd12,32'd6,32'd9,32'd6,32'd12,32'd4,32'd20,32'd15,32'd6,32'd6,32'd6,32'd6,32'd6,32'd10,32'd6,32'd4,32'd6,32'd6,32'd6,32'd18,32'd18,32'd6,32'd6,32'd24,32'd16,32'd19,32'd19,32'd10,32'd10,32'd24,32'd6,32'd6,32'd6,32'd8,32'd6,32'd19,32'd4,32'd6,32'd6,32'd12,32'd12,32'd8,32'd10,32'd4,32'd6,32'd6,32'd22,32'd4,32'd10,32'd15,32'd14,32'd18,32'd8,32'd6,32'd18,32'd4,32'd4,32'd4,32'd6,32'd6,32'd18,32'd9,32'd18,32'd8,32'd8,32'd14,32'd7,32'd9,32'd19,32'd6,32'd4,32'd3,32'd4,32'd10,32'd4,32'd12,32'd4,32'd4,32'd4,32'd10,32'd18,32'd18,32'd18,32'd9,32'd18,32'd6,32'd20,32'd6,32'd6,32'd9,32'd18,32'd19,32'd23,32'd10,32'd24,32'd6,32'd6,32'd6,32'd6,32'd8,32'd8,32'd4,32'd10,32'd6,32'd20,32'd4,32'd4,32'd18,32'd7,32'd8,32'd4,32'd6,32'd6,32'd4,32'd6,32'd18,32'd6,32'd19,32'd23,32'd9,32'd12,32'd22,32'd12,32'd24,32'd9,32'd10,32'd14,32'd10,32'd6,32'd8,32'd12,32'd24,32'd20,32'd9,32'd3,32'd4,32'd12,32'd8,32'd7,32'd14,32'd9,32'd24,32'd16,32'd16,32'd9,32'd4,32'd4,32'd6,32'd4,32'd10,32'd8,32'd21,32'd10,32'd19,32'd20,32'd6,32'd24,32'd4,32'd18,32'd10,32'd10,32'd12,32'd8,32'd6,32'd6,32'd10,32'd10,32'd12,32'd18,32'd6,32'd6,32'd6,32'd12,32'd18,32'd4,32'd10,32'd18,32'd16,32'd21,32'd12,32'd19,32'd8,32'd5,32'd6,32'd9,32'd10,32'd10,32'd18,32'd6,32'd6,32'd16,32'd6,32'd6,32'd6,32'd6,32'd4,32'd4,32'd18,32'd6,32'd20,32'd12,32'd3,32'd15,32'd9,32'd9,32'd4,32'd6,32'd6,32'd6,32'd6,32'd6,32'd18,32'd22,32'd21,32'd9,32'd18,32'd6,32'd5,32'd10,32'd12,32'd13,32'd21,32'd6,32'd20,32'd4,32'd8,32'd8,32'd9,32'd9,32'd20,32'd24,32'd20,32'd20,32'd18,32'd6,32'd18,32'd9,32'd14,32'd14,32'd9,32'd19,32'd20,32'd12,32'd5,32'd3,32'd14,32'd14,32'd18,32'd10,32'd6,32'd6,32'd9,32'd12,32'd16,32'd10,32'd3,32'd3,32'd15,32'd9,32'd15,32'd18,32'd16,32'd12,32'd6,32'd21,32'd6,32'd6,32'd12,32'd18,32'd5,32'd5,32'd17,32'd12,32'd4,32'd4,32'd3,32'd24,32'd18,32'd12,32'd15,32'd12,32'd6,32'd6,32'd13,32'd8,32'd20,32'd14,32'd12,32'd12,32'd12,32'd4,32'd6,32'd6,32'd9,32'd9,32'd6,32'd6,32'd12,32'd12,32'd6,32'd6,32'd16,32'd3,32'd4,32'd8,32'd6,32'd6,32'd9,32'd14,32'd10,32'd10,32'd18,32'd10,32'd6,32'd6,32'd6,32'd24,32'd15,32'd15,32'd18,32'd10,32'd9,32'd18,32'd10,32'd16,32'd12,32'd12,32'd6,32'd10,32'd9,32'd22,32'd24,32'd9,32'd24,32'd18,32'd18,32'd16,32'd12,32'd12,32'd6,32'd6,32'd8,32'd15,32'd14,32'd9,32'd6,32'd4,32'd6,32'd6,32'd18,32'd6,32'd4,32'd10,32'd14,32'd5,32'd8,32'd9,32'd12,32'd5,32'd10,32'd6,32'd10,32'd4,32'd3,32'd18,32'd8,32'd3,32'd18,32'd18,32'd9,32'd9,32'd24,32'd19,32'd9,32'd18,32'd24,32'd18,32'd18,32'd14,32'd12,32'd12,32'd4,32'd14,32'd16,32'd5,32'd6,32'd21,32'd6,32'd16,32'd14,32'd6,32'd4,32'd6,32'd4,32'd12,32'd14,32'd3,32'd9,32'd6,32'd6,32'd6,32'd6,32'd6,32'd6,32'd6,32'd9,32'd6,32'd6,32'd6,32'd15,32'd20,32'd6,32'd18,32'd5,32'd16,32'd6,32'd12,32'd17,32'd6,32'd18,32'd10,32'd19,32'd9,32'd6,32'd4,32'd4,32'd12,32'd21,32'd8,32'd24,32'd21,32'd14,32'd8,32'd24,32'd11,32'd11,32'd18,32'd9,32'd6,32'd8,32'd23,32'd9,32'd5,32'd5,32'd10,32'd6,32'd6,32'd18,32'd6,32'd6,32'd6,32'd18,32'd12,32'd12,32'd6,32'd18,32'd6,32'd6,32'd6,32'd22,32'd18,32'd22,32'd12,32'd12,32'd3,32'd6,32'd22,32'd21,32'd10,32'd18,32'd8,32'd8,32'd10,32'd12,32'd9,32'd22,32'd12,32'd12,32'd10,32'd18,32'd16,32'd4,32'd5,32'd18,32'd4,32'd19,32'd8,32'd3,32'd6,32'd8,32'd7,32'd6,32'd6,32'd6,32'd8,32'd22,32'd16,32'd16,32'd10,32'd6,32'd10,32'd10,32'd10,32'd11,32'd6,32'd6,32'd18,32'd6,32'd6,32'd6,32'd10,32'd10,32'd4,32'd18,32'd15,32'd18,32'd2,32'd2,32'd9,32'd18,32'd6,32'd4,32'd6,32'd23,32'd7,32'd17,32'd20,32'd6,32'd9,32'd9,32'd5,32'd4,32'd16,32'd9,32'd12,32'd24,32'd8,32'd6,32'd24,32'd8,32'd6,32'd12,32'd9,32'd9,32'd6,32'd6,32'd15,32'd9,32'd20,32'd7,32'd12,32'd9,32'd18,32'd14,32'd18,32'd4,32'd6,32'd6,32'd18,32'd9,32'd19,32'd9,32'd2,32'd8,32'd4,32'd4,32'd6,32'd9,32'd20,32'd8,32'd14,32'd6,32'd16,32'd18,32'd4,32'd24,32'd8,32'd4,32'd5,32'd10,32'd20,32'd12,32'd6,32'd6,32'd9,32'd21,32'd10,32'd12,32'd6,32'd12,32'd8,32'd4,32'd4,32'd18,32'd10,32'd9,32'd9,32'd19,32'd6,32'd7,32'd7,32'd6,32'd10,32'd4,32'd16,32'd20,32'd24,32'd9,32'd9,32'd18,32'd9,32'd24,32'd9,32'd12,32'd17,32'd14,32'd12,32'd6,32'd6,32'd4,32'd18,32'd9,32'd7,32'd9,32'd6,32'd12,32'd12,32'd12,32'd22,32'd18,32'd18,32'd8,32'd6,32'd12,32'd12,32'd24,32'd8,32'd8,32'd24,32'd7,32'd5,32'd8,32'd8,32'd8,32'd8,32'd9,32'd8,32'd16,32'd18,32'd16,32'd8,32'd4,32'd4,32'd6,32'd11,32'd6,32'd6,32'd4,32'd12,32'd10,32'd12,32'd10,32'd10,32'd8,32'd12,32'd12,32'd9,32'd21,32'd5,32'd12,32'd12,32'd10,32'd10,32'd22,32'd18,32'd4,32'd6,32'd6,32'd6,32'd4,32'd6,32'd12,32'd10,32'd3,32'd4,32'd12,32'd4,32'd12,32'd20,32'd6,32'd6,32'd6,32'd6,32'd4,32'd24,32'd12,32'd21,32'd9,32'd22,32'd18,32'd18,32'd6,32'd24,32'd24,32'd6,32'd6,32'd6,32'd9,32'd16,32'd6,32'd6,32'd22,32'd18,32'd9,32'd9,32'd12,32'd6,32'd6,32'd6,32'd16,32'd6,32'd4,32'd10,32'd2,32'd2,32'd2,32'd19,32'd4,32'd4,32'd6,32'd4,32'd6,32'd12,32'd10,32'd6,32'd12,32'd20,32'd5,32'd6,32'd8,32'd10,32'd24,32'd2,32'd22,32'd10,32'd12,32'd4,32'd4,32'd6,32'd9,32'd6,32'd18,32'd6,32'd10,32'd6,32'd6,32'd10,32'd10,32'd9,32'd18,32'd6,32'd6,32'd6,32'd6,32'd5,32'd5,32'd6,32'd24,32'd6,32'd8,32'd9,32'd6,32'd12,32'd9,32'd8,32'd8,32'd12,32'd6,32'd15,32'd3,32'd12,32'd20,32'd12,32'd9,32'd6,32'd6,32'd12,32'd9,32'd4,32'd6,32'd12,32'd12,32'd6,32'd18,32'd9,32'd6,32'd18,32'd18,32'd6,32'd20,32'd18,32'd12,32'd7,32'd18,32'd6,32'd6,32'd2,32'd2,32'd2,32'd2,32'd24,32'd12,32'd6,32'd6,32'd5,32'd5,32'd6,32'd6,32'd6,32'd8,32'd8,32'd8,32'd13,32'd18,32'd9,32'd6,32'd6,32'd6,32'd6,32'd6,32'd9,32'd10,32'd11,32'd7,32'd22,32'd6,32'd19,32'd18,32'd10,32'd20,32'd20,32'd12,32'd22,32'd8,32'd18,32'd12,32'd6,32'd6,32'd8,32'd8,32'd12,32'd4,32'd6,32'd8,32'd6,32'd8,32'd15,32'd8,32'd9,32'd18,32'd23,32'd9,32'd18,32'd9,32'd6,32'd6,32'd6,32'd6,32'd6,32'd24,32'd6,32'd6,32'd22,32'd6,32'd18,32'd20,32'd20,32'd6,32'd6,32'd6,32'd18,32'd18,32'd6,32'd4,32'd20,32'd18,32'd9,32'd6,32'd6,32'd6,32'd4,32'd10,32'd18,32'd20,32'd9,32'd4,32'd3,32'd18,32'd5,32'd24,32'd15,32'd4,32'd4,32'd8,32'd24,32'd8,32'd8,32'd12,32'd12,32'd12,32'd15,32'd9,32'd12,32'd12,32'd11,32'd18,32'd10,32'd4,32'd10,32'd4,32'd8,32'd9,32'd9,32'd9,32'd9,32'd15,32'd9,32'd6,32'd6,32'd6,32'd6,32'd12,32'd12,32'd6,32'd20,32'd20,32'd14,32'd16,32'd6,32'd6,32'd12,32'd15,32'd9,32'd4,32'd19,32'd12,32'd10,32'd18,32'd24,32'd6,32'd6,32'd6,32'd6,32'd6,32'd18,32'd6,32'd6,32'd9,32'd12,32'd14,32'd21,32'd9,32'd20,32'd6,32'd6,32'd14,32'd14,32'd12,32'd9,32'd24,32'd22,32'd7,32'd21,32'd9,32'd7,32'd2,32'd2,32'd6,32'd6,32'd18,32'd8,32'd18,32'd6,32'd18,32'd21,32'd22,32'd6,32'd6,32'd6,32'd15,32'd6,32'd19,32'd18,32'd18,32'd18,32'd9,32'd9,32'd9,32'd9,32'd6,32'd8,32'd16,32'd5,32'd6,32'd9,32'd20,32'd6,32'd12,32'd12,32'd14,32'd10,32'd6,32'd6,32'd4,32'd6,32'd14,32'd7,32'd6,32'd9,32'd4,32'd4,32'd6,32'd24,32'd6,32'd6,32'd4,32'd4,32'd6,32'd6,32'd8,32'd4,32'd20,32'd19,32'd4,32'd9,32'd6,32'd14,32'd6,32'd21,32'd4,32'd10,32'd19,32'd16,32'd14,32'd20,32'd6,32'd22,32'd11,32'd24,32'd9,32'd24,32'd10,32'd10,32'd9,32'd12,32'd4,32'd9,32'd9,32'd9,32'd6,32'd6,32'd4,32'd10,32'd6,32'd9,32'd14,32'd14,32'd6,32'd9,32'd6,32'd9,32'd24,32'd10,32'd9,32'd9,32'd21,32'd6,32'd13,32'd6,32'd9,32'd14,32'd24,32'd9,32'd18,32'd9,32'd19,32'd9,32'd6,32'd22,32'd8,32'd5,32'd4,32'd14,32'd8,32'd8,32'd6,32'd18,32'd24,32'd6,32'd20,32'd20,32'd6,32'd18,32'd18,32'd19,32'd6,32'd3,32'd10,32'd3,32'd3,32'd4,32'd12,32'd3,32'd6,32'd3,32'd6,32'd6,32'd4,32'd4,32'd4,32'd12,32'd16,32'd7,32'd18,32'd9,32'd22,32'd8,32'd9,32'd14,32'd6,32'd6,32'd19,32'd21,32'd6,32'd8,32'd21,32'd11,32'd12,32'd6,32'd6,32'd8,32'd15,32'd4,32'd9,32'd16,32'd18,32'd19,32'd6,32'd6,32'd9,32'd9,32'd4,32'd4,32'd9,32'd18,32'd12,32'd12,32'd6,32'd4,32'd24,32'd13,32'd24,32'd19,32'd5,32'd8,32'd8,32'd8,32'd24,32'd8,32'd12,32'd6,32'd21,32'd23,32'd10,32'd5,32'd5,32'd3,32'd6,32'd16,32'd9,32'd8,32'd8,32'd6,32'd12,32'd12,32'd4,32'd20,32'd14,32'd10,32'd8,32'd4,32'd8,32'd6,32'd8,32'd6,32'd16,32'd10,32'd10,32'd6,32'd22,32'd14,32'd9,32'd12,32'd18,32'd8,32'd9,32'd7,32'd19,32'd15,32'd9,32'd6,32'd18,32'd4,32'd4,32'd20,32'd16,32'd6,32'd6,32'd6,32'd6,32'd15,32'd6,32'd4,32'd4,32'd12,32'd11,32'd6,32'd18,32'd10,32'd24,32'd9,32'd18,32'd9,32'd14,32'd16,32'd8,32'd9,32'd6,32'd10,32'd10,32'd14,32'd22,32'd13,32'd20,32'd11,32'd18,32'd4,32'd4,32'd9,32'd11,32'd4,32'd18,32'd14,32'd19,32'd6,32'd12,32'd21,32'd12,32'd18,32'd18,32'd9,32'd9,32'd6,32'd10,32'd12,32'd6,32'd23,32'd12,32'd6,32'd4,32'd6,32'd6,32'd4,32'd7,32'd16,32'd21,32'd6,32'd6,32'd8,32'd6,32'd12,32'd8,32'd4,32'd16,32'd16,32'd6,32'd8,32'd16,32'd6,32'd20,32'd6,32'd22,32'd19,32'd9,32'd9,32'd24,32'd4,32'd4,32'd6,32'd12,32'd18,32'd9,32'd18,32'd8,32'd18,32'd6,32'd10,32'd21,32'd5,32'd6,32'd9,32'd12,32'd9,32'd8,32'd4,32'd9,32'd9,32'd20,32'd12,32'd6,32'd9,32'd4,32'd10,32'd9,32'd18,32'd24,32'd9,32'd8,32'd12,32'd10,32'd10,32'd8,32'd6,32'd18,32'd16,32'd6,32'd16,32'd3,32'd18,32'd6,32'd6,32'd6,32'd6,32'd22,32'd18,32'd12,32'd10,32'd11,32'd3,32'd21,32'd8,32'd6,32'd6,32'd5,32'd6,32'd6,32'd18,32'd9,32'd9,32'd18,32'd24,32'd18,32'd24,32'd6,32'd6,32'd9,32'd9,32'd18,32'd8,32'd23,32'd12,32'd10,32'd21,32'd8,32'd9,32'd9,32'd20,32'd9,32'd9,32'd9,32'd10,32'd8,32'd11,32'd19,32'd23,32'd12,32'd6,32'd6,32'd12,32'd8,32'd8,32'd5,32'd5,32'd18,32'd24,32'd14,32'd3,32'd8,32'd6,32'd20,32'd18,32'd4,32'd6,32'd4,32'd4,32'd4,32'd18,32'd4,32'd18,32'd12,32'd9,32'd19,32'd4,32'd6,32'd6,32'd8,32'd9,32'd6,32'd4,32'd4,32'd12,32'd18,32'd9,32'd6,32'd6,32'd8,32'd6,32'd22,32'd9,32'd7,32'd4,32'd22,32'd7,32'd8,32'd12,32'd18,32'd9,32'd14,32'd3,32'd3,32'd14,32'd14,32'd18,32'd17,32'd4,32'd4,32'd24,32'd12,32'd10,32'd6,32'd6,32'd4,32'd4,32'd22,32'd20,32'd4,32'd18,32'd6,32'd19,32'd9,32'd14,32'd12,32'd9,32'd16,32'd12,32'd20,32'd8,32'd8,32'd12,32'd20,32'd6,32'd12,32'd12,32'd12,32'd21,32'd10,32'd8,32'd8,32'd6,32'd6,32'd6,32'd6,32'd6,32'd6,32'd15,32'd15,32'd3,32'd14,32'd5,32'd9,32'd9,32'd8,32'd18,32'd18,32'd6,32'd3,32'd9,32'd3,32'd6,32'd9,32'd6,32'd6,32'd4,32'd6,32'd10,32'd10,32'd3,32'd12,32'd18,32'd23,32'd9,32'd18,32'd18,32'd18,32'd24,32'd16,32'd10,32'd19,32'd14,32'd9,32'd4,32'd8,32'd12,32'd10,32'd4,32'd10,32'd6,32'd10,32'd20,32'd4,32'd6,32'd6,32'd10,32'd11,32'd6,32'd6,32'd10,32'd6,32'd24,32'd6,32'd6,32'd14,32'd18,32'd6,32'd6,32'd4,32'd14,32'd12,32'd15,32'd24,32'd10,32'd10,32'd10,32'd3,32'd24,32'd8,32'd18,32'd6,32'd4,32'd10,32'd8,32'd9,32'd8,32'd6,32'd6,32'd6,32'd6,32'd9,32'd9,32'd14,32'd14,32'd3,32'd14,32'd3,32'd9,32'd6,32'd6,32'd9,32'd9,32'd12,32'd18,32'd4,32'd4,32'd6,32'd6,32'd18,32'd3,32'd8,32'd9,32'd6,32'd18,32'd6,32'd16,32'd4,32'd4,32'd24,32'd11,32'd8,32'd8,32'd16,32'd8,32'd6,32'd6,32'd4,32'd24,32'd18,32'd18,32'd12,32'd2,32'd12,32'd6,32'd6,32'd6,32'd24,32'd9,32'd4,32'd3,32'd8,32'd9,32'd6,32'd3,32'd12,32'd6,32'd10,32'd10,32'd10,32'd16,32'd6,32'd6,32'd6,32'd21,32'd18,32'd6,32'd9,32'd9,32'd9,32'd9,32'd6,32'd9,32'd10,32'd15,32'd8,32'd4,32'd6,32'd21,32'd18,32'd23,32'd24,32'd12,32'd11,32'd5,32'd4,32'd5,32'd21,32'd6,32'd6,32'd4,32'd7,32'd8,32'd14,32'd9,32'd6,32'd6,32'd15,32'd2,32'd10,32'd6,32'd9,32'd6,32'd6,32'd10,32'd24,32'd4,32'd6,32'd6,32'd6,32'd2,32'd9,32'd6,32'd6,32'd21,32'd18,32'd16,32'd16,32'd18,32'd24,32'd10,32'd10,32'd24,32'd6,32'd11,32'd22,32'd18,32'd24,32'd14,32'd22,32'd7,32'd12,32'd18,32'd24,32'd22,32'd15,32'd14,32'd11,32'd18,32'd18,32'd6,32'd6,32'd6,32'd18,32'd4,32'd4,32'd6,32'd6,32'd19,32'd9,32'd6,32'd6,32'd9,32'd6,32'd11,32'd6,32'd18,32'd9,32'd4,32'd4,32'd9,32'd9,32'd21,32'd9,32'd10,32'd10,32'd10,32'd4,32'd12,32'd19,32'd6,32'd6,32'd5,32'd5,32'd24,32'd6,32'd12,32'd18,32'd6,32'd6,32'd6,32'd18,32'd3,32'd16,32'd18,32'd18,32'd10,32'd24,32'd3,32'd24,32'd18,32'd6,32'd15,32'd9,32'd13,32'd11,32'd17,32'd21,32'd9,32'd18,32'd6,32'd14,32'd4,32'd9,32'd6,32'd6,32'd6,32'd10,32'd10,32'd19,32'd19,32'd9,32'd9,32'd6,32'd6,32'd6,32'd6,32'd6,32'd8,32'd18,32'd16,32'd22,32'd10,32'd18,32'd6,32'd4,32'd4,32'd10,32'd9,32'd3,32'd9,32'd6,32'd9,32'd13,32'd9,32'd6,32'd6,32'd12,32'd18,32'd6,32'd6,32'd15,32'd6,32'd6,32'd6,32'd6,32'd6,32'd6,32'd19,32'd20,32'd18,32'd3,32'd5,32'd8,32'd14,32'd12,32'd12,32'd24,32'd6,32'd18,32'd5,32'd22,32'd6,32'd20,32'd9,32'd6,32'd18,32'd3,32'd3,32'd6,32'd19,32'd18,32'd3,32'd5,32'd6,32'd6,32'd9,32'd6,32'd6,32'd6,32'd6,32'd6,32'd10,32'd6,32'd6,32'd16,32'd6,32'd13,32'd24,32'd6,32'd6,32'd3,32'd10,32'd4,32'd8,32'd24,32'd18,32'd9,32'd9,32'd9,32'd9,32'd2,32'd2,32'd6,32'd2,32'd6,32'd10,32'd8,32'd12,32'd6,32'd12,32'd6,32'd6,32'd9,32'd4,32'd13,32'd3,32'd6,32'd6,32'd6,32'd5,32'd24,32'd5,32'd6,32'd10,32'd12,32'd6,32'd6,32'd7,32'd16,32'd10,32'd20,32'd6,32'd10,32'd10,32'd18,32'd24,32'd15,32'd22,32'd24,32'd5,32'd21,32'd15,32'd2,32'd2,32'd14,32'd18,32'd18,32'd18,32'd6,32'd10,32'd15,32'd10,32'd16,32'd15,32'd15,32'd18,32'd14,32'd9,32'd6,32'd6,32'd4,32'd4,32'd24,32'd6,32'd16,32'd6,32'd18,32'd6,32'd12,32'd4,32'd9,32'd6,32'd22,32'd22,32'd7,32'd22,32'd20,32'd14,32'd6,32'd19,32'd4,32'd19,32'd18,32'd4,32'd5,32'd18,32'd9,32'd6,32'd6,32'd14,32'd12,32'd18,32'd8,32'd18,32'd9,32'd9,32'd3,32'd2,32'd2,32'd2,32'd2,32'd20,32'd22,32'd24,32'd11,32'd6,32'd6,32'd8,32'd22,32'd18,32'd12,32'd6,32'd10,32'd9,32'd9,32'd20,32'd9,32'd16,32'd9,32'd10,32'd6,32'd18,32'd24,32'd3,32'd10,32'd9,32'd9,32'd8,32'd3,32'd17,32'd6,32'd19,32'd8,32'd6,32'd6,32'd6,32'd6,32'd6,32'd17,32'd22,32'd6,32'd9,32'd12,32'd24,32'd5,32'd12,32'd12,32'd15,32'd11,32'd22,32'd19,32'd4,32'd12,32'd6,32'd18,32'd8,32'd18,32'd12,32'd10,32'd14,32'd18,32'd18,32'd20,32'd12,32'd6,32'd9,32'd9,32'd6,32'd6,32'd12,32'd12,32'd6,32'd6,32'd8,32'd20,32'd4,32'd4,32'd6,32'd18,32'd22,32'd18,32'd10,32'd10,32'd8,32'd4,32'd18,32'd6,32'd4,32'd4,32'd15,32'd4,32'd24,32'd6,32'd16,32'd24,32'd12,32'd18,32'd6,32'd6,32'd6,32'd6,32'd6,32'd12,32'd14,32'd8,32'd9,32'd9,32'd7,32'd14,32'd20,32'd18,32'd4,32'd16,32'd18,32'd9,32'd6,32'd12,32'd16,32'd3,32'd8,32'd24,32'd4,32'd4,32'd12,32'd18,32'd24,32'd12,32'd12,32'd6,32'd4,32'd18,32'd14,32'd4,32'd4,32'd19,32'd4,32'd6,32'd6,32'd22,32'd4,32'd6,32'd20,32'd4,32'd21,32'd14,32'd24,32'd6,32'd6,32'd13,32'd18,32'd3,32'd6,32'd5,32'd15,32'd24,32'd14,32'd10,32'd6,32'd24,32'd6,32'd4,32'd6,32'd6,32'd9,32'd14,32'd14,32'd6,32'd24,32'd19,32'd12,32'd12,32'd7,32'd4,32'd12,32'd12,32'd4,32'd9,32'd18,32'd12,32'd12}
`define RECTANGLE1_HEIGHTS {32'd22,32'd8,32'd20,32'd6,32'd6,32'd6,32'd6,32'd3,32'd3,32'd2,32'd6,32'd10,32'd6,32'd12,32'd12,32'd3,32'd4,32'd6,32'd8,32'd15,32'd15,32'd9,32'd4,32'd21,32'd9,32'd12,32'd12,32'd15,32'd15,32'd8,32'd8,32'd12,32'd12,32'd20,32'd4,32'd14,32'd14,32'd14,32'd15,32'd8,32'd3,32'd4,32'd12,32'd9,32'd9,32'd18,32'd6,32'd6,32'd22,32'd12,32'd6,32'd18,32'd18,32'd6,32'd18,32'd6,32'd3,32'd10,32'd3,32'd15,32'd6,32'd4,32'd6,32'd3,32'd3,32'd9,32'd6,32'd9,32'd9,32'd6,32'd6,32'd9,32'd9,32'd9,32'd10,32'd4,32'd3,32'd9,32'd9,32'd9,32'd18,32'd6,32'd9,32'd3,32'd6,32'd6,32'd6,32'd9,32'd10,32'd18,32'd18,32'd6,32'd4,32'd6,32'd2,32'd14,32'd14,32'd7,32'd8,32'd6,32'd11,32'd17,32'd17,32'd10,32'd3,32'd3,32'd3,32'd18,32'd18,32'd3,32'd18,32'd10,32'd10,32'd10,32'd10,32'd6,32'd18,32'd10,32'd10,32'd19,32'd19,32'd15,32'd12,32'd4,32'd15,32'd9,32'd12,32'd3,32'd2,32'd6,32'd6,32'd6,32'd6,32'd12,32'd12,32'd8,32'd8,32'd4,32'd6,32'd4,32'd3,32'd18,32'd18,32'd16,32'd19,32'd6,32'd3,32'd6,32'd3,32'd6,32'd6,32'd13,32'd6,32'd12,32'd9,32'd6,32'd4,32'd10,32'd3,32'd3,32'd18,32'd6,32'd6,32'd14,32'd14,32'd4,32'd3,32'd9,32'd9,32'd10,32'd10,32'd18,32'd3,32'd6,32'd2,32'd9,32'd8,32'd11,32'd3,32'd10,32'd2,32'd3,32'd5,32'd14,32'd6,32'd15,32'd15,32'd9,32'd9,32'd6,32'd2,32'd3,32'd18,32'd6,32'd6,32'd6,32'd8,32'd5,32'd6,32'd9,32'd12,32'd8,32'd6,32'd6,32'd6,32'd8,32'd6,32'd12,32'd16,32'd9,32'd20,32'd20,32'd22,32'd22,32'd14,32'd14,32'd16,32'd16,32'd16,32'd4,32'd8,32'd4,32'd3,32'd10,32'd6,32'd3,32'd2,32'd8,32'd24,32'd24,32'd13,32'd12,32'd15,32'd4,32'd22,32'd22,32'd9,32'd10,32'd8,32'd6,32'd12,32'd12,32'd20,32'd6,32'd9,32'd6,32'd7,32'd5,32'd6,32'd5,32'd5,32'd6,32'd16,32'd16,32'd19,32'd18,32'd4,32'd8,32'd8,32'd10,32'd9,32'd9,32'd6,32'd6,32'd12,32'd4,32'd14,32'd14,32'd6,32'd5,32'd10,32'd14,32'd6,32'd24,32'd3,32'd3,32'd22,32'd6,32'd9,32'd12,32'd8,32'd9,32'd6,32'd6,32'd16,32'd10,32'd10,32'd6,32'd7,32'd7,32'd9,32'd3,32'd18,32'd18,32'd19,32'd5,32'd6,32'd6,32'd18,32'd23,32'd20,32'd4,32'd9,32'd9,32'd6,32'd6,32'd9,32'd24,32'd15,32'd24,32'd10,32'd3,32'd3,32'd7,32'd12,32'd12,32'd4,32'd8,32'd9,32'd4,32'd8,32'd4,32'd8,32'd16,32'd7,32'd6,32'd2,32'd5,32'd10,32'd10,32'd10,32'd10,32'd18,32'd8,32'd5,32'd7,32'd9,32'd10,32'd9,32'd12,32'd12,32'd9,32'd3,32'd2,32'd14,32'd6,32'd12,32'd6,32'd6,32'd12,32'd24,32'd24,32'd9,32'd12,32'd6,32'd7,32'd15,32'd6,32'd13,32'd6,32'd6,32'd6,32'd7,32'd3,32'd6,32'd3,32'd6,32'd6,32'd20,32'd20,32'd6,32'd9,32'd18,32'd6,32'd12,32'd18,32'd20,32'd20,32'd3,32'd3,32'd9,32'd3,32'd12,32'd3,32'd8,32'd12,32'd9,32'd6,32'd6,32'd3,32'd3,32'd6,32'd6,32'd6,32'd9,32'd3,32'd6,32'd6,32'd3,32'd12,32'd6,32'd4,32'd6,32'd18,32'd6,32'd7,32'd6,32'd4,32'd14,32'd5,32'd9,32'd20,32'd9,32'd6,32'd15,32'd6,32'd4,32'd3,32'd8,32'd12,32'd12,32'd12,32'd8,32'd7,32'd7,32'd9,32'd9,32'd10,32'd7,32'd5,32'd5,32'd5,32'd9,32'd14,32'd6,32'd19,32'd5,32'd6,32'd7,32'd9,32'd7,32'd19,32'd7,32'd6,32'd7,32'd3,32'd12,32'd8,32'd3,32'd6,32'd4,32'd12,32'd24,32'd6,32'd6,32'd4,32'd4,32'd20,32'd22,32'd12,32'd12,32'd7,32'd12,32'd2,32'd14,32'd18,32'd6,32'd14,32'd12,32'd20,32'd18,32'd18,32'd12,32'd14,32'd8,32'd12,32'd12,32'd8,32'd8,32'd6,32'd18,32'd9,32'd9,32'd22,32'd22,32'd4,32'd6,32'd4,32'd9,32'd6,32'd6,32'd2,32'd6,32'd20,32'd5,32'd9,32'd9,32'd9,32'd9,32'd3,32'd4,32'd10,32'd15,32'd6,32'd6,32'd10,32'd6,32'd8,32'd18,32'd6,32'd2,32'd19,32'd19,32'd6,32'd3,32'd6,32'd9,32'd18,32'd6,32'd4,32'd12,32'd10,32'd6,32'd15,32'd4,32'd6,32'd8,32'd12,32'd12,32'd20,32'd20,32'd6,32'd5,32'd9,32'd20,32'd3,32'd19,32'd9,32'd20,32'd3,32'd3,32'd4,32'd4,32'd20,32'd20,32'd15,32'd15,32'd8,32'd6,32'd6,32'd19,32'd7,32'd7,32'd24,32'd24,32'd6,32'd14,32'd9,32'd20,32'd9,32'd9,32'd14,32'd18,32'd4,32'd24,32'd22,32'd22,32'd3,32'd3,32'd6,32'd6,32'd4,32'd6,32'd12,32'd12,32'd18,32'd9,32'd9,32'd9,32'd12,32'd16,32'd8,32'd9,32'd6,32'd9,32'd9,32'd4,32'd16,32'd6,32'd2,32'd4,32'd10,32'd10,32'd9,32'd10,32'd14,32'd6,32'd3,32'd15,32'd3,32'd9,32'd15,32'd3,32'd22,32'd22,32'd6,32'd10,32'd4,32'd3,32'd12,32'd8,32'd19,32'd4,32'd4,32'd4,32'd6,32'd4,32'd4,32'd9,32'd9,32'd12,32'd12,32'd12,32'd12,32'd9,32'd8,32'd10,32'd21,32'd10,32'd6,32'd7,32'd9,32'd6,32'd6,32'd4,32'd4,32'd9,32'd16,32'd14,32'd8,32'd12,32'd18,32'd20,32'd20,32'd3,32'd6,32'd4,32'd8,32'd12,32'd18,32'd12,32'd6,32'd23,32'd6,32'd6,32'd12,32'd6,32'd4,32'd5,32'd6,32'd10,32'd15,32'd4,32'd12,32'd8,32'd8,32'd9,32'd10,32'd14,32'd15,32'd3,32'd6,32'd18,32'd18,32'd12,32'd9,32'd8,32'd8,32'd9,32'd5,32'd9,32'd9,32'd20,32'd24,32'd10,32'd10,32'd16,32'd16,32'd6,32'd6,32'd6,32'd3,32'd3,32'd13,32'd2,32'd6,32'd6,32'd10,32'd4,32'd12,32'd18,32'd5,32'd7,32'd5,32'd7,32'd5,32'd10,32'd10,32'd18,32'd6,32'd10,32'd9,32'd6,32'd18,32'd3,32'd18,32'd3,32'd3,32'd4,32'd4,32'd6,32'd3,32'd21,32'd10,32'd3,32'd3,32'd10,32'd11,32'd3,32'd3,32'd9,32'd10,32'd13,32'd3,32'd18,32'd8,32'd3,32'd6,32'd14,32'd4,32'd15,32'd13,32'd6,32'd20,32'd9,32'd6,32'd10,32'd10,32'd12,32'd5,32'd12,32'd3,32'd18,32'd3,32'd9,32'd14,32'd5,32'd4,32'd3,32'd18,32'd3,32'd15,32'd9,32'd3,32'd3,32'd3,32'd20,32'd9,32'd6,32'd9,32'd14,32'd9,32'd3,32'd6,32'd11,32'd11,32'd9,32'd13,32'd13,32'd10,32'd16,32'd10,32'd9,32'd9,32'd9,32'd2,32'd3,32'd9,32'd15,32'd5,32'd9,32'd3,32'd3,32'd6,32'd6,32'd4,32'd9,32'd8,32'd8,32'd22,32'd8,32'd3,32'd10,32'd6,32'd6,32'd6,32'd14,32'd12,32'd16,32'd18,32'd12,32'd10,32'd3,32'd10,32'd6,32'd7,32'd12,32'd8,32'd6,32'd9,32'd6,32'd20,32'd20,32'd18,32'd9,32'd9,32'd8,32'd6,32'd4,32'd6,32'd6,32'd8,32'd6,32'd6,32'd4,32'd9,32'd20,32'd19,32'd20,32'd8,32'd20,32'd3,32'd20,32'd9,32'd9,32'd10,32'd9,32'd5,32'd5,32'd7,32'd3,32'd14,32'd6,32'd9,32'd9,32'd6,32'd2,32'd3,32'd8,32'd4,32'd3,32'd16,32'd16,32'd16,32'd16,32'd12,32'd12,32'd15,32'd4,32'd7,32'd4,32'd22,32'd22,32'd4,32'd9,32'd12,32'd22,32'd9,32'd9,32'd12,32'd9,32'd3,32'd21,32'd12,32'd6,32'd6,32'd6,32'd4,32'd5,32'd3,32'd6,32'd8,32'd14,32'd24,32'd6,32'd14,32'd5,32'd4,32'd2,32'd6,32'd19,32'd13,32'd5,32'd10,32'd9,32'd4,32'd6,32'd4,32'd14,32'd6,32'd6,32'd13,32'd13,32'd10,32'd9,32'd4,32'd8,32'd14,32'd6,32'd8,32'd6,32'd9,32'd6,32'd10,32'd3,32'd4,32'd4,32'd6,32'd8,32'd9,32'd9,32'd6,32'd6,32'd6,32'd6,32'd8,32'd8,32'd9,32'd6,32'd3,32'd10,32'd14,32'd3,32'd8,32'd8,32'd6,32'd3,32'd8,32'd12,32'd12,32'd4,32'd6,32'd8,32'd3,32'd12,32'd11,32'd6,32'd6,32'd9,32'd9,32'd9,32'd18,32'd18,32'd14,32'd9,32'd4,32'd6,32'd18,32'd6,32'd4,32'd4,32'd9,32'd14,32'd20,32'd20,32'd9,32'd9,32'd3,32'd2,32'd3,32'd4,32'd6,32'd9,32'd8,32'd6,32'd5,32'd9,32'd3,32'd6,32'd2,32'd10,32'd5,32'd5,32'd7,32'd7,32'd8,32'd2,32'd6,32'd6,32'd4,32'd9,32'd4,32'd7,32'd18,32'd12,32'd6,32'd3,32'd3,32'd6,32'd12,32'd21,32'd6,32'd6,32'd2,32'd9,32'd9,32'd9,32'd13,32'd3,32'd8,32'd8,32'd18,32'd18,32'd11,32'd6,32'd6,32'd5,32'd9,32'd6,32'd12,32'd3,32'd12,32'd12,32'd5,32'd2,32'd8,32'd8,32'd4,32'd6,32'd9,32'd14,32'd18,32'd5,32'd3,32'd5,32'd12,32'd4,32'd9,32'd18,32'd9,32'd10,32'd3,32'd9,32'd6,32'd6,32'd7,32'd9,32'd13,32'd13,32'd6,32'd6,32'd17,32'd17,32'd20,32'd20,32'd14,32'd14,32'd12,32'd18,32'd14,32'd6,32'd12,32'd12,32'd7,32'd6,32'd8,32'd9,32'd9,32'd6,32'd12,32'd9,32'd12,32'd4,32'd6,32'd6,32'd3,32'd9,32'd6,32'd3,32'd6,32'd9,32'd6,32'd6,32'd9,32'd4,32'd6,32'd4,32'd8,32'd6,32'd22,32'd5,32'd9,32'd6,32'd10,32'd4,32'd12,32'd12,32'd10,32'd9,32'd8,32'd4,32'd11,32'd18,32'd9,32'd9,32'd3,32'd9,32'd10,32'd4,32'd24,32'd12,32'd10,32'd4,32'd10,32'd12,32'd9,32'd14,32'd12,32'd10,32'd23,32'd3,32'd6,32'd23,32'd3,32'd2,32'd4,32'd4,32'd2,32'd2,32'd6,32'd3,32'd21,32'd21,32'd10,32'd6,32'd4,32'd8,32'd15,32'd6,32'd16,32'd8,32'd9,32'd4,32'd9,32'd12,32'd4,32'd9,32'd9,32'd9,32'd20,32'd6,32'd12,32'd16,32'd6,32'd6,32'd9,32'd9,32'd16,32'd16,32'd9,32'd9,32'd6,32'd9,32'd9,32'd9,32'd10,32'd3,32'd6,32'd3,32'd12,32'd6,32'd13,32'd11,32'd9,32'd12,32'd12,32'd10,32'd2,32'd6,32'd12,32'd10,32'd10,32'd6,32'd3,32'd5,32'd3,32'd3,32'd6,32'd8,32'd6,32'd6,32'd6,32'd3,32'd4,32'd9,32'd12,32'd15,32'd6,32'd8,32'd8,32'd8,32'd9,32'd9,32'd2,32'd13,32'd9,32'd12,32'd3,32'd6,32'd4,32'd13,32'd3,32'd9,32'd9,32'd9,32'd6,32'd4,32'd4,32'd18,32'd18,32'd12,32'd22,32'd16,32'd6,32'd9,32'd6,32'd10,32'd10,32'd7,32'd5,32'd6,32'd4,32'd3,32'd6,32'd8,32'd3,32'd4,32'd15,32'd12,32'd3,32'd13,32'd2,32'd10,32'd12,32'd12,32'd10,32'd9,32'd9,32'd18,32'd12,32'd10,32'd14,32'd3,32'd3,32'd8,32'd6,32'd7,32'd7,32'd4,32'd6,32'd6,32'd6,32'd2,32'd6,32'd16,32'd16,32'd18,32'd4,32'd11,32'd3,32'd6,32'd10,32'd24,32'd24,32'd6,32'd2,32'd13,32'd9,32'd9,32'd2,32'd6,32'd16,32'd12,32'd9,32'd12,32'd12,32'd8,32'd10,32'd4,32'd6,32'd8,32'd6,32'd10,32'd6,32'd4,32'd10,32'd9,32'd6,32'd6,32'd6,32'd9,32'd6,32'd4,32'd6,32'd3,32'd8,32'd6,32'd6,32'd3,32'd6,32'd3,32'd15,32'd9,32'd9,32'd5,32'd6,32'd3,32'd6,32'd18,32'd10,32'd11,32'd11,32'd9,32'd6,32'd3,32'd10,32'd6,32'd9,32'd6,32'd3,32'd9,32'd6,32'd14,32'd9,32'd18,32'd4,32'd6,32'd6,32'd7,32'd9,32'd9,32'd5,32'd6,32'd3,32'd6,32'd13,32'd10,32'd9,32'd9,32'd2,32'd6,32'd4,32'd4,32'd8,32'd12,32'd10,32'd10,32'd8,32'd4,32'd15,32'd12,32'd6,32'd6,32'd6,32'd4,32'd3,32'd10,32'd3,32'd9,32'd21,32'd8,32'd6,32'd10,32'd9,32'd9,32'd16,32'd4,32'd6,32'd12,32'd6,32'd9,32'd6,32'd6,32'd9,32'd3,32'd2,32'd3,32'd10,32'd9,32'd12,32'd9,32'd6,32'd16,32'd11,32'd10,32'd9,32'd8,32'd14,32'd14,32'd20,32'd20,32'd6,32'd20,32'd12,32'd12,32'd8,32'd18,32'd21,32'd21,32'd16,32'd12,32'd14,32'd14,32'd18,32'd6,32'd8,32'd5,32'd8,32'd8,32'd12,32'd12,32'd4,32'd6,32'd2,32'd15,32'd16,32'd16,32'd5,32'd5,32'd4,32'd6,32'd10,32'd16,32'd14,32'd14,32'd9,32'd9,32'd8,32'd5,32'd18,32'd13,32'd4,32'd13,32'd6,32'd3,32'd9,32'd9,32'd9,32'd12,32'd15,32'd4,32'd6,32'd3,32'd6,32'd4,32'd3,32'd3,32'd23,32'd4,32'd3,32'd23,32'd9,32'd9,32'd4,32'd6,32'd6,32'd6,32'd6,32'd3,32'd6,32'd6,32'd6,32'd9,32'd9,32'd9,32'd8,32'd9,32'd9,32'd8,32'd18,32'd18,32'd18,32'd3,32'd17,32'd17,32'd6,32'd17,32'd8,32'd9,32'd4,32'd6,32'd8,32'd9,32'd8,32'd14,32'd10,32'd4,32'd4,32'd20,32'd3,32'd5,32'd18,32'd11,32'd11,32'd6,32'd7,32'd9,32'd3,32'd7,32'd4,32'd11,32'd12,32'd8,32'd8,32'd6,32'd6,32'd9,32'd9,32'd6,32'd6,32'd8,32'd8,32'd14,32'd12,32'd9,32'd10,32'd7,32'd9,32'd6,32'd10,32'd14,32'd14,32'd8,32'd12,32'd4,32'd24,32'd6,32'd3,32'd6,32'd6,32'd9,32'd9,32'd6,32'd6,32'd10,32'd6,32'd9,32'd6,32'd14,32'd4,32'd6,32'd9,32'd3,32'd3,32'd12,32'd3,32'd5,32'd12,32'd8,32'd14,32'd12,32'd12,32'd20,32'd20,32'd19,32'd19,32'd4,32'd8,32'd15,32'd9,32'd15,32'd15,32'd12,32'd12,32'd9,32'd7,32'd12,32'd12,32'd14,32'd3,32'd6,32'd23,32'd9,32'd6,32'd12,32'd9,32'd7,32'd8,32'd9,32'd12,32'd4,32'd9,32'd3,32'd3,32'd8,32'd12,32'd18,32'd6,32'd8,32'd10,32'd6,32'd6,32'd19,32'd14,32'd10,32'd10,32'd4,32'd18,32'd9,32'd10,32'd12,32'd10,32'd6,32'd10,32'd6,32'd3,32'd6,32'd6,32'd3,32'd6,32'd9,32'd9,32'd9,32'd9,32'd10,32'd6,32'd9,32'd9,32'd9,32'd9,32'd2,32'd2,32'd3,32'd9,32'd11,32'd11,32'd22,32'd22,32'd12,32'd12,32'd4,32'd2,32'd6,32'd9,32'd9,32'd9,32'd18,32'd6,32'd3,32'd2,32'd8,32'd9,32'd12,32'd3,32'd16,32'd6,32'd9,32'd21,32'd10,32'd10,32'd11,32'd6,32'd6,32'd9,32'd6,32'd13,32'd16,32'd4,32'd6,32'd10,32'd6,32'd2,32'd6,32'd10,32'd6,32'd16,32'd10,32'd6,32'd6,32'd6,32'd6,32'd22,32'd6,32'd12,32'd12,32'd16,32'd9,32'd8,32'd8,32'd9,32'd6,32'd4,32'd6,32'd6,32'd9,32'd9,32'd7,32'd4,32'd6,32'd20,32'd3,32'd3,32'd4,32'd4,32'd4,32'd9,32'd9,32'd13,32'd15,32'd11,32'd2,32'd6,32'd6,32'd6,32'd4,32'd8,32'd15,32'd8,32'd10,32'd9,32'd9,32'd6,32'd6,32'd8,32'd4,32'd16,32'd3,32'd9,32'd3,32'd6,32'd9,32'd18,32'd18,32'd9,32'd9,32'd3,32'd9,32'd3,32'd9,32'd3,32'd12,32'd4,32'd9,32'd11,32'd11,32'd6,32'd11,32'd2,32'd3,32'd3,32'd3,32'd6,32'd6,32'd6,32'd6,32'd10,32'd9,32'd6,32'd14,32'd9,32'd6,32'd8,32'd10,32'd12,32'd6,32'd14,32'd4,32'd9,32'd9,32'd10,32'd9,32'd3,32'd9,32'd9,32'd6,32'd20,32'd21,32'd13,32'd21,32'd6,32'd6,32'd10,32'd10,32'd9,32'd9,32'd8,32'd13,32'd3,32'd2,32'd21,32'd9,32'd9,32'd9,32'd6,32'd3,32'd15,32'd4,32'd3,32'd6,32'd14,32'd4,32'd18,32'd4,32'd4,32'd6,32'd6,32'd4,32'd8,32'd8,32'd8,32'd6,32'd10,32'd6,32'd4,32'd4,32'd16,32'd9,32'd9,32'd4,32'd20,32'd17,32'd10,32'd10,32'd6,32'd4,32'd9,32'd6,32'd3,32'd8,32'd7,32'd6,32'd3,32'd12,32'd4,32'd9,32'd6,32'd4,32'd3,32'd4,32'd3,32'd4,32'd3,32'd4,32'd6,32'd6,32'd14,32'd12,32'd15,32'd6,32'd5,32'd5,32'd6,32'd3,32'd8,32'd6,32'd4,32'd4,32'd9,32'd4,32'd3,32'd3,32'd12,32'd18,32'd5,32'd12,32'd19,32'd9,32'd4,32'd19,32'd9,32'd19,32'd9,32'd9,32'd10,32'd10,32'd9,32'd5,32'd4,32'd9,32'd3,32'd6,32'd4,32'd9,32'd6,32'd14,32'd14,32'd14,32'd3,32'd2,32'd12,32'd12,32'd3,32'd6,32'd8,32'd9,32'd9,32'd5,32'd12,32'd14,32'd6,32'd6,32'd4,32'd3,32'd8,32'd8,32'd19,32'd19,32'd9,32'd9,32'd6,32'd3,32'd6,32'd8,32'd9,32'd11,32'd3,32'd8,32'd9,32'd2,32'd8,32'd10,32'd16,32'd16,32'd4,32'd16,32'd6,32'd9,32'd3,32'd18,32'd6,32'd14,32'd14,32'd18,32'd8,32'd12,32'd6,32'd16,32'd16,32'd7,32'd4,32'd10,32'd16,32'd2,32'd14,32'd6,32'd16,32'd9,32'd12,32'd12,32'd14,32'd9,32'd6,32'd10,32'd10,32'd9,32'd6,32'd14,32'd4,32'd6,32'd3,32'd12,32'd6,32'd16,32'd2,32'd6,32'd6,32'd9,32'd7,32'd13,32'd13,32'd3,32'd9,32'd10,32'd10,32'd10,32'd9,32'd10,32'd9,32'd18,32'd10,32'd22,32'd6,32'd16,32'd3,32'd6,32'd3,32'd6,32'd2,32'd6,32'd6,32'd6,32'd10,32'd6,32'd9,32'd4,32'd4,32'd3,32'd15,32'd4,32'd3,32'd4,32'd3,32'd23,32'd23,32'd6,32'd4,32'd9,32'd4,32'd4,32'd2,32'd14,32'd6,32'd3,32'd6,32'd13,32'd13,32'd6,32'd6,32'd12,32'd4,32'd5,32'd12,32'd3,32'd5,32'd10,32'd16,32'd14,32'd9,32'd14,32'd6,32'd6,32'd3,32'd6,32'd9,32'd12,32'd9,32'd6,32'd10,32'd12,32'd8,32'd6,32'd14,32'd9,32'd6,32'd10,32'd3,32'd6,32'd12,32'd3,32'd6,32'd6,32'd4,32'd9,32'd9,32'd9,32'd5,32'd3,32'd6,32'd2,32'd6,32'd2,32'd15,32'd6,32'd6,32'd12,32'd9,32'd6,32'd5,32'd8,32'd12,32'd18,32'd4,32'd9,32'd3,32'd4,32'd9,32'd6,32'd12,32'd4,32'd6,32'd4,32'd3,32'd8,32'd10,32'd5,32'd4,32'd4,32'd5,32'd9,32'd4,32'd4,32'd10,32'd20,32'd14,32'd8,32'd14,32'd9,32'd9,32'd8,32'd22,32'd4,32'd3,32'd8,32'd12,32'd12,32'd6,32'd9,32'd11,32'd8,32'd8,32'd9,32'd10,32'd3,32'd6,32'd6,32'd3,32'd4,32'd3,32'd6,32'd6,32'd6,32'd4,32'd4,32'd3,32'd10,32'd4,32'd4,32'd14,32'd6,32'd5,32'd10,32'd18,32'd8,32'd6,32'd6,32'd9,32'd4,32'd5,32'd4,32'd3,32'd3,32'd12,32'd11,32'd9,32'd12,32'd18,32'd18,32'd12,32'd12,32'd2,32'd10,32'd14,32'd12,32'd8,32'd12,32'd3,32'd3,32'd11,32'd10,32'd18,32'd18,32'd9,32'd14,32'd12,32'd3,32'd9,32'd7,32'd3,32'd15,32'd12,32'd12,32'd9,32'd6,32'd17,32'd10,32'd11,32'd6,32'd2,32'd12,32'd9,32'd12,32'd18,32'd17,32'd4,32'd4,32'd8,32'd15,32'd4,32'd8,32'd5,32'd8,32'd9,32'd4,32'd4,32'd18,32'd18,32'd6,32'd6,32'd8,32'd6,32'd15,32'd10,32'd6,32'd12,32'd6,32'd9,32'd19,32'd23,32'd18,32'd3,32'd3,32'd18,32'd2,32'd9,32'd3,32'd6,32'd12,32'd5,32'd4,32'd6,32'd5,32'd13,32'd10,32'd10,32'd6,32'd6,32'd9,32'd6,32'd6,32'd6,32'd6,32'd6,32'd10,32'd10,32'd9,32'd7,32'd14,32'd14,32'd6,32'd6,32'd20,32'd20,32'd19,32'd6,32'd12,32'd8,32'd6,32'd10,32'd4,32'd3,32'd9,32'd19,32'd6,32'd19,32'd9,32'd6,32'd9,32'd9,32'd9,32'd12,32'd6,32'd6,32'd22,32'd3,32'd3,32'd10,32'd6,32'd3,32'd3,32'd5,32'd11,32'd18,32'd8,32'd8,32'd9,32'd4,32'd16,32'd10,32'd6,32'd4,32'd9,32'd9,32'd11,32'd6,32'd3,32'd15,32'd9,32'd9,32'd4,32'd12,32'd7,32'd6,32'd6,32'd7,32'd3,32'd6,32'd6,32'd18,32'd3,32'd6,32'd7,32'd10,32'd6,32'd6,32'd4,32'd3,32'd9,32'd8,32'd8,32'd20,32'd4,32'd10,32'd3,32'd9,32'd18,32'd12,32'd12,32'd21,32'd9,32'd15,32'd15,32'd9,32'd14,32'd6,32'd6,32'd15,32'd15,32'd12,32'd12,32'd18,32'd4,32'd17,32'd17,32'd6,32'd6,32'd4,32'd9,32'd9,32'd9,32'd11,32'd11,32'd3,32'd18,32'd10,32'd6,32'd9,32'd3,32'd9,32'd8,32'd16,32'd16,32'd9,32'd6,32'd14,32'd14,32'd15,32'd14,32'd22,32'd9,32'd9,32'd4,32'd3,32'd8,32'd8,32'd21,32'd12,32'd12,32'd10,32'd9,32'd3,32'd6,32'd9,32'd18,32'd10,32'd7,32'd9,32'd18,32'd6,32'd10,32'd5,32'd5,32'd16,32'd10,32'd9,32'd9,32'd6,32'd6,32'd3,32'd9,32'd6,32'd6,32'd6,32'd6,32'd16,32'd6,32'd6,32'd12,32'd10,32'd15,32'd12,32'd6,32'd3,32'd6,32'd5,32'd5,32'd9,32'd8,32'd10,32'd12,32'd3,32'd13,32'd9,32'd18,32'd12,32'd6,32'd3,32'd7,32'd9,32'd10,32'd6,32'd18,32'd14,32'd9,32'd15,32'd14,32'd9,32'd6,32'd14,32'd12,32'd14,32'd24,32'd24,32'd20,32'd6,32'd11,32'd24,32'd10,32'd3,32'd6,32'd6,32'd3,32'd4,32'd10,32'd10,32'd6,32'd6,32'd8,32'd2,32'd4,32'd16,32'd3,32'd6,32'd12,32'd9,32'd4,32'd24,32'd2,32'd4,32'd6,32'd12,32'd3,32'd3,32'd9,32'd9,32'd10,32'd7,32'd9,32'd9,32'd9,32'd9,32'd2,32'd4,32'd9,32'd9,32'd6,32'd9,32'd14,32'd11,32'd5,32'd6,32'd14,32'd14,32'd6,32'd6,32'd4,32'd6,32'd12,32'd12,32'd7,32'd19,32'd6,32'd9,32'd17,32'd9,32'd12,32'd12,32'd4,32'd9,32'd7,32'd21,32'd9,32'd10,32'd9,32'd4,32'd12,32'd9,32'd9,32'd3,32'd6,32'd3,32'd12,32'd4,32'd3,32'd9,32'd4,32'd6,32'd6,32'd18,32'd4,32'd23,32'd6,32'd3,32'd9,32'd8,32'd12,32'd12,32'd9,32'd12,32'd12,32'd12,32'd6,32'd3,32'd3,32'd6,32'd6,32'd12,32'd12,32'd9,32'd9,32'd20,32'd14,32'd22,32'd6,32'd4,32'd9,32'd3,32'd9,32'd19,32'd19,32'd4,32'd6,32'd14,32'd6,32'd15,32'd6,32'd6,32'd6,32'd9,32'd9,32'd6,32'd2,32'd9,32'd9,32'd6,32'd9,32'd18,32'd18,32'd12,32'd14,32'd9,32'd6,32'd2,32'd8,32'd16,32'd14,32'd10,32'd12,32'd5,32'd9,32'd4,32'd10,32'd3,32'd10,32'd16,32'd12,32'd16,32'd6,32'd14,32'd9,32'd18,32'd18,32'd9,32'd3,32'd3,32'd16,32'd8,32'd10,32'd7,32'd4,32'd15,32'd15,32'd9,32'd9,32'd9,32'd4,32'd9,32'd9,32'd4,32'd9,32'd4,32'd2,32'd12,32'd10,32'd19,32'd12,32'd10,32'd12,32'd19,32'd4,32'd6,32'd6,32'd4,32'd4,32'd23,32'd21,32'd9,32'd20,32'd9,32'd12,32'd21,32'd3,32'd9,32'd6,32'd9,32'd9,32'd6,32'd9,32'd6,32'd16,32'd6,32'd6,32'd12,32'd12,32'd5,32'd12,32'd14,32'd6,32'd10,32'd14,32'd13,32'd15,32'd9,32'd6,32'd4,32'd16,32'd4,32'd4,32'd3,32'd19,32'd9,32'd8,32'd6,32'd18,32'd4,32'd10,32'd18,32'd18,32'd6,32'd4,32'd3,32'd3,32'd9,32'd14,32'd10,32'd6,32'd4,32'd9,32'd4,32'd4,32'd6,32'd6,32'd9,32'd9,32'd13,32'd13,32'd14,32'd9,32'd6,32'd9,32'd3,32'd15,32'd12,32'd10,32'd6,32'd11,32'd4,32'd4,32'd9,32'd3,32'd2,32'd12,32'd9,32'd18,32'd9,32'd2,32'd3,32'd9,32'd8,32'd9,32'd16,32'd16,32'd6,32'd6,32'd4,32'd3,32'd18,32'd3,32'd4,32'd6,32'd18,32'd22,32'd22,32'd24,32'd24,32'd17,32'd12,32'd4,32'd6,32'd6,32'd6,32'd8,32'd3,32'd3,32'd6,32'd9,32'd6,32'd6,32'd6,32'd4,32'd6,32'd4,32'd6,32'd16,32'd6,32'd14,32'd8,32'd14,32'd18,32'd11,32'd11,32'd10,32'd14,32'd6,32'd12,32'd6,32'd16,32'd22,32'd22,32'd7,32'd8,32'd10,32'd9,32'd15,32'd6,32'd6,32'd4,32'd4,32'd12,32'd6,32'd6,32'd10,32'd4,32'd13,32'd2,32'd14,32'd18,32'd6,32'd6,32'd8,32'd3,32'd12,32'd12,32'd10,32'd24,32'd12,32'd2,32'd3,32'd10,32'd6,32'd6,32'd9,32'd9,32'd6,32'd6,32'd6,32'd9,32'd9,32'd6,32'd10,32'd10,32'd15,32'd3,32'd3,32'd2,32'd4,32'd6,32'd10,32'd10,32'd2,32'd12,32'd9,32'd9,32'd4,32'd9,32'd3,32'd6,32'd12,32'd6,32'd9,32'd4,32'd9,32'd9,32'd9,32'd9,32'd9,32'd5,32'd14,32'd10,32'd6,32'd6,32'd9,32'd12,32'd14,32'd2,32'd20,32'd12,32'd3,32'd6,32'd12,32'd6,32'd6,32'd14,32'd12,32'd23,32'd13,32'd13,32'd6,32'd6,32'd5,32'd6,32'd9,32'd9,32'd11,32'd2,32'd14,32'd9,32'd9,32'd3,32'd9,32'd11,32'd9,32'd19,32'd13,32'd13,32'd10,32'd10,32'd12,32'd12,32'd15,32'd15,32'd15,32'd6,32'd3,32'd12,32'd10,32'd14,32'd6,32'd3,32'd12,32'd6,32'd9,32'd13,32'd11,32'd9,32'd10,32'd10,32'd6,32'd9,32'd10,32'd15,32'd3,32'd12,32'd7,32'd6,32'd6,32'd10,32'd6,32'd16,32'd19,32'd6,32'd9,32'd7,32'd9}
`define RECTANGLE1_WEIGHTS {32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168,32'd4294967168}
`define RECTANGLE2_XS {32'd12,32'd0,32'd17,32'd3,32'd12,32'd0,32'd15,32'd0,32'd3,32'd0,32'd15,32'd1,32'd15,32'd0,32'd21,32'd12,32'd0,32'd0,32'd16,32'd3,32'd13,32'd3,32'd13,32'd10,32'd14,32'd2,32'd6,32'd5,32'd15,32'd1,32'd18,32'd0,32'd20,32'd5,32'd12,32'd3,32'd18,32'd2,32'd11,32'd9,32'd5,32'd5,32'd11,32'd8,32'd14,32'd9,32'd14,32'd4,32'd5,32'd12,32'd9,32'd8,32'd14,32'd10,32'd12,32'd2,32'd6,32'd9,32'd5,32'd8,32'd8,32'd1,32'd9,32'd0,32'd5,32'd1,32'd12,32'd1,32'd10,32'd1,32'd8,32'd4,32'd4,32'd5,32'd12,32'd6,32'd0,32'd1,32'd9,32'd10,32'd12,32'd12,32'd12,32'd0,32'd7,32'd1,32'd14,32'd1,32'd11,32'd11,32'd12,32'd0,32'd12,32'd5,32'd6,32'd3,32'd18,32'd10,32'd12,32'd4,32'd8,32'd6,32'd12,32'd7,32'd2,32'd0,32'd6,32'd9,32'd12,32'd0,32'd12,32'd0,32'd15,32'd6,32'd14,32'd5,32'd12,32'd3,32'd17,32'd7,32'd16,32'd10,32'd4,32'd3,32'd4,32'd5,32'd12,32'd0,32'd5,32'd0,32'd14,32'd0,32'd15,32'd0,32'd19,32'd2,32'd17,32'd7,32'd18,32'd0,32'd3,32'd1,32'd21,32'd4,32'd20,32'd0,32'd6,32'd0,32'd0,32'd0,32'd18,32'd12,32'd11,32'd7,32'd6,32'd5,32'd9,32'd4,32'd6,32'd0,32'd11,32'd10,32'd9,32'd0,32'd17,32'd5,32'd3,32'd10,32'd10,32'd2,32'd20,32'd6,32'd6,32'd2,32'd5,32'd9,32'd9,32'd11,32'd2,32'd2,32'd5,32'd10,32'd8,32'd8,32'd13,32'd3,32'd16,32'd10,32'd11,32'd4,32'd5,32'd9,32'd11,32'd4,32'd15,32'd3,32'd12,32'd5,32'd10,32'd6,32'd9,32'd19,32'd9,32'd8,32'd0,32'd13,32'd3,32'd12,32'd12,32'd11,32'd4,32'd16,32'd5,32'd17,32'd2,32'd20,32'd3,32'd18,32'd7,32'd10,32'd8,32'd15,32'd2,32'd3,32'd7,32'd2,32'd2,32'd10,32'd6,32'd17,32'd9,32'd12,32'd10,32'd13,32'd8,32'd15,32'd11,32'd12,32'd4,32'd12,32'd0,32'd12,32'd4,32'd11,32'd8,32'd11,32'd12,32'd7,32'd9,32'd11,32'd8,32'd8,32'd2,32'd20,32'd2,32'd21,32'd0,32'd10,32'd8,32'd12,32'd0,32'd16,32'd1,32'd6,32'd3,32'd9,32'd3,32'd14,32'd10,32'd7,32'd1,32'd14,32'd5,32'd17,32'd0,32'd6,32'd10,32'd16,32'd10,32'd12,32'd9,32'd6,32'd0,32'd15,32'd3,32'd10,32'd4,32'd11,32'd10,32'd7,32'd9,32'd9,32'd3,32'd20,32'd1,32'd15,32'd0,32'd8,32'd1,32'd17,32'd2,32'd13,32'd0,32'd18,32'd3,32'd15,32'd7,32'd16,32'd8,32'd16,32'd4,32'd3,32'd0,32'd10,32'd6,32'd13,32'd9,32'd18,32'd7,32'd14,32'd7,32'd7,32'd3,32'd14,32'd10,32'd12,32'd10,32'd6,32'd5,32'd15,32'd1,32'd19,32'd9,32'd11,32'd10,32'd9,32'd7,32'd12,32'd10,32'd12,32'd3,32'd11,32'd0,32'd0,32'd0,32'd4,32'd8,32'd5,32'd7,32'd11,32'd9,32'd13,32'd9,32'd12,32'd3,32'd13,32'd9,32'd12,32'd10,32'd12,32'd9,32'd12,32'd11,32'd5,32'd5,32'd9,32'd1,32'd14,32'd2,32'd18,32'd0,32'd16,32'd7,32'd18,32'd0,32'd15,32'd0,32'd21,32'd7,32'd11,32'd12,32'd7,32'd7,32'd10,32'd8,32'd15,32'd8,32'd14,32'd0,32'd6,32'd0,32'd14,32'd0,32'd14,32'd0,32'd3,32'd8,32'd13,32'd8,32'd12,32'd4,32'd13,32'd6,32'd4,32'd3,32'd18,32'd8,32'd2,32'd4,32'd10,32'd5,32'd3,32'd5,32'd8,32'd9,32'd3,32'd15,32'd0,32'd4,32'd7,32'd13,32'd0,32'd18,32'd6,32'd15,32'd3,32'd18,32'd8,32'd18,32'd4,32'd16,32'd6,32'd11,32'd6,32'd9,32'd12,32'd16,32'd6,32'd18,32'd6,32'd18,32'd11,32'd18,32'd1,32'd18,32'd3,32'd12,32'd10,32'd6,32'd1,32'd8,32'd6,32'd15,32'd0,32'd15,32'd2,32'd13,32'd1,32'd7,32'd8,32'd12,32'd9,32'd12,32'd2,32'd12,32'd10,32'd12,32'd9,32'd14,32'd5,32'd4,32'd4,32'd12,32'd9,32'd12,32'd6,32'd15,32'd4,32'd15,32'd5,32'd11,32'd8,32'd11,32'd5,32'd17,32'd7,32'd0,32'd2,32'd17,32'd2,32'd10,32'd3,32'd14,32'd2,32'd9,32'd6,32'd13,32'd10,32'd12,32'd2,32'd12,32'd6,32'd10,32'd5,32'd16,32'd5,32'd3,32'd3,32'd0,32'd0,32'd1,32'd9,32'd13,32'd2,32'd4,32'd3,32'd12,32'd10,32'd6,32'd7,32'd12,32'd6,32'd15,32'd9,32'd6,32'd4,32'd12,32'd5,32'd16,32'd1,32'd15,32'd11,32'd11,32'd7,32'd15,32'd8,32'd13,32'd2,32'd14,32'd0,32'd10,32'd11,32'd7,32'd0,32'd22,32'd0,32'd19,32'd3,32'd12,32'd8,32'd9,32'd8,32'd13,32'd8,32'd15,32'd11,32'd12,32'd7,32'd22,32'd3,32'd14,32'd7,32'd13,32'd11,32'd15,32'd1,32'd21,32'd0,32'd6,32'd2,32'd13,32'd0,32'd14,32'd4,32'd17,32'd6,32'd12,32'd5,32'd14,32'd6,32'd9,32'd2,32'd12,32'd3,32'd13,32'd0,32'd7,32'd6,32'd8,32'd0,32'd13,32'd7,32'd17,32'd12,32'd17,32'd0,32'd11,32'd1,32'd7,32'd0,32'd11,32'd10,32'd5,32'd2,32'd20,32'd3,32'd19,32'd6,32'd8,32'd4,32'd7,32'd20,32'd5,32'd10,32'd3,32'd11,32'd5,32'd14,32'd10,32'd12,32'd2,32'd19,32'd6,32'd15,32'd10,32'd15,32'd9,32'd9,32'd8,32'd0,32'd9,32'd10,32'd9,32'd12,32'd0,32'd13,32'd9,32'd17,32'd7,32'd12,32'd10,32'd14,32'd5,32'd12,32'd2,32'd8,32'd6,32'd12,32'd9,32'd3,32'd0,32'd0,32'd6,32'd10,32'd0,32'd4,32'd7,32'd14,32'd6,32'd16,32'd3,32'd4,32'd4,32'd3,32'd5,32'd16,32'd5,32'd17,32'd12,32'd10,32'd11,32'd0,32'd4,32'd16,32'd3,32'd10,32'd7,32'd12,32'd7,32'd10,32'd6,32'd16,32'd3,32'd12,32'd9,32'd13,32'd8,32'd13,32'd2,32'd13,32'd0,32'd6,32'd0,32'd10,32'd1,32'd15,32'd2,32'd11,32'd0,32'd5,32'd10,32'd13,32'd10,32'd13,32'd10,32'd13,32'd7,32'd13,32'd1,32'd15,32'd0,32'd9,32'd7,32'd21,32'd3,32'd21,32'd7,32'd11,32'd7,32'd10,32'd0,32'd6,32'd12,32'd12,32'd2,32'd4,32'd0,32'd13,32'd0,32'd5,32'd5,32'd20,32'd2,32'd0,32'd7,32'd5,32'd2,32'd7,32'd7,32'd14,32'd5,32'd10,32'd4,32'd12,32'd1,32'd16,32'd2,32'd18,32'd9,32'd12,32'd5,32'd2,32'd9,32'd6,32'd10,32'd1,32'd12,32'd5,32'd0,32'd21,32'd2,32'd10,32'd11,32'd9,32'd9,32'd6,32'd4,32'd12,32'd10,32'd11,32'd5,32'd10,32'd2,32'd9,32'd3,32'd18,32'd7,32'd18,32'd3,32'd7,32'd9,32'd11,32'd0,32'd18,32'd2,32'd6,32'd0,32'd11,32'd3,32'd8,32'd4,32'd1,32'd4,32'd0,32'd14,32'd0,32'd14,32'd6,32'd12,32'd8,32'd12,32'd0,32'd13,32'd7,32'd11,32'd2,32'd13,32'd8,32'd12,32'd10,32'd16,32'd10,32'd1,32'd0,32'd14,32'd9,32'd13,32'd0,32'd10,32'd8,32'd14,32'd9,32'd13,32'd10,32'd12,32'd4,32'd9,32'd0,32'd15,32'd0,32'd16,32'd5,32'd17,32'd7,32'd3,32'd2,32'd13,32'd2,32'd13,32'd1,32'd13,32'd12,32'd13,32'd2,32'd20,32'd4,32'd9,32'd6,32'd12,32'd7,32'd6,32'd0,32'd4,32'd3,32'd15,32'd1,32'd6,32'd1,32'd1,32'd7,32'd0,32'd5,32'd17,32'd6,32'd16,32'd1,32'd19,32'd0,32'd7,32'd12,32'd14,32'd7,32'd15,32'd3,32'd14,32'd1,32'd15,32'd4,32'd18,32'd11,32'd11,32'd9,32'd9,32'd1,32'd1,32'd0,32'd9,32'd1,32'd11,32'd12,32'd12,32'd7,32'd14,32'd6,32'd11,32'd1,32'd11,32'd0,32'd4,32'd10,32'd12,32'd10,32'd11,32'd8,32'd10,32'd11,32'd12,32'd0,32'd13,32'd3,32'd11,32'd8,32'd14,32'd9,32'd10,32'd11,32'd10,32'd8,32'd14,32'd1,32'd14,32'd0,32'd0,32'd8,32'd6,32'd1,32'd13,32'd1,32'd9,32'd3,32'd15,32'd0,32'd14,32'd1,32'd14,32'd3,32'd15,32'd6,32'd12,32'd9,32'd15,32'd4,32'd6,32'd4,32'd9,32'd1,32'd3,32'd4,32'd19,32'd1,32'd9,32'd6,32'd7,32'd1,32'd20,32'd11,32'd12,32'd12,32'd13,32'd9,32'd13,32'd5,32'd17,32'd3,32'd14,32'd2,32'd12,32'd8,32'd7,32'd1,32'd12,32'd2,32'd14,32'd2,32'd20,32'd7,32'd15,32'd0,32'd1,32'd8,32'd11,32'd8,32'd15,32'd6,32'd10,32'd10,32'd6,32'd7,32'd9,32'd11,32'd13,32'd8,32'd12,32'd7,32'd14,32'd1,32'd0,32'd1,32'd13,32'd0,32'd11,32'd1,32'd14,32'd5,32'd6,32'd1,32'd5,32'd1,32'd12,32'd0,32'd21,32'd0,32'd17,32'd0,32'd8,32'd9,32'd13,32'd8,32'd7,32'd4,32'd14,32'd6,32'd15,32'd8,32'd14,32'd6,32'd6,32'd8,32'd18,32'd4,32'd2,32'd2,32'd17,32'd4,32'd6,32'd3,32'd16,32'd0,32'd14,32'd11,32'd10,32'd6,32'd8,32'd6,32'd16,32'd3,32'd6,32'd8,32'd10,32'd5,32'd12,32'd0,32'd5,32'd0,32'd12,32'd9,32'd16,32'd2,32'd20,32'd0,32'd15,32'd4,32'd18,32'd4,32'd16,32'd5,32'd17,32'd12,32'd18,32'd10,32'd13,32'd4,32'd17,32'd7,32'd13,32'd7,32'd11,32'd2,32'd14,32'd0,32'd13,32'd9,32'd12,32'd4,32'd9,32'd3,32'd14,32'd2,32'd5,32'd0,32'd8,32'd2,32'd16,32'd11,32'd7,32'd1,32'd12,32'd0,32'd14,32'd0,32'd9,32'd9,32'd13,32'd10,32'd7,32'd9,32'd12,32'd7,32'd8,32'd5,32'd15,32'd9,32'd12,32'd7,32'd15,32'd3,32'd15,32'd10,32'd7,32'd11,32'd10,32'd1,32'd15,32'd1,32'd11,32'd2,32'd17,32'd7,32'd10,32'd10,32'd6,32'd6,32'd13,32'd3,32'd6,32'd0,32'd15,32'd0,32'd4,32'd0,32'd6,32'd8,32'd12,32'd3,32'd12,32'd12,32'd15,32'd10,32'd13,32'd4,32'd16,32'd4,32'd3,32'd11,32'd4,32'd5,32'd14,32'd12,32'd14,32'd9,32'd7,32'd4,32'd14,32'd6,32'd9,32'd0,32'd14,32'd3,32'd19,32'd6,32'd16,32'd7,32'd16,32'd11,32'd11,32'd9,32'd2,32'd3,32'd9,32'd8,32'd5,32'd4,32'd10,32'd3,32'd10,32'd3,32'd7,32'd3,32'd10,32'd9,32'd7,32'd10,32'd1,32'd9,32'd6,32'd0,32'd1,32'd10,32'd6,32'd12,32'd0,32'd13,32'd0,32'd8,32'd4,32'd16,32'd0,32'd14,32'd5,32'd14,32'd5,32'd12,32'd11,32'd6,32'd11,32'd11,32'd0,32'd4,32'd9,32'd7,32'd9,32'd5,32'd10,32'd12,32'd5,32'd2,32'd3,32'd12,32'd0,32'd18,32'd9,32'd9,32'd0,32'd2,32'd0,32'd15,32'd9,32'd11,32'd11,32'd10,32'd10,32'd1,32'd11,32'd17,32'd5,32'd6,32'd4,32'd11,32'd9,32'd5,32'd8,32'd3,32'd1,32'd12,32'd1,32'd19,32'd0,32'd15,32'd7,32'd20,32'd3,32'd13,32'd9,32'd7,32'd5,32'd16,32'd8,32'd11,32'd10,32'd13,32'd0,32'd18,32'd3,32'd18,32'd8,32'd14,32'd12,32'd9,32'd11,32'd9,32'd9,32'd9,32'd9,32'd14,32'd6,32'd4,32'd10,32'd13,32'd9,32'd1,32'd8,32'd4,32'd2,32'd14,32'd4,32'd11,32'd8,32'd10,32'd4,32'd11,32'd5,32'd0,32'd0,32'd13,32'd8,32'd20,32'd3,32'd15,32'd0,32'd15,32'd0,32'd17,32'd4,32'd15,32'd2,32'd9,32'd0,32'd15,32'd2,32'd9,32'd1,32'd13,32'd8,32'd14,32'd7,32'd9,32'd0,32'd12,32'd12,32'd12,32'd10,32'd12,32'd10,32'd12,32'd2,32'd17,32'd5,32'd13,32'd3,32'd3,32'd2,32'd12,32'd8,32'd20,32'd4,32'd13,32'd2,32'd15,32'd3,32'd11,32'd0,32'd9,32'd7,32'd7,32'd13,32'd10,32'd14,32'd10,32'd12,32'd12,32'd12,32'd3,32'd12,32'd1,32'd19,32'd0,32'd17,32'd9,32'd7,32'd10,32'd12,32'd2,32'd0,32'd0,32'd8,32'd2,32'd11,32'd12,32'd8,32'd6,32'd4,32'd3,32'd15,32'd10,32'd12,32'd7,32'd12,32'd7,32'd9,32'd7,32'd12,32'd0,32'd18,32'd2,32'd1,32'd1,32'd6,32'd4,32'd18,32'd1,32'd6,32'd0,32'd14,32'd8,32'd0,32'd4,32'd10,32'd5,32'd15,32'd1,32'd19,32'd10,32'd19,32'd4,32'd3,32'd2,32'd14,32'd3,32'd17,32'd4,32'd7,32'd8,32'd13,32'd9,32'd13,32'd6,32'd14,32'd0,32'd19,32'd8,32'd12,32'd12,32'd15,32'd1,32'd10,32'd4,32'd16,32'd5,32'd14,32'd12,32'd12,32'd9,32'd17,32'd1,32'd20,32'd10,32'd11,32'd10,32'd14,32'd7,32'd10,32'd12,32'd13,32'd1,32'd2,32'd11,32'd13,32'd8,32'd10,32'd10,32'd0,32'd2,32'd9,32'd0,32'd12,32'd0,32'd3,32'd5,32'd8,32'd8,32'd17,32'd4,32'd14,32'd6,32'd5,32'd0,32'd18,32'd1,32'd3,32'd1,32'd14,32'd3,32'd14,32'd10,32'd14,32'd2,32'd12,32'd12,32'd12,32'd7,32'd15,32'd11,32'd5,32'd4,32'd18,32'd3,32'd18,32'd8,32'd10,32'd7,32'd9,32'd6,32'd2,32'd4,32'd17,32'd6,32'd7,32'd8,32'd1,32'd2,32'd7,32'd12,32'd8,32'd14,32'd9,32'd11,32'd10,32'd5,32'd12,32'd7,32'd11,32'd10,32'd5,32'd14,32'd2,32'd3,32'd0,32'd18,32'd1,32'd17,32'd0,32'd19,32'd6,32'd8,32'd4,32'd14,32'd10,32'd12,32'd6,32'd9,32'd1,32'd19,32'd1,32'd9,32'd8,32'd12,32'd6,32'd3,32'd5,32'd9,32'd5,32'd13,32'd2,32'd11,32'd0,32'd12,32'd10,32'd13,32'd7,32'd13,32'd2,32'd18,32'd3,32'd4,32'd9,32'd4,32'd11,32'd7,32'd6,32'd3,32'd2,32'd20,32'd1,32'd22,32'd8,32'd15,32'd0,32'd17,32'd1,32'd18,32'd3,32'd16,32'd4,32'd17,32'd3,32'd8,32'd0,32'd19,32'd5,32'd4,32'd0,32'd11,32'd10,32'd14,32'd3,32'd16,32'd5,32'd17,32'd4,32'd13,32'd1,32'd14,32'd0,32'd6,32'd0,32'd13,32'd0,32'd14,32'd0,32'd20,32'd1,32'd12,32'd12,32'd14,32'd7,32'd13,32'd11,32'd12,32'd10,32'd13,32'd8,32'd13,32'd8,32'd13,32'd0,32'd5,32'd0,32'd15,32'd0,32'd15,32'd5,32'd17,32'd9,32'd12,32'd2,32'd0,32'd0,32'd17,32'd0,32'd18,32'd1,32'd2,32'd0,32'd13,32'd2,32'd20,32'd0,32'd15,32'd6,32'd10,32'd0,32'd3,32'd9,32'd13,32'd7,32'd15,32'd1,32'd7,32'd8,32'd4,32'd8,32'd11,32'd6,32'd9,32'd9,32'd8,32'd4,32'd10,32'd10,32'd0,32'd0,32'd0,32'd16,32'd3,32'd12,32'd11,32'd10,32'd7,32'd16,32'd0,32'd7,32'd12,32'd8,32'd10,32'd7,32'd3,32'd14,32'd0,32'd15,32'd0,32'd15,32'd4,32'd15,32'd3,32'd15,32'd4,32'd12,32'd8,32'd12,32'd9,32'd12,32'd1,32'd16,32'd0,32'd18,32'd0,32'd12,32'd7,32'd8,32'd10,32'd4,32'd11,32'd9,32'd12,32'd8,32'd8,32'd14,32'd2,32'd20,32'd2,32'd6,32'd8,32'd13,32'd9,32'd6,32'd12,32'd9,32'd5,32'd13,32'd0,32'd18,32'd5,32'd12,32'd5,32'd13,32'd0,32'd2,32'd0,32'd3,32'd3,32'd17,32'd8,32'd15,32'd11,32'd11,32'd3,32'd16,32'd3,32'd14,32'd0,32'd9,32'd1,32'd18,32'd6,32'd16,32'd9,32'd16,32'd1,32'd5,32'd1,32'd5,32'd2,32'd13,32'd0,32'd15,32'd9,32'd16,32'd3,32'd10,32'd9,32'd15,32'd1,32'd13,32'd6,32'd18,32'd5,32'd14,32'd10,32'd12,32'd12,32'd11,32'd12,32'd16,32'd9,32'd8,32'd2,32'd20,32'd3,32'd8,32'd4,32'd14,32'd8,32'd14,32'd4,32'd14,32'd1,32'd19,32'd2,32'd3,32'd8,32'd15,32'd11,32'd6,32'd6,32'd2,32'd0,32'd7,32'd2,32'd4,32'd5,32'd2,32'd9,32'd12,32'd5,32'd12,32'd0,32'd12,32'd2,32'd17,32'd9,32'd11,32'd5,32'd13,32'd3,32'd12,32'd3,32'd12,32'd12,32'd7,32'd3,32'd11,32'd1,32'd16,32'd9,32'd12,32'd4,32'd8,32'd8,32'd17,32'd6,32'd11,32'd8,32'd9,32'd5,32'd14,32'd6,32'd5,32'd0,32'd12,32'd1,32'd12,32'd2,32'd12,32'd0,32'd12,32'd7,32'd10,32'd10,32'd5,32'd9,32'd11,32'd11,32'd5,32'd8,32'd10,32'd0,32'd14,32'd5,32'd12,32'd2,32'd3,32'd11,32'd12,32'd11,32'd11,32'd7,32'd10,32'd12,32'd16,32'd3,32'd16,32'd3,32'd15,32'd10,32'd12,32'd11,32'd7,32'd12,32'd16,32'd0,32'd9,32'd1,32'd15,32'd0,32'd14,32'd1,32'd20,32'd2,32'd2,32'd1,32'd12,32'd0,32'd13,32'd5,32'd14,32'd7,32'd11,32'd1,32'd10,32'd9,32'd6,32'd9,32'd5,32'd8,32'd13,32'd3,32'd18,32'd2,32'd20,32'd0,32'd6,32'd0,32'd12,32'd10,32'd20,32'd0,32'd6,32'd8,32'd4,32'd5,32'd8,32'd0,32'd20,32'd8,32'd20,32'd3,32'd11,32'd8,32'd1,32'd7,32'd2,32'd17,32'd7,32'd9,32'd1,32'd11,32'd6,32'd14,32'd12,32'd6,32'd1,32'd18,32'd2,32'd12,32'd7,32'd14,32'd10,32'd12,32'd9,32'd20,32'd0,32'd12,32'd5,32'd14,32'd11,32'd12,32'd5,32'd13,32'd4,32'd6,32'd0,32'd9,32'd8,32'd5,32'd3,32'd8,32'd1,32'd9,32'd9,32'd13,32'd2,32'd4,32'd9,32'd13,32'd11,32'd12,32'd9,32'd18,32'd9,32'd10,32'd5,32'd7,32'd2,32'd3,32'd0,32'd0,32'd10,32'd6,32'd4,32'd5,32'd3,32'd12,32'd4,32'd12,32'd11,32'd8,32'd10,32'd1,32'd5,32'd2,32'd0,32'd5,32'd3,32'd19,32'd5,32'd13,32'd9,32'd9,32'd5,32'd5,32'd5,32'd16,32'd0,32'd16,32'd6,32'd12,32'd7,32'd14,32'd7,32'd13,32'd4,32'd15,32'd0,32'd10,32'd11,32'd18,32'd7,32'd11,32'd6,32'd13,32'd2,32'd10,32'd5,32'd18,32'd0,32'd12,32'd6,32'd12,32'd9,32'd5,32'd2,32'd14,32'd2,32'd14,32'd10,32'd4,32'd8,32'd12,32'd0,32'd14,32'd0,32'd12,32'd2,32'd20,32'd2,32'd10,32'd0,32'd11,32'd3,32'd8,32'd2,32'd11,32'd7,32'd9,32'd4,32'd7,32'd14,32'd9,32'd14,32'd7,32'd11,32'd2,32'd8,32'd1,32'd6,32'd1,32'd12,32'd9,32'd11,32'd1,32'd9,32'd8,32'd14,32'd3,32'd11,32'd7,32'd12,32'd12,32'd15,32'd8,32'd5,32'd11,32'd4,32'd10,32'd9,32'd8,32'd12,32'd11,32'd11,32'd0,32'd12,32'd11,32'd18,32'd6,32'd15,32'd1,32'd13,32'd8,32'd12,32'd8,32'd12,32'd10,32'd6,32'd0,32'd15,32'd1,32'd12,32'd2,32'd12,32'd8,32'd13,32'd0,32'd15,32'd0,32'd17,32'd0,32'd12,32'd7,32'd10,32'd5,32'd16,32'd5,32'd13,32'd1,32'd15,32'd4,32'd12,32'd4,32'd13,32'd1,32'd1,32'd0,32'd11,32'd9,32'd18,32'd0,32'd20,32'd0,32'd19,32'd1,32'd12,32'd5,32'd13,32'd8,32'd9,32'd0,32'd4,32'd11,32'd12,32'd10,32'd12,32'd2,32'd3,32'd10,32'd3,32'd3,32'd14,32'd1,32'd10,32'd2,32'd16,32'd0,32'd15,32'd3,32'd20,32'd2,32'd16,32'd2,32'd15,32'd9,32'd20,32'd8,32'd19,32'd1,32'd8,32'd5,32'd15,32'd0,32'd12,32'd5,32'd10,32'd2,32'd4,32'd10,32'd6,32'd17,32'd3,32'd14,32'd2,32'd4,32'd8,32'd10,32'd0,32'd13,32'd0,32'd20,32'd3,32'd19,32'd0,32'd1,32'd2,32'd22,32'd3,32'd18,32'd2,32'd12,32'd3,32'd11,32'd1,32'd13,32'd12,32'd2,32'd2,32'd18,32'd0,32'd2,32'd8,32'd18,32'd9,32'd9,32'd1,32'd8,32'd9,32'd11,32'd11,32'd12,32'd4,32'd17,32'd8,32'd13,32'd6,32'd13,32'd8,32'd14,32'd0,32'd15,32'd10,32'd17,32'd7,32'd5,32'd0,32'd15,32'd6,32'd15,32'd5,32'd15,32'd9,32'd13,32'd12,32'd13,32'd1,32'd14,32'd7,32'd6,32'd3,32'd1,32'd1,32'd5,32'd1,32'd3,32'd8,32'd5,32'd5,32'd3,32'd5,32'd8,32'd7,32'd12,32'd6,32'd14,32'd10,32'd10,32'd5,32'd13,32'd0,32'd11,32'd6,32'd16,32'd6,32'd7,32'd8,32'd13,32'd4,32'd13,32'd8,32'd13,32'd3,32'd9,32'd3,32'd18,32'd3,32'd11,32'd5,32'd10,32'd3,32'd8,32'd7,32'd2,32'd17,32'd1,32'd12,32'd3,32'd3,32'd0,32'd12,32'd6,32'd11,32'd3,32'd15,32'd8,32'd14,32'd11,32'd14,32'd0,32'd15,32'd0,32'd10,32'd10,32'd5,32'd6,32'd8,32'd5,32'd17,32'd0,32'd15,32'd6,32'd4,32'd3,32'd19,32'd3,32'd19,32'd3,32'd15,32'd2,32'd8,32'd3,32'd6,32'd0,32'd13,32'd9,32'd13,32'd8,32'd10,32'd0,32'd20,32'd3,32'd20,32'd8,32'd13,32'd12,32'd12,32'd3,32'd3,32'd6,32'd14,32'd6,32'd14,32'd9,32'd13,32'd0,32'd15,32'd12,32'd22,32'd7,32'd11,32'd8,32'd22,32'd5,32'd18,32'd5,32'd14,32'd2,32'd12,32'd0,32'd18,32'd9,32'd3,32'd2,32'd19,32'd0,32'd15,32'd1,32'd14,32'd9,32'd14,32'd0,32'd10,32'd8,32'd10,32'd2,32'd3,32'd9,32'd1,32'd8,32'd10,32'd6,32'd8,32'd10,32'd5,32'd9,32'd6,32'd16,32'd10,32'd12,32'd11,32'd6,32'd6,32'd14,32'd10,32'd14,32'd12,32'd17,32'd2,32'd18,32'd2,32'd14,32'd5,32'd8,32'd6,32'd19,32'd7,32'd15,32'd1,32'd12,32'd9,32'd15,32'd0,32'd6,32'd3,32'd13,32'd0,32'd12,32'd0,32'd19,32'd0,32'd14,32'd6,32'd2,32'd3,32'd12,32'd12,32'd12,32'd4,32'd6,32'd10,32'd8,32'd0,32'd5,32'd5,32'd10,32'd1,32'd6,32'd8,32'd14,32'd9,32'd9,32'd8,32'd14,32'd1,32'd17,32'd0,32'd9,32'd0,32'd18,32'd7,32'd18,32'd6,32'd20,32'd8,32'd14,32'd9,32'd13,32'd10,32'd9,32'd8,32'd12,32'd6,32'd13,32'd5,32'd20,32'd3,32'd3,32'd3,32'd11,32'd5,32'd14,32'd8,32'd10,32'd6,32'd12,32'd11,32'd11,32'd12,32'd6,32'd16,32'd4,32'd5,32'd7,32'd14,32'd0,32'd16,32'd8,32'd12,32'd9,32'd13,32'd0,32'd6,32'd1,32'd6,32'd7,32'd15,32'd8,32'd12,32'd4,32'd12,32'd7,32'd16,32'd1,32'd20,32'd6,32'd14,32'd2,32'd4,32'd0,32'd15,32'd3,32'd18,32'd5,32'd17,32'd0,32'd14,32'd1,32'd12,32'd1,32'd14,32'd1,32'd18,32'd9,32'd13,32'd9,32'd15,32'd8,32'd11,32'd5,32'd15,32'd3,32'd15,32'd10,32'd12,32'd6,32'd5,32'd0,32'd18,32'd3,32'd18,32'd0,32'd21,32'd9,32'd16,32'd10,32'd3,32'd2,32'd9,32'd7,32'd11,32'd4,32'd5,32'd10,32'd6,32'd8,32'd12,32'd3,32'd10,32'd1,32'd15,32'd1,32'd12,32'd8,32'd9,32'd10,32'd13,32'd11,32'd5,32'd2,32'd14,32'd7,32'd9,32'd8,32'd15,32'd8,32'd14,32'd9,32'd13,32'd10,32'd8,32'd0,32'd18,32'd0,32'd9,32'd4,32'd0,32'd2,32'd16,32'd6,32'd12,32'd12,32'd9,32'd8,32'd9,32'd0,32'd8,32'd0,32'd15,32'd8,32'd15,32'd0,32'd15,32'd0,32'd7,32'd8,32'd7,32'd9,32'd6,32'd9,32'd12,32'd10,32'd13,32'd1,32'd14,32'd6,32'd12,32'd3,32'd15,32'd8,32'd10,32'd4,32'd7,32'd3,32'd17,32'd11,32'd15,32'd3,32'd14,32'd1,32'd20,32'd10,32'd9,32'd11,32'd8,32'd4,32'd12,32'd0,32'd10,32'd8,32'd10,32'd10,32'd13,32'd4,32'd12,32'd0,32'd3,32'd9,32'd12,32'd5,32'd7,32'd4,32'd14,32'd5,32'd12,32'd2,32'd13,32'd10,32'd13,32'd9,32'd13,32'd0,32'd13,32'd1,32'd18,32'd3,32'd18,32'd6,32'd11,32'd10,32'd11,32'd0,32'd13,32'd2,32'd1,32'd0,32'd13,32'd2,32'd5,32'd2,32'd5,32'd2,32'd20,32'd9,32'd5,32'd4,32'd10,32'd10,32'd6,32'd6,32'd0,32'd13,32'd3,32'd13,32'd6,32'd18,32'd9,32'd14,32'd9,32'd14,32'd12,32'd13,32'd0,32'd7,32'd9,32'd12,32'd9,32'd1,32'd0,32'd7,32'd8,32'd8,32'd8,32'd13,32'd1,32'd13,32'd12,32'd13,32'd7,32'd14,32'd10,32'd8,32'd7,32'd8,32'd3,32'd18,32'd5,32'd14,32'd2,32'd9,32'd2,32'd16,32'd3,32'd18,32'd3,32'd18,32'd9,32'd4,32'd0,32'd9,32'd10,32'd6,32'd8,32'd19,32'd4,32'd16,32'd5,32'd8,32'd12,32'd3,32'd8,32'd10,32'd3,32'd3,32'd6,32'd4,32'd4,32'd14,32'd5,32'd3,32'd2,32'd2,32'd9,32'd12,32'd0,32'd8,32'd8,32'd14,32'd0,32'd17,32'd8,32'd14,32'd4,32'd12,32'd2,32'd20,32'd5,32'd6,32'd1,32'd6,32'd0,32'd7,32'd6,32'd10,32'd1,32'd9,32'd11,32'd11,32'd9,32'd11,32'd8,32'd11,32'd4,32'd8,32'd6,32'd9,32'd10,32'd12,32'd9,32'd11,32'd9,32'd10,32'd5,32'd15,32'd1,32'd14,32'd3,32'd5,32'd1,32'd3,32'd2,32'd4,32'd1,32'd15,32'd8,32'd6,32'd3,32'd14,32'd1,32'd8,32'd3,32'd19,32'd2,32'd4,32'd8,32'd10,32'd6,32'd0,32'd17,32'd1,32'd12,32'd10,32'd12,32'd0,32'd12,32'd2,32'd20,32'd11,32'd20,32'd2,32'd2,32'd10,32'd2,32'd5,32'd8,32'd4,32'd18,32'd5,32'd9,32'd6,32'd11,32'd9,32'd5,32'd8,32'd5,32'd7,32'd11,32'd8,32'd20,32'd4,32'd12,32'd9,32'd16,32'd5,32'd5,32'd9,32'd8,32'd1,32'd10,32'd6,32'd4,32'd11,32'd5,32'd6,32'd5,32'd8,32'd3,32'd10,32'd6}
`define RECTANGLE2_YS {32'd1,32'd17,32'd2,32'd19,32'd19,32'd19,32'd19,32'd14,32'd16,32'd19,32'd19,32'd6,32'd19,32'd12,32'd12,32'd20,32'd16,32'd18,32'd14,32'd13,32'd13,32'd13,32'd13,32'd8,32'd15,32'd15,32'd15,32'd13,32'd13,32'd13,32'd13,32'd8,32'd8,32'd0,32'd20,32'd1,32'd1,32'd0,32'd14,32'd13,32'd9,32'd11,32'd1,32'd0,32'd0,32'd9,32'd9,32'd2,32'd13,32'd1,32'd2,32'd14,32'd14,32'd5,32'd6,32'd6,32'd8,32'd8,32'd5,32'd11,32'd17,32'd20,32'd19,32'd17,32'd18,32'd17,32'd4,32'd8,32'd8,32'd9,32'd7,32'd7,32'd7,32'd5,32'd9,32'd16,32'd4,32'd3,32'd4,32'd0,32'd6,32'd5,32'd0,32'd1,32'd9,32'd10,32'd9,32'd13,32'd12,32'd2,32'd2,32'd13,32'd13,32'd10,32'd13,32'd10,32'd10,32'd14,32'd12,32'd13,32'd12,32'd3,32'd3,32'd0,32'd6,32'd6,32'd15,32'd12,32'd12,32'd15,32'd12,32'd8,32'd8,32'd4,32'd5,32'd11,32'd12,32'd14,32'd14,32'd4,32'd4,32'd3,32'd12,32'd2,32'd5,32'd6,32'd5,32'd19,32'd19,32'd16,32'd16,32'd16,32'd16,32'd0,32'd0,32'd16,32'd16,32'd20,32'd18,32'd21,32'd22,32'd6,32'd6,32'd6,32'd0,32'd2,32'd8,32'd7,32'd7,32'd11,32'd11,32'd11,32'd7,32'd9,32'd4,32'd6,32'd9,32'd11,32'd17,32'd17,32'd12,32'd11,32'd11,32'd7,32'd7,32'd4,32'd3,32'd5,32'd5,32'd3,32'd3,32'd0,32'd1,32'd8,32'd12,32'd15,32'd19,32'd13,32'd2,32'd6,32'd11,32'd20,32'd16,32'd13,32'd6,32'd14,32'd14,32'd6,32'd6,32'd2,32'd4,32'd9,32'd12,32'd16,32'd18,32'd14,32'd16,32'd1,32'd5,32'd7,32'd7,32'd1,32'd2,32'd16,32'd15,32'd5,32'd4,32'd7,32'd0,32'd6,32'd2,32'd2,32'd0,32'd0,32'd0,32'd0,32'd8,32'd8,32'd4,32'd9,32'd2,32'd8,32'd8,32'd7,32'd8,32'd9,32'd19,32'd19,32'd0,32'd0,32'd0,32'd7,32'd7,32'd7,32'd0,32'd0,32'd1,32'd11,32'd7,32'd19,32'd6,32'd6,32'd3,32'd2,32'd17,32'd2,32'd8,32'd6,32'd3,32'd6,32'd6,32'd20,32'd8,32'd8,32'd3,32'd2,32'd1,32'd2,32'd2,32'd9,32'd10,32'd10,32'd13,32'd13,32'd2,32'd10,32'd8,32'd8,32'd7,32'd6,32'd6,32'd6,32'd13,32'd0,32'd19,32'd6,32'd1,32'd9,32'd15,32'd7,32'd14,32'd10,32'd12,32'd12,32'd16,32'd19,32'd14,32'd15,32'd13,32'd13,32'd4,32'd10,32'd1,32'd1,32'd4,32'd12,32'd6,32'd10,32'd15,32'd0,32'd1,32'd7,32'd8,32'd8,32'd9,32'd14,32'd4,32'd0,32'd0,32'd0,32'd4,32'd18,32'd18,32'd6,32'd7,32'd7,32'd16,32'd4,32'd0,32'd19,32'd12,32'd8,32'd9,32'd5,32'd6,32'd8,32'd12,32'd1,32'd0,32'd0,32'd14,32'd14,32'd6,32'd7,32'd11,32'd0,32'd0,32'd6,32'd0,32'd7,32'd9,32'd0,32'd16,32'd2,32'd3,32'd19,32'd13,32'd9,32'd17,32'd13,32'd0,32'd0,32'd7,32'd7,32'd6,32'd0,32'd1,32'd11,32'd2,32'd6,32'd1,32'd1,32'd2,32'd1,32'd15,32'd15,32'd15,32'd15,32'd4,32'd4,32'd9,32'd0,32'd3,32'd9,32'd6,32'd3,32'd1,32'd1,32'd20,32'd20,32'd6,32'd7,32'd8,32'd20,32'd17,32'd8,32'd2,32'd15,32'd20,32'd17,32'd17,32'd15,32'd18,32'd18,32'd5,32'd11,32'd11,32'd11,32'd1,32'd9,32'd14,32'd7,32'd0,32'd12,32'd0,32'd1,32'd20,32'd14,32'd1,32'd6,32'd3,32'd0,32'd4,32'd9,32'd6,32'd6,32'd9,32'd22,32'd1,32'd0,32'd0,32'd1,32'd15,32'd10,32'd10,32'd15,32'd15,32'd6,32'd17,32'd7,32'd7,32'd11,32'd0,32'd5,32'd1,32'd4,32'd7,32'd8,32'd17,32'd4,32'd17,32'd3,32'd17,32'd14,32'd17,32'd15,32'd12,32'd7,32'd7,32'd9,32'd9,32'd10,32'd0,32'd17,32'd17,32'd13,32'd13,32'd1,32'd13,32'd13,32'd13,32'd5,32'd10,32'd8,32'd4,32'd4,32'd5,32'd10,32'd14,32'd14,32'd12,32'd5,32'd10,32'd8,32'd9,32'd6,32'd6,32'd11,32'd11,32'd8,32'd10,32'd1,32'd16,32'd1,32'd1,32'd18,32'd19,32'd12,32'd11,32'd17,32'd4,32'd22,32'd20,32'd14,32'd9,32'd11,32'd8,32'd8,32'd8,32'd12,32'd2,32'd5,32'd7,32'd0,32'd0,32'd1,32'd8,32'd6,32'd9,32'd2,32'd5,32'd0,32'd0,32'd17,32'd15,32'd20,32'd8,32'd6,32'd2,32'd4,32'd13,32'd5,32'd2,32'd7,32'd7,32'd12,32'd6,32'd10,32'd10,32'd1,32'd1,32'd10,32'd19,32'd10,32'd1,32'd11,32'd0,32'd13,32'd2,32'd2,32'd11,32'd19,32'd7,32'd4,32'd4,32'd13,32'd13,32'd16,32'd5,32'd6,32'd5,32'd12,32'd12,32'd0,32'd0,32'd1,32'd0,32'd9,32'd4,32'd9,32'd9,32'd9,32'd6,32'd20,32'd0,32'd2,32'd2,32'd17,32'd17,32'd20,32'd20,32'd20,32'd17,32'd9,32'd9,32'd6,32'd8,32'd17,32'd9,32'd10,32'd14,32'd19,32'd17,32'd18,32'd18,32'd6,32'd10,32'd12,32'd18,32'd1,32'd13,32'd11,32'd9,32'd5,32'd9,32'd17,32'd2,32'd8,32'd8,32'd22,32'd6,32'd12,32'd16,32'd0,32'd0,32'd6,32'd3,32'd10,32'd1,32'd11,32'd12,32'd2,32'd15,32'd3,32'd4,32'd19,32'd20,32'd20,32'd15,32'd15,32'd12,32'd12,32'd10,32'd10,32'd6,32'd16,32'd12,32'd3,32'd11,32'd8,32'd8,32'd0,32'd6,32'd12,32'd12,32'd16,32'd0,32'd2,32'd14,32'd9,32'd8,32'd11,32'd10,32'd10,32'd8,32'd10,32'd20,32'd5,32'd11,32'd9,32'd9,32'd10,32'd0,32'd15,32'd15,32'd14,32'd16,32'd16,32'd16,32'd18,32'd10,32'd14,32'd14,32'd10,32'd1,32'd1,32'd0,32'd10,32'd0,32'd8,32'd7,32'd9,32'd0,32'd0,32'd4,32'd0,32'd2,32'd2,32'd6,32'd5,32'd0,32'd0,32'd4,32'd0,32'd5,32'd5,32'd1,32'd1,32'd17,32'd17,32'd18,32'd19,32'd19,32'd4,32'd11,32'd18,32'd19,32'd10,32'd3,32'd11,32'd11,32'd8,32'd6,32'd8,32'd8,32'd8,32'd8,32'd8,32'd5,32'd18,32'd11,32'd16,32'd17,32'd4,32'd8,32'd4,32'd21,32'd21,32'd14,32'd14,32'd9,32'd7,32'd3,32'd0,32'd17,32'd17,32'd0,32'd4,32'd2,32'd7,32'd4,32'd0,32'd2,32'd11,32'd10,32'd5,32'd6,32'd8,32'd8,32'd16,32'd9,32'd5,32'd6,32'd3,32'd6,32'd18,32'd14,32'd14,32'd12,32'd6,32'd8,32'd1,32'd12,32'd18,32'd15,32'd2,32'd2,32'd2,32'd2,32'd4,32'd4,32'd2,32'd6,32'd20,32'd7,32'd7,32'd1,32'd6,32'd0,32'd0,32'd6,32'd6,32'd3,32'd14,32'd2,32'd2,32'd1,32'd1,32'd3,32'd12,32'd14,32'd19,32'd15,32'd15,32'd15,32'd23,32'd18,32'd6,32'd11,32'd1,32'd3,32'd7,32'd7,32'd14,32'd14,32'd8,32'd8,32'd12,32'd12,32'd12,32'd12,32'd20,32'd4,32'd19,32'd19,32'd16,32'd1,32'd1,32'd8,32'd6,32'd2,32'd9,32'd11,32'd16,32'd14,32'd3,32'd5,32'd0,32'd16,32'd4,32'd9,32'd1,32'd1,32'd6,32'd5,32'd11,32'd7,32'd16,32'd0,32'd4,32'd4,32'd4,32'd4,32'd16,32'd9,32'd1,32'd1,32'd0,32'd1,32'd16,32'd1,32'd21,32'd1,32'd14,32'd14,32'd6,32'd2,32'd10,32'd10,32'd12,32'd19,32'd10,32'd17,32'd18,32'd18,32'd19,32'd19,32'd18,32'd4,32'd3,32'd3,32'd0,32'd0,32'd5,32'd5,32'd0,32'd0,32'd8,32'd7,32'd10,32'd7,32'd1,32'd1,32'd12,32'd10,32'd14,32'd1,32'd0,32'd0,32'd6,32'd14,32'd19,32'd8,32'd10,32'd7,32'd7,32'd14,32'd13,32'd3,32'd6,32'd1,32'd8,32'd5,32'd0,32'd19,32'd10,32'd3,32'd16,32'd22,32'd7,32'd2,32'd2,32'd3,32'd3,32'd17,32'd1,32'd1,32'd0,32'd4,32'd6,32'd7,32'd4,32'd4,32'd5,32'd5,32'd8,32'd10,32'd10,32'd2,32'd19,32'd9,32'd4,32'd2,32'd19,32'd20,32'd21,32'd21,32'd18,32'd5,32'd16,32'd16,32'd17,32'd17,32'd15,32'd9,32'd11,32'd11,32'd15,32'd18,32'd18,32'd11,32'd11,32'd1,32'd5,32'd1,32'd5,32'd6,32'd0,32'd8,32'd1,32'd16,32'd20,32'd17,32'd18,32'd1,32'd13,32'd1,32'd5,32'd5,32'd0,32'd0,32'd6,32'd6,32'd5,32'd18,32'd19,32'd6,32'd8,32'd8,32'd15,32'd16,32'd1,32'd7,32'd2,32'd2,32'd0,32'd0,32'd18,32'd11,32'd20,32'd4,32'd10,32'd0,32'd16,32'd12,32'd5,32'd7,32'd1,32'd10,32'd15,32'd10,32'd12,32'd12,32'd12,32'd12,32'd12,32'd9,32'd10,32'd10,32'd8,32'd17,32'd17,32'd12,32'd12,32'd14,32'd14,32'd8,32'd9,32'd8,32'd13,32'd2,32'd13,32'd13,32'd3,32'd4,32'd0,32'd0,32'd0,32'd7,32'd4,32'd5,32'd9,32'd9,32'd0,32'd9,32'd6,32'd13,32'd15,32'd8,32'd3,32'd4,32'd12,32'd3,32'd0,32'd19,32'd20,32'd20,32'd6,32'd2,32'd3,32'd0,32'd1,32'd14,32'd15,32'd0,32'd6,32'd11,32'd0,32'd8,32'd7,32'd10,32'd16,32'd10,32'd11,32'd11,32'd10,32'd0,32'd1,32'd1,32'd8,32'd8,32'd0,32'd0,32'd2,32'd2,32'd0,32'd0,32'd12,32'd0,32'd3,32'd9,32'd10,32'd10,32'd13,32'd6,32'd6,32'd17,32'd10,32'd14,32'd12,32'd0,32'd8,32'd5,32'd10,32'd4,32'd7,32'd5,32'd9,32'd6,32'd7,32'd6,32'd18,32'd18,32'd15,32'd8,32'd18,32'd19,32'd20,32'd18,32'd0,32'd8,32'd1,32'd6,32'd3,32'd7,32'd2,32'd2,32'd2,32'd4,32'd8,32'd3,32'd3,32'd6,32'd15,32'd15,32'd22,32'd15,32'd19,32'd19,32'd0,32'd5,32'd2,32'd3,32'd4,32'd7,32'd3,32'd9,32'd12,32'd12,32'd0,32'd17,32'd3,32'd0,32'd18,32'd16,32'd16,32'd16,32'd4,32'd4,32'd17,32'd19,32'd0,32'd0,32'd6,32'd6,32'd7,32'd15,32'd10,32'd6,32'd0,32'd20,32'd16,32'd2,32'd6,32'd10,32'd22,32'd16,32'd6,32'd16,32'd2,32'd8,32'd10,32'd15,32'd10,32'd5,32'd3,32'd16,32'd1,32'd1,32'd0,32'd0,32'd18,32'd0,32'd0,32'd6,32'd6,32'd1,32'd0,32'd21,32'd14,32'd11,32'd0,32'd0,32'd3,32'd0,32'd12,32'd7,32'd15,32'd1,32'd12,32'd12,32'd19,32'd18,32'd11,32'd15,32'd2,32'd2,32'd18,32'd20,32'd9,32'd13,32'd13,32'd18,32'd20,32'd18,32'd6,32'd7,32'd13,32'd13,32'd13,32'd6,32'd0,32'd4,32'd18,32'd10,32'd15,32'd12,32'd2,32'd2,32'd4,32'd0,32'd19,32'd14,32'd14,32'd3,32'd7,32'd2,32'd1,32'd0,32'd0,32'd7,32'd11,32'd4,32'd9,32'd8,32'd4,32'd2,32'd2,32'd7,32'd11,32'd9,32'd10,32'd15,32'd18,32'd1,32'd1,32'd3,32'd7,32'd7,32'd11,32'd3,32'd22,32'd13,32'd7,32'd0,32'd13,32'd15,32'd0,32'd2,32'd0,32'd10,32'd5,32'd21,32'd21,32'd6,32'd4,32'd9,32'd9,32'd7,32'd13,32'd5,32'd5,32'd6,32'd5,32'd1,32'd1,32'd0,32'd7,32'd1,32'd21,32'd13,32'd2,32'd0,32'd0,32'd10,32'd23,32'd1,32'd3,32'd0,32'd10,32'd10,32'd12,32'd8,32'd9,32'd9,32'd9,32'd8,32'd7,32'd5,32'd9,32'd2,32'd17,32'd13,32'd18,32'd14,32'd13,32'd18,32'd18,32'd19,32'd19,32'd6,32'd5,32'd2,32'd19,32'd18,32'd17,32'd8,32'd19,32'd17,32'd9,32'd6,32'd11,32'd0,32'd0,32'd8,32'd16,32'd3,32'd2,32'd1,32'd3,32'd3,32'd3,32'd6,32'd2,32'd3,32'd5,32'd6,32'd9,32'd19,32'd7,32'd4,32'd1,32'd13,32'd4,32'd11,32'd4,32'd8,32'd18,32'd3,32'd6,32'd11,32'd0,32'd7,32'd5,32'd5,32'd4,32'd5,32'd1,32'd1,32'd4,32'd4,32'd4,32'd4,32'd4,32'd1,32'd5,32'd5,32'd19,32'd5,32'd7,32'd5,32'd12,32'd13,32'd2,32'd18,32'd12,32'd11,32'd7,32'd4,32'd9,32'd6,32'd8,32'd11,32'd15,32'd15,32'd4,32'd15,32'd13,32'd14,32'd15,32'd15,32'd8,32'd8,32'd11,32'd11,32'd11,32'd22,32'd3,32'd8,32'd2,32'd3,32'd2,32'd2,32'd2,32'd18,32'd16,32'd17,32'd8,32'd8,32'd4,32'd4,32'd2,32'd4,32'd14,32'd10,32'd5,32'd1,32'd10,32'd10,32'd8,32'd10,32'd9,32'd9,32'd6,32'd6,32'd16,32'd12,32'd16,32'd16,32'd10,32'd0,32'd1,32'd2,32'd19,32'd14,32'd6,32'd6,32'd3,32'd3,32'd20,32'd17,32'd4,32'd0,32'd0,32'd0,32'd3,32'd10,32'd15,32'd3,32'd0,32'd1,32'd7,32'd2,32'd18,32'd2,32'd7,32'd0,32'd6,32'd13,32'd7,32'd7,32'd18,32'd10,32'd18,32'd16,32'd17,32'd18,32'd1,32'd20,32'd21,32'd1,32'd18,32'd18,32'd18,32'd14,32'd7,32'd7,32'd9,32'd8,32'd14,32'd14,32'd14,32'd18,32'd7,32'd18,32'd9,32'd0,32'd6,32'd11,32'd13,32'd13,32'd9,32'd19,32'd4,32'd4,32'd0,32'd4,32'd11,32'd5,32'd12,32'd20,32'd7,32'd3,32'd15,32'd0,32'd7,32'd10,32'd2,32'd4,32'd21,32'd12,32'd0,32'd12,32'd12,32'd11,32'd1,32'd4,32'd19,32'd6,32'd8,32'd11,32'd11,32'd3,32'd3,32'd5,32'd5,32'd5,32'd5,32'd6,32'd6,32'd12,32'd12,32'd7,32'd6,32'd9,32'd4,32'd8,32'd15,32'd9,32'd16,32'd9,32'd10,32'd15,32'd18,32'd16,32'd0,32'd5,32'd3,32'd19,32'd17,32'd13,32'd13,32'd12,32'd0,32'd7,32'd12,32'd7,32'd13,32'd7,32'd14,32'd14,32'd7,32'd7,32'd7,32'd12,32'd22,32'd18,32'd13,32'd14,32'd13,32'd11,32'd11,32'd1,32'd1,32'd1,32'd1,32'd2,32'd15,32'd12,32'd7,32'd10,32'd10,32'd8,32'd8,32'd1,32'd2,32'd0,32'd0,32'd9,32'd18,32'd18,32'd1,32'd0,32'd16,32'd16,32'd17,32'd12,32'd10,32'd10,32'd10,32'd7,32'd9,32'd12,32'd17,32'd16,32'd6,32'd6,32'd18,32'd9,32'd14,32'd9,32'd12,32'd5,32'd10,32'd8,32'd8,32'd7,32'd6,32'd5,32'd8,32'd0,32'd8,32'd7,32'd8,32'd16,32'd16,32'd17,32'd16,32'd18,32'd19,32'd0,32'd0,32'd0,32'd6,32'd2,32'd8,32'd10,32'd6,32'd3,32'd10,32'd11,32'd3,32'd1,32'd0,32'd2,32'd2,32'd0,32'd0,32'd5,32'd8,32'd10,32'd1,32'd7,32'd0,32'd0,32'd0,32'd4,32'd17,32'd10,32'd4,32'd6,32'd6,32'd11,32'd21,32'd14,32'd1,32'd7,32'd9,32'd19,32'd13,32'd3,32'd5,32'd5,32'd12,32'd2,32'd10,32'd7,32'd18,32'd1,32'd0,32'd9,32'd22,32'd6,32'd17,32'd8,32'd0,32'd0,32'd17,32'd17,32'd14,32'd14,32'd11,32'd14,32'd8,32'd8,32'd0,32'd6,32'd5,32'd5,32'd8,32'd8,32'd20,32'd18,32'd18,32'd8,32'd13,32'd4,32'd9,32'd17,32'd10,32'd15,32'd8,32'd7,32'd13,32'd2,32'd0,32'd0,32'd0,32'd0,32'd2,32'd5,32'd11,32'd11,32'd5,32'd7,32'd12,32'd1,32'd13,32'd4,32'd5,32'd5,32'd16,32'd6,32'd5,32'd19,32'd3,32'd8,32'd6,32'd19,32'd20,32'd6,32'd0,32'd0,32'd8,32'd11,32'd8,32'd6,32'd11,32'd2,32'd13,32'd0,32'd2,32'd5,32'd2,32'd2,32'd15,32'd2,32'd2,32'd1,32'd17,32'd17,32'd18,32'd18,32'd15,32'd15,32'd13,32'd6,32'd6,32'd8,32'd3,32'd15,32'd10,32'd13,32'd6,32'd8,32'd5,32'd16,32'd5,32'd6,32'd5,32'd5,32'd21,32'd15,32'd0,32'd18,32'd4,32'd0,32'd2,32'd2,32'd8,32'd8,32'd5,32'd5,32'd17,32'd17,32'd11,32'd0,32'd16,32'd23,32'd7,32'd11,32'd1,32'd7,32'd0,32'd11,32'd14,32'd3,32'd4,32'd5,32'd9,32'd11,32'd15,32'd1,32'd2,32'd4,32'd8,32'd0,32'd16,32'd16,32'd4,32'd5,32'd12,32'd1,32'd19,32'd19,32'd8,32'd15,32'd7,32'd8,32'd4,32'd7,32'd9,32'd9,32'd15,32'd19,32'd16,32'd7,32'd15,32'd10,32'd10,32'd8,32'd10,32'd13,32'd22,32'd16,32'd16,32'd2,32'd1,32'd19,32'd18,32'd19,32'd19,32'd19,32'd8,32'd5,32'd9,32'd11,32'd7,32'd2,32'd12,32'd12,32'd15,32'd6,32'd2,32'd15,32'd1,32'd1,32'd5,32'd13,32'd8,32'd8,32'd3,32'd3,32'd7,32'd7,32'd0,32'd5,32'd3,32'd0,32'd3,32'd1,32'd18,32'd18,32'd1,32'd1,32'd6,32'd6,32'd3,32'd17,32'd16,32'd13,32'd1,32'd17,32'd14,32'd6,32'd10,32'd10,32'd3,32'd3,32'd0,32'd1,32'd14,32'd14,32'd5,32'd0,32'd0,32'd12,32'd11,32'd10,32'd0,32'd8,32'd20,32'd12,32'd11,32'd11,32'd0,32'd0,32'd3,32'd3,32'd16,32'd18,32'd8,32'd11,32'd6,32'd3,32'd1,32'd4,32'd12,32'd2,32'd11,32'd17,32'd8,32'd8,32'd19,32'd8,32'd18,32'd6,32'd1,32'd9,32'd7,32'd16,32'd16,32'd0,32'd9,32'd5,32'd9,32'd4,32'd4,32'd12,32'd11,32'd11,32'd16,32'd12,32'd6,32'd12,32'd4,32'd0,32'd10,32'd18,32'd10,32'd10,32'd6,32'd5,32'd5,32'd0,32'd16,32'd8,32'd15,32'd16,32'd5,32'd11,32'd16,32'd14,32'd11,32'd11,32'd20,32'd14,32'd1,32'd0,32'd0,32'd12,32'd11,32'd14,32'd14,32'd9,32'd5,32'd7,32'd11,32'd6,32'd12,32'd13,32'd8,32'd5,32'd19,32'd19,32'd2,32'd6,32'd4,32'd5,32'd9,32'd6,32'd3,32'd12,32'd4,32'd7,32'd7,32'd4,32'd9,32'd5,32'd17,32'd5,32'd17,32'd1,32'd1,32'd0,32'd5,32'd0,32'd18,32'd6,32'd11,32'd14,32'd16,32'd7,32'd16,32'd11,32'd11,32'd6,32'd6,32'd0,32'd4,32'd10,32'd0,32'd13,32'd11,32'd14,32'd16,32'd8,32'd7,32'd11,32'd9,32'd3,32'd21,32'd12,32'd11,32'd0,32'd7,32'd6,32'd2,32'd7,32'd20,32'd12,32'd8,32'd16,32'd12,32'd14,32'd3,32'd13,32'd5,32'd16,32'd15,32'd18,32'd1,32'd2,32'd2,32'd3,32'd7,32'd18,32'd0,32'd1,32'd20,32'd3,32'd0,32'd8,32'd0,32'd11,32'd10,32'd9,32'd11,32'd10,32'd2,32'd7,32'd21,32'd4,32'd6,32'd18,32'd16,32'd6,32'd18,32'd19,32'd17,32'd20,32'd21,32'd12,32'd10,32'd11,32'd10,32'd10,32'd4,32'd0,32'd5,32'd2,32'd4,32'd13,32'd7,32'd10,32'd3,32'd0,32'd0,32'd6,32'd11,32'd11,32'd8,32'd8,32'd13,32'd11,32'd9,32'd9,32'd5,32'd12,32'd12,32'd6,32'd8,32'd18,32'd17,32'd17,32'd17,32'd0,32'd5,32'd3,32'd11,32'd11,32'd18,32'd18,32'd17,32'd10,32'd8,32'd19,32'd0,32'd4,32'd2,32'd11,32'd0,32'd10,32'd14,32'd16,32'd9,32'd10,32'd13,32'd19,32'd16,32'd3,32'd5,32'd13,32'd6,32'd5,32'd6,32'd6,32'd9,32'd9,32'd12,32'd0,32'd9,32'd16,32'd17,32'd13,32'd17,32'd17,32'd4,32'd5,32'd5,32'd5,32'd0,32'd9,32'd6,32'd7,32'd11,32'd8,32'd6,32'd7,32'd12,32'd12,32'd16,32'd17,32'd3,32'd0,32'd1,32'd10,32'd23,32'd11,32'd0,32'd0,32'd11,32'd3,32'd4,32'd20,32'd11,32'd11,32'd14,32'd11,32'd1,32'd3,32'd3,32'd12,32'd12,32'd5,32'd5,32'd6,32'd6,32'd5,32'd14,32'd14,32'd19,32'd3,32'd0,32'd7,32'd2,32'd3,32'd0,32'd2,32'd10,32'd19,32'd2,32'd8,32'd13,32'd7,32'd4,32'd5,32'd5,32'd21,32'd6,32'd9,32'd11,32'd14,32'd14,32'd5,32'd9,32'd11,32'd5,32'd2,32'd2,32'd20,32'd20,32'd4,32'd4,32'd4,32'd4,32'd2,32'd2,32'd10,32'd10,32'd4,32'd4,32'd5,32'd6,32'd10,32'd9,32'd8,32'd4,32'd10,32'd22,32'd6,32'd5,32'd8,32'd5,32'd11,32'd10,32'd0,32'd0,32'd6,32'd3,32'd20,32'd19,32'd2,32'd8,32'd8,32'd14,32'd15,32'd18,32'd17,32'd3,32'd11,32'd2,32'd0,32'd20,32'd5,32'd10,32'd12,32'd8,32'd6,32'd3,32'd2,32'd17,32'd7,32'd20,32'd1,32'd7,32'd0,32'd0,32'd17,32'd8,32'd11,32'd11,32'd14,32'd11,32'd20,32'd11,32'd0,32'd12,32'd2,32'd0,32'd6,32'd19,32'd16,32'd5,32'd10,32'd0,32'd3,32'd16,32'd16,32'd2,32'd12,32'd14,32'd15,32'd3,32'd6,32'd7,32'd13,32'd0,32'd3,32'd6,32'd6,32'd7,32'd6,32'd2,32'd2,32'd12,32'd12,32'd8,32'd8,32'd11,32'd19,32'd0,32'd0,32'd4,32'd4,32'd11,32'd15,32'd1,32'd1,32'd5,32'd5,32'd6,32'd11,32'd13,32'd16,32'd15,32'd17,32'd12,32'd5,32'd1,32'd1,32'd7,32'd17,32'd10,32'd10,32'd9,32'd10,32'd2,32'd1,32'd5,32'd13,32'd1,32'd4,32'd5,32'd3,32'd10,32'd1,32'd6,32'd7,32'd3,32'd2,32'd6,32'd0,32'd12,32'd8,32'd0,32'd0,32'd11,32'd3,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd20,32'd17,32'd18,32'd3,32'd11,32'd11,32'd20,32'd20,32'd14,32'd20,32'd19,32'd7,32'd12,32'd7,32'd5,32'd8,32'd21,32'd12,32'd0,32'd6,32'd3,32'd8,32'd8,32'd8,32'd2,32'd0,32'd17,32'd6,32'd13,32'd7,32'd7,32'd3,32'd0,32'd6,32'd5,32'd6,32'd2,32'd2,32'd2,32'd7,32'd0,32'd15,32'd5,32'd7,32'd7,32'd0,32'd0,32'd14,32'd5,32'd4,32'd0,32'd18,32'd17,32'd15,32'd15,32'd18,32'd1,32'd0,32'd0,32'd9,32'd8,32'd7,32'd11,32'd13,32'd0,32'd20,32'd2,32'd16,32'd11,32'd15,32'd0,32'd1,32'd6,32'd6,32'd12,32'd18,32'd18,32'd0,32'd0,32'd17,32'd9,32'd11,32'd11,32'd17,32'd17,32'd23,32'd6,32'd7,32'd7,32'd8,32'd7,32'd12,32'd3,32'd8,32'd17,32'd0,32'd0,32'd2,32'd14,32'd20,32'd2,32'd7,32'd7,32'd16,32'd4,32'd18,32'd4,32'd1,32'd6,32'd11,32'd11,32'd2,32'd5,32'd8,32'd1,32'd15,32'd8,32'd6,32'd7,32'd11,32'd6,32'd3,32'd13,32'd19,32'd4,32'd16,32'd14,32'd8,32'd15,32'd7,32'd17,32'd17,32'd6,32'd11,32'd1,32'd17,32'd10,32'd6,32'd4,32'd7,32'd9,32'd17,32'd1,32'd1,32'd0,32'd17,32'd14,32'd15,32'd14,32'd14,32'd12,32'd12,32'd0,32'd0,32'd4,32'd7,32'd0,32'd6,32'd13,32'd16,32'd22,32'd12,32'd1,32'd1,32'd12,32'd14,32'd13,32'd8,32'd5,32'd14,32'd8,32'd14,32'd0,32'd0,32'd2,32'd11,32'd5,32'd5,32'd20,32'd5,32'd6,32'd6,32'd9,32'd6,32'd6,32'd14,32'd4,32'd7,32'd14,32'd13,32'd14,32'd12,32'd6,32'd7,32'd2,32'd14,32'd22,32'd19,32'd2,32'd5,32'd3,32'd19,32'd1,32'd3,32'd4,32'd4,32'd0,32'd19,32'd18,32'd13,32'd17,32'd19,32'd10,32'd4,32'd3,32'd3,32'd0,32'd0,32'd7,32'd7,32'd15,32'd15,32'd14,32'd11,32'd11,32'd12,32'd0,32'd0,32'd0,32'd9,32'd6,32'd7,32'd0,32'd10,32'd16,32'd16,32'd10,32'd10,32'd0,32'd3,32'd6,32'd2,32'd4,32'd8,32'd10,32'd7,32'd6,32'd20,32'd2,32'd2,32'd0,32'd1,32'd14,32'd14,32'd16,32'd16,32'd1,32'd11,32'd17,32'd8,32'd2,32'd8,32'd14,32'd2,32'd1,32'd11,32'd3,32'd17,32'd15,32'd8,32'd7,32'd7,32'd21,32'd0,32'd3,32'd1,32'd2,32'd14,32'd20,32'd7,32'd0,32'd0,32'd6,32'd16,32'd11,32'd7,32'd6,32'd9,32'd14,32'd8,32'd6,32'd15,32'd20,32'd18,32'd18,32'd19,32'd7,32'd6,32'd0,32'd0,32'd4,32'd0,32'd5,32'd8,32'd16,32'd6,32'd10,32'd7,32'd1,32'd7,32'd12,32'd12,32'd11,32'd3,32'd2,32'd5,32'd1,32'd12,32'd0,32'd23,32'd1,32'd0,32'd19,32'd3,32'd4,32'd13,32'd5,32'd11,32'd2,32'd18,32'd4,32'd19,32'd16,32'd16,32'd6,32'd1,32'd1,32'd0,32'd0,32'd0,32'd4,32'd13,32'd12,32'd11,32'd11,32'd11,32'd11,32'd11,32'd5,32'd3,32'd20,32'd0,32'd0,32'd1,32'd0,32'd3,32'd0,32'd0,32'd15,32'd10,32'd14,32'd14,32'd15,32'd8,32'd8,32'd6,32'd14,32'd17,32'd13,32'd12,32'd7,32'd0,32'd0,32'd1,32'd1,32'd5,32'd4,32'd12,32'd20,32'd5,32'd10,32'd2,32'd5,32'd16,32'd16,32'd12,32'd11,32'd8,32'd3,32'd1,32'd6,32'd0,32'd19,32'd17,32'd15,32'd5,32'd5,32'd6,32'd0,32'd9,32'd11,32'd19,32'd8,32'd18,32'd16,32'd0,32'd0,32'd8,32'd8,32'd10,32'd0,32'd12,32'd16,32'd4,32'd4,32'd4,32'd17,32'd2,32'd19,32'd16,32'd8,32'd12,32'd12,32'd23,32'd18,32'd6,32'd6,32'd13,32'd6,32'd20,32'd6,32'd11,32'd0,32'd3,32'd8,32'd6,32'd6,32'd0,32'd6,32'd3,32'd0,32'd5,32'd6,32'd17,32'd17,32'd17,32'd12,32'd5,32'd1,32'd1,32'd10,32'd18,32'd17,32'd13,32'd8,32'd12,32'd14,32'd11,32'd1,32'd3,32'd3,32'd17,32'd12,32'd1,32'd5,32'd7,32'd7,32'd13,32'd11,32'd5,32'd1,32'd1,32'd7,32'd1,32'd3,32'd4,32'd5,32'd2,32'd1,32'd13,32'd1,32'd16,32'd6,32'd8,32'd1,32'd1,32'd8,32'd21,32'd12,32'd5,32'd13,32'd11,32'd3,32'd13,32'd20,32'd6,32'd6,32'd0,32'd5,32'd8,32'd5,32'd11,32'd3,32'd11,32'd14,32'd2,32'd12,32'd4,32'd8,32'd3,32'd19,32'd11,32'd13,32'd5,32'd20,32'd12,32'd4,32'd7}
`define RECTANGLE2_WIDTHS {32'd3,32'd24,32'd1,32'd9,32'd9,32'd9,32'd9,32'd18,32'd19,32'd18,32'd9,32'd11,32'd9,32'd3,32'd3,32'd6,32'd12,32'd11,32'd5,32'd8,32'd8,32'd17,32'd9,32'd3,32'd7,32'd16,32'd16,32'd4,32'd4,32'd5,32'd5,32'd4,32'd4,32'd2,32'd9,32'd3,32'd3,32'd3,32'd4,32'd6,32'd19,32'd13,32'd2,32'd2,32'd2,32'd5,32'd8,32'd12,32'd17,32'd9,32'd5,32'd2,32'd2,32'd3,32'd2,32'd9,32'd6,32'd5,32'd18,32'd8,32'd8,32'd11,32'd9,32'd18,32'd18,32'd10,32'd12,32'd13,32'd13,32'd16,32'd9,32'd14,32'd16,32'd13,32'd4,32'd9,32'd24,32'd18,32'd6,32'd2,32'd2,32'd3,32'd2,32'd18,32'd16,32'd9,32'd8,32'd6,32'd2,32'd1,32'd1,32'd9,32'd9,32'd10,32'd18,32'd3,32'd3,32'd4,32'd6,32'd16,32'd8,32'd6,32'd6,32'd7,32'd22,32'd18,32'd18,32'd3,32'd3,32'd18,32'd3,32'd9,32'd9,32'd6,32'd4,32'd6,32'd3,32'd4,32'd4,32'd1,32'd1,32'd6,32'd8,32'd16,32'd19,32'd7,32'd9,32'd18,32'd18,32'd10,32'd10,32'd9,32'd9,32'd5,32'd5,32'd5,32'd5,32'd9,32'd6,32'd9,32'd18,32'd2,32'd2,32'd6,32'd1,32'd10,32'd18,32'd10,32'd24,32'd6,32'd6,32'd11,32'd13,32'd3,32'd12,32'd6,32'd15,32'd9,32'd18,32'd18,32'd3,32'd5,32'd5,32'd7,32'd7,32'd13,32'd20,32'd4,32'd4,32'd2,32'd2,32'd1,32'd18,32'd15,32'd18,32'd6,32'd6,32'd2,32'd20,32'd2,32'd18,32'd10,32'd8,32'd3,32'd7,32'd5,32'd5,32'd2,32'd2,32'd6,32'd19,32'd6,32'd7,32'd6,32'd6,32'd12,32'd6,32'd4,32'd4,32'd12,32'd3,32'd5,32'd3,32'd9,32'd10,32'd8,32'd9,32'd3,32'd3,32'd2,32'd4,32'd4,32'd2,32'd2,32'd2,32'd2,32'd3,32'd3,32'd3,32'd7,32'd6,32'd9,32'd19,32'd19,32'd9,32'd20,32'd18,32'd5,32'd1,32'd1,32'd9,32'd3,32'd4,32'd9,32'd1,32'd1,32'd2,32'd4,32'd6,32'd11,32'd7,32'd5,32'd8,32'd3,32'd6,32'd3,32'd3,32'd6,32'd3,32'd4,32'd4,32'd11,32'd2,32'd2,32'd1,32'd1,32'd9,32'd6,32'd5,32'd12,32'd8,32'd8,32'd17,32'd17,32'd3,32'd13,32'd7,32'd7,32'd3,32'd6,32'd4,32'd5,32'd5,32'd3,32'd19,32'd7,32'd2,32'd7,32'd2,32'd3,32'd5,32'd12,32'd9,32'd9,32'd5,32'd4,32'd4,32'd3,32'd7,32'd7,32'd5,32'd6,32'd1,32'd1,32'd1,32'd4,32'd10,32'd10,32'd2,32'd3,32'd6,32'd9,32'd6,32'd6,32'd9,32'd9,32'd6,32'd4,32'd4,32'd4,32'd2,32'd18,32'd18,32'd6,32'd5,32'd5,32'd6,32'd5,32'd6,32'd5,32'd5,32'd5,32'd8,32'd4,32'd3,32'd10,32'd9,32'd6,32'd4,32'd4,32'd4,32'd4,32'd3,32'd3,32'd4,32'd7,32'd2,32'd2,32'd2,32'd3,32'd14,32'd2,32'd18,32'd24,32'd9,32'd17,32'd5,32'd18,32'd9,32'd5,32'd2,32'd2,32'd2,32'd3,32'd16,32'd3,32'd6,32'd6,32'd2,32'd7,32'd3,32'd3,32'd3,32'd18,32'd9,32'd6,32'd9,32'd9,32'd4,32'd4,32'd6,32'd2,32'd2,32'd6,32'd6,32'd2,32'd3,32'd3,32'd6,32'd6,32'd2,32'd6,32'd2,32'd6,32'd8,32'd2,32'd2,32'd9,32'd9,32'd18,32'd18,32'd9,32'd10,32'd10,32'd6,32'd19,32'd3,32'd3,32'd8,32'd5,32'd10,32'd9,32'd6,32'd17,32'd3,32'd3,32'd6,32'd22,32'd4,32'd4,32'd7,32'd4,32'd14,32'd3,32'd6,32'd9,32'd9,32'd19,32'd8,32'd5,32'd3,32'd3,32'd5,32'd3,32'd3,32'd3,32'd3,32'd4,32'd3,32'd4,32'd4,32'd4,32'd2,32'd6,32'd7,32'd10,32'd4,32'd11,32'd3,32'd11,32'd3,32'd1,32'd3,32'd10,32'd3,32'd18,32'd2,32'd3,32'd18,32'd9,32'd10,32'd6,32'd9,32'd9,32'd9,32'd9,32'd9,32'd1,32'd10,32'd4,32'd4,32'd3,32'd6,32'd18,32'd11,32'd1,32'd3,32'd3,32'd8,32'd7,32'd16,32'd2,32'd6,32'd3,32'd7,32'd3,32'd3,32'd5,32'd5,32'd6,32'd3,32'd2,32'd8,32'd2,32'd2,32'd9,32'd24,32'd10,32'd6,32'd12,32'd5,32'd18,32'd8,32'd2,32'd6,32'd3,32'd2,32'd2,32'd2,32'd19,32'd10,32'd7,32'd4,32'd3,32'd3,32'd2,32'd18,32'd16,32'd24,32'd9,32'd22,32'd2,32'd2,32'd9,32'd20,32'd10,32'd2,32'd2,32'd13,32'd9,32'd4,32'd11,32'd9,32'd5,32'd12,32'd6,32'd5,32'd3,32'd3,32'd8,32'd8,32'd3,32'd5,32'd7,32'd8,32'd7,32'd2,32'd2,32'd7,32'd24,32'd6,32'd7,32'd5,32'd2,32'd2,32'd5,32'd5,32'd5,32'd3,32'd3,32'd6,32'd3,32'd3,32'd1,32'd1,32'd9,32'd5,32'd6,32'd2,32'd7,32'd6,32'd5,32'd2,32'd8,32'd1,32'd2,32'd2,32'd18,32'd18,32'd9,32'd9,32'd9,32'd9,32'd3,32'd3,32'd2,32'd2,32'd6,32'd6,32'd7,32'd6,32'd15,32'd6,32'd6,32'd7,32'd6,32'd10,32'd8,32'd8,32'd19,32'd9,32'd5,32'd4,32'd2,32'd4,32'd24,32'd3,32'd18,32'd10,32'd18,32'd2,32'd4,32'd19,32'd2,32'd2,32'd3,32'd2,32'd12,32'd8,32'd5,32'd3,32'd1,32'd5,32'd10,32'd14,32'd9,32'd5,32'd5,32'd2,32'd2,32'd3,32'd3,32'd3,32'd3,32'd2,32'd5,32'd2,32'd6,32'd8,32'd24,32'd6,32'd2,32'd3,32'd11,32'd11,32'd9,32'd2,32'd6,32'd3,32'd6,32'd5,32'd2,32'd7,32'd7,32'd20,32'd10,32'd9,32'd12,32'd3,32'd19,32'd5,32'd24,32'd1,32'd9,32'd19,32'd16,32'd9,32'd9,32'd4,32'd8,32'd4,32'd16,32'd16,32'd18,32'd3,32'd3,32'd2,32'd4,32'd5,32'd4,32'd7,32'd24,32'd4,32'd4,32'd3,32'd2,32'd5,32'd5,32'd2,32'd6,32'd2,32'd2,32'd2,32'd2,32'd2,32'd2,32'd3,32'd3,32'd9,32'd9,32'd9,32'd18,32'd18,32'd4,32'd18,32'd9,32'd11,32'd2,32'd11,32'd14,32'd4,32'd4,32'd3,32'd4,32'd3,32'd4,32'd4,32'd4,32'd2,32'd9,32'd4,32'd11,32'd10,32'd2,32'd18,32'd2,32'd6,32'd6,32'd7,32'd7,32'd6,32'd7,32'd10,32'd9,32'd18,32'd18,32'd4,32'd2,32'd24,32'd18,32'd10,32'd4,32'd2,32'd24,32'd8,32'd15,32'd18,32'd10,32'd3,32'd5,32'd4,32'd4,32'd7,32'd1,32'd6,32'd6,32'd4,32'd4,32'd3,32'd4,32'd5,32'd20,32'd3,32'd18,32'd2,32'd11,32'd7,32'd15,32'd19,32'd2,32'd18,32'd4,32'd2,32'd6,32'd9,32'd9,32'd6,32'd2,32'd3,32'd2,32'd6,32'd2,32'd20,32'd15,32'd3,32'd3,32'd2,32'd3,32'd2,32'd10,32'd6,32'd4,32'd6,32'd6,32'd6,32'd18,32'd18,32'd2,32'd6,32'd8,32'd16,32'd19,32'd19,32'd10,32'd10,32'd24,32'd6,32'd6,32'd6,32'd8,32'd6,32'd19,32'd2,32'd6,32'd6,32'd12,32'd6,32'd4,32'd5,32'd2,32'd3,32'd2,32'd22,32'd4,32'd10,32'd5,32'd7,32'd9,32'd4,32'd2,32'd9,32'd2,32'd2,32'd2,32'd2,32'd2,32'd6,32'd9,32'd9,32'd8,32'd8,32'd14,32'd7,32'd9,32'd19,32'd2,32'd2,32'd1,32'd2,32'd5,32'd2,32'd6,32'd2,32'd2,32'd2,32'd5,32'd6,32'd6,32'd6,32'd3,32'd18,32'd3,32'd20,32'd6,32'd6,32'd9,32'd18,32'd19,32'd23,32'd10,32'd24,32'd2,32'd2,32'd2,32'd2,32'd4,32'd4,32'd4,32'd5,32'd3,32'd10,32'd2,32'd2,32'd9,32'd7,32'd8,32'd2,32'd2,32'd2,32'd2,32'd2,32'd6,32'd6,32'd19,32'd23,32'd9,32'd12,32'd11,32'd4,32'd12,32'd3,32'd5,32'd7,32'd5,32'd6,32'd4,32'd4,32'd12,32'd10,32'd3,32'd1,32'd2,32'd4,32'd4,32'd7,32'd7,32'd3,32'd12,32'd8,32'd8,32'd3,32'd2,32'd2,32'd2,32'd2,32'd5,32'd4,32'd7,32'd10,32'd19,32'd10,32'd6,32'd24,32'd4,32'd18,32'd10,32'd10,32'd6,32'd4,32'd6,32'd6,32'd10,32'd10,32'd12,32'd9,32'd6,32'd6,32'd3,32'd4,32'd6,32'd4,32'd10,32'd18,32'd16,32'd7,32'd6,32'd19,32'd4,32'd5,32'd3,32'd9,32'd10,32'd10,32'd18,32'd3,32'd2,32'd8,32'd3,32'd2,32'd2,32'd2,32'd2,32'd2,32'd9,32'd6,32'd10,32'd6,32'd3,32'd15,32'd9,32'd9,32'd2,32'd3,32'd2,32'd2,32'd2,32'd2,32'd18,32'd22,32'd7,32'd9,32'd6,32'd2,32'd5,32'd10,32'd4,32'd13,32'd7,32'd3,32'd10,32'd2,32'd4,32'd4,32'd3,32'd3,32'd10,32'd12,32'd10,32'd10,32'd9,32'd6,32'd18,32'd3,32'd14,32'd14,32'd9,32'd19,32'd20,32'd12,32'd5,32'd1,32'd7,32'd7,32'd18,32'd10,32'd2,32'd2,32'd3,32'd6,32'd8,32'd5,32'd3,32'd3,32'd5,32'd3,32'd5,32'd9,32'd8,32'd6,32'd3,32'd21,32'd2,32'd3,32'd4,32'd18,32'd5,32'd5,32'd17,32'd6,32'd2,32'd2,32'd1,32'd8,32'd6,32'd4,32'd15,32'd12,32'd2,32'd6,32'd13,32'd4,32'd20,32'd14,32'd12,32'd12,32'd4,32'd2,32'd2,32'd2,32'd9,32'd9,32'd2,32'd2,32'd4,32'd4,32'd2,32'd2,32'd8,32'd1,32'd2,32'd4,32'd3,32'd3,32'd3,32'd7,32'd5,32'd10,32'd18,32'd10,32'd3,32'd2,32'd2,32'd12,32'd15,32'd15,32'd18,32'd10,32'd9,32'd18,32'd10,32'd16,32'd6,32'd6,32'd2,32'd5,32'd9,32'd11,32'd24,32'd9,32'd12,32'd6,32'd6,32'd8,32'd4,32'd6,32'd3,32'd3,32'd4,32'd15,32'd14,32'd9,32'd2,32'd2,32'd2,32'd2,32'd18,32'd2,32'd4,32'd10,32'd7,32'd5,32'd4,32'd9,32'd6,32'd5,32'd10,32'd3,32'd10,32'd4,32'd1,32'd18,32'd8,32'd1,32'd18,32'd18,32'd9,32'd9,32'd24,32'd19,32'd9,32'd18,32'd8,32'd6,32'd9,32'd7,32'd6,32'd6,32'd4,32'd7,32'd8,32'd5,32'd6,32'd21,32'd2,32'd16,32'd14,32'd6,32'd2,32'd6,32'd2,32'd12,32'd7,32'd3,32'd3,32'd3,32'd6,32'd6,32'd2,32'd2,32'd2,32'd2,32'd9,32'd2,32'd2,32'd2,32'd5,32'd20,32'd3,32'd6,32'd5,32'd16,32'd3,32'd4,32'd17,32'd2,32'd9,32'd5,32'd19,32'd3,32'd6,32'd4,32'd4,32'd6,32'd7,32'd4,32'd12,32'd21,32'd14,32'd8,32'd12,32'd11,32'd11,32'd18,32'd9,32'd6,32'd8,32'd23,32'd9,32'd5,32'd5,32'd5,32'd2,32'd2,32'd18,32'd2,32'd2,32'd6,32'd18,32'd4,32'd6,32'd3,32'd18,32'd2,32'd2,32'd6,32'd22,32'd18,32'd11,32'd6,32'd6,32'd3,32'd6,32'd11,32'd21,32'd10,32'd9,32'd4,32'd4,32'd5,32'd4,32'd3,32'd11,32'd6,32'd6,32'd5,32'd18,32'd16,32'd4,32'd5,32'd18,32'd2,32'd19,32'd4,32'd3,32'd3,32'd4,32'd7,32'd2,32'd2,32'd3,32'd4,32'd11,32'd8,32'd8,32'd5,32'd3,32'd5,32'd5,32'd5,32'd11,32'd6,32'd6,32'd18,32'd6,32'd2,32'd2,32'd5,32'd5,32'd2,32'd6,32'd5,32'd6,32'd1,32'd1,32'd3,32'd18,32'd2,32'd2,32'd2,32'd23,32'd7,32'd17,32'd20,32'd6,32'd9,32'd9,32'd5,32'd4,32'd16,32'd3,32'd6,32'd24,32'd4,32'd3,32'd8,32'd4,32'd6,32'd6,32'd9,32'd9,32'd6,32'd6,32'd15,32'd9,32'd20,32'd7,32'd6,32'd9,32'd18,32'd14,32'd18,32'd4,32'd2,32'd2,32'd6,32'd9,32'd19,32'd3,32'd1,32'd4,32'd2,32'd2,32'd2,32'd3,32'd20,32'd4,32'd7,32'd6,32'd16,32'd18,32'd2,32'd12,32'd8,32'd2,32'd5,32'd10,32'd10,32'd6,32'd3,32'd2,32'd9,32'd7,32'd10,32'd6,32'd3,32'd4,32'd4,32'd2,32'd2,32'd9,32'd10,32'd9,32'd9,32'd19,32'd3,32'd7,32'd7,32'd6,32'd10,32'd4,32'd8,32'd20,32'd24,32'd9,32'd9,32'd18,32'd9,32'd12,32'd9,32'd12,32'd17,32'd14,32'd6,32'd2,32'd2,32'd2,32'd6,32'd3,32'd7,32'd9,32'd2,32'd6,32'd6,32'd12,32'd22,32'd18,32'd18,32'd4,32'd6,32'd6,32'd12,32'd12,32'd4,32'd4,32'd24,32'd7,32'd5,32'd4,32'd4,32'd4,32'd4,32'd3,32'd4,32'd16,32'd18,32'd8,32'd4,32'd4,32'd4,32'd3,32'd11,32'd3,32'd3,32'd2,32'd6,32'd5,32'd4,32'd5,32'd5,32'd4,32'd6,32'd6,32'd9,32'd21,32'd5,32'd4,32'd4,32'd5,32'd5,32'd11,32'd9,32'd2,32'd3,32'd3,32'd3,32'd2,32'd2,32'd4,32'd5,32'd1,32'd2,32'd6,32'd2,32'd6,32'd20,32'd2,32'd2,32'd2,32'd6,32'd4,32'd24,32'd6,32'd7,32'd9,32'd11,32'd18,32'd18,32'd2,32'd8,32'd8,32'd2,32'd6,32'd6,32'd9,32'd16,32'd6,32'd6,32'd22,32'd18,32'd9,32'd9,32'd12,32'd6,32'd2,32'd6,32'd8,32'd2,32'd2,32'd5,32'd2,32'd2,32'd2,32'd19,32'd2,32'd2,32'd3,32'd2,32'd3,32'd4,32'd10,32'd6,32'd6,32'd20,32'd5,32'd3,32'd4,32'd10,32'd8,32'd1,32'd22,32'd5,32'd4,32'd2,32'd2,32'd3,32'd3,32'd2,32'd18,32'd3,32'd5,32'd3,32'd3,32'd5,32'd5,32'd9,32'd18,32'd6,32'd6,32'd6,32'd6,32'd5,32'd5,32'd3,32'd8,32'd6,32'd4,32'd3,32'd2,32'd12,32'd9,32'd4,32'd4,32'd6,32'd6,32'd5,32'd1,32'd4,32'd20,32'd12,32'd9,32'd6,32'd6,32'd12,32'd3,32'd4,32'd3,32'd4,32'd6,32'd3,32'd9,32'd9,32'd6,32'd18,32'd18,32'd3,32'd20,32'd9,32'd12,32'd7,32'd18,32'd2,32'd2,32'd1,32'd1,32'd1,32'd1,32'd12,32'd6,32'd6,32'd6,32'd5,32'd5,32'd3,32'd3,32'd2,32'd4,32'd4,32'd4,32'd13,32'd18,32'd9,32'd2,32'd2,32'd6,32'd6,32'd6,32'd3,32'd5,32'd11,32'd7,32'd11,32'd6,32'd19,32'd18,32'd5,32'd10,32'd10,32'd6,32'd11,32'd4,32'd9,32'd6,32'd3,32'd3,32'd4,32'd4,32'd6,32'd2,32'd2,32'd4,32'd3,32'd4,32'd5,32'd4,32'd9,32'd18,32'd23,32'd9,32'd18,32'd9,32'd2,32'd2,32'd2,32'd2,32'd2,32'd24,32'd6,32'd6,32'd22,32'd6,32'd18,32'd20,32'd20,32'd2,32'd2,32'd2,32'd9,32'd9,32'd3,32'd4,32'd10,32'd18,32'd3,32'd2,32'd2,32'd2,32'd2,32'd10,32'd6,32'd20,32'd3,32'd2,32'd3,32'd6,32'd5,32'd8,32'd15,32'd4,32'd4,32'd4,32'd12,32'd8,32'd8,32'd12,32'd6,32'd6,32'd5,32'd9,32'd6,32'd6,32'd11,32'd9,32'd10,32'd4,32'd10,32'd2,32'd4,32'd9,32'd9,32'd9,32'd9,32'd15,32'd9,32'd6,32'd6,32'd2,32'd2,32'd4,32'd4,32'd2,32'd10,32'd10,32'd7,32'd8,32'd6,32'd6,32'd4,32'd5,32'd9,32'd4,32'd19,32'd6,32'd5,32'd9,32'd8,32'd2,32'd2,32'd2,32'd2,32'd2,32'd18,32'd3,32'd3,32'd3,32'd6,32'd7,32'd7,32'd3,32'd10,32'd6,32'd6,32'd7,32'd7,32'd6,32'd9,32'd12,32'd22,32'd7,32'd21,32'd9,32'd7,32'd1,32'd1,32'd2,32'd2,32'd18,32'd8,32'd18,32'd2,32'd18,32'd7,32'd11,32'd6,32'd2,32'd2,32'd5,32'd2,32'd19,32'd18,32'd18,32'd18,32'd9,32'd9,32'd9,32'd9,32'd2,32'd8,32'd16,32'd5,32'd6,32'd9,32'd10,32'd2,32'd6,32'd6,32'd7,32'd10,32'd3,32'd2,32'd2,32'd3,32'd7,32'd7,32'd2,32'd9,32'd2,32'd2,32'd2,32'd8,32'd6,32'd6,32'd2,32'd2,32'd6,32'd6,32'd8,32'd2,32'd20,32'd19,32'd4,32'd9,32'd2,32'd14,32'd3,32'd21,32'd4,32'd10,32'd19,32'd16,32'd14,32'd20,32'd6,32'd11,32'd11,32'd12,32'd9,32'd12,32'd5,32'd5,32'd3,32'd4,32'd4,32'd3,32'd9,32'd9,32'd3,32'd2,32'd2,32'd5,32'd3,32'd3,32'd7,32'd7,32'd6,32'd9,32'd6,32'd9,32'd8,32'd5,32'd3,32'd3,32'd7,32'd6,32'd13,32'd6,32'd9,32'd14,32'd24,32'd9,32'd18,32'd9,32'd19,32'd9,32'd6,32'd11,32'd4,32'd5,32'd4,32'd14,32'd4,32'd4,32'd3,32'd18,32'd8,32'd3,32'd10,32'd10,32'd2,32'd9,32'd18,32'd19,32'd2,32'd1,32'd5,32'd3,32'd1,32'd2,32'd6,32'd1,32'd2,32'd1,32'd6,32'd6,32'd2,32'd2,32'd2,32'd6,32'd8,32'd7,32'd18,32'd9,32'd11,32'd8,32'd9,32'd7,32'd3,32'd3,32'd19,32'd21,32'd3,32'd4,32'd21,32'd11,32'd6,32'd2,32'd2,32'd4,32'd15,32'd4,32'd3,32'd16,32'd6,32'd19,32'd3,32'd3,32'd3,32'd3,32'd2,32'd2,32'd9,32'd18,32'd6,32'd6,32'd2,32'd2,32'd24,32'd13,32'd8,32'd19,32'd5,32'd8,32'd4,32'd4,32'd8,32'd4,32'd6,32'd2,32'd7,32'd23,32'd10,32'd5,32'd5,32'd1,32'd3,32'd8,32'd3,32'd4,32'd4,32'd3,32'd12,32'd6,32'd4,32'd20,32'd7,32'd10,32'd4,32'd2,32'd4,32'd6,32'd4,32'd6,32'd8,32'd5,32'd5,32'd2,32'd11,32'd7,32'd9,32'd4,32'd18,32'd8,32'd9,32'd7,32'd19,32'd15,32'd9,32'd6,32'd6,32'd2,32'd2,32'd20,32'd16,32'd2,32'd2,32'd2,32'd2,32'd5,32'd6,32'd4,32'd4,32'd12,32'd11,32'd3,32'd18,32'd10,32'd24,32'd3,32'd18,32'd9,32'd14,32'd8,32'd4,32'd3,32'd2,32'd5,32'd5,32'd7,32'd11,32'd13,32'd20,32'd11,32'd18,32'd2,32'd2,32'd3,32'd11,32'd2,32'd6,32'd14,32'd19,32'd6,32'd4,32'd21,32'd4,32'd6,32'd6,32'd3,32'd3,32'd2,32'd10,32'd4,32'd2,32'd23,32'd4,32'd2,32'd4,32'd3,32'd2,32'd4,32'd7,32'd16,32'd7,32'd3,32'd6,32'd4,32'd2,32'd6,32'd4,32'd4,32'd16,32'd8,32'd3,32'd8,32'd8,32'd2,32'd20,32'd3,32'd11,32'd19,32'd9,32'd9,32'd12,32'd2,32'd2,32'd2,32'd4,32'd18,32'd3,32'd18,32'd8,32'd18,32'd2,32'd10,32'd7,32'd5,32'd2,32'd3,32'd4,32'd3,32'd4,32'd4,32'd9,32'd9,32'd20,32'd12,32'd6,32'd3,32'd4,32'd10,32'd9,32'd6,32'd8,32'd3,32'd4,32'd4,32'd5,32'd5,32'd4,32'd2,32'd6,32'd16,32'd2,32'd16,32'd3,32'd6,32'd3,32'd2,32'd2,32'd6,32'd22,32'd6,32'd6,32'd5,32'd11,32'd3,32'd21,32'd8,32'd2,32'd6,32'd5,32'd2,32'd2,32'd18,32'd9,32'd9,32'd18,32'd12,32'd18,32'd12,32'd3,32'd3,32'd9,32'd9,32'd18,32'd4,32'd23,32'd12,32'd5,32'd7,32'd4,32'd3,32'd3,32'd10,32'd9,32'd9,32'd9,32'd5,32'd4,32'd11,32'd19,32'd23,32'd6,32'd2,32'd2,32'd6,32'd4,32'd4,32'd5,32'd5,32'd18,32'd12,32'd7,32'd3,32'd8,32'd6,32'd20,32'd18,32'd2,32'd2,32'd2,32'd2,32'd2,32'd9,32'd4,32'd18,32'd12,32'd3,32'd19,32'd4,32'd6,32'd6,32'd8,32'd9,32'd2,32'd2,32'd2,32'd6,32'd18,32'd9,32'd2,32'd3,32'd8,32'd2,32'd22,32'd9,32'd7,32'd4,32'd22,32'd7,32'd4,32'd4,32'd18,32'd9,32'd14,32'd1,32'd1,32'd7,32'd7,32'd9,32'd17,32'd4,32'd4,32'd12,32'd6,32'd10,32'd2,32'd3,32'd2,32'd2,32'd22,32'd20,32'd2,32'd18,32'd6,32'd19,32'd3,32'd7,32'd4,32'd9,32'd8,32'd6,32'd10,32'd4,32'd4,32'd6,32'd20,32'd6,32'd6,32'd6,32'd6,32'd21,32'd10,32'd4,32'd4,32'd2,32'd3,32'd3,32'd3,32'd3,32'd3,32'd5,32'd5,32'd1,32'd7,32'd5,32'd3,32'd3,32'd4,32'd6,32'd18,32'd6,32'd1,32'd9,32'd1,32'd3,32'd3,32'd2,32'd2,32'd2,32'd2,32'd10,32'd10,32'd1,32'd6,32'd18,32'd23,32'd9,32'd18,32'd18,32'd9,32'd8,32'd8,32'd5,32'd19,32'd14,32'd9,32'd4,32'd4,32'd6,32'd5,32'd2,32'd10,32'd3,32'd10,32'd20,32'd4,32'd2,32'd2,32'd10,32'd11,32'd3,32'd3,32'd10,32'd3,32'd8,32'd3,32'd3,32'd14,32'd18,32'd3,32'd3,32'd4,32'd14,32'd4,32'd15,32'd8,32'd10,32'd5,32'd5,32'd1,32'd12,32'd4,32'd18,32'd6,32'd2,32'd5,32'd8,32'd3,32'd4,32'd2,32'd2,32'd2,32'd2,32'd9,32'd9,32'd14,32'd14,32'd3,32'd14,32'd3,32'd9,32'd2,32'd2,32'd9,32'd9,32'd12,32'd9,32'd2,32'd2,32'd2,32'd2,32'd18,32'd3,32'd4,32'd9,32'd6,32'd18,32'd6,32'd8,32'd2,32'd2,32'd8,32'd11,32'd4,32'd4,32'd16,32'd4,32'd2,32'd2,32'd2,32'd12,32'd18,32'd18,32'd12,32'd1,32'd12,32'd2,32'd2,32'd2,32'd24,32'd9,32'd2,32'd1,32'd4,32'd3,32'd2,32'd1,32'd6,32'd3,32'd5,32'd5,32'd5,32'd8,32'd6,32'd6,32'd6,32'd21,32'd18,32'd2,32'd9,32'd9,32'd9,32'd9,32'd6,32'd9,32'd10,32'd5,32'd8,32'd4,32'd2,32'd21,32'd6,32'd23,32'd8,32'd4,32'd11,32'd5,32'd4,32'd5,32'd7,32'd2,32'd6,32'd2,32'd7,32'd4,32'd7,32'd3,32'd2,32'd2,32'd5,32'd1,32'd5,32'd2,32'd3,32'd3,32'd2,32'd10,32'd8,32'd2,32'd3,32'd2,32'd2,32'd2,32'd3,32'd2,32'd2,32'd21,32'd18,32'd8,32'd8,32'd18,32'd12,32'd5,32'd5,32'd24,32'd6,32'd11,32'd22,32'd9,32'd12,32'd7,32'd11,32'd7,32'd12,32'd9,32'd8,32'd22,32'd15,32'd7,32'd11,32'd18,32'd18,32'd2,32'd2,32'd6,32'd6,32'd2,32'd2,32'd6,32'd6,32'd19,32'd9,32'd6,32'd6,32'd9,32'd6,32'd11,32'd2,32'd6,32'd9,32'd2,32'd2,32'd3,32'd9,32'd7,32'd3,32'd5,32'd5,32'd5,32'd2,32'd6,32'd19,32'd3,32'd2,32'd5,32'd5,32'd8,32'd2,32'd6,32'd9,32'd2,32'd2,32'd2,32'd6,32'd3,32'd16,32'd18,32'd6,32'd10,32'd24,32'd3,32'd8,32'd6,32'd6,32'd5,32'd9,32'd13,32'd11,32'd17,32'd7,32'd9,32'd6,32'd2,32'd14,32'd4,32'd9,32'd6,32'd3,32'd3,32'd5,32'd10,32'd19,32'd19,32'd9,32'd9,32'd3,32'd3,32'd2,32'd2,32'd3,32'd4,32'd9,32'd8,32'd11,32'd10,32'd18,32'd6,32'd2,32'd2,32'd5,32'd9,32'd3,32'd3,32'd3,32'd9,32'd13,32'd9,32'd2,32'd2,32'd12,32'd18,32'd6,32'd6,32'd15,32'd6,32'd3,32'd3,32'd2,32'd3,32'd2,32'd19,32'd20,32'd6,32'd3,32'd5,32'd4,32'd14,32'd4,32'd12,32'd8,32'd2,32'd18,32'd5,32'd11,32'd3,32'd10,32'd9,32'd2,32'd6,32'd1,32'd1,32'd2,32'd19,32'd18,32'd3,32'd5,32'd6,32'd3,32'd9,32'd2,32'd2,32'd2,32'd2,32'd2,32'd5,32'd6,32'd6,32'd16,32'd6,32'd13,32'd24,32'd3,32'd2,32'd1,32'd5,32'd2,32'd8,32'd8,32'd6,32'd9,32'd9,32'd9,32'd9,32'd1,32'd1,32'd6,32'd1,32'd6,32'd10,32'd8,32'd6,32'd2,32'd12,32'd3,32'd3,32'd3,32'd2,32'd13,32'd3,32'd6,32'd6,32'd3,32'd5,32'd8,32'd5,32'd3,32'd10,32'd6,32'd3,32'd2,32'd7,32'd16,32'd10,32'd10,32'd3,32'd5,32'd5,32'd9,32'd8,32'd15,32'd11,32'd12,32'd5,32'd7,32'd5,32'd1,32'd1,32'd7,32'd9,32'd18,32'd18,32'd2,32'd5,32'd5,32'd10,32'd16,32'd5,32'd5,32'd9,32'd7,32'd9,32'd2,32'd2,32'd2,32'd2,32'd12,32'd2,32'd8,32'd6,32'd18,32'd6,32'd12,32'd4,32'd3,32'd2,32'd11,32'd11,32'd7,32'd22,32'd20,32'd7,32'd2,32'd19,32'd2,32'd19,32'd18,32'd2,32'd5,32'd18,32'd3,32'd6,32'd3,32'd14,32'd6,32'd18,32'd4,32'd18,32'd9,32'd9,32'd1,32'd1,32'd1,32'd1,32'd1,32'd10,32'd11,32'd12,32'd11,32'd3,32'd3,32'd4,32'd22,32'd18,32'd12,32'd2,32'd10,32'd3,32'd3,32'd10,32'd3,32'd8,32'd3,32'd5,32'd6,32'd9,32'd8,32'd3,32'd10,32'd3,32'd3,32'd4,32'd3,32'd17,32'd6,32'd19,32'd4,32'd3,32'd3,32'd3,32'd3,32'd2,32'd17,32'd22,32'd6,32'd3,32'd12,32'd8,32'd5,32'd4,32'd4,32'd5,32'd11,32'd11,32'd19,32'd2,32'd4,32'd3,32'd18,32'd8,32'd18,32'd6,32'd5,32'd7,32'd9,32'd9,32'd20,32'd6,32'd2,32'd9,32'd9,32'd2,32'd2,32'd6,32'd6,32'd3,32'd2,32'd4,32'd10,32'd2,32'd2,32'd3,32'd18,32'd22,32'd18,32'd10,32'd10,32'd8,32'd4,32'd18,32'd6,32'd2,32'd2,32'd5,32'd2,32'd8,32'd3,32'd16,32'd8,32'd12,32'd6,32'd2,32'd2,32'd2,32'd2,32'd6,32'd4,32'd7,32'd4,32'd9,32'd9,32'd7,32'd14,32'd10,32'd18,32'd2,32'd16,32'd18,32'd9,32'd6,32'd12,32'd8,32'd3,32'd8,32'd8,32'd2,32'd2,32'd6,32'd18,32'd8,32'd4,32'd12,32'd6,32'd2,32'd18,32'd7,32'd2,32'd2,32'd19,32'd2,32'd2,32'd2,32'd11,32'd2,32'd2,32'd10,32'd2,32'd21,32'd7,32'd8,32'd3,32'd3,32'd13,32'd6,32'd3,32'd2,32'd5,32'd15,32'd8,32'd14,32'd10,32'd2,32'd8,32'd2,32'd2,32'd2,32'd2,32'd3,32'd14,32'd14,32'd6,32'd8,32'd19,32'd4,32'd12,32'd7,32'd4,32'd12,32'd12,32'd2,32'd9,32'd18,32'd4,32'd12}
`define RECTANGLE2_HEIGHTS {32'd11,32'd4,32'd20,32'd2,32'd2,32'd2,32'd2,32'd1,32'd1,32'd1,32'd2,32'd5,32'd2,32'd6,32'd6,32'd3,32'd4,32'd3,32'd4,32'd5,32'd5,32'd3,32'd2,32'd7,32'd3,32'd4,32'd4,32'd5,32'd5,32'd4,32'd4,32'd6,32'd6,32'd10,32'd2,32'd7,32'd7,32'd7,32'd5,32'd4,32'd1,32'd2,32'd12,32'd9,32'd9,32'd9,32'd3,32'd2,32'd11,32'd12,32'd6,32'd9,32'd9,32'd6,32'd9,32'd3,32'd3,32'd5,32'd1,32'd5,32'd3,32'd2,32'd2,32'd1,32'd1,32'd3,32'd3,32'd3,32'd3,32'd2,32'd2,32'd3,32'd3,32'd3,32'd5,32'd2,32'd1,32'd3,32'd3,32'd9,32'd9,32'd6,32'd9,32'd1,32'd2,32'd2,32'd3,32'd3,32'd10,32'd18,32'd18,32'd2,32'd2,32'd2,32'd1,32'd7,32'd7,32'd7,32'd4,32'd3,32'd11,32'd17,32'd17,32'd10,32'd1,32'd1,32'd1,32'd6,32'd6,32'd1,32'd6,32'd5,32'd5,32'd5,32'd5,32'd3,32'd6,32'd5,32'd5,32'd19,32'd19,32'd15,32'd12,32'd2,32'd5,32'd3,32'd6,32'd1,32'd1,32'd2,32'd2,32'd2,32'd2,32'd6,32'd6,32'd4,32'd4,32'd2,32'd3,32'd2,32'd1,32'd9,32'd9,32'd8,32'd19,32'd2,32'd1,32'd2,32'd1,32'd3,32'd3,32'd13,32'd2,32'd6,32'd3,32'd3,32'd2,32'd5,32'd1,32'd1,32'd6,32'd6,32'd6,32'd7,32'd7,32'd2,32'd1,32'd9,32'd9,32'd10,32'd10,32'd18,32'd1,32'd2,32'd1,32'd3,32'd4,32'd11,32'd1,32'd10,32'd1,32'd3,32'd5,32'd7,32'd3,32'd5,32'd5,32'd9,32'd9,32'd3,32'd1,32'd3,32'd9,32'd3,32'd3,32'd2,32'd4,32'd5,32'd6,32'd3,32'd6,32'd4,32'd6,32'd2,32'd2,32'd4,32'd3,32'd6,32'd16,32'd9,32'd20,32'd20,32'd22,32'd22,32'd14,32'd14,32'd16,32'd16,32'd16,32'd4,32'd8,32'd2,32'd1,32'd5,32'd2,32'd1,32'd1,32'd4,32'd24,32'd24,32'd13,32'd6,32'd5,32'd2,32'd22,32'd22,32'd9,32'd5,32'd4,32'd2,32'd4,32'd6,32'd10,32'd6,32'd3,32'd6,32'd7,32'd5,32'd6,32'd5,32'd5,32'd2,32'd16,32'd16,32'd19,32'd18,32'd2,32'd8,32'd8,32'd5,32'd3,32'd3,32'd3,32'd3,32'd6,32'd2,32'd7,32'd7,32'd6,32'd5,32'd5,32'd7,32'd6,32'd24,32'd1,32'd3,32'd22,32'd3,32'd9,32'd6,32'd4,32'd3,32'd2,32'd2,32'd8,32'd5,32'd5,32'd6,32'd7,32'd7,32'd9,32'd3,32'd18,32'd18,32'd19,32'd5,32'd3,32'd2,32'd9,32'd23,32'd10,32'd2,32'd3,32'd3,32'd3,32'd2,32'd9,32'd24,32'd15,32'd24,32'd10,32'd1,32'd1,32'd7,32'd6,32'd6,32'd4,32'd4,32'd9,32'd4,32'd4,32'd4,32'd4,32'd8,32'd7,32'd3,32'd2,32'd5,32'd5,32'd5,32'd5,32'd5,32'd9,32'd8,32'd5,32'd7,32'd9,32'd10,32'd9,32'd6,32'd6,32'd9,32'd1,32'd1,32'd7,32'd2,32'd4,32'd2,32'd2,32'd4,32'd24,32'd24,32'd9,32'd6,32'd3,32'd7,32'd15,32'd3,32'd13,32'd3,32'd6,32'd6,32'd7,32'd1,32'd2,32'd3,32'd2,32'd2,32'd10,32'd10,32'd3,32'd9,32'd9,32'd3,32'd4,32'd9,32'd10,32'd10,32'd3,32'd3,32'd9,32'd3,32'd12,32'd3,32'd4,32'd12,32'd9,32'd2,32'd2,32'd1,32'd1,32'd2,32'd2,32'd2,32'd3,32'd1,32'd6,32'd6,32'd3,32'd6,32'd2,32'd2,32'd3,32'd6,32'd6,32'd7,32'd3,32'd2,32'd14,32'd5,32'd3,32'd10,32'd3,32'd6,32'd5,32'd2,32'd2,32'd1,32'd8,32'd6,32'd6,32'd6,32'd4,32'd7,32'd7,32'd9,32'd9,32'd5,32'd7,32'd5,32'd5,32'd5,32'd9,32'd7,32'd6,32'd19,32'd5,32'd3,32'd7,32'd3,32'd7,32'd19,32'd7,32'd2,32'd7,32'd1,32'd12,32'd8,32'd1,32'd3,32'd2,32'd4,32'd12,32'd2,32'd2,32'd2,32'd2,32'd20,32'd11,32'd6,32'd6,32'd7,32'd4,32'd1,32'd7,32'd18,32'd6,32'd7,32'd6,32'd10,32'd6,32'd9,32'd4,32'd7,32'd4,32'd6,32'd6,32'd4,32'd4,32'd3,32'd6,32'd9,32'd3,32'd11,32'd11,32'd2,32'd2,32'd2,32'd3,32'd2,32'd6,32'd1,32'd3,32'd10,32'd5,32'd9,32'd9,32'd9,32'd9,32'd1,32'd2,32'd5,32'd5,32'd6,32'd6,32'd10,32'd2,32'd4,32'd9,32'd2,32'd1,32'd19,32'd19,32'd2,32'd1,32'd2,32'd9,32'd9,32'd2,32'd2,32'd6,32'd5,32'd2,32'd5,32'd2,32'd3,32'd4,32'd6,32'd6,32'd10,32'd10,32'd6,32'd5,32'd9,32'd10,32'd3,32'd19,32'd9,32'd10,32'd1,32'd3,32'd4,32'd4,32'd10,32'd10,32'd5,32'd5,32'd4,32'd6,32'd6,32'd19,32'd7,32'd7,32'd24,32'd24,32'd6,32'd7,32'd3,32'd10,32'd3,32'd3,32'd7,32'd9,32'd4,32'd24,32'd11,32'd11,32'd1,32'd1,32'd2,32'd2,32'd2,32'd2,32'd6,32'd6,32'd9,32'd9,32'd3,32'd3,32'd4,32'd8,32'd4,32'd3,32'd3,32'd3,32'd3,32'd2,32'd8,32'd6,32'd1,32'd2,32'd5,32'd5,32'd9,32'd5,32'd7,32'd6,32'd1,32'd5,32'd1,32'd9,32'd5,32'd1,32'd22,32'd22,32'd6,32'd10,32'd2,32'd3,32'd4,32'd8,32'd19,32'd4,32'd2,32'd2,32'd2,32'd4,32'd4,32'd9,32'd9,32'd6,32'd6,32'd6,32'd6,32'd9,32'd4,32'd10,32'd21,32'd10,32'd2,32'd7,32'd9,32'd6,32'd3,32'd2,32'd2,32'd9,32'd8,32'd7,32'd4,32'd12,32'd9,32'd10,32'd10,32'd1,32'd2,32'd2,32'd4,32'd6,32'd9,32'd4,32'd2,32'd23,32'd2,32'd2,32'd4,32'd2,32'd2,32'd5,32'd3,32'd5,32'd5,32'd2,32'd4,32'd8,32'd8,32'd9,32'd5,32'd14,32'd15,32'd3,32'd2,32'd18,32'd18,32'd6,32'd9,32'd8,32'd8,32'd9,32'd5,32'd9,32'd9,32'd10,32'd24,32'd10,32'd10,32'd16,32'd16,32'd2,32'd2,32'd2,32'd1,32'd1,32'd13,32'd1,32'd2,32'd2,32'd10,32'd2,32'd6,32'd6,32'd5,32'd7,32'd5,32'd7,32'd5,32'd5,32'd5,32'd9,32'd2,32'd5,32'd3,32'd2,32'd9,32'd1,32'd9,32'd3,32'd3,32'd4,32'd4,32'd3,32'd3,32'd21,32'd5,32'd1,32'd1,32'd5,32'd11,32'd1,32'd1,32'd3,32'd5,32'd13,32'd1,32'd9,32'd4,32'd1,32'd2,32'd7,32'd4,32'd5,32'd13,32'd3,32'd20,32'd3,32'd3,32'd5,32'd5,32'd6,32'd5,32'd4,32'd1,32'd6,32'd1,32'd9,32'd14,32'd5,32'd2,32'd1,32'd9,32'd1,32'd15,32'd9,32'd3,32'd3,32'd3,32'd10,32'd9,32'd6,32'd9,32'd7,32'd9,32'd1,32'd2,32'd11,32'd11,32'd9,32'd13,32'd13,32'd5,32'd8,32'd5,32'd3,32'd3,32'd3,32'd1,32'd1,32'd9,32'd5,32'd5,32'd3,32'd1,32'd1,32'd2,32'd2,32'd2,32'd3,32'd4,32'd4,32'd11,32'd4,32'd1,32'd10,32'd3,32'd3,32'd2,32'd7,32'd6,32'd8,32'd9,32'd6,32'd10,32'd1,32'd5,32'd2,32'd7,32'd6,32'd4,32'd6,32'd9,32'd3,32'd10,32'd10,32'd9,32'd9,32'd9,32'd8,32'd2,32'd2,32'd3,32'd3,32'd4,32'd3,32'd2,32'd2,32'd9,32'd10,32'd19,32'd10,32'd4,32'd10,32'd3,32'd10,32'd9,32'd9,32'd5,32'd9,32'd5,32'd5,32'd7,32'd1,32'd7,32'd3,32'd3,32'd3,32'd2,32'd1,32'd1,32'd4,32'd2,32'd1,32'd16,32'd16,32'd16,32'd16,32'd6,32'd6,32'd5,32'd4,32'd7,32'd2,32'd11,32'd11,32'd2,32'd3,32'd6,32'd11,32'd9,32'd9,32'd12,32'd9,32'd3,32'd7,32'd4,32'd2,32'd2,32'd2,32'd2,32'd5,32'd3,32'd6,32'd4,32'd7,32'd12,32'd3,32'd7,32'd5,32'd2,32'd2,32'd6,32'd19,32'd13,32'd5,32'd5,32'd3,32'd4,32'd6,32'd2,32'd7,32'd3,32'd6,32'd13,32'd13,32'd10,32'd9,32'd4,32'd8,32'd14,32'd2,32'd4,32'd3,32'd3,32'd2,32'd5,32'd1,32'd2,32'd2,32'd3,32'd8,32'd3,32'd3,32'd2,32'd2,32'd2,32'd3,32'd4,32'd4,32'd9,32'd6,32'd3,32'd5,32'd7,32'd1,32'd4,32'd8,32'd3,32'd1,32'd8,32'd4,32'd6,32'd2,32'd2,32'd4,32'd1,32'd6,32'd11,32'd3,32'd6,32'd9,32'd9,32'd9,32'd9,32'd9,32'd7,32'd3,32'd2,32'd3,32'd6,32'd2,32'd2,32'd2,32'd9,32'd7,32'd20,32'd20,32'd9,32'd9,32'd1,32'd1,32'd3,32'd2,32'd6,32'd9,32'd4,32'd2,32'd5,32'd3,32'd3,32'd6,32'd2,32'd10,32'd5,32'd5,32'd7,32'd7,32'd4,32'd2,32'd3,32'd3,32'd2,32'd3,32'd2,32'd7,32'd6,32'd4,32'd2,32'd1,32'd1,32'd2,32'd4,32'd21,32'd3,32'd3,32'd1,32'd3,32'd9,32'd9,32'd13,32'd3,32'd4,32'd4,32'd6,32'd6,32'd11,32'd6,32'd6,32'd5,32'd9,32'd3,32'd6,32'd1,32'd12,32'd6,32'd5,32'd1,32'd4,32'd4,32'd2,32'd3,32'd9,32'd14,32'd18,32'd5,32'd3,32'd5,32'd4,32'd2,32'd9,32'd6,32'd3,32'd5,32'd1,32'd3,32'd2,32'd2,32'd7,32'd9,32'd13,32'd13,32'd2,32'd2,32'd17,32'd17,32'd20,32'd20,32'd14,32'd14,32'd12,32'd18,32'd14,32'd6,32'd6,32'd6,32'd7,32'd3,32'd4,32'd3,32'd3,32'd2,32'd6,32'd9,32'd12,32'd2,32'd2,32'd2,32'd1,32'd3,32'd3,32'd1,32'd2,32'd3,32'd3,32'd3,32'd9,32'd4,32'd2,32'd2,32'd4,32'd2,32'd11,32'd5,32'd9,32'd3,32'd10,32'd4,32'd12,32'd12,32'd5,32'd3,32'd4,32'd2,32'd11,32'd9,32'd9,32'd9,32'd1,32'd9,32'd5,32'd2,32'd24,32'd4,32'd5,32'd2,32'd5,32'd6,32'd3,32'd7,32'd4,32'd5,32'd23,32'd1,32'd3,32'd23,32'd1,32'd1,32'd2,32'd2,32'd1,32'd1,32'd2,32'd1,32'd21,32'd21,32'd5,32'd3,32'd4,32'd4,32'd5,32'd3,32'd8,32'd4,32'd3,32'd2,32'd9,32'd6,32'd2,32'd3,32'd9,32'd3,32'd20,32'd2,32'd6,32'd8,32'd6,32'd6,32'd3,32'd3,32'd16,32'd16,32'd9,32'd9,32'd2,32'd9,32'd9,32'd9,32'd10,32'd1,32'd6,32'd3,32'd6,32'd3,32'd13,32'd11,32'd3,32'd12,32'd12,32'd5,32'd1,32'd6,32'd4,32'd5,32'd5,32'd3,32'd3,32'd5,32'd3,32'd1,32'd2,32'd4,32'd3,32'd2,32'd2,32'd1,32'd2,32'd3,32'd6,32'd5,32'd2,32'd4,32'd4,32'd4,32'd9,32'd9,32'd1,32'd13,32'd9,32'd4,32'd1,32'd6,32'd4,32'd13,32'd1,32'd9,32'd9,32'd3,32'd2,32'd2,32'd2,32'd9,32'd9,32'd6,32'd11,32'd8,32'd2,32'd3,32'd3,32'd10,32'd10,32'd7,32'd5,32'd6,32'd4,32'd3,32'd3,32'd4,32'd1,32'd2,32'd5,32'd4,32'd1,32'd13,32'd1,32'd5,32'd6,32'd6,32'd5,32'd3,32'd9,32'd18,32'd6,32'd5,32'd7,32'd3,32'd3,32'd4,32'd6,32'd7,32'd7,32'd4,32'd2,32'd3,32'd3,32'd1,32'd3,32'd16,32'd16,32'd18,32'd4,32'd11,32'd3,32'd6,32'd10,32'd24,32'd24,32'd6,32'd1,32'd13,32'd9,32'd9,32'd1,32'd3,32'd8,32'd4,32'd3,32'd4,32'd4,32'd4,32'd5,32'd2,32'd6,32'd4,32'd3,32'd5,32'd6,32'd4,32'd5,32'd3,32'd3,32'd2,32'd2,32'd3,32'd3,32'd2,32'd2,32'd1,32'd4,32'd3,32'd2,32'd1,32'd2,32'd1,32'd5,32'd9,32'd9,32'd5,32'd2,32'd1,32'd6,32'd18,32'd5,32'd11,32'd11,32'd9,32'd6,32'd1,32'd5,32'd3,32'd3,32'd2,32'd1,32'd9,32'd3,32'd7,32'd9,32'd6,32'd2,32'd3,32'd3,32'd7,32'd9,32'd3,32'd5,32'd2,32'd3,32'd6,32'd13,32'd5,32'd9,32'd9,32'd2,32'd2,32'd2,32'd2,32'd4,32'd6,32'd5,32'd5,32'd4,32'd2,32'd5,32'd6,32'd3,32'd2,32'd2,32'd2,32'd1,32'd5,32'd3,32'd3,32'd7,32'd4,32'd2,32'd5,32'd9,32'd9,32'd16,32'd4,32'd6,32'd6,32'd2,32'd9,32'd3,32'd3,32'd3,32'd1,32'd1,32'd1,32'd5,32'd3,32'd6,32'd3,32'd3,32'd8,32'd11,32'd5,32'd3,32'd4,32'd7,32'd7,32'd10,32'd10,32'd6,32'd10,32'd4,32'd4,32'd4,32'd9,32'd7,32'd7,32'd8,32'd6,32'd7,32'd7,32'd9,32'd3,32'd4,32'd5,32'd4,32'd4,32'd6,32'd6,32'd4,32'd2,32'd1,32'd5,32'd16,32'd16,32'd5,32'd5,32'd4,32'd3,32'd10,32'd8,32'd7,32'd7,32'd9,32'd9,32'd8,32'd5,32'd18,32'd13,32'd4,32'd13,32'd3,32'd1,32'd9,32'd9,32'd9,32'd6,32'd5,32'd2,32'd3,32'd3,32'd2,32'd2,32'd1,32'd1,32'd23,32'd4,32'd3,32'd23,32'd3,32'd3,32'd2,32'd3,32'd3,32'd3,32'd2,32'd1,32'd2,32'd2,32'd2,32'd3,32'd9,32'd3,32'd4,32'd9,32'd9,32'd4,32'd9,32'd9,32'd9,32'd1,32'd17,32'd17,32'd6,32'd17,32'd8,32'd9,32'd2,32'd3,32'd4,32'd3,32'd4,32'd7,32'd5,32'd2,32'd4,32'd20,32'd1,32'd5,32'd18,32'd11,32'd11,32'd6,32'd7,32'd9,32'd1,32'd7,32'd4,32'd11,32'd12,32'd4,32'd4,32'd2,32'd2,32'd3,32'd3,32'd3,32'd3,32'd4,32'd4,32'd14,32'd12,32'd3,32'd5,32'd7,32'd9,32'd2,32'd5,32'd7,32'd7,32'd4,32'd6,32'd4,32'd24,32'd6,32'd1,32'd3,32'd2,32'd3,32'd3,32'd3,32'd6,32'd5,32'd6,32'd9,32'd3,32'd7,32'd2,32'd2,32'd3,32'd1,32'd1,32'd6,32'd1,32'd5,32'd4,32'd4,32'd7,32'd12,32'd12,32'd20,32'd20,32'd19,32'd19,32'd2,32'd4,32'd5,32'd3,32'd5,32'd5,32'd6,32'd6,32'd9,32'd7,32'd6,32'd6,32'd7,32'd1,32'd2,32'd23,32'd9,32'd3,32'd4,32'd3,32'd7,32'd4,32'd3,32'd4,32'd2,32'd3,32'd1,32'd1,32'd4,32'd6,32'd9,32'd3,32'd4,32'd5,32'd3,32'd3,32'd19,32'd7,32'd5,32'd5,32'd4,32'd9,32'd9,32'd5,32'd12,32'd5,32'd6,32'd5,32'd2,32'd1,32'd2,32'd2,32'd1,32'd2,32'd9,32'd9,32'd9,32'd9,32'd10,32'd2,32'd3,32'd3,32'd3,32'd3,32'd1,32'd1,32'd1,32'd9,32'd11,32'd11,32'd11,32'd11,32'd6,32'd6,32'd2,32'd1,32'd6,32'd9,32'd9,32'd9,32'd9,32'd2,32'd3,32'd1,32'd8,32'd9,32'd6,32'd3,32'd8,32'd6,32'd3,32'd7,32'd5,32'd5,32'd11,32'd3,32'd3,32'd3,32'd3,32'd13,32'd16,32'd2,32'd3,32'd5,32'd2,32'd2,32'd2,32'd5,32'd2,32'd16,32'd5,32'd2,32'd2,32'd2,32'd2,32'd11,32'd2,32'd4,32'd4,32'd16,32'd9,32'd8,32'd8,32'd9,32'd3,32'd2,32'd3,32'd3,32'd3,32'd3,32'd7,32'd4,32'd2,32'd10,32'd1,32'd3,32'd4,32'd4,32'd4,32'd9,32'd9,32'd13,32'd15,32'd11,32'd1,32'd6,32'd6,32'd6,32'd4,32'd8,32'd15,32'd8,32'd5,32'd3,32'd3,32'd3,32'd3,32'd4,32'd2,32'd8,32'd1,32'd3,32'd1,32'd2,32'd3,32'd18,32'd18,32'd9,32'd9,32'd1,32'd3,32'd1,32'd9,32'd1,32'd12,32'd2,32'd3,32'd11,32'd11,32'd6,32'd11,32'd1,32'd1,32'd1,32'd1,32'd2,32'd2,32'd2,32'd2,32'd10,32'd3,32'd2,32'd7,32'd3,32'd2,32'd4,32'd10,32'd6,32'd3,32'd7,32'd2,32'd9,32'd9,32'd10,32'd9,32'd3,32'd3,32'd9,32'd2,32'd20,32'd21,32'd13,32'd21,32'd3,32'd3,32'd10,32'd10,32'd3,32'd3,32'd4,32'd13,32'd1,32'd1,32'd7,32'd3,32'd9,32'd3,32'd6,32'd1,32'd5,32'd2,32'd1,32'd3,32'd7,32'd2,32'd9,32'd2,32'd2,32'd3,32'd2,32'd2,32'd4,32'd4,32'd8,32'd6,32'd5,32'd6,32'd2,32'd2,32'd8,32'd9,32'd9,32'd4,32'd10,32'd17,32'd5,32'd5,32'd3,32'd2,32'd3,32'd2,32'd3,32'd4,32'd7,32'd6,32'd3,32'd4,32'd2,32'd3,32'd2,32'd2,32'd1,32'd2,32'd1,32'd2,32'd1,32'd2,32'd3,32'd3,32'd7,32'd4,32'd5,32'd2,32'd5,32'd5,32'd6,32'd1,32'd8,32'd6,32'd2,32'd2,32'd9,32'd2,32'd1,32'd1,32'd12,32'd18,32'd5,32'd6,32'd19,32'd9,32'd4,32'd19,32'd9,32'd19,32'd3,32'd3,32'd10,32'd10,32'd9,32'd5,32'd4,32'd3,32'd1,32'd2,32'd2,32'd3,32'd2,32'd7,32'd7,32'd7,32'd1,32'd1,32'd6,32'd6,32'd1,32'd2,32'd4,32'd9,32'd9,32'd5,32'd6,32'd7,32'd6,32'd2,32'd4,32'd1,32'd8,32'd8,32'd19,32'd19,32'd9,32'd9,32'd2,32'd1,32'd3,32'd4,32'd9,32'd11,32'd1,32'd4,32'd9,32'd1,32'd4,32'd5,32'd8,32'd8,32'd4,32'd8,32'd3,32'd9,32'd3,32'd6,32'd3,32'd7,32'd7,32'd18,32'd8,32'd6,32'd6,32'd8,32'd8,32'd7,32'd2,32'd5,32'd8,32'd1,32'd7,32'd2,32'd8,32'd9,32'd6,32'd6,32'd7,32'd3,32'd3,32'd5,32'd5,32'd9,32'd3,32'd7,32'd2,32'd6,32'd1,32'd4,32'd2,32'd8,32'd1,32'd2,32'd2,32'd3,32'd7,32'd13,32'd13,32'd1,32'd3,32'd10,32'd10,32'd10,32'd9,32'd10,32'd3,32'd6,32'd5,32'd11,32'd2,32'd8,32'd1,32'd2,32'd1,32'd6,32'd1,32'd2,32'd3,32'd3,32'd5,32'd6,32'd9,32'd4,32'd4,32'd3,32'd15,32'd2,32'd1,32'd2,32'd1,32'd23,32'd23,32'd6,32'd2,32'd9,32'd4,32'd2,32'd1,32'd7,32'd6,32'd1,32'd6,32'd13,32'd13,32'd6,32'd6,32'd12,32'd2,32'd5,32'd12,32'd1,32'd5,32'd10,32'd8,32'd7,32'd9,32'd7,32'd3,32'd3,32'd3,32'd6,32'd3,32'd6,32'd9,32'd3,32'd5,32'd6,32'd4,32'd3,32'd7,32'd3,32'd3,32'd10,32'd1,32'd6,32'd6,32'd1,32'd2,32'd2,32'd2,32'd9,32'd9,32'd9,32'd5,32'd1,32'd6,32'd1,32'd3,32'd1,32'd15,32'd2,32'd6,32'd4,32'd9,32'd6,32'd5,32'd8,32'd6,32'd6,32'd2,32'd3,32'd1,32'd2,32'd3,32'd6,32'd6,32'd2,32'd2,32'd4,32'd3,32'd8,32'd5,32'd5,32'd4,32'd4,32'd5,32'd9,32'd4,32'd2,32'd10,32'd10,32'd7,32'd8,32'd7,32'd9,32'd9,32'd4,32'd11,32'd4,32'd3,32'd4,32'd4,32'd6,32'd2,32'd3,32'd11,32'd4,32'd4,32'd9,32'd10,32'd1,32'd2,32'd2,32'd1,32'd2,32'd1,32'd3,32'd6,32'd6,32'd2,32'd2,32'd1,32'd5,32'd2,32'd2,32'd7,32'd6,32'd5,32'd10,32'd18,32'd4,32'd2,32'd2,32'd3,32'd4,32'd5,32'd2,32'd1,32'd1,32'd6,32'd11,32'd9,32'd6,32'd9,32'd9,32'd4,32'd4,32'd1,32'd5,32'd7,32'd6,32'd4,32'd4,32'd1,32'd1,32'd11,32'd10,32'd18,32'd18,32'd9,32'd14,32'd6,32'd1,32'd3,32'd7,32'd1,32'd5,32'd4,32'd4,32'd3,32'd2,32'd17,32'd10,32'd11,32'd3,32'd1,32'd6,32'd9,32'd6,32'd9,32'd17,32'd2,32'd2,32'd4,32'd5,32'd2,32'd4,32'd5,32'd8,32'd3,32'd2,32'd2,32'd18,32'd18,32'd3,32'd3,32'd4,32'd3,32'd5,32'd5,32'd3,32'd6,32'd2,32'd9,32'd19,32'd23,32'd9,32'd1,32'd1,32'd9,32'd1,32'd3,32'd1,32'd6,32'd6,32'd5,32'd2,32'd3,32'd5,32'd13,32'd5,32'd5,32'd3,32'd2,32'd3,32'd3,32'd6,32'd6,32'd2,32'd2,32'd10,32'd10,32'd9,32'd7,32'd7,32'd7,32'd6,32'd6,32'd20,32'd20,32'd19,32'd3,32'd4,32'd8,32'd6,32'd5,32'd4,32'd1,32'd3,32'd19,32'd2,32'd19,32'd9,32'd6,32'd9,32'd9,32'd9,32'd12,32'd2,32'd2,32'd22,32'd3,32'd1,32'd5,32'd2,32'd1,32'd1,32'd5,32'd11,32'd18,32'd8,32'd4,32'd3,32'd2,32'd8,32'd5,32'd3,32'd4,32'd9,32'd3,32'd11,32'd2,32'd1,32'd5,32'd9,32'd9,32'd2,32'd4,32'd7,32'd6,32'd2,32'd7,32'd3,32'd6,32'd6,32'd6,32'd1,32'd6,32'd7,32'd5,32'd3,32'd6,32'd2,32'd3,32'd3,32'd4,32'd4,32'd20,32'd2,32'd5,32'd1,32'd3,32'd9,32'd6,32'd4,32'd21,32'd9,32'd15,32'd15,32'd9,32'd14,32'd2,32'd2,32'd5,32'd5,32'd6,32'd6,32'd6,32'd2,32'd17,32'd17,32'd2,32'd2,32'd2,32'd9,32'd9,32'd9,32'd11,32'd11,32'd1,32'd6,32'd5,32'd2,32'd3,32'd1,32'd3,32'd4,32'd16,32'd16,32'd9,32'd3,32'd7,32'd7,32'd5,32'd7,32'd22,32'd9,32'd9,32'd2,32'd1,32'd4,32'd4,32'd21,32'd6,32'd12,32'd10,32'd9,32'd1,32'd2,32'd9,32'd18,32'd5,32'd7,32'd9,32'd18,32'd3,32'd10,32'd5,32'd5,32'd8,32'd5,32'd3,32'd3,32'd3,32'd2,32'd1,32'd9,32'd2,32'd2,32'd2,32'd2,32'd8,32'd2,32'd2,32'd12,32'd5,32'd5,32'd12,32'd2,32'd3,32'd2,32'd5,32'd5,32'd3,32'd4,32'd5,32'd4,32'd3,32'd13,32'd3,32'd9,32'd6,32'd6,32'd3,32'd7,32'd9,32'd10,32'd6,32'd18,32'd7,32'd9,32'd15,32'd7,32'd9,32'd2,32'd14,32'd12,32'd7,32'd24,32'd24,32'd10,32'd6,32'd11,32'd24,32'd5,32'd1,32'd3,32'd3,32'd1,32'd2,32'd5,32'd5,32'd2,32'd3,32'd4,32'd1,32'd2,32'd8,32'd3,32'd3,32'd4,32'd3,32'd4,32'd24,32'd1,32'd2,32'd3,32'd6,32'd1,32'd1,32'd9,32'd9,32'd5,32'd7,32'd9,32'd9,32'd3,32'd3,32'd1,32'd2,32'd3,32'd3,32'd2,32'd3,32'd7,32'd11,32'd5,32'd2,32'd14,32'd14,32'd6,32'd2,32'd4,32'd6,32'd6,32'd6,32'd7,32'd19,32'd3,32'd3,32'd17,32'd9,32'd4,32'd4,32'd4,32'd9,32'd7,32'd21,32'd9,32'd10,32'd9,32'd4,32'd6,32'd3,32'd3,32'd3,32'd2,32'd1,32'd6,32'd4,32'd3,32'd3,32'd4,32'd2,32'd2,32'd6,32'd2,32'd23,32'd2,32'd3,32'd9,32'd4,32'd6,32'd6,32'd3,32'd6,32'd6,32'd6,32'd2,32'd1,32'd1,32'd2,32'd2,32'd6,32'd6,32'd9,32'd9,32'd10,32'd7,32'd11,32'd3,32'd2,32'd3,32'd1,32'd3,32'd19,32'd19,32'd4,32'd2,32'd7,32'd6,32'd15,32'd2,32'd2,32'd2,32'd9,32'd9,32'd2,32'd1,32'd3,32'd3,32'd2,32'd3,32'd9,32'd9,32'd12,32'd14,32'd9,32'd2,32'd1,32'd8,32'd8,32'd7,32'd5,32'd4,32'd5,32'd3,32'd4,32'd10,32'd1,32'd5,32'd8,32'd6,32'd8,32'd3,32'd14,32'd9,32'd18,32'd18,32'd9,32'd1,32'd1,32'd8,32'd4,32'd5,32'd7,32'd2,32'd15,32'd15,32'd9,32'd9,32'd9,32'd4,32'd3,32'd3,32'd2,32'd3,32'd2,32'd1,32'd6,32'd10,32'd19,32'd6,32'd10,32'd6,32'd19,32'd4,32'd2,32'd2,32'd2,32'd2,32'd23,32'd21,32'd3,32'd20,32'd3,32'd4,32'd7,32'd3,32'd9,32'd2,32'd9,32'd9,32'd6,32'd9,32'd2,32'd8,32'd3,32'd3,32'd6,32'd4,32'd5,32'd4,32'd14,32'd2,32'd5,32'd14,32'd13,32'd5,32'd3,32'd2,32'd2,32'd8,32'd4,32'd4,32'd3,32'd19,32'd3,32'd4,32'd3,32'd9,32'd4,32'd10,32'd18,32'd18,32'd3,32'd2,32'd1,32'd1,32'd9,32'd7,32'd10,32'd2,32'd2,32'd9,32'd4,32'd2,32'd3,32'd2,32'd9,32'd9,32'd13,32'd13,32'd7,32'd9,32'd3,32'd3,32'd1,32'd5,32'd6,32'd5,32'd6,32'd11,32'd2,32'd2,32'd3,32'd1,32'd1,32'd6,32'd9,32'd6,32'd9,32'd1,32'd1,32'd9,32'd4,32'd3,32'd16,32'd8,32'd6,32'd3,32'd4,32'd1,32'd9,32'd1,32'd2,32'd2,32'd18,32'd22,32'd22,32'd24,32'd24,32'd17,32'd6,32'd2,32'd2,32'd6,32'd6,32'd8,32'd1,32'd1,32'd2,32'd9,32'd2,32'd6,32'd6,32'd2,32'd6,32'd4,32'd6,32'd8,32'd3,32'd14,32'd8,32'd7,32'd9,32'd11,32'd11,32'd5,32'd7,32'd2,32'd4,32'd2,32'd16,32'd22,32'd22,32'd7,32'd8,32'd10,32'd3,32'd5,32'd3,32'd6,32'd2,32'd4,32'd4,32'd6,32'd6,32'd10,32'd2,32'd13,32'd1,32'd14,32'd18,32'd6,32'd3,32'd4,32'd1,32'd6,32'd6,32'd5,32'd24,32'd6,32'd1,32'd3,32'd10,32'd2,32'd2,32'd9,32'd9,32'd3,32'd3,32'd6,32'd9,32'd9,32'd3,32'd10,32'd10,32'd15,32'd1,32'd1,32'd1,32'd2,32'd2,32'd5,32'd5,32'd1,32'd6,32'd9,32'd9,32'd4,32'd9,32'd3,32'd6,32'd4,32'd6,32'd3,32'd4,32'd9,32'd9,32'd9,32'd9,32'd3,32'd5,32'd7,32'd5,32'd2,32'd2,32'd3,32'd4,32'd7,32'd1,32'd20,32'd6,32'd1,32'd2,32'd6,32'd2,32'd3,32'd7,32'd4,32'd23,32'd13,32'd13,32'd3,32'd2,32'd5,32'd6,32'd3,32'd3,32'd11,32'd1,32'd7,32'd9,32'd9,32'd1,32'd9,32'd11,32'd9,32'd19,32'd13,32'd13,32'd10,32'd10,32'd4,32'd6,32'd15,32'd15,32'd15,32'd2,32'd3,32'd6,32'd10,32'd7,32'd3,32'd3,32'd6,32'd2,32'd9,32'd13,32'd11,32'd9,32'd10,32'd10,32'd6,32'd3,32'd5,32'd5,32'd3,32'd4,32'd7,32'd2,32'd3,32'd5,32'd3,32'd8,32'd19,32'd2,32'd3,32'd7,32'd3}
`define RECTANGLE2_WEIGHTS {32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd256,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd384,32'd256,32'd384,32'd256,32'd256,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd256,32'd384,32'd384,32'd384,32'd384,32'd384,32'd256,32'd256,32'd256,32'd256,32'd256,32'd384,32'd384,32'd384,32'd384}
`define RECTANGLE3_XS {32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd3,32'd18,32'd0,32'd0,32'd11,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd13,32'd4,32'd16,32'd7,32'd3,32'd6,32'd15,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd6,32'd12,32'd10,32'd11,32'd0,32'd7,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd14,32'd7,32'd12,32'd0,32'd12,32'd0,32'd0,32'd3,32'd19,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd5,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd8,32'd10,32'd0,32'd0,32'd7,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd10,32'd7,32'd0,32'd0,32'd5,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd8,32'd4,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd8,32'd0,32'd13,32'd0,32'd0,32'd12,32'd0,32'd11,32'd10,32'd0,32'd2,32'd0,32'd0,32'd9,32'd11,32'd5,32'd15,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd14,32'd6,32'd0,32'd9,32'd12,32'd0,32'd13,32'd3,32'd18,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd4,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd12,32'd10,32'd3,32'd13,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd6,32'd0,32'd0,32'd11,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd1,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd5,32'd9,32'd12,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd7,32'd15,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd9,32'd7,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd2,32'd20,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd20,32'd0,32'd0,32'd12,32'd11,32'd0,32'd0,32'd3,32'd19,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd7,32'd14,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd12,32'd13,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd16,32'd9,32'd12,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd1,32'd11,32'd0,32'd0,32'd11,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd9,32'd3,32'd0,32'd0,32'd0,32'd0,32'd19,32'd0,32'd19,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd3,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd10,32'd6,32'd14,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd19,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd12,32'd7,32'd12,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd9,32'd0,32'd0,32'd5,32'd11,32'd11,32'd12,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd11,32'd6,32'd11,32'd0,32'd11,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd15,32'd0,32'd0,32'd0,32'd4,32'd9,32'd13,32'd12,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd12,32'd7,32'd11,32'd0,32'd5,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd12,32'd5,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd17,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd7,32'd15,32'd12,32'd0,32'd12,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd11,32'd3,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd7,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd14,32'd0,32'd6,32'd12,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd10,32'd0,32'd0,32'd0,32'd1,32'd0,32'd0,32'd12,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd7,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd5,32'd0,32'd9,32'd0,32'd6,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd1,32'd6,32'd12,32'd0,32'd0,32'd11,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd4,32'd15,32'd0,32'd0,32'd0,32'd17,32'd7,32'd2,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd4,32'd0,32'd0,32'd16,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd12,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd7,32'd0,32'd12,32'd10,32'd0,32'd0,32'd0,32'd0,32'd9,32'd11,32'd5,32'd15,32'd0,32'd15,32'd0,32'd0,32'd10,32'd10,32'd0,32'd0,32'd7,32'd0,32'd11,32'd10,32'd11,32'd7,32'd11,32'd0,32'd5,32'd14,32'd12,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd14,32'd4,32'd17,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd1,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd14,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd5,32'd15,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd10,32'd4,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd11,32'd0,32'd0,32'd0,32'd0,32'd7,32'd14,32'd0,32'd0,32'd4,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd5,32'd3,32'd10,32'd8,32'd11,32'd16,32'd10,32'd6,32'd0,32'd11,32'd11,32'd9,32'd0,32'd10,32'd0,32'd9,32'd0,32'd9,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd6,32'd9,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd10,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd11,32'd9,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd12,32'd5,32'd11,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd12,32'd12,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd1,32'd0,32'd0,32'd0,32'd0,32'd7,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd6,32'd0,32'd8,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd1,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd4,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd7,32'd4,32'd17,32'd0,32'd0,32'd4,32'd8,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd16,32'd0,32'd16,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd10,32'd10,32'd0,32'd0,32'd7,32'd0,32'd0,32'd5,32'd0,32'd10,32'd0,32'd8,32'd0,32'd16,32'd0,32'd4,32'd10,32'd9,32'd0,32'd1,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd12,32'd8,32'd0,32'd0,32'd10,32'd11,32'd0,32'd6,32'd0,32'd0,32'd0,32'd1,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd12,32'd4,32'd16,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd17,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd7,32'd11,32'd0,32'd0,32'd0,32'd12,32'd7,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd20,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd5,32'd0,32'd0,32'd6,32'd14,32'd6,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd12,32'd0,32'd0,32'd7,32'd0,32'd0,32'd10,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd4,32'd16,32'd0,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd7,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd5,32'd0,32'd0,32'd5,32'd14,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd1,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd8,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd17,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd15,32'd0,32'd0,32'd3,32'd10,32'd10,32'd4,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd18,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd12,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd17,32'd0,32'd0,32'd0,32'd0,32'd0,32'd1,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd3,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd2,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd9,32'd12,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd11,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd11,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0}
`define RECTANGLE3_YS {32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd18,32'd18,32'd0,32'd0,32'd21,32'd18,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd17,32'd17,32'd14,32'd14,32'd10,32'd22,32'd8,32'd8,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd22,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd17,32'd17,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd13,32'd9,32'd10,32'd14,32'd0,32'd19,32'd19,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd20,32'd20,32'd0,32'd21,32'd0,32'd0,32'd15,32'd15,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd9,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd16,32'd11,32'd0,32'd0,32'd12,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd15,32'd15,32'd0,32'd0,32'd11,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd19,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd11,32'd9,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd13,32'd0,32'd8,32'd0,32'd0,32'd16,32'd0,32'd13,32'd13,32'd0,32'd11,32'd0,32'd0,32'd5,32'd5,32'd19,32'd19,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd14,32'd12,32'd0,32'd12,32'd12,32'd0,32'd12,32'd11,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd9,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd6,32'd6,32'd7,32'd19,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd12,32'd0,32'd0,32'd15,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd17,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd13,32'd12,32'd12,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd12,32'd12,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd11,32'd11,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd14,32'd14,32'd0,32'd0,32'd20,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd14,32'd0,32'd0,32'd16,32'd15,32'd0,32'd0,32'd13,32'd13,32'd0,32'd0,32'd0,32'd0,32'd22,32'd0,32'd15,32'd15,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd16,32'd14,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd18,32'd18,32'd16,32'd16,32'd0,32'd20,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd14,32'd0,32'd0,32'd10,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd17,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd21,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd13,32'd14,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd5,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd21,32'd19,32'd19,32'd18,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd7,32'd16,32'd15,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd4,32'd0,32'd0,32'd12,32'd11,32'd11,32'd15,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd11,32'd20,32'd11,32'd0,32'd11,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd17,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd9,32'd12,32'd12,32'd14,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd12,32'd12,32'd12,32'd0,32'd17,32'd0,32'd18,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd2,32'd11,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd15,32'd15,32'd12,32'd0,32'd21,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd16,32'd0,32'd13,32'd13,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd16,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd9,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd16,32'd16,32'd0,32'd9,32'd10,32'd0,32'd0,32'd0,32'd18,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd21,32'd21,32'd0,32'd0,32'd0,32'd21,32'd0,32'd0,32'd11,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd9,32'd0,32'd0,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd9,32'd0,32'd19,32'd0,32'd9,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd9,32'd9,32'd0,32'd0,32'd12,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd21,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd18,32'd0,32'd6,32'd18,32'd0,32'd0,32'd0,32'd6,32'd15,32'd12,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd18,32'd0,32'd0,32'd18,32'd0,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd9,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd11,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd11,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd8,32'd0,32'd5,32'd10,32'd0,32'd0,32'd0,32'd0,32'd15,32'd15,32'd14,32'd14,32'd0,32'd14,32'd0,32'd0,32'd9,32'd10,32'd0,32'd0,32'd16,32'd0,32'd16,32'd16,32'd15,32'd9,32'd20,32'd0,32'd20,32'd20,32'd16,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd20,32'd0,32'd8,32'd7,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd21,32'd0,32'd0,32'd18,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd7,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd16,32'd17,32'd19,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd16,32'd14,32'd16,32'd0,32'd0,32'd0,32'd0,32'd18,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd19,32'd0,32'd0,32'd0,32'd0,32'd14,32'd14,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd20,32'd12,32'd15,32'd21,32'd13,32'd19,32'd12,32'd15,32'd0,32'd17,32'd13,32'd13,32'd0,32'd15,32'd0,32'd13,32'd0,32'd13,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd11,32'd11,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd18,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd4,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd22,32'd21,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd19,32'd9,32'd9,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd12,32'd11,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd7,32'd0,32'd2,32'd20,32'd20,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd16,32'd0,32'd0,32'd0,32'd14,32'd0,32'd14,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd13,32'd17,32'd17,32'd0,32'd0,32'd6,32'd7,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd16,32'd16,32'd0,32'd16,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd12,32'd12,32'd0,32'd0,32'd16,32'd0,32'd0,32'd13,32'd0,32'd12,32'd0,32'd16,32'd0,32'd17,32'd0,32'd9,32'd10,32'd10,32'd0,32'd19,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd9,32'd7,32'd0,32'd0,32'd15,32'd15,32'd0,32'd15,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd11,32'd15,32'd15,32'd0,32'd0,32'd0,32'd5,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd9,32'd9,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd9,32'd0,32'd0,32'd19,32'd19,32'd8,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd20,32'd20,32'd0,32'd14,32'd19,32'd0,32'd0,32'd15,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd18,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd17,32'd17,32'd0,32'd17,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd17,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd8,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd14,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd18,32'd18,32'd0,32'd3,32'd5,32'd5,32'd0,32'd0,32'd0,32'd0,32'd15,32'd8,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd13,32'd0,32'd0,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd7,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd18,32'd18,32'd0,32'd0,32'd14,32'd14,32'd11,32'd9,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd19,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd11,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd19,32'd0,32'd0,32'd0,32'd0,32'd0,32'd17,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd18,32'd0,32'd0,32'd0,32'd16,32'd0,32'd0,32'd0,32'd0,32'd0,32'd20,32'd21,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd14,32'd14,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd13,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd11,32'd11,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd11,32'd0,32'd0,32'd0,32'd19,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd11,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd15,32'd0,32'd0,32'd0,32'd0,32'd0,32'd20,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0}
`define RECTANGLE3_WIDTHS {32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd3,32'd3,32'd0,32'd0,32'd11,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd5,32'd4,32'd4,32'd2,32'd9,32'd3,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd9,32'd6,32'd4,32'd6,32'd0,32'd4,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd5,32'd5,32'd5,32'd0,32'd6,32'd0,32'd0,32'd2,32'd2,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd8,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd4,32'd6,32'd0,32'd0,32'd5,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd7,32'd7,32'd0,32'd0,32'd4,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd6,32'd9,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd5,32'd0,32'd5,32'd0,32'd0,32'd5,32'd0,32'd8,32'd4,32'd0,32'd10,32'd0,32'd0,32'd4,32'd4,32'd4,32'd4,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd6,32'd0,32'd2,32'd6,32'd0,32'd2,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd9,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd5,32'd3,32'd3,32'd5,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd9,32'd0,32'd0,32'd9,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd7,32'd3,32'd3,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd2,32'd2,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd8,32'd8,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd2,32'd2,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd2,32'd0,32'd0,32'd5,32'd2,32'd0,32'd0,32'd2,32'd2,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd3,32'd3,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd5,32'd4,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd3,32'd3,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd11,32'd0,32'd0,32'd6,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd2,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd9,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd6,32'd4,32'd4,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd4,32'd5,32'd2,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd9,32'd0,32'd0,32'd9,32'd2,32'd2,32'd2,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd2,32'd5,32'd2,32'd0,32'd2,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd0,32'd0,32'd0,32'd10,32'd2,32'd2,32'd9,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd5,32'd7,32'd5,32'd0,32'd4,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd12,32'd8,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd2,32'd2,32'd9,32'd0,32'd10,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd10,32'd10,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd3,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd7,32'd5,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd12,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd6,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd7,32'd0,32'd6,32'd0,32'd7,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd6,32'd6,32'd0,32'd0,32'd11,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd3,32'd4,32'd0,32'd0,32'd0,32'd3,32'd4,32'd11,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd4,32'd0,32'd0,32'd4,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd7,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd10,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd6,32'd0,32'd12,32'd4,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd4,32'd4,32'd0,32'd4,32'd0,32'd0,32'd8,32'd4,32'd0,32'd0,32'd3,32'd0,32'd3,32'd3,32'd2,32'd6,32'd5,32'd0,32'd5,32'd5,32'd4,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd3,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd3,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd3,32'd9,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd6,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd4,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd5,32'd10,32'd10,32'd6,32'd11,32'd4,32'd9,32'd6,32'd0,32'd3,32'd4,32'd4,32'd0,32'd2,32'd0,32'd4,32'd0,32'd4,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd9,32'd3,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd10,32'd7,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd7,32'd7,32'd6,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd6,32'd6,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd12,32'd0,32'd12,32'd5,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd3,32'd0,32'd7,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd10,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd7,32'd3,32'd3,32'd0,32'd0,32'd3,32'd4,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd0,32'd4,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd4,32'd4,32'd0,32'd0,32'd6,32'd0,32'd0,32'd7,32'd0,32'd4,32'd0,32'd4,32'd0,32'd4,32'd0,32'd8,32'd5,32'd5,32'd0,32'd11,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd6,32'd4,32'd0,32'd0,32'd8,32'd3,32'd0,32'd8,32'd0,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd6,32'd4,32'd4,32'd0,32'd0,32'd0,32'd12,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd7,32'd9,32'd0,32'd0,32'd0,32'd12,32'd6,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd8,32'd0,32'd0,32'd4,32'd4,32'd6,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd5,32'd0,32'd12,32'd4,32'd0,32'd0,32'd2,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd0,32'd4,32'd0,32'd0,32'd0,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd5,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd8,32'd0,32'd12,32'd5,32'd5,32'd0,32'd0,32'd0,32'd0,32'd9,32'd12,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd5,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd3,32'd4,32'd9,32'd8,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd3,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd9,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd12,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd11,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd12,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd5,32'd7,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd4,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0}
`define RECTANGLE3_HEIGHTS {32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd6,32'd6,32'd0,32'd0,32'd3,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd6,32'd6,32'd10,32'd2,32'd7,32'd7,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd5,32'd5,32'd5,32'd3,32'd0,32'd5,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd4,32'd4,32'd0,32'd3,32'd0,32'd0,32'd9,32'd9,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd4,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd5,32'd4,32'd0,32'd0,32'd6,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd7,32'd7,32'd0,32'd0,32'd5,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd10,32'd2,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd4,32'd0,32'd0,32'd4,32'd0,32'd4,32'd8,32'd0,32'd3,32'd0,32'd0,32'd5,32'd5,32'd5,32'd5,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd10,32'd3,32'd0,32'd9,32'd3,32'd0,32'd9,32'd10,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd2,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd6,32'd6,32'd6,32'd4,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd12,32'd0,32'd0,32'd2,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd4,32'd6,32'd6,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd11,32'd11,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd10,32'd10,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd10,32'd10,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd10,32'd0,32'd0,32'd7,32'd9,32'd0,32'd0,32'd11,32'd11,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd6,32'd6,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd5,32'd5,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd6,32'd6,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd2,32'd0,32'd0,32'd8,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd5,32'd9,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd5,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd3,32'd5,32'd5,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd6,32'd8,32'd9,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd4,32'd0,32'd0,32'd3,32'd10,32'd10,32'd9,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd10,32'd0,32'd10,32'd4,32'd10,32'd0,32'd10,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd2,32'd11,32'd11,32'd2,32'd0,32'd0,32'd11,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd4,32'd7,32'd12,32'd0,32'd7,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd2,32'd7,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd9,32'd9,32'd7,32'd0,32'd2,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd3,32'd3,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd6,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd3,32'd4,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd11,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd5,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd3,32'd0,32'd4,32'd0,32'd3,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd9,32'd9,32'd0,32'd0,32'd8,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd6,32'd5,32'd0,32'd0,32'd0,32'd6,32'd5,32'd7,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd5,32'd0,32'd0,32'd5,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd3,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd6,32'd0,32'd3,32'd8,32'd0,32'd0,32'd0,32'd0,32'd7,32'd7,32'd10,32'd10,32'd0,32'd10,32'd0,32'd0,32'd4,32'd9,32'd0,32'd0,32'd8,32'd0,32'd7,32'd7,32'd9,32'd3,32'd4,32'd0,32'd4,32'd4,32'd6,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd8,32'd7,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd7,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd7,32'd7,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd7,32'd2,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd4,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd4,32'd6,32'd9,32'd3,32'd4,32'd5,32'd3,32'd3,32'd0,32'd7,32'd5,32'd5,32'd0,32'd9,32'd0,32'd5,32'd0,32'd5,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd11,32'd11,32'd6,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd3,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd2,32'd3,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd3,32'd3,32'd4,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd6,32'd3,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd3,32'd0,32'd2,32'd4,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd10,32'd0,32'd5,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd2,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd7,32'd7,32'd7,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd8,32'd0,32'd8,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd8,32'd8,32'd0,32'd0,32'd5,32'd0,32'd0,32'd7,32'd0,32'd8,32'd0,32'd6,32'd0,32'd7,32'd0,32'd3,32'd5,32'd5,32'd0,32'd3,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd3,32'd5,32'd0,32'd0,32'd3,32'd7,32'd0,32'd3,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd6,32'd9,32'd9,32'd0,32'd0,32'd0,32'd5,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd4,32'd0,32'd0,32'd0,32'd3,32'd6,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd3,32'd0,32'd0,32'd5,32'd5,32'd3,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd4,32'd0,32'd2,32'd5,32'd0,32'd0,32'd9,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd4,32'd0,32'd0,32'd0,32'd0,32'd7,32'd7,32'd0,32'd7,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd8,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd2,32'd5,32'd5,32'd0,32'd0,32'd0,32'd0,32'd2,32'd8,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd0,32'd0,32'd10,32'd7,32'd11,32'd3,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd8,32'd6,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd4,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd2,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd2,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd9,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd2,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd2,32'd0,32'd0,32'd0,32'd8,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd5,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd6,32'd5,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd3,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd5,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd3,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd7,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd6,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0}
`define RECTANGLE3_WEIGHTS {32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd256,32'd256,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd256,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd256,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd256,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0}
`define FEATURE_THRESHOLD {32'd4294967293,32'd10,32'd0,32'd4294967294,32'd7,32'd3,32'd4294967291,32'd2,32'd0,32'd4294967295,32'd4294967294,32'd9,32'd2,32'd4294967289,32'd4,32'd4294967291,32'd14,32'd6,32'd0,32'd6,32'd4294967292,32'd4294967294,32'd0,32'd10,32'd3,32'd1,32'd4294967276,32'd4294967293,32'd4294967291,32'd5,32'd4294967287,32'd5,32'd4294967291,32'd6,32'd4294967292,32'd1,32'd4294967295,32'd3,32'd1,32'd4294967295,32'd1,32'd0,32'd4294967294,32'd3,32'd4294967293,32'd4294967289,32'd4294967289,32'd1,32'd18,32'd4294967266,32'd10,32'd2,32'd4294967291,32'd0,32'd2,32'd4,32'd4294967293,32'd4294967288,32'd2,32'd4294967292,32'd0,32'd0,32'd1,32'd1,32'd1,32'd2,32'd9,32'd2,32'd4294967282,32'd3,32'd0,32'd4294967283,32'd4294967266,32'd4294967286,32'd4294967294,32'd0,32'd4294967294,32'd4294967285,32'd1,32'd4,32'd4294967295,32'd3,32'd4,32'd4294967295,32'd4294967293,32'd1,32'd7,32'd4294967294,32'd5,32'd1,32'd2,32'd4,32'd4294967293,32'd3,32'd1,32'd4294967290,32'd4,32'd0,32'd2,32'd4294967288,32'd16,32'd4294967282,32'd4294967266,32'd36,32'd4294967294,32'd2,32'd1,32'd4294967292,32'd1,32'd4294967295,32'd4294967293,32'd4294967285,32'd4294967281,32'd4294967294,32'd4294967293,32'd3,32'd4294967291,32'd2,32'd4294967292,32'd4294967295,32'd2,32'd4294967281,32'd4294967282,32'd5,32'd14,32'd1,32'd4294967287,32'd1,32'd4294967294,32'd1,32'd4294967291,32'd4294967293,32'd1,32'd4294967286,32'd8,32'd4294967293,32'd3,32'd1,32'd4294967294,32'd1,32'd0,32'd6,32'd4294967293,32'd4294967285,32'd0,32'd6,32'd4294967294,32'd4294967289,32'd4294967295,32'd4294967294,32'd8,32'd54,32'd4294967285,32'd4294967292,32'd4294967291,32'd4294967292,32'd4294967291,32'd7,32'd2,32'd4294967294,32'd4294967293,32'd0,32'd0,32'd21,32'd2,32'd6,32'd4294967295,32'd1,32'd4294967295,32'd1,32'd4294967291,32'd4294967295,32'd4294967295,32'd4294967294,32'd4294967295,32'd0,32'd4294967293,32'd4294967292,32'd4294967295,32'd4294967293,32'd0,32'd4294967295,32'd20,32'd3,32'd6,32'd1,32'd7,32'd4294967294,32'd5,32'd2,32'd0,32'd6,32'd4294967286,32'd0,32'd2,32'd4294967295,32'd0,32'd3,32'd2,32'd4294967284,32'd0,32'd4,32'd4294967292,32'd1,32'd3,32'd6,32'd4294967293,32'd7,32'd2,32'd1,32'd7,32'd11,32'd11,32'd16,32'd4294967291,32'd1,32'd4294967274,32'd4294967288,32'd12,32'd1,32'd4294967292,32'd4294967287,32'd1,32'd25,32'd1,32'd1,32'd4294967295,32'd4294967292,32'd4294967295,32'd4294967294,32'd41,32'd4294967295,32'd4294967292,32'd4294967295,32'd4294967294,32'd4,32'd3,32'd2,32'd4,32'd8,32'd10,32'd6,32'd4294967287,32'd3,32'd5,32'd10,32'd4294967291,32'd11,32'd0,32'd4,32'd4294967294,32'd0,32'd7,32'd4294967293,32'd2,32'd0,32'd4294967295,32'd4294967291,32'd12,32'd4294967286,32'd9,32'd4294967285,32'd2,32'd10,32'd2,32'd11,32'd9,32'd4294967280,32'd4294967294,32'd4294967291,32'd1,32'd4294967295,32'd4294967293,32'd4294967266,32'd1,32'd3,32'd4294967293,32'd6,32'd3,32'd4294967292,32'd4294967295,32'd15,32'd4294967295,32'd0,32'd10,32'd5,32'd1,32'd0,32'd11,32'd20,32'd4294967292,32'd4294967292,32'd0,32'd0,32'd2,32'd4294967292,32'd4294967293,32'd0,32'd6,32'd4,32'd17,32'd4294967295,32'd4294967292,32'd2,32'd4294967290,32'd4294967294,32'd28,32'd47,32'd0,32'd4294967285,32'd4294967295,32'd1,32'd4294967294,32'd14,32'd2,32'd4,32'd3,32'd4294967295,32'd4294967293,32'd4,32'd1,32'd4294967293,32'd4294967289,32'd4294967295,32'd4294967293,32'd4294967293,32'd5,32'd4,32'd8,32'd4294967293,32'd5,32'd4294967292,32'd4,32'd6,32'd4294967294,32'd4294967287,32'd4294967292,32'd4,32'd4294967294,32'd1,32'd4294967286,32'd6,32'd1,32'd0,32'd4294967280,32'd5,32'd7,32'd4,32'd4294967294,32'd4294967287,32'd4294967293,32'd7,32'd4294967294,32'd4294967295,32'd7,32'd1,32'd4294967285,32'd4294967294,32'd4,32'd4,32'd4,32'd0,32'd4294967294,32'd4294967295,32'd4294967294,32'd4294967286,32'd4294967292,32'd8,32'd4294967285,32'd4294967280,32'd4294967295,32'd4294967294,32'd4294967295,32'd4294967294,32'd3,32'd0,32'd4294967291,32'd8,32'd6,32'd4294967293,32'd3,32'd4294967290,32'd4294967295,32'd6,32'd0,32'd0,32'd4294967292,32'd2,32'd4294967294,32'd1,32'd4294967294,32'd4294967294,32'd4294967292,32'd3,32'd4294967291,32'd4294967295,32'd1,32'd0,32'd19,32'd3,32'd4294967293,32'd4294967294,32'd4294967294,32'd10,32'd4294967292,32'd3,32'd0,32'd4294967295,32'd5,32'd4,32'd3,32'd14,32'd4294967289,32'd1,32'd9,32'd3,32'd6,32'd1,32'd4294967276,32'd4294967292,32'd0,32'd7,32'd1,32'd4,32'd4294967281,32'd4294967280,32'd4294967283,32'd4294967291,32'd4294967290,32'd7,32'd1,32'd9,32'd5,32'd4294967292,32'd30,32'd4294967280,32'd4294967292,32'd4294967291,32'd4294967281,32'd14,32'd1,32'd4294967295,32'd4294967292,32'd4,32'd10,32'd1,32'd4294967291,32'd12,32'd1,32'd5,32'd4294967294,32'd4294967291,32'd29,32'd1,32'd4294967293,32'd2,32'd3,32'd4294967294,32'd4294967287,32'd4294967294,32'd3,32'd2,32'd4294967295,32'd1,32'd4294967287,32'd0,32'd4294967295,32'd5,32'd4294967289,32'd4294967285,32'd38,32'd0,32'd4294967289,32'd4294967289,32'd5,32'd2,32'd4294967295,32'd1,32'd4294967292,32'd4294967293,32'd4294967295,32'd2,32'd4294967294,32'd2,32'd4294967294,32'd4294967294,32'd4294967285,32'd4294967294,32'd0,32'd3,32'd4294967292,32'd0,32'd1,32'd7,32'd19,32'd8,32'd4294967293,32'd3,32'd4,32'd3,32'd4294967294,32'd4294967290,32'd4294967293,32'd4294967289,32'd4294967286,32'd4294967293,32'd2,32'd14,32'd85,32'd4294967294,32'd0,32'd4294967293,32'd5,32'd0,32'd4294967295,32'd4,32'd4294967291,32'd4294967295,32'd0,32'd4294967295,32'd4294967294,32'd4294967284,32'd4,32'd4294967286,32'd4294967290,32'd4294967294,32'd4294967292,32'd1,32'd8,32'd4294967266,32'd37,32'd1,32'd1,32'd4294967280,32'd4294967267,32'd4294967294,32'd4294967294,32'd4294967290,32'd0,32'd2,32'd4294967294,32'd4294967290,32'd3,32'd4294967290,32'd6,32'd4294967293,32'd4294967293,32'd4294967293,32'd4294967294,32'd4294967294,32'd26,32'd0,32'd1,32'd4294967295,32'd2,32'd4294967287,32'd4294967288,32'd4294967295,32'd4294967290,32'd2,32'd4,32'd4,32'd4294967294,32'd12,32'd4294967294,32'd7,32'd7,32'd4294967295,32'd1,32'd4294967294,32'd3,32'd4294967293,32'd0,32'd5,32'd4294967295,32'd0,32'd4294967294,32'd4294967291,32'd4294967291,32'd4294967293,32'd2,32'd4294967290,32'd4294967289,32'd2,32'd4294967288,32'd4294967291,32'd1,32'd4294967286,32'd4294967287,32'd0,32'd4294967292,32'd4294967292,32'd5,32'd4,32'd4294967288,32'd4294967287,32'd5,32'd2,32'd4294967295,32'd0,32'd3,32'd5,32'd0,32'd4294967291,32'd4294967290,32'd5,32'd4,32'd3,32'd13,32'd3,32'd4294967294,32'd4294967292,32'd9,32'd4294967288,32'd4,32'd2,32'd11,32'd4294967283,32'd5,32'd3,32'd3,32'd4294967289,32'd1,32'd7,32'd5,32'd4294967293,32'd0,32'd20,32'd4294967259,32'd5,32'd4294967283,32'd4294967292,32'd4294967294,32'd4294967294,32'd2,32'd2,32'd4294967292,32'd0,32'd4294967293,32'd4294967292,32'd14,32'd1,32'd23,32'd4294967278,32'd1,32'd4294967294,32'd1,32'd4294967291,32'd4294967292,32'd66,32'd4294967291,32'd9,32'd2,32'd4294967295,32'd4294967284,32'd4294967278,32'd2,32'd0,32'd12,32'd4294967292,32'd1,32'd2,32'd0,32'd4294967291,32'd4294967287,32'd4294967290,32'd1,32'd5,32'd8,32'd4294967287,32'd5,32'd4294967287,32'd26,32'd4294967255,32'd4294967294,32'd3,32'd13,32'd4294967289,32'd4294967295,32'd14,32'd4294967293,32'd4294967294,32'd1,32'd11,32'd4294967295,32'd4,32'd4294967295,32'd5,32'd0,32'd1,32'd4294967295,32'd1,32'd4294967295,32'd11,32'd1,32'd4294967293,32'd4,32'd1,32'd4294967294,32'd4294967289,32'd2,32'd3,32'd4294967294,32'd7,32'd9,32'd4294967284,32'd2,32'd6,32'd4294967290,32'd2,32'd4294967293,32'd4294967287,32'd4294967295,32'd4294967289,32'd4294967294,32'd4294967294,32'd5,32'd4294967284,32'd4294967290,32'd6,32'd0,32'd4294967294,32'd68,32'd9,32'd2,32'd4294967295,32'd4,32'd4294967291,32'd4294967294,32'd4294967294,32'd4294967290,32'd2,32'd5,32'd4,32'd4294967295,32'd10,32'd4294967295,32'd4294967295,32'd4,32'd4294967289,32'd4294967295,32'd4294967294,32'd4294967294,32'd4294967295,32'd4294967287,32'd1,32'd4294967291,32'd2,32'd3,32'd4294967292,32'd4,32'd4294967295,32'd4294967292,32'd1,32'd4,32'd4294967256,32'd4294967287,32'd6,32'd1,32'd4294967292,32'd0,32'd19,32'd8,32'd5,32'd11,32'd13,32'd4294967291,32'd4294967294,32'd5,32'd0,32'd4294967288,32'd4294967293,32'd1,32'd4294967294,32'd7,32'd4294967289,32'd1,32'd7,32'd4294967290,32'd0,32'd1,32'd4294967294,32'd4294967293,32'd3,32'd2,32'd4294967295,32'd4294967295,32'd2,32'd4,32'd24,32'd6,32'd2,32'd4294967293,32'd4,32'd4,32'd4294967288,32'd4294967289,32'd0,32'd4294967292,32'd4294967294,32'd0,32'd4294967295,32'd3,32'd0,32'd5,32'd0,32'd13,32'd4294967292,32'd6,32'd4294967295,32'd0,32'd2,32'd0,32'd9,32'd4294967294,32'd4294967292,32'd2,32'd8,32'd6,32'd4294967291,32'd4294967287,32'd5,32'd4294967292,32'd3,32'd4,32'd0,32'd4294967281,32'd2,32'd4294967292,32'd4294967294,32'd15,32'd4294967283,32'd4294967294,32'd3,32'd7,32'd4294967288,32'd2,32'd2,32'd0,32'd4294967293,32'd4294967295,32'd4294967291,32'd5,32'd1,32'd4294967288,32'd4294967294,32'd4294967286,32'd4294967281,32'd4294967274,32'd4294967294,32'd3,32'd6,32'd4294967294,32'd4294967295,32'd4294967294,32'd3,32'd0,32'd2,32'd25,32'd6,32'd2,32'd6,32'd4294967295,32'd0,32'd4,32'd4294967288,32'd8,32'd6,32'd6,32'd4294967291,32'd5,32'd4294967288,32'd4294967295,32'd4294967295,32'd2,32'd13,32'd4294967287,32'd0,32'd4294967288,32'd1,32'd4,32'd6,32'd4294967280,32'd4294967295,32'd4294967294,32'd4294967291,32'd4294967294,32'd4294967294,32'd9,32'd7,32'd4294967295,32'd4294967294,32'd4294967281,32'd4294967290,32'd0,32'd4294967289,32'd4294967295,32'd4294967294,32'd9,32'd4294967294,32'd1,32'd4294967294,32'd13,32'd4294967290,32'd4294967295,32'd4294967290,32'd0,32'd4294967291,32'd6,32'd4294967290,32'd4294967294,32'd4294967295,32'd2,32'd4294967295,32'd2,32'd4294967295,32'd4294967291,32'd53,32'd3,32'd4294967294,32'd4,32'd3,32'd1,32'd4294967295,32'd4294967295,32'd2,32'd4294967294,32'd4294967294,32'd0,32'd4294967294,32'd2,32'd2,32'd2,32'd0,32'd4294967289,32'd4294967295,32'd4294967294,32'd0,32'd4294967292,32'd4294967292,32'd1,32'd6,32'd4294967294,32'd10,32'd41,32'd4294967289,32'd1,32'd4294967290,32'd4294967288,32'd4294967293,32'd4294967295,32'd2,32'd3,32'd1,32'd4294967293,32'd4294967293,32'd4294967290,32'd2,32'd4294967295,32'd4294967294,32'd4294967294,32'd4294967295,32'd0,32'd9,32'd4294967292,32'd2,32'd4294967293,32'd4294967290,32'd4294967293,32'd4294967293,32'd4294967291,32'd2,32'd4294967295,32'd4294967291,32'd4294967289,32'd4294967293,32'd4,32'd4294967295,32'd1,32'd10,32'd4294967295,32'd11,32'd4294967293,32'd0,32'd0,32'd3,32'd4294967282,32'd7,32'd1,32'd4294967294,32'd0,32'd4294967293,32'd1,32'd4294967294,32'd4294967286,32'd3,32'd8,32'd4294967287,32'd4294967286,32'd5,32'd1,32'd1,32'd4,32'd2,32'd4294967280,32'd4294967294,32'd4294967294,32'd4294967294,32'd4294967283,32'd3,32'd4294967294,32'd4294967292,32'd2,32'd4294967295,32'd4294967291,32'd3,32'd2,32'd3,32'd3,32'd4294967288,32'd4294967294,32'd13,32'd5,32'd4294967279,32'd4294967295,32'd4294967285,32'd0,32'd33,32'd6,32'd4294967292,32'd5,32'd4294967286,32'd4294967292,32'd4294967291,32'd0,32'd4294967295,32'd4294967287,32'd0,32'd4294967294,32'd1,32'd1,32'd4294967295,32'd11,32'd4294967291,32'd4294967289,32'd8,32'd0,32'd4294967294,32'd4294967282,32'd4294967271,32'd4294967292,32'd1,32'd4294967293,32'd4294967295,32'd4,32'd4294967285,32'd0,32'd2,32'd2,32'd4294967289,32'd4294967294,32'd4294967295,32'd0,32'd4294967285,32'd4294967278,32'd4294967293,32'd4294967295,32'd4294967278,32'd0,32'd4294967294,32'd2,32'd5,32'd5,32'd6,32'd3,32'd2,32'd4294967291,32'd14,32'd4294967293,32'd4294967289,32'd4294967293,32'd6,32'd4,32'd4,32'd0,32'd1,32'd8,32'd4,32'd1,32'd4294967288,32'd4294967290,32'd2,32'd4294967289,32'd4294967290,32'd4,32'd1,32'd3,32'd10,32'd4294967293,32'd4294967255,32'd7,32'd22,32'd2,32'd7,32'd4294967295,32'd1,32'd0,32'd0,32'd2,32'd4294967290,32'd4294967295,32'd4294967295,32'd4294967294,32'd4294967295,32'd7,32'd0,32'd0,32'd4,32'd1,32'd44,32'd1,32'd4294967293,32'd3,32'd4294967289,32'd0,32'd4294967291,32'd11,32'd2,32'd4,32'd4294967293,32'd2,32'd10,32'd4294967293,32'd1,32'd0,32'd0,32'd4294967293,32'd1,32'd4294967295,32'd4294967295,32'd1,32'd4294967295,32'd24,32'd5,32'd4294967292,32'd6,32'd2,32'd4294967293,32'd6,32'd4294967282,32'd4294967295,32'd2,32'd1,32'd6,32'd4294967287,32'd3,32'd4294967295,32'd3,32'd4294967291,32'd4294967294,32'd4294967293,32'd9,32'd4294967289,32'd1,32'd3,32'd4,32'd2,32'd1,32'd2,32'd4294967294,32'd4294967295,32'd4294967295,32'd4294967293,32'd4,32'd2,32'd14,32'd4294967295,32'd4294967291,32'd8,32'd1,32'd8,32'd5,32'd7,32'd9,32'd4294967294,32'd28,32'd4294967291,32'd4294967295,32'd4294967293,32'd3,32'd0,32'd4294967289,32'd4294967294,32'd4294967286,32'd4294967294,32'd17,32'd4294967295,32'd0,32'd5,32'd4294967293,32'd4294967292,32'd11,32'd1,32'd0,32'd4294967291,32'd1,32'd8,32'd4,32'd4294967291,32'd4294967294,32'd4294967294,32'd4,32'd4294967295,32'd4294967294,32'd1,32'd2,32'd12,32'd1,32'd4294967295,32'd4,32'd0,32'd2,32'd4294967291,32'd4294967291,32'd4294967291,32'd6,32'd7,32'd4294967290,32'd20,32'd25,32'd0,32'd9,32'd14,32'd0,32'd1,32'd4294967292,32'd4294967292,32'd6,32'd4294967294,32'd0,32'd6,32'd4294967285,32'd0,32'd4294967295,32'd4294967295,32'd0,32'd6,32'd1,32'd4294967291,32'd0,32'd3,32'd4294967293,32'd4,32'd4294967295,32'd5,32'd1,32'd2,32'd2,32'd5,32'd2,32'd2,32'd4294967280,32'd6,32'd4294967286,32'd3,32'd0,32'd2,32'd4294967290,32'd4294967295,32'd4294967292,32'd4294967293,32'd4294967290,32'd4294967294,32'd4294967293,32'd4294967290,32'd4,32'd9,32'd4294967295,32'd4294967293,32'd4294967293,32'd4294967284,32'd4294967291,32'd4294967295,32'd2,32'd3,32'd4294967295,32'd4,32'd0,32'd3,32'd1,32'd9,32'd4294967281,32'd4294967281,32'd4294967290,32'd4294967291,32'd13,32'd4294967292,32'd0,32'd5,32'd7,32'd4294967290,32'd4294967294,32'd4294967292,32'd1,32'd4294967287,32'd4294967290,32'd4294967294,32'd3,32'd3,32'd4294967289,32'd3,32'd3,32'd1,32'd4294967295,32'd4294967295,32'd4294967290,32'd0,32'd3,32'd4294967294,32'd4294967286,32'd2,32'd2,32'd4294967294,32'd4294967292,32'd12,32'd1,32'd1,32'd4294967292,32'd4294967295,32'd4294967292,32'd0,32'd0,32'd4294967294,32'd6,32'd4294967295,32'd4294967290,32'd2,32'd4294967293,32'd4294967293,32'd2,32'd4294967291,32'd4294967291,32'd4,32'd4294967290,32'd5,32'd0,32'd4294967294,32'd1,32'd3,32'd4,32'd1,32'd16,32'd4294967292,32'd6,32'd4294967292,32'd8,32'd1,32'd0,32'd0,32'd4294967292,32'd3,32'd2,32'd4294967295,32'd6,32'd4294967295,32'd13,32'd0,32'd7,32'd4294967293,32'd4294967288,32'd4294967289,32'd11,32'd11,32'd3,32'd3,32'd4,32'd4294967294,32'd14,32'd4294967290,32'd22,32'd12,32'd1,32'd3,32'd6,32'd6,32'd4294967292,32'd4294967293,32'd4294967295,32'd4,32'd1,32'd4294967290,32'd0,32'd4294967295,32'd4294967293,32'd2,32'd0,32'd0,32'd4294967295,32'd4294967293,32'd4294967286,32'd13,32'd5,32'd4294967293,32'd4294967287,32'd4294967291,32'd2,32'd4294967292,32'd4294967291,32'd4294967279,32'd4294967291,32'd3,32'd5,32'd4294967281,32'd1,32'd29,32'd4294967289,32'd4294967293,32'd15,32'd22,32'd1,32'd4294967291,32'd1,32'd9,32'd4294967294,32'd4294967294,32'd4294967295,32'd4,32'd2,32'd4294967293,32'd4294967292,32'd8,32'd3,32'd2,32'd4294967294,32'd1,32'd23,32'd4294967287,32'd1,32'd15,32'd4294967281,32'd4,32'd4294967294,32'd4294967286,32'd5,32'd4294967294,32'd3,32'd0,32'd6,32'd2,32'd1,32'd4,32'd4294967291,32'd4294967294,32'd4294967293,32'd4294967295,32'd4294967292,32'd4,32'd4294967294,32'd4294967293,32'd4294967291,32'd0,32'd4,32'd12,32'd3,32'd4294967292,32'd4294967294,32'd4294967295,32'd9,32'd20,32'd4294967293,32'd4294967294,32'd4294967293,32'd0,32'd4294967295,32'd4294967288,32'd4294967293,32'd5,32'd4,32'd4294967294,32'd4294967294,32'd4294967293,32'd1,32'd4294967295,32'd4294967293,32'd4294967290,32'd4294967288,32'd4294967294,32'd4294967293,32'd4294967292,32'd3,32'd4294967293,32'd4294967292,32'd0,32'd3,32'd12,32'd4294967289,32'd2,32'd1,32'd0,32'd0,32'd0,32'd4294967294,32'd4,32'd0,32'd4294967295,32'd4294967295,32'd2,32'd18,32'd2,32'd5,32'd12,32'd21,32'd1,32'd4294967291,32'd4294967293,32'd4294967292,32'd4294967295,32'd4294967295,32'd4294967293,32'd2,32'd4294967288,32'd12,32'd4294967295,32'd0,32'd4294967293,32'd2,32'd7,32'd2,32'd4294967293,32'd4294967293,32'd4294967294,32'd3,32'd7,32'd4294967278,32'd3,32'd4294967292,32'd7,32'd4294967290,32'd0,32'd4294967281,32'd4294967287,32'd4294967288,32'd1,32'd4,32'd10,32'd5,32'd6,32'd3,32'd4294967291,32'd3,32'd4294967295,32'd4294967287,32'd4294967293,32'd4294967294,32'd10,32'd4294967293,32'd3,32'd5,32'd4294967293,32'd6,32'd3,32'd4294967294,32'd4294967294,32'd1,32'd4,32'd0,32'd14,32'd0,32'd4294967291,32'd4294967284,32'd4294967283,32'd4294967294,32'd4294967295,32'd2,32'd0,32'd4294967294,32'd2,32'd3,32'd11,32'd4294967290,32'd2,32'd4294967292,32'd4,32'd4294967289,32'd1,32'd3,32'd3,32'd4294967292,32'd6,32'd1,32'd4,32'd1,32'd4,32'd0,32'd4294967292,32'd3,32'd4294967295,32'd4,32'd4294967294,32'd3,32'd4294967294,32'd3,32'd4294967295,32'd1,32'd4294967292,32'd4294967284,32'd10,32'd1,32'd4294967285,32'd4294967293,32'd5,32'd3,32'd7,32'd4294967290,32'd2,32'd1,32'd8,32'd1,32'd3,32'd4294967291,32'd1,32'd6,32'd12,32'd2,32'd1,32'd1,32'd4294967290,32'd2,32'd4294967294,32'd3,32'd4294967295,32'd4294967295,32'd4294967294,32'd3,32'd1,32'd0,32'd5,32'd12,32'd4294967280,32'd7,32'd0,32'd4294967295,32'd4294967295,32'd4,32'd4294967289,32'd4294967291,32'd4294967258,32'd4294967292,32'd4294967294,32'd4294967289,32'd1,32'd0,32'd7,32'd4294967293,32'd4294967294,32'd4294967293,32'd4294967291,32'd4294967295,32'd7,32'd0,32'd4294967293,32'd1,32'd1,32'd7,32'd2,32'd28,32'd4294967286,32'd4294967291,32'd6,32'd1,32'd42,32'd4294967294,32'd3,32'd11,32'd0,32'd14,32'd29,32'd4294967294,32'd1,32'd7,32'd4,32'd4294967294,32'd4294967293,32'd4294967293,32'd4294967294,32'd12,32'd0,32'd4294967294,32'd4294967294,32'd4294967294,32'd1,32'd54,32'd4294967293,32'd5,32'd9,32'd0,32'd6,32'd6,32'd14,32'd0,32'd4294967293,32'd4294967293,32'd3,32'd4294967293,32'd5,32'd4,32'd4294967293,32'd8,32'd4294967293,32'd4294967283,32'd0,32'd4294967294,32'd4294967290,32'd4294967286,32'd24,32'd3,32'd4294967293,32'd4294967290,32'd3,32'd2,32'd0,32'd4294967293,32'd0,32'd4294967292,32'd4294967290,32'd17,32'd4294967287,32'd2,32'd4294967286,32'd3,32'd8,32'd4294967292,32'd3,32'd5,32'd2,32'd27,32'd4294967295,32'd4294967289,32'd0,32'd4294967294,32'd9,32'd4294967295,32'd4294967294,32'd4294967293,32'd1,32'd2,32'd4294967282,32'd0,32'd4294967292,32'd1,32'd4294967285,32'd4294967294,32'd2,32'd4294967292,32'd4294967295,32'd4294967294,32'd4294967292,32'd0,32'd4294967295,32'd4294967295,32'd1,32'd4294967294,32'd4294967291,32'd4294967293,32'd3,32'd4294967291,32'd4294967284,32'd4294967288,32'd8,32'd1,32'd4294967292,32'd2,32'd4294967292,32'd4,32'd4294967295,32'd4294967292,32'd0,32'd0,32'd4294967293,32'd2,32'd0,32'd4294967293,32'd3,32'd4294967293,32'd4294967294,32'd4294967290,32'd4294967293,32'd2,32'd58,32'd4294967294,32'd4294967293,32'd2,32'd3,32'd4294967291,32'd3,32'd1,32'd3,32'd0,32'd0,32'd4294967288,32'd1,32'd1,32'd4294967279,32'd1,32'd3,32'd4294967291,32'd4294967291,32'd4294967294,32'd6,32'd5,32'd1,32'd4294967284,32'd2,32'd7,32'd6,32'd4294967291,32'd4294967290,32'd1,32'd4294967292,32'd3,32'd5,32'd4294967294,32'd13,32'd2,32'd4294967293,32'd4294967290,32'd2,32'd5,32'd4294967292,32'd1,32'd4294967293,32'd7,32'd10,32'd1,32'd0,32'd4,32'd4294967295,32'd4294967289,32'd4294967292,32'd2,32'd7,32'd13,32'd4294967295,32'd4294967295,32'd1,32'd1,32'd4294967293,32'd2,32'd5,32'd1,32'd4294967293,32'd1,32'd2,32'd4294967295,32'd4294967293,32'd4294967291,32'd7,32'd4294967292,32'd1,32'd4294967291,32'd4294967295,32'd4294967295,32'd2,32'd4294967282,32'd4294967290,32'd4294967293,32'd4294967287,32'd4294967293,32'd3,32'd4294967295,32'd1,32'd4294967294,32'd4294967291,32'd4294967293,32'd4294967295,32'd4294967295,32'd1,32'd4,32'd2,32'd1,32'd4294967293,32'd3,32'd4294967292,32'd4,32'd0,32'd0,32'd1,32'd10,32'd3,32'd1,32'd1,32'd3,32'd4294967292,32'd3,32'd4294967295,32'd5,32'd14,32'd2,32'd0,32'd3,32'd7,32'd4294967295,32'd4294967291,32'd3,32'd4294967293,32'd1,32'd4294967293,32'd4294967291,32'd0,32'd5,32'd4294967294,32'd4,32'd0,32'd0,32'd4,32'd4294967287,32'd4,32'd3,32'd4294967290,32'd1,32'd4294967295,32'd4294967294,32'd4294967292,32'd5,32'd4,32'd4294967295,32'd7,32'd4294967279,32'd4294967295,32'd1,32'd4294967288,32'd4294967292,32'd4294967287,32'd20,32'd4294967291,32'd1,32'd3,32'd7,32'd2,32'd4294967292,32'd10,32'd11,32'd4294967294,32'd6,32'd4294967284,32'd10,32'd4294967295,32'd4294967282,32'd7,32'd0,32'd4,32'd4294967294,32'd3,32'd4294967285,32'd3,32'd4294967295,32'd3,32'd6,32'd4294967285,32'd4294967291,32'd8,32'd2,32'd2,32'd4294967293,32'd0,32'd6,32'd4,32'd4294967293,32'd4294967290,32'd1,32'd0,32'd1,32'd6,32'd1,32'd4294967294,32'd1,32'd5,32'd4294967290,32'd0,32'd4294967294,32'd4294967294,32'd4294967293,32'd4294967292,32'd4294967290,32'd2,32'd4294967295,32'd16,32'd4294967295,32'd7,32'd2,32'd15,32'd0,32'd4294967290,32'd1,32'd3,32'd4294967295,32'd4294967295,32'd0,32'd4294967292,32'd14,32'd8,32'd4294967293,32'd2,32'd3,32'd4294967294,32'd4294967294,32'd4294967293,32'd4294967245,32'd5,32'd4294967295,32'd2,32'd1,32'd4294967289,32'd3,32'd0,32'd4294967288,32'd0,32'd4294967292,32'd4,32'd0,32'd2,32'd12,32'd4294967295,32'd4294967290,32'd20,32'd15,32'd4294967294,32'd4294967286,32'd4294967291,32'd3,32'd11,32'd3,32'd4294967294,32'd1,32'd4294967293,32'd1,32'd4294967293,32'd4294967294,32'd4294967294,32'd4294967294,32'd13,32'd10,32'd4294967294,32'd6,32'd5,32'd6,32'd4,32'd4294967291,32'd0,32'd4294967293,32'd3,32'd4294967295,32'd2,32'd4294967293,32'd4294967291,32'd1,32'd0,32'd13,32'd0,32'd2,32'd4294967294,32'd4,32'd3,32'd4294967292,32'd4294967291,32'd0,32'd4294967294,32'd5,32'd0,32'd0,32'd0,32'd2,32'd4294967293,32'd15,32'd4,32'd4294967293,32'd4294967291,32'd0,32'd4294967293,32'd7,32'd4294967289,32'd4294967294,32'd4294967289,32'd0,32'd2,32'd4294967295,32'd4,32'd4,32'd6,32'd0,32'd6,32'd4294967294,32'd8,32'd4294967290,32'd4294967295,32'd4294967294,32'd4294967289,32'd4294967295,32'd4294967292,32'd4294967293,32'd1,32'd5,32'd15,32'd0,32'd4294967280,32'd4294967294,32'd7,32'd3,32'd5,32'd70,32'd12,32'd4294967295,32'd4294967294,32'd4294967285,32'd0,32'd3,32'd10,32'd4294967290,32'd0,32'd4,32'd4,32'd2,32'd4294967294,32'd4294967293,32'd7,32'd4294967295,32'd4,32'd1,32'd3,32'd0,32'd4294967291,32'd4294967294,32'd3,32'd1,32'd6,32'd4294967289,32'd4294967295,32'd7,32'd4294967290,32'd1,32'd2,32'd17,32'd4294967285,32'd4294967293,32'd1,32'd4294967289,32'd4294967293,32'd4294967293,32'd3,32'd1,32'd4294967293,32'd4294967287,32'd7,32'd4294967295,32'd4294967289,32'd4294967285,32'd4294967289,32'd4294967293,32'd4294967294,32'd4294967295,32'd4294967279,32'd11,32'd4294967292,32'd0,32'd6,32'd0,32'd4294967295,32'd4294967293,32'd6,32'd4294967295,32'd8,32'd4294967293,32'd27,32'd4294967295,32'd1,32'd2,32'd4294967294,32'd1,32'd4294967288,32'd4294967295,32'd16,32'd4294967291,32'd4294967292,32'd4294967288,32'd4294967289,32'd3,32'd1,32'd0,32'd4294967293,32'd3,32'd1,32'd1,32'd4,32'd4294967294,32'd0,32'd1,32'd2,32'd4294967295,32'd1,32'd4,32'd4,32'd6,32'd0,32'd4,32'd1,32'd2,32'd4294967294,32'd5,32'd4,32'd6,32'd2,32'd4,32'd5,32'd10,32'd4294967294,32'd2,32'd21,32'd2,32'd6,32'd3,32'd4294967294,32'd4294967289,32'd1,32'd4,32'd2,32'd4294967294,32'd4294967284,32'd3,32'd1,32'd3,32'd4294967290,32'd24,32'd4294967290,32'd3,32'd4294967293,32'd4294967287,32'd9,32'd4294967295,32'd4294967287,32'd4294967289,32'd4,32'd1,32'd1,32'd12,32'd4294967294,32'd1,32'd4294967289,32'd10,32'd0,32'd1,32'd9,32'd4294967275,32'd4294967293,32'd8,32'd5,32'd5,32'd6,32'd4294967288,32'd11,32'd0,32'd4,32'd2,32'd0,32'd4294967294,32'd5,32'd4294967294,32'd4294967292,32'd4294967292,32'd2,32'd4294967295,32'd4294967293,32'd4294967293,32'd2,32'd4294967291,32'd2,32'd2,32'd4294967294,32'd1,32'd2,32'd4294967287,32'd4294967273,32'd29,32'd2,32'd4294967284,32'd7,32'd0,32'd4294967292,32'd3,32'd3,32'd3,32'd0,32'd4294967288,32'd4294967290,32'd4294967294,32'd4294967295,32'd4294967291,32'd4294967294,32'd4294967293,32'd4294967295,32'd4294967294,32'd2,32'd0,32'd4294967294,32'd4294967292,32'd12,32'd2,32'd4294967293,32'd4294967293,32'd4294967295,32'd4294967291,32'd3,32'd4294967295,32'd0,32'd2,32'd3,32'd12,32'd4,32'd4294967294,32'd2,32'd4294967293,32'd4294967294,32'd1,32'd4294967295,32'd7,32'd4294967294,32'd3,32'd1,32'd4294967281,32'd6,32'd4294967295,32'd4294967283,32'd4294967294,32'd4294967295,32'd4294967294,32'd2,32'd18,32'd1,32'd4,32'd2,32'd2,32'd0,32'd7,32'd1,32'd4294967293,32'd3,32'd1,32'd24,32'd0,32'd4294967292,32'd4294967291,32'd4294967292,32'd1,32'd1,32'd1,32'd1,32'd2,32'd4294967295,32'd7,32'd4294967290,32'd4294967294,32'd4294967293,32'd4294967280,32'd4294967290,32'd4294967290,32'd4294967280,32'd4294967282,32'd4294967290,32'd4294967290,32'd0,32'd2,32'd4,32'd0,32'd3,32'd4294967284,32'd1,32'd4294967292,32'd4294967291,32'd0,32'd4294967295,32'd4294967295,32'd4,32'd4294967293,32'd3,32'd4294967292,32'd7,32'd4,32'd4294967293,32'd4,32'd2,32'd4294967290,32'd8,32'd4294967295,32'd6,32'd4294967292,32'd4,32'd1,32'd4294967289,32'd4294967295,32'd4294967292,32'd4294967295,32'd1,32'd4,32'd5,32'd0,32'd4294967293,32'd4294967293,32'd9,32'd4294967294,32'd4294967288,32'd4294967291,32'd4294967292,32'd5,32'd2,32'd26,32'd3,32'd5,32'd4294967292,32'd4294967295,32'd5,32'd4294967293,32'd4294967293,32'd4294967294,32'd2,32'd8,32'd4294967293,32'd4294967293,32'd6,32'd4294967293,32'd4294967292,32'd2,32'd4294967295,32'd4294967284,32'd4294967291,32'd4,32'd1,32'd5,32'd4294967293,32'd35,32'd0,32'd1,32'd4294967288,32'd4294967278,32'd6,32'd4294967291,32'd4294967295,32'd4294967285,32'd4294967293,32'd4294967294,32'd4294967291,32'd4294967291,32'd4294967295,32'd4294967294,32'd3,32'd4294967288,32'd4294967287,32'd4294967293,32'd1,32'd1,32'd4294967294,32'd23,32'd4294967290,32'd4294967292,32'd4294967287,32'd15,32'd12,32'd4294967259,32'd0,32'd3,32'd4294967291,32'd13,32'd1,32'd4294967294,32'd4294967293,32'd2,32'd4294967286,32'd4294967284,32'd0,32'd0,32'd2,32'd4294967292,32'd0,32'd4294967293,32'd4294967291,32'd6,32'd4294967295,32'd4294967291,32'd4294967288,32'd4294967292,32'd12,32'd1,32'd4294967295,32'd4294967295,32'd5,32'd4294967295,32'd11,32'd4294967290,32'd1,32'd2,32'd4294967290,32'd4,32'd1,32'd2,32'd7,32'd3,32'd2,32'd4,32'd18,32'd4294967294,32'd4294967290,32'd36,32'd3,32'd1,32'd4294967295,32'd13,32'd1,32'd4,32'd0,32'd4294967286,32'd4294967292,32'd4,32'd4294967295,32'd4294967287,32'd4294967286,32'd2,32'd10,32'd4294967294,32'd4294967295,32'd21,32'd1,32'd42,32'd4294967293,32'd7,32'd5,32'd12,32'd0,32'd4294967286,32'd4294967292,32'd4294967294,32'd4,32'd7,32'd1,32'd4294967295,32'd4294967295,32'd4294967292,32'd4294967290,32'd4294967292,32'd4294967290,32'd4294967294,32'd0,32'd5,32'd4294967294,32'd4294967270,32'd5,32'd2,32'd4294967285,32'd0,32'd6,32'd4294967294,32'd3,32'd1,32'd4294967292,32'd3,32'd5,32'd8,32'd3,32'd4294967295,32'd4294967294,32'd3,32'd5,32'd0,32'd1,32'd4,32'd4,32'd0,32'd4294967291,32'd4294967292,32'd5,32'd4294967295,32'd6,32'd3,32'd2,32'd4294967295,32'd18,32'd4294967292,32'd2,32'd2,32'd4,32'd2,32'd4294967284,32'd17,32'd4294967290,32'd0,32'd7,32'd19,32'd4294967294,32'd4294967277,32'd4294967292,32'd4294967288,32'd4294967290,32'd4294967295,32'd0,32'd4294967295,32'd1,32'd2,32'd4294967292,32'd0,32'd4294967293,32'd4294967292,32'd4294967293,32'd4294967294,32'd4294967288,32'd4294967294,32'd4294967292,32'd4294967293,32'd0,32'd4294967293,32'd4294967291,32'd4294967295,32'd4294967293,32'd1,32'd3,32'd4,32'd4294967294,32'd4294967295,32'd4294967291,32'd4294967294,32'd4294967294,32'd4294967267,32'd4294967289,32'd1,32'd1,32'd0,32'd5,32'd4294967295,32'd3,32'd4294967290,32'd4294967294,32'd5,32'd4294967295,32'd4294967283,32'd4294967293,32'd4294967295,32'd0,32'd0,32'd8,32'd5,32'd0,32'd0,32'd4294967293,32'd0,32'd4294967291,32'd4294967295,32'd2,32'd4294967287,32'd4294967289,32'd5,32'd4294967294,32'd2,32'd6,32'd2,32'd2,32'd6,32'd2,32'd4294967294,32'd4294967292,32'd4294967293,32'd8,32'd4294967288,32'd4294967269,32'd17,32'd4294967287,32'd4294967291,32'd7,32'd6,32'd16,32'd4294967295,32'd4294967295,32'd2,32'd4294967293,32'd3,32'd4294967294,32'd4294967295,32'd7,32'd6,32'd0,32'd3,32'd4294967288,32'd4294967291,32'd4294967293,32'd2,32'd4294967293,32'd4294967294,32'd4294967295,32'd4294967295,32'd4294967295,32'd4294967282,32'd4,32'd4294967295,32'd4294967289,32'd0,32'd4294967291,32'd4294967291,32'd0,32'd4,32'd1,32'd3,32'd4,32'd1,32'd1,32'd0,32'd1,32'd1,32'd8,32'd4294967292,32'd0,32'd4294967295,32'd4294967291,32'd4294967294,32'd3,32'd2,32'd3,32'd1,32'd4,32'd4,32'd1,32'd4294967282,32'd0,32'd2,32'd1,32'd1,32'd4294967295,32'd2,32'd1,32'd4294967294,32'd30,32'd9,32'd4294967292,32'd2,32'd0,32'd3,32'd4294967290,32'd2,32'd4294967295,32'd3,32'd0,32'd1,32'd4294967292,32'd4294967288,32'd4294967293,32'd5,32'd4294967290,32'd4294967292,32'd8,32'd4294967295,32'd23,32'd4294967273,32'd4294967294,32'd7,32'd3,32'd5,32'd4294967294,32'd4294967292,32'd0,32'd5,32'd1,32'd8,32'd4294967287,32'd4294967290,32'd4,32'd3,32'd4294967294,32'd0,32'd4,32'd0,32'd2,32'd2,32'd12,32'd4,32'd4294967290,32'd4294967290,32'd9,32'd0,32'd15,32'd0,32'd3,32'd4294967286,32'd4294967293,32'd4294967290,32'd0,32'd4294967295,32'd0,32'd4294967294,32'd4294967291,32'd33,32'd11,32'd0,32'd2,32'd4294967292,32'd4294967294,32'd2,32'd4294967293,32'd4294967293,32'd4294967294,32'd4294967291,32'd1,32'd3,32'd4294967292,32'd4294967292,32'd3,32'd4,32'd10,32'd4294967295,32'd4294967294,32'd0,32'd4294967293,32'd4294967295,32'd4294967295,32'd4,32'd0,32'd4,32'd1,32'd4294967293,32'd1,32'd1,32'd11,32'd0,32'd10,32'd24,32'd5,32'd4294967287,32'd4294967294,32'd4294967295,32'd4294967293,32'd2,32'd0,32'd7,32'd6,32'd4294967295,32'd3,32'd3,32'd4294967292,32'd3,32'd4294967279,32'd0,32'd4294967291,32'd4294967288,32'd4294967295,32'd4294967291,32'd4,32'd4294967295,32'd2,32'd4294967291,32'd1,32'd4294967260,32'd3,32'd2,32'd1,32'd1,32'd19,32'd2,32'd4294967288,32'd4294967290,32'd3,32'd0,32'd4294967286,32'd4,32'd0,32'd4294967295,32'd5,32'd2,32'd2,32'd48,32'd4294967291,32'd4294967289,32'd15,32'd0,32'd11,32'd4294967290,32'd4294967287,32'd6,32'd6,32'd4294967295,32'd4,32'd0,32'd2,32'd2,32'd4,32'd9,32'd12,32'd1,32'd2,32'd4294967278,32'd4294967293,32'd2,32'd4294967295,32'd4294967295,32'd2,32'd1,32'd4294967294,32'd5,32'd12,32'd3,32'd3,32'd4294967293,32'd1,32'd4294967294,32'd0,32'd13,32'd2,32'd1,32'd3,32'd2,32'd4294967292}
`define FEATURE_ABOVE {32'd0,32'd215,32'd28,32'd4294967292,32'd4294967157,32'd4294967181,32'd15,32'd111,32'd44,32'd4294967275,32'd23,32'd4294967183,32'd4294967265,32'd4294967276,32'd88,32'd4294967273,32'd4294967230,32'd81,32'd27,32'd4294967243,32'd18,32'd4294967293,32'd4294967291,32'd75,32'd4294967241,32'd35,32'd16,32'd4294967273,32'd10,32'd4294967189,32'd15,32'd60,32'd10,32'd202,32'd19,32'd4294967237,32'd4294967284,32'd51,32'd4294967264,32'd8,32'd85,32'd4294967288,32'd7,32'd4294967159,32'd20,32'd4294967272,32'd11,32'd15,32'd51,32'd4294967277,32'd4294967268,32'd4294967231,32'd15,32'd0,32'd86,32'd38,32'd25,32'd4294967288,32'd71,32'd4294967278,32'd4294967258,32'd23,32'd40,32'd43,32'd62,32'd4294967220,32'd4294967184,32'd92,32'd10,32'd4294967178,32'd4294967249,32'd10,32'd10,32'd4294967276,32'd26,32'd37,32'd22,32'd4294967278,32'd33,32'd4294967122,32'd4294967289,32'd76,32'd4294967184,32'd4294967291,32'd0,32'd19,32'd200,32'd4294967293,32'd4294967163,32'd34,32'd54,32'd4294967167,32'd9,32'd4294967237,32'd4294967212,32'd4294967274,32'd53,32'd4294967249,32'd36,32'd4294967276,32'd46,32'd4294967269,32'd9,32'd56,32'd4,32'd51,32'd59,32'd4294967293,32'd4294967293,32'd4294967266,32'd18,32'd4294967273,32'd11,32'd4294967256,32'd4294967295,32'd4294967121,32'd17,32'd19,32'd8,32'd0,32'd4294967229,32'd4294967275,32'd0,32'd53,32'd4294967201,32'd45,32'd22,32'd40,32'd8,32'd4294967215,32'd16,32'd4294967292,32'd4294967230,32'd4294967271,32'd116,32'd4294967270,32'd50,32'd16,32'd4294967295,32'd4294967208,32'd40,32'd140,32'd4294967294,32'd4294967292,32'd41,32'd4294967113,32'd4294967284,32'd4294967290,32'd4294967283,32'd4294967289,32'd4294967054,32'd229,32'd18,32'd4294967268,32'd7,32'd4294967270,32'd18,32'd4294967237,32'd105,32'd4294967272,32'd26,32'd4294967250,32'd4294967284,32'd4294967086,32'd32,32'd122,32'd25,32'd7,32'd24,32'd27,32'd4294967292,32'd4294967294,32'd25,32'd4294967216,32'd21,32'd40,32'd24,32'd4294967290,32'd28,32'd4294967263,32'd25,32'd4294967258,32'd109,32'd4294967186,32'd115,32'd18,32'd4294967279,32'd4294967265,32'd95,32'd4294967205,32'd33,32'd4294967194,32'd21,32'd4294967196,32'd52,32'd4294967257,32'd4294967215,32'd54,32'd28,32'd4294967237,32'd4294967245,32'd82,32'd4294967288,32'd44,32'd4294967177,32'd62,32'd3,32'd4294967218,32'd34,32'd36,32'd24,32'd41,32'd4294967106,32'd4294967024,32'd4294967269,32'd54,32'd4294967288,32'd5,32'd122,32'd24,32'd4294967272,32'd14,32'd49,32'd150,32'd4294967158,32'd71,32'd4294967275,32'd17,32'd1,32'd21,32'd4294967188,32'd4294967288,32'd3,32'd4294967294,32'd4294967291,32'd4294967094,32'd57,32'd4294967245,32'd90,32'd4294967090,32'd4294967025,32'd4294967174,32'd4294967270,32'd4294967290,32'd167,32'd4294967041,32'd4294967276,32'd4294966934,32'd6,32'd34,32'd4294967266,32'd26,32'd4294967178,32'd4294967290,32'd56,32'd46,32'd0,32'd6,32'd43,32'd5,32'd4294967115,32'd14,32'd4294967231,32'd314,32'd4294967214,32'd4294966679,32'd4294967154,32'd16,32'd4294967274,32'd21,32'd10,32'd4294967283,32'd4294967267,32'd15,32'd27,32'd36,32'd4294967289,32'd4294967251,32'd4294967172,32'd7,32'd35,32'd134,32'd0,32'd25,32'd191,32'd4294967179,32'd14,32'd4294967288,32'd80,32'd306,32'd4294967273,32'd22,32'd9,32'd33,32'd60,32'd7,32'd4294967264,32'd35,32'd84,32'd37,32'd325,32'd4294967295,32'd4294967294,32'd4294967260,32'd4294967275,32'd23,32'd4294967113,32'd4294967053,32'd9,32'd1,32'd6,32'd66,32'd4294967267,32'd4294967255,32'd4294967197,32'd4294967232,32'd34,32'd4294967259,32'd4294967268,32'd45,32'd4294967230,32'd29,32'd4294967272,32'd4294967273,32'd4294967277,32'd31,32'd57,32'd79,32'd4294967049,32'd23,32'd79,32'd0,32'd66,32'd46,32'd4294967262,32'd7,32'd4294967291,32'd77,32'd4294967291,32'd4294967277,32'd4294967290,32'd4294967104,32'd38,32'd42,32'd4294967291,32'd4294967218,32'd4294967125,32'd4294967188,32'd4294967256,32'd11,32'd4294967293,32'd4294967176,32'd4294967257,32'd4294967288,32'd128,32'd39,32'd4294967273,32'd27,32'd45,32'd83,32'd4294967211,32'd29,32'd4294967271,32'd24,32'd4294967264,32'd20,32'd4294967290,32'd4294963456,32'd4294967272,32'd10,32'd4,32'd31,32'd4294967237,32'd24,32'd4294967203,32'd4294967268,32'd4294967267,32'd88,32'd53,32'd6,32'd69,32'd16,32'd4294967254,32'd62,32'd4294967226,32'd4294967289,32'd4294967291,32'd4294967261,32'd4294967294,32'd78,32'd4294967268,32'd20,32'd4294967291,32'd4294967227,32'd4294967292,32'd24,32'd4294967191,32'd4294967252,32'd92,32'd4294967234,32'd4294967265,32'd4294967288,32'd4,32'd44,32'd4294967264,32'd57,32'd36,32'd4294967211,32'd55,32'd58,32'd50,32'd394,32'd8,32'd4294967231,32'd4294967128,32'd67,32'd4294967096,32'd27,32'd7,32'd3,32'd26,32'd138,32'd35,32'd47,32'd14,32'd4294967288,32'd16,32'd4294967277,32'd8,32'd4294967183,32'd28,32'd175,32'd4294967173,32'd1,32'd116,32'd4294967263,32'd4,32'd3,32'd14,32'd83,32'd41,32'd4294967267,32'd4,32'd4294967114,32'd4294967195,32'd76,32'd18,32'd160,32'd54,32'd79,32'd22,32'd4294967277,32'd89,32'd4294967217,32'd20,32'd4294967151,32'd4294967186,32'd4294967271,32'd4294967287,32'd7,32'd4294967273,32'd20,32'd9,32'd65,32'd29,32'd4294967255,32'd2,32'd4294967138,32'd18,32'd4294967270,32'd4294967155,32'd11,32'd12,32'd4294967288,32'd98,32'd145,32'd4294967285,32'd1,32'd14,32'd4294967293,32'd4294967295,32'd4294967175,32'd4294967290,32'd4294967225,32'd20,32'd4294967271,32'd17,32'd3,32'd26,32'd118,32'd7,32'd4294967255,32'd39,32'd89,32'd4294966893,32'd75,32'd17,32'd53,32'd64,32'd4294967160,32'd26,32'd4294967265,32'd32,32'd4294967274,32'd11,32'd4294967295,32'd4294967129,32'd188,32'd4294966845,32'd4294967295,32'd37,32'd4294967290,32'd4294967236,32'd4294967238,32'd4294967290,32'd4294967186,32'd9,32'd4294967262,32'd39,32'd4,32'd23,32'd4294967270,32'd4294967242,32'd4294967294,32'd0,32'd4294967278,32'd0,32'd8,32'd4294967206,32'd4294967288,32'd4294963456,32'd4294967246,32'd31,32'd4294967271,32'd16,32'd1,32'd24,32'd4294967291,32'd4294967281,32'd4294967198,32'd21,32'd4294967271,32'd4294967218,32'd4294967274,32'd112,32'd1,32'd26,32'd4294967275,32'd3,32'd4294967257,32'd91,32'd4294967243,32'd4294967275,32'd4294967294,32'd4294967233,32'd4294967270,32'd22,32'd4294967251,32'd4,32'd52,32'd70,32'd4294967176,32'd4294967289,32'd129,32'd22,32'd140,32'd94,32'd4294967266,32'd76,32'd4294967295,32'd4294967254,32'd4294967271,32'd4294967272,32'd4294967130,32'd30,32'd18,32'd4294967294,32'd4294967294,32'd5,32'd4294967274,32'd4294967225,32'd0,32'd20,32'd33,32'd16,32'd4294967292,32'd29,32'd4294967292,32'd4294967291,32'd12,32'd17,32'd4294967295,32'd4294967224,32'd126,32'd17,32'd4294967242,32'd4294967228,32'd205,32'd4294967258,32'd23,32'd57,32'd4294967182,32'd67,32'd4294967259,32'd4294967277,32'd82,32'd75,32'd50,32'd78,32'd38,32'd4294967260,32'd7,32'd111,32'd12,32'd73,32'd4294967282,32'd4294967108,32'd15,32'd4294967099,32'd4294967232,32'd59,32'd10,32'd25,32'd4294967127,32'd59,32'd8,32'd4294967243,32'd53,32'd4294967277,32'd4294967006,32'd4294967287,32'd18,32'd4294967269,32'd4294967293,32'd4294967201,32'd4294967210,32'd4294967287,32'd4294967281,32'd4294967295,32'd4,32'd130,32'd4294967275,32'd119,32'd15,32'd72,32'd21,32'd22,32'd4294967292,32'd4294967290,32'd4294967094,32'd4294967291,32'd4294967215,32'd4294967194,32'd4294967290,32'd4294967287,32'd6,32'd48,32'd4294967219,32'd293,32'd5,32'd4294967227,32'd50,32'd4294967227,32'd8,32'd4294967278,32'd8,32'd15,32'd4294967218,32'd61,32'd18,32'd4294967190,32'd24,32'd4294967165,32'd15,32'd3,32'd4294967110,32'd65,32'd8,32'd4294967260,32'd68,32'd4294967293,32'd21,32'd24,32'd4294967150,32'd4294967255,32'd97,32'd9,32'd4294967269,32'd4294967225,32'd4294967260,32'd10,32'd58,32'd4294967269,32'd4294967248,32'd9,32'd23,32'd4294967189,32'd42,32'd4294967292,32'd19,32'd4294967253,32'd4294967280,32'd4294967274,32'd4294967239,32'd95,32'd16,32'd4294967164,32'd4294967044,32'd4294967274,32'd4294967193,32'd4294967291,32'd22,32'd4294967244,32'd11,32'd4294967264,32'd2,32'd32,32'd11,32'd4294967260,32'd38,32'd7,32'd26,32'd197,32'd4294967201,32'd97,32'd4294967294,32'd70,32'd21,32'd4294967292,32'd1,32'd4294967276,32'd50,32'd75,32'd4294967114,32'd4294967254,32'd103,32'd4294967266,32'd4294967239,32'd210,32'd8,32'd4294967263,32'd30,32'd4294967259,32'd3,32'd4294967288,32'd41,32'd4294967273,32'd66,32'd4294967172,32'd4,32'd110,32'd30,32'd4294967293,32'd85,32'd4294967132,32'd4,32'd4294967272,32'd95,32'd4294967197,32'd0,32'd4294967254,32'd4294967148,32'd122,32'd66,32'd4294967079,32'd4294967087,32'd4294967250,32'd1,32'd4294967176,32'd32,32'd0,32'd1,32'd4294967166,32'd4294967288,32'd60,32'd2,32'd4294967193,32'd86,32'd4294967269,32'd30,32'd4294967209,32'd27,32'd3,32'd4294967226,32'd4294967183,32'd4294967261,32'd4294967261,32'd40,32'd33,32'd88,32'd51,32'd63,32'd5,32'd4294967143,32'd4294967230,32'd4294967290,32'd3,32'd0,32'd12,32'd4294967252,32'd25,32'd4294967267,32'd4294967225,32'd18,32'd4294967223,32'd25,32'd139,32'd4294967294,32'd4294967209,32'd4294967259,32'd4294967279,32'd38,32'd30,32'd420,32'd24,32'd4294967273,32'd4294967270,32'd89,32'd94,32'd4294967289,32'd11,32'd4294966996,32'd18,32'd83,32'd54,32'd10,32'd18,32'd4294967202,32'd17,32'd2,32'd4294966721,32'd4294967276,32'd21,32'd85,32'd4294967195,32'd4294967275,32'd4294967282,32'd70,32'd36,32'd4294967269,32'd5,32'd4294967273,32'd4294967203,32'd4294967240,32'd15,32'd4294967252,32'd6,32'd4294967289,32'd15,32'd4294967264,32'd89,32'd142,32'd4294967273,32'd8,32'd26,32'd4294967196,32'd37,32'd105,32'd4294967155,32'd124,32'd4294967224,32'd4294967187,32'd34,32'd13,32'd4294967286,32'd4294967274,32'd211,32'd4294967205,32'd4294966969,32'd4294967276,32'd110,32'd4294967287,32'd4294967291,32'd6,32'd33,32'd243,32'd15,32'd11,32'd8,32'd11,32'd4294967167,32'd44,32'd19,32'd4294967273,32'd4294967264,32'd4294967291,32'd0,32'd2,32'd4294967258,32'd4294967224,32'd18,32'd2,32'd17,32'd4294967263,32'd29,32'd4294967270,32'd7,32'd0,32'd104,32'd4294967272,32'd57,32'd4294967289,32'd4294967115,32'd4294967288,32'd4294967288,32'd4294967273,32'd24,32'd4294967290,32'd4294967258,32'd4294967273,32'd6,32'd6,32'd4294967241,32'd4294967248,32'd71,32'd2,32'd19,32'd4294967090,32'd4294967266,32'd4294967255,32'd75,32'd4294967212,32'd44,32'd7,32'd3,32'd4294967184,32'd23,32'd4294967268,32'd28,32'd6,32'd4294967254,32'd4294967191,32'd4294967244,32'd4294967253,32'd7,32'd4294967292,32'd11,32'd18,32'd5,32'd4294967265,32'd29,32'd4294967238,32'd20,32'd77,32'd159,32'd4294967289,32'd51,32'd4294967270,32'd18,32'd4294967265,32'd38,32'd27,32'd4294967170,32'd54,32'd4294967291,32'd4294967294,32'd23,32'd94,32'd4294967276,32'd4294967293,32'd21,32'd9,32'd32,32'd4294967177,32'd21,32'd4294967202,32'd4294967289,32'd4294967295,32'd4294967269,32'd0,32'd17,32'd53,32'd4294967248,32'd4294967262,32'd4294967292,32'd3,32'd4294967168,32'd4294967258,32'd40,32'd62,32'd27,32'd4294967165,32'd16,32'd4294967208,32'd18,32'd38,32'd4294967243,32'd78,32'd4294967260,32'd4294967260,32'd4294967278,32'd0,32'd4294967258,32'd4294967265,32'd15,32'd43,32'd110,32'd4294967277,32'd11,32'd4294967151,32'd4294967275,32'd65,32'd63,32'd0,32'd8,32'd4294967293,32'd4294967293,32'd4294967271,32'd15,32'd4294967243,32'd2,32'd4294967294,32'd4294967272,32'd4294967294,32'd9,32'd4294967151,32'd4294967273,32'd42,32'd4294967256,32'd4294967273,32'd2,32'd4294966862,32'd48,32'd4294967278,32'd4294967292,32'd4294967293,32'd2,32'd4294967134,32'd4294967210,32'd4294967295,32'd4294966998,32'd4294967289,32'd20,32'd4294967266,32'd32,32'd4294967258,32'd14,32'd4294967243,32'd28,32'd16,32'd54,32'd0,32'd69,32'd4294967270,32'd5,32'd144,32'd21,32'd4294967293,32'd16,32'd4294967277,32'd22,32'd41,32'd6,32'd4294967294,32'd4294967292,32'd4294967278,32'd41,32'd34,32'd64,32'd4294967291,32'd4294967293,32'd10,32'd35,32'd4294967266,32'd6,32'd4294967295,32'd27,32'd4294967269,32'd30,32'd4294967291,32'd4294967288,32'd4294967123,32'd4294967253,32'd89,32'd55,32'd34,32'd19,32'd54,32'd19,32'd4294967275,32'd20,32'd182,32'd4294967216,32'd4294967228,32'd26,32'd50,32'd4294967232,32'd39,32'd65,32'd4294967288,32'd4294967288,32'd35,32'd11,32'd4294967287,32'd4294967205,32'd4294967217,32'd4294967219,32'd99,32'd20,32'd4294967287,32'd4294967262,32'd51,32'd49,32'd4294967240,32'd28,32'd8,32'd29,32'd10,32'd24,32'd4,32'd19,32'd4294967252,32'd0,32'd4,32'd4294967164,32'd15,32'd33,32'd4294967169,32'd52,32'd119,32'd54,32'd4294967256,32'd4294967263,32'd4294967294,32'd4294967272,32'd4294967276,32'd4294967080,32'd4294967295,32'd4294967168,32'd4294967289,32'd117,32'd151,32'd18,32'd66,32'd48,32'd4294967219,32'd20,32'd4294967208,32'd24,32'd6,32'd74,32'd4294967257,32'd42,32'd4294967206,32'd4294967293,32'd4294967068,32'd35,32'd4294967274,32'd124,32'd4294967293,32'd4294967290,32'd4294967182,32'd37,32'd65,32'd19,32'd4294967148,32'd4294967287,32'd107,32'd21,32'd0,32'd4294967254,32'd4294967051,32'd18,32'd29,32'd103,32'd4294967184,32'd4294967165,32'd34,32'd70,32'd3,32'd26,32'd4294967251,32'd26,32'd4294967137,32'd66,32'd4294967158,32'd32,32'd4294967268,32'd91,32'd4294967170,32'd59,32'd70,32'd56,32'd78,32'd4294967272,32'd105,32'd4294967291,32'd4294967287,32'd4294967290,32'd4294967278,32'd4,32'd18,32'd4294967271,32'd16,32'd4294967265,32'd4294967011,32'd4294967293,32'd4294967285,32'd4294967198,32'd4294967292,32'd4294967288,32'd4294966687,32'd56,32'd42,32'd4294967292,32'd39,32'd4294967202,32'd4294967209,32'd4294967279,32'd7,32'd4294967262,32'd4294967235,32'd4294967272,32'd4,32'd20,32'd4294967237,32'd4294967079,32'd4294967244,32'd4294967267,32'd48,32'd3,32'd74,32'd4294967289,32'd17,32'd4294967277,32'd4294967096,32'd69,32'd18,32'd267,32'd369,32'd4294967242,32'd73,32'd4294967165,32'd4294967262,32'd61,32'd4294967295,32'd4294967274,32'd41,32'd1,32'd4294967274,32'd62,32'd1,32'd4294967253,32'd0,32'd5,32'd32,32'd79,32'd4294967269,32'd7,32'd29,32'd4294967156,32'd19,32'd79,32'd4294967279,32'd95,32'd53,32'd4294967218,32'd4294967235,32'd101,32'd69,32'd4294967209,32'd18,32'd43,32'd12,32'd86,32'd36,32'd4294967238,32'd19,32'd1,32'd18,32'd4294967295,32'd11,32'd4294967270,32'd20,32'd4294967291,32'd4294967251,32'd61,32'd22,32'd4294967277,32'd1,32'd4294967290,32'd4,32'd4294967292,32'd4294967218,32'd41,32'd4294967280,32'd69,32'd29,32'd4294967178,32'd49,32'd4294967042,32'd21,32'd4,32'd4,32'd4294967266,32'd82,32'd3,32'd4294967261,32'd115,32'd77,32'd4294967291,32'd4294967270,32'd4294967266,32'd32,32'd4294967265,32'd6,32'd4,32'd49,32'd4294967186,32'd12,32'd4294967175,32'd4294967265,32'd18,32'd31,32'd4294967261,32'd22,32'd4,32'd4294967217,32'd4294967265,32'd17,32'd60,32'd32,32'd4,32'd19,32'd4294967157,32'd66,32'd4294967203,32'd18,32'd4294967262,32'd29,32'd13,32'd34,32'd4294967263,32'd4294967180,32'd1,32'd20,32'd54,32'd4294967286,32'd3,32'd103,32'd4294967271,32'd29,32'd4294967191,32'd5,32'd23,32'd30,32'd12,32'd53,32'd65,32'd78,32'd28,32'd77,32'd4294967221,32'd64,32'd10,32'd4294967233,32'd67,32'd9,32'd27,32'd4294967267,32'd39,32'd4294967218,32'd22,32'd33,32'd4294967281,32'd4294967115,32'd27,32'd4294967063,32'd0,32'd4294967291,32'd25,32'd93,32'd4294967121,32'd4294967204,32'd100,32'd4294967022,32'd19,32'd4294966976,32'd9,32'd4294967207,32'd126,32'd4294967154,32'd50,32'd4294967058,32'd4294967145,32'd4294967295,32'd0,32'd4294967259,32'd4294967205,32'd51,32'd17,32'd6,32'd27,32'd4294967277,32'd4294967210,32'd4,32'd33,32'd4294967250,32'd28,32'd4294967295,32'd98,32'd4294967199,32'd2,32'd4294967277,32'd4294967274,32'd4294967189,32'd22,32'd4294967266,32'd14,32'd4294967261,32'd47,32'd4294967188,32'd9,32'd25,32'd139,32'd4294967270,32'd2,32'd4294967168,32'd4294967099,32'd21,32'd23,32'd43,32'd1280,32'd4294967255,32'd4294967289,32'd5,32'd45,32'd44,32'd0,32'd4294967293,32'd4294967179,32'd45,32'd4294967247,32'd4294967274,32'd4294967247,32'd4294967155,32'd2,32'd11,32'd4294967024,32'd4294967273,32'd4294967215,32'd4294967289,32'd16,32'd74,32'd4294967288,32'd4294967197,32'd41,32'd4294967204,32'd48,32'd4294967219,32'd129,32'd4294967292,32'd22,32'd4294967269,32'd31,32'd4294967274,32'd4294967165,32'd4294967255,32'd30,32'd2,32'd4294967248,32'd58,32'd4294967125,32'd4294967159,32'd22,32'd4294967265,32'd4294967289,32'd4294967145,32'd133,32'd4294967262,32'd19,32'd6,32'd26,32'd4294967258,32'd0,32'd4294967294,32'd4294967233,32'd4294967117,32'd4294967284,32'd2,32'd20,32'd4294967219,32'd28,32'd4294967266,32'd19,32'd4294967272,32'd28,32'd4294967269,32'd23,32'd4294967193,32'd22,32'd0,32'd57,32'd50,32'd4294967179,32'd4294967272,32'd54,32'd4294967211,32'd31,32'd15,32'd35,32'd31,32'd35,32'd4294967208,32'd4294967222,32'd4294967215,32'd51,32'd98,32'd63,32'd4294967025,32'd250,32'd4294967236,32'd4294967215,32'd16,32'd4294967294,32'd18,32'd4294967268,32'd4,32'd4294967270,32'd4294967242,32'd4294967277,32'd4294967156,32'd11,32'd35,32'd4294967270,32'd52,32'd4294967010,32'd4294967259,32'd4294967295,32'd9,32'd2,32'd4294967268,32'd64,32'd4294967293,32'd69,32'd1,32'd62,32'd17,32'd4294967229,32'd17,32'd4294967274,32'd4,32'd14,32'd4294967209,32'd200,32'd4294967104,32'd4294967176,32'd4294967145,32'd4294967290,32'd126,32'd3,32'd14,32'd4294967276,32'd24,32'd4294967047,32'd25,32'd4294967249,32'd4294967216,32'd4294967261,32'd4294966921,32'd4294967155,32'd24,32'd4294967262,32'd85,32'd4294967153,32'd37,32'd93,32'd32,32'd4294967267,32'd26,32'd4294967288,32'd4294967295,32'd4294967267,32'd101,32'd4294967252,32'd20,32'd4294967213,32'd54,32'd4294967187,32'd21,32'd15,32'd10,32'd4294967156,32'd15,32'd31,32'd90,32'd56,32'd4294967288,32'd4294967238,32'd90,32'd4294967126,32'd38,32'd4294967149,32'd4294967262,32'd4,32'd4294967259,32'd4294967263,32'd4294967199,32'd4294967270,32'd32,32'd4294967261,32'd73,32'd4294967293,32'd77,32'd4294967269,32'd23,32'd76,32'd37,32'd4294967272,32'd4294967292,32'd128,32'd4294967200,32'd79,32'd18,32'd4294967147,32'd4294967282,32'd4294967039,32'd62,32'd44,32'd18,32'd20,32'd348,32'd4294967133,32'd4294967231,32'd4294967187,32'd79,32'd0,32'd4294967162,32'd4294967269,32'd4294967210,32'd10,32'd30,32'd4294967295,32'd67,32'd39,32'd4294967200,32'd4294967170,32'd4294966789,32'd4294967277,32'd4294967153,32'd5,32'd29,32'd2,32'd4294967151,32'd4294967270,32'd4294967290,32'd4294967291,32'd4294967282,32'd4294967239,32'd23,32'd53,32'd42,32'd151,32'd20,32'd5,32'd26,32'd4294967270,32'd4294967256,32'd4294967141,32'd35,32'd4294967247,32'd40,32'd29,32'd97,32'd4294967132,32'd116,32'd4294967210,32'd4294967270,32'd4294967087,32'd41,32'd4294967164,32'd5,32'd4294967274,32'd68,32'd4294967275,32'd70,32'd4294967131,32'd4294967268,32'd4294967285,32'd102,32'd4294967116,32'd4294967260,32'd4294967294,32'd3,32'd4294967247,32'd4294967061,32'd32,32'd1,32'd22,32'd0,32'd4294967276,32'd4294967060,32'd20,32'd99,32'd160,32'd15,32'd102,32'd52,32'd4294967194,32'd4294967247,32'd29,32'd0,32'd55,32'd4294967269,32'd4294967194,32'd4294967188,32'd0,32'd4294967158,32'd4294967291,32'd4294967289,32'd4294967281,32'd1,32'd16,32'd4294967272,32'd159,32'd4294967151,32'd20,32'd4294967268,32'd75,32'd33,32'd33,32'd0,32'd4294967265,32'd4294967273,32'd22,32'd144,32'd2,32'd22,32'd4,32'd4294967205,32'd4294967158,32'd4294967293,32'd79,32'd90,32'd4294967240,32'd4294966979,32'd4294967277,32'd4294967292,32'd45,32'd0,32'd4294967155,32'd1,32'd18,32'd4294967272,32'd59,32'd142,32'd15,32'd9,32'd22,32'd35,32'd4,32'd2,32'd4294967238,32'd4294967294,32'd27,32'd4294967251,32'd24,32'd17,32'd25,32'd4294967264,32'd103,32'd5,32'd19,32'd4294967293,32'd4294967207,32'd4294967292,32'd19,32'd4294967274,32'd105,32'd16,32'd20,32'd54,32'd20,32'd4294967183,32'd36,32'd8,32'd4294967269,32'd8,32'd4,32'd71,32'd34,32'd4294967261,32'd4294967247,32'd4294967293,32'd4294967276,32'd4294967268,32'd4294967283,32'd39,32'd93,32'd4294967254,32'd0,32'd4294967172,32'd4294967207,32'd5,32'd4294967207,32'd13,32'd110,32'd46,32'd4294967243,32'd3,32'd22,32'd53,32'd4294967258,32'd75,32'd4294967195,32'd4294967272,32'd8,32'd4294967292,32'd100,32'd4294967242,32'd25,32'd4294967294,32'd4294967243,32'd156,32'd4294967208,32'd4294967295,32'd20,32'd28,32'd3,32'd39,32'd44,32'd4294967277,32'd4294966697,32'd4294967148,32'd16,32'd4294967273,32'd4294967251,32'd214,32'd26,32'd26,32'd26,32'd4294967076,32'd4294967136,32'd132,32'd4294967293,32'd4294967070,32'd4294967259,32'd4294967263,32'd22,32'd34,32'd95,32'd4294967045,32'd33,32'd4294967257,32'd4294967265,32'd56,32'd4,32'd4294967158,32'd4294966947,32'd80,32'd18,32'd66,32'd4294967245,32'd11,32'd4294967288,32'd1,32'd81,32'd5,32'd54,32'd4294967294,32'd4294967289,32'd4294967256,32'd68,32'd4294967269,32'd15,32'd4294967293,32'd15,32'd0,32'd4294967118,32'd4294967252,32'd105,32'd4294967272,32'd14,32'd1,32'd4294967274,32'd2,32'd71,32'd59,32'd4294967231,32'd28,32'd17,32'd4294967184,32'd22,32'd4294967135,32'd31,32'd12,32'd43,32'd119,32'd4294967250,32'd50,32'd53,32'd4294967168,32'd25,32'd4294967167,32'd4294967263,32'd123,32'd4294966977,32'd4294967147,32'd43,32'd69,32'd4294967069,32'd4294967263,32'd18,32'd58,32'd30,32'd4294967206,32'd20,32'd4294967294,32'd4294967262,32'd4294967151,32'd4294967236,32'd32,32'd38,32'd4294967229,32'd4294967224,32'd4294967263,32'd42,32'd76,32'd5,32'd4294967198,32'd4294967281,32'd4294967294,32'd27,32'd93,32'd116,32'd10,32'd91,32'd4294967263,32'd24,32'd8,32'd29,32'd4294967253,32'd7,32'd141,32'd4294967270,32'd55,32'd74,32'd73,32'd39,32'd4294967207,32'd248,32'd122,32'd4294967295,32'd206,32'd4294967292,32'd158,32'd4294967230,32'd17,32'd275,32'd24,32'd78,32'd3,32'd4294967053,32'd20,32'd30,32'd4294967249,32'd4294967157,32'd4294967139,32'd4294967289,32'd4294967295,32'd4294967052,32'd73,32'd60,32'd0,32'd4,32'd4294967169,32'd4294967213,32'd23,32'd4294967269,32'd48,32'd4,32'd51,32'd4294967162,32'd33,32'd4294967277,32'd48,32'd4294967125,32'd1,32'd7,32'd20,32'd4294967290,32'd8,32'd4294967294,32'd20,32'd31,32'd2,32'd4294967128,32'd22,32'd4294967173,32'd4294967231,32'd70,32'd4294967200,32'd4294967274,32'd63,32'd4294967168,32'd28,32'd4294967271,32'd27,32'd4294967275,32'd4294967020,32'd163,32'd31,32'd25,32'd46,32'd5,32'd26,32'd4294967268,32'd6,32'd149,32'd4294967286,32'd4294967210,32'd75,32'd4294967271,32'd48,32'd29,32'd14,32'd17,32'd4294967291,32'd184,32'd27,32'd4294967230,32'd4294967237,32'd4294967258,32'd2,32'd71,32'd53,32'd4294967243,32'd19,32'd4294967293,32'd4294967246,32'd4294967102,32'd4294967205,32'd4294967292,32'd4294967258,32'd4294967295,32'd4294967275,32'd4294967259,32'd2,32'd1,32'd6,32'd129,32'd79,32'd4294967266,32'd4294967157,32'd99,32'd118,32'd80,32'd23,32'd4294967234,32'd4294967285,32'd4294967136,32'd4294967265,32'd4294967184,32'd25,32'd4294967293,32'd4294967203,32'd4294967230,32'd4294967124,32'd44,32'd4294967239,32'd6,32'd4294967112,32'd91,32'd1,32'd4294967264,32'd31,32'd4294967260,32'd4294967158,32'd34,32'd34,32'd24,32'd46,32'd4294967210,32'd90,32'd66,32'd4294967271,32'd2,32'd4294967243,32'd0,32'd4294967118,32'd22,32'd4294967295,32'd7,32'd27,32'd112,32'd16,32'd73,32'd4294967154,32'd4294966968,32'd4294967239,32'd68,32'd4294967259,32'd117,32'd4294967293,32'd4294967289,32'd4,32'd12,32'd4294967252,32'd20,32'd4294967266,32'd52,32'd71,32'd76,32'd4294967248,32'd21,32'd4294967258,32'd4294966981,32'd4294967183,32'd98,32'd4294967082,32'd4294967200,32'd6,32'd23,32'd4294967276,32'd27,32'd4294967153,32'd149,32'd4294967292,32'd27,32'd4294967175,32'd75,32'd50,32'd4294967292,32'd4294967295,32'd4294967043,32'd4294967257,32'd4294967174,32'd56,32'd4294967243,32'd4294967236,32'd19,32'd0,32'd4294967205,32'd66,32'd4294967137,32'd4294967294,32'd0,32'd4294967139,32'd4294967294,32'd18,32'd48,32'd4294967099,32'd8,32'd4294967293,32'd4294967219,32'd4294967269,32'd24,32'd4294967267,32'd4294967234,32'd42,32'd21,32'd4294967294,32'd4294966967,32'd4294967245,32'd24,32'd4294967269,32'd4294967294,32'd7,32'd30,32'd4294967294,32'd21,32'd4294967098,32'd23,32'd4294967205,32'd4294967140,32'd51,32'd4294967287,32'd4294967274,32'd137,32'd6,32'd4294967144,32'd4294967267,32'd132,32'd4294967248,32'd77,32'd4294967260,32'd4294967277,32'd49,32'd25,32'd3,32'd4294967170,32'd2,32'd19,32'd4294967267,32'd4,32'd67,32'd4294967269,32'd4294967239,32'd24,32'd4294967097,32'd61,32'd4294967229,32'd74,32'd16,32'd47,32'd26,32'd15,32'd4294967205,32'd25,32'd87,32'd57,32'd73,32'd10,32'd4294967270,32'd4294967184,32'd4294967257,32'd4294967260,32'd67,32'd49,32'd201,32'd4294967216,32'd4294967189,32'd4294967195,32'd4294967164,32'd4294967255,32'd69,32'd4294967090,32'd50,32'd152,32'd4294967091,32'd4294967272,32'd9,32'd99,32'd4294967233,32'd93,32'd2,32'd4294967291,32'd43,32'd4294967200,32'd69,32'd0,32'd89,32'd4294967274,32'd52,32'd4294967258,32'd26,32'd94,32'd4294967275,32'd4294967275,32'd8,32'd4294967204,32'd50,32'd18,32'd4294967130,32'd4294967273,32'd46,32'd4294967291,32'd269,32'd4294967228,32'd4294967247,32'd38,32'd4,32'd4294967292,32'd190,32'd4294967194,32'd72,32'd69,32'd18,32'd4294967143,32'd55,32'd4294967139,32'd4294967212,32'd4294967200,32'd21,32'd68,32'd2,32'd4294967292,32'd17,32'd76,32'd4294967285,32'd4294967294,32'd21,32'd4294967147,32'd25,32'd143,32'd4294967248,32'd6,32'd92,32'd141,32'd4294967291,32'd4294967264,32'd99,32'd27,32'd25,32'd74,32'd33,32'd6,32'd4294967206,32'd72,32'd67,32'd7,32'd23,32'd4294967268,32'd22,32'd6,32'd28,32'd8,32'd28,32'd4294967229,32'd4294967236,32'd4294967173,32'd4294967279,32'd4294967252,32'd20,32'd94,32'd4294967206,32'd4294967260,32'd27,32'd15,32'd4294967292,32'd67,32'd42,32'd4294967153,32'd40,32'd72,32'd129,32'd74,32'd4294967262,32'd48,32'd4294967272,32'd28,32'd24,32'd4294967287,32'd4294967049,32'd4294967284,32'd4294967165,32'd26,32'd4294967270,32'd50,32'd4294967238,32'd15,32'd4294967270,32'd4294967274,32'd3,32'd4294967261,32'd4294967182,32'd25,32'd91,32'd4294967256,32'd17,32'd43,32'd4294967113,32'd32,32'd0,32'd4294967252,32'd3,32'd105,32'd22,32'd5,32'd4294967269,32'd2,32'd53,32'd33,32'd40,32'd86,32'd4294967197,32'd4294967289,32'd4294967074,32'd4294967294,32'd3,32'd25,32'd4294967266,32'd20,32'd4294967261,32'd12,32'd4294967272,32'd4294967295,32'd6,32'd4294967287,32'd104,32'd4294967104,32'd14,32'd61,32'd4294967269,32'd4294967217,32'd0,32'd19,32'd4294967229,32'd4294967279,32'd4,32'd4294967218,32'd4294967264,32'd127,32'd1,32'd96,32'd4294967018,32'd3,32'd4294966955,32'd59,32'd4294967266,32'd125,32'd4294967228,32'd4294967204,32'd5,32'd4294967159,32'd29,32'd26,32'd4294967254,32'd4294967294,32'd8,32'd33,32'd4294967121,32'd4294967188,32'd4294967208,32'd24,32'd6,32'd4294967229,32'd9,32'd26,32'd4294967261,32'd4294967239,32'd68,32'd37,32'd168,32'd74,32'd82,32'd3,32'd4294967268,32'd195,32'd0,32'd3,32'd32,32'd56,32'd4294967238,32'd4294967295,32'd31,32'd4294967086,32'd20,32'd4294967272,32'd35,32'd4294967270,32'd19,32'd4294967268,32'd62,32'd33,32'd4294967110,32'd4294967267,32'd98,32'd4294967247,32'd52,32'd4294967295,32'd15,32'd102,32'd8,32'd4294967247,32'd18,32'd4294967239,32'd4294967290,32'd4294967293,32'd20,32'd4294967253,32'd34,32'd76,32'd4,32'd3,32'd2,32'd4294967210,32'd37,32'd7,32'd4294967140,32'd4294967270,32'd31,32'd4294967295,32'd146,32'd138,32'd4294967294,32'd19,32'd160,32'd4294967268,32'd4294967208,32'd102,32'd4294967288,32'd2,32'd4294967205,32'd4294967291,32'd27,32'd4294967228,32'd4294967261,32'd4294967167,32'd26,32'd4294967227,32'd4294967283,32'd3,32'd4294967085,32'd4294967204,32'd33,32'd1,32'd4294967279,32'd4294967090,32'd4294967245,32'd13,32'd26,32'd4294967108,32'd4294967269,32'd77,32'd17,32'd4294967160,32'd4294967172,32'd4294967254,32'd102,32'd47,32'd49,32'd94,32'd95,32'd52,32'd68,32'd140,32'd4294967263,32'd36,32'd98,32'd4294967162,32'd29,32'd4294967292,32'd4294966949,32'd40,32'd118,32'd30,32'd4294967292,32'd20,32'd4294966996,32'd4294967253,32'd4294967259,32'd19,32'd130,32'd4294967075,32'd9,32'd4294967254,32'd4294967000,32'd32,32'd66,32'd22,32'd4294967160,32'd156,32'd139,32'd4294967258,32'd4294967293,32'd26,32'd4294967250,32'd130,32'd4294967137,32'd4294967213,32'd4294967262,32'd4294967281,32'd4294967293,32'd16,32'd4294967265,32'd6,32'd10,32'd43,32'd90,32'd4294967276,32'd2,32'd156,32'd4294967158,32'd19,32'd34,32'd4294967204,32'd9,32'd4294967244,32'd4294967206,32'd20,32'd4294967169,32'd110,32'd104,32'd4294967200,32'd4294967192,32'd35,32'd4294967122,32'd4294967111,32'd32,32'd48,32'd4294967091,32'd4294967241,32'd32,32'd23,32'd4294967256,32'd121,32'd4294967235,32'd108,32'd86,32'd4294967192,32'd16,32'd4294967075,32'd8,32'd4294967209,32'd58,32'd37,32'd51,32'd4294967217,32'd142,32'd19,32'd42,32'd4294967102,32'd4294967132,32'd4294967273,32'd0,32'd21,32'd4294967292,32'd4294967294,32'd4294967252,32'd4294967283,32'd5,32'd83,32'd196,32'd20,32'd4294967213,32'd40,32'd0,32'd24,32'd4294967242,32'd20,32'd5,32'd19,32'd4294967262,32'd41,32'd5,32'd21,32'd4294967234,32'd4,32'd8,32'd4294967076,32'd135,32'd25,32'd7,32'd31,32'd4294967260,32'd4294967269,32'd4294967264,32'd25,32'd4294967161,32'd91,32'd16,32'd4294967144,32'd8,32'd4294967012,32'd0,32'd24,32'd4294967103,32'd4294967229,32'd4294967295,32'd29,32'd4294967239,32'd56,32'd25,32'd4294967159,32'd4294967118,32'd49,32'd4294967224,32'd30,32'd4294967184,32'd22,32'd4294967221,32'd33,32'd4294967247,32'd34,32'd91,32'd4294967206,32'd65,32'd115,32'd74,32'd38,32'd105,32'd4294967198,32'd8,32'd4294967285,32'd1,32'd4294967053,32'd4294967268,32'd4294967290,32'd157,32'd29,32'd7,32'd4294967137,32'd48,32'd4294967098,32'd9,32'd23,32'd60,32'd31,32'd4294967081,32'd4294967282,32'd4294967247,32'd4294967104,32'd58,32'd4294967189,32'd133,32'd4294967294,32'd4294967255,32'd30,32'd65,32'd25,32'd4294967247,32'd4294967272,32'd13,32'd30,32'd5,32'd4294967082,32'd4294967236,32'd21,32'd55,32'd44,32'd6,32'd4294967237,32'd4294967132,32'd66,32'd4294967028,32'd4294967126,32'd23,32'd4294967171,32'd18,32'd4294967237,32'd76,32'd53,32'd4294967262,32'd4294967236,32'd24,32'd4294967283,32'd29,32'd39,32'd76,32'd4294967136,32'd64,32'd63,32'd122,32'd87,32'd16,32'd48,32'd4294967103,32'd72,32'd81,32'd8,32'd4294967186,32'd4294967161,32'd27,32'd103,32'd4294967213,32'd0,32'd57,32'd4294967227,32'd4294967163,32'd5,32'd4294967168,32'd8,32'd82,32'd4294967223,32'd63,32'd5,32'd17,32'd7,32'd4294967190,32'd4294967255,32'd31,32'd4294967098,32'd4294967273,32'd106,32'd4294967289,32'd15,32'd4294967208,32'd61,32'd79,32'd4294967230,32'd29,32'd4294967206,32'd4294967126,32'd25,32'd134,32'd4294967256,32'd4294967273,32'd146,32'd109,32'd4294967232,32'd46,32'd46,32'd68,32'd82,32'd71,32'd134,32'd4294967220,32'd4294967263,32'd4294967294,32'd66,32'd31,32'd68,32'd39,32'd4294967134,32'd30,32'd4294967261,32'd32,32'd4294967214,32'd4294967274,32'd4294967222,32'd4294967277,32'd12,32'd126,32'd4294967025,32'd50,32'd68,32'd2,32'd16,32'd100,32'd9,32'd25,32'd10,32'd18,32'd4294967210,32'd4294967189,32'd4294967254,32'd38,32'd109,32'd156,32'd168,32'd4294967268,32'd10,32'd87,32'd9,32'd4294967204,32'd20,32'd4294967091,32'd4294967229,32'd4294967105,32'd69,32'd6,32'd4294967173,32'd59,32'd162,32'd48,32'd95,32'd180,32'd139,32'd27,32'd4294967251,32'd4294967290,32'd5,32'd91,32'd35,32'd4294967134,32'd4294967150,32'd4294967261,32'd4294966991,32'd4294967135,32'd13,32'd50,32'd7,32'd81,32'd4294967258,32'd32,32'd4294967247,32'd23,32'd4294967087,32'd4294967181,32'd4294967124,32'd30,32'd35,32'd4294967278,32'd122,32'd150,32'd75,32'd66,32'd177,32'd98,32'd4294967159,32'd13,32'd138,32'd30,32'd36,32'd4294966957,32'd51,32'd4294967240,32'd4294966917,32'd123,32'd120,32'd197,32'd4294967289,32'd4294967257,32'd164,32'd30,32'd4294967096,32'd20,32'd4294967237,32'd155,32'd186,32'd4294967124,32'd135,32'd54,32'd106,32'd4294967092,32'd128,32'd188,32'd4294967102,32'd99,32'd146,32'd4294967228,32'd4294967271,32'd174,32'd4294967258,32'd4294967211,32'd119,32'd69,32'd58,32'd4294967017,32'd221,32'd90,32'd151,32'd4294967095,32'd109,32'd57,32'd56,32'd4294967056,32'd161,32'd151,32'd136,32'd170,32'd4294967012}
`define FEATURE_BELOW {32'd62,32'd4294967279,32'd4294967272,32'd4294967194,32'd14,32'd4294967290,32'd4294967218,32'd4294967276,32'd4294967289,32'd83,32'd4294967239,32'd4294967290,32'd25,32'd96,32'd9,32'd90,32'd24,32'd4294967273,32'd4294967291,32'd10,32'd4294967261,32'd4294967198,32'd33,32'd4294967274,32'd21,32'd4294967268,32'd4294967266,32'd82,32'd149,32'd4294967292,32'd4294967170,32'd4294967273,32'd43,32'd4294967279,32'd4294967169,32'd4,32'd33,32'd4294967272,32'd27,32'd4294967250,32'd5,32'd4294967146,32'd101,32'd4294967288,32'd4294967229,32'd47,32'd108,32'd4294967255,32'd4,32'd151,32'd17,32'd3,32'd4294967242,32'd4294967216,32'd0,32'd4294967269,32'd4294967247,32'd4294967105,32'd2,32'd156,32'd28,32'd4294967258,32'd4294967288,32'd4294967267,32'd4294967292,32'd4294967295,32'd20,32'd4294967275,32'd54,32'd4294967291,32'd28,32'd4294967236,32'd151,32'd100,32'd4294967250,32'd4294967266,32'd4294967196,32'd210,32'd4294967256,32'd4294967289,32'd57,32'd4294967272,32'd19,32'd4294967188,32'd36,32'd4294967251,32'd11,32'd4294967202,32'd20,32'd4294967263,32'd4,32'd4294967290,32'd69,32'd5,32'd18,32'd92,32'd7,32'd10,32'd4294967289,32'd122,32'd4294967287,32'd50,32'd89,32'd4294967271,32'd95,32'd4294967269,32'd3,32'd4294967176,32'd25,32'd42,32'd4294967272,32'd105,32'd150,32'd36,32'd44,32'd4294967288,32'd4294967225,32'd4294967253,32'd103,32'd4294967211,32'd18,32'd116,32'd65,32'd4294967265,32'd21,32'd4294967268,32'd4294967203,32'd4294967266,32'd129,32'd2,32'd4294967209,32'd4294967177,32'd25,32'd84,32'd7,32'd83,32'd4294967292,32'd4294967253,32'd81,32'd4294967295,32'd4294967274,32'd4294967275,32'd67,32'd4294967185,32'd4294967286,32'd4294967289,32'd66,32'd4294967118,32'd57,32'd4294967115,32'd15,32'd4294967278,32'd4294967202,32'd50,32'd149,32'd68,32'd4294967135,32'd9,32'd4,32'd74,32'd4294967241,32'd23,32'd30,32'd4294967289,32'd4294967284,32'd4294967274,32'd4294967224,32'd4294967228,32'd4294967261,32'd4294967254,32'd102,32'd4294967195,32'd4294967232,32'd3,32'd4294967226,32'd4294967262,32'd4294967195,32'd4294967111,32'd4294967228,32'd42,32'd4294967244,32'd37,32'd2,32'd2,32'd4,32'd4294967239,32'd17,32'd62,32'd4294967288,32'd5,32'd4294967232,32'd4,32'd4294967232,32'd5,32'd4294967266,32'd48,32'd12,32'd4294967244,32'd4294967177,32'd80,32'd13,32'd5,32'd4294967100,32'd0,32'd4294967291,32'd6,32'd4294967232,32'd16,32'd4294967255,32'd4294967273,32'd4294967261,32'd2,32'd4294967288,32'd16,32'd44,32'd4294967291,32'd4294967085,32'd59,32'd4294967277,32'd4294967294,32'd57,32'd4294966600,32'd4294967271,32'd9,32'd4294967290,32'd2,32'd103,32'd4294967182,32'd4294967227,32'd4294967231,32'd4294967292,32'd30,32'd4294967237,32'd46,32'd4294967181,32'd15,32'd4294967271,32'd29,32'd4294967275,32'd15,32'd4294967286,32'd20,32'd42,32'd26,32'd4294967278,32'd14,32'd117,32'd15,32'd4294967240,32'd4294967293,32'd42,32'd4294967281,32'd4294967292,32'd53,32'd4294967270,32'd4294967286,32'd4294967227,32'd74,32'd4294967268,32'd114,32'd4294967288,32'd4294967053,32'd5,32'd11,32'd4294967294,32'd15,32'd4294967290,32'd4294967215,32'd100,32'd4294967231,32'd4294967241,32'd25,32'd38,32'd4294967069,32'd4294967263,32'd3,32'd4294967158,32'd17,32'd4294967290,32'd46,32'd4294967261,32'd4,32'd4294967205,32'd4294967269,32'd4294967277,32'd21,32'd4294967251,32'd32,32'd4294967272,32'd13,32'd107,32'd4294967187,32'd4294967242,32'd4294967295,32'd4294967271,32'd57,32'd37,32'd4294967276,32'd4294967273,32'd4294967287,32'd4294967279,32'd36,32'd4294967192,32'd23,32'd125,32'd4294967222,32'd4294967289,32'd17,32'd4294967233,32'd85,32'd4294967241,32'd4294967291,32'd45,32'd24,32'd4294967294,32'd18,32'd4294967264,32'd42,32'd44,32'd2,32'd4,32'd4294967240,32'd66,32'd27,32'd139,32'd4294967250,32'd4294967269,32'd4294967294,32'd4294967287,32'd4294967259,32'd4294967272,32'd83,32'd4294967270,32'd1,32'd36,32'd94,32'd4294967168,32'd4294967292,32'd4294967180,32'd25,32'd4294967163,32'd18,32'd4294967265,32'd4294967275,32'd4294967170,32'd23,32'd4294967290,32'd19,32'd24,32'd302,32'd4294967189,32'd17,32'd32,32'd30,32'd4294967274,32'd4294967275,32'd96,32'd4294967227,32'd4294967265,32'd4294967294,32'd2,32'd4294967275,32'd75,32'd4294967262,32'd52,32'd4294967123,32'd4294967123,32'd14,32'd107,32'd165,32'd4294967215,32'd4294967229,32'd11,32'd4294967232,32'd1,32'd32,32'd68,32'd5,32'd4294967264,32'd43,32'd4294967269,32'd4294967116,32'd37,32'd4294967291,32'd5,32'd34,32'd4294967146,32'd21,32'd4294967186,32'd4294967288,32'd61,32'd4294967260,32'd4294967114,32'd19,32'd4294967143,32'd4294967168,32'd7,32'd36,32'd4294967268,32'd32,32'd86,32'd60,32'd4294967195,32'd4294967251,32'd97,32'd4294967265,32'd4294967234,32'd33,32'd4294967236,32'd4294967235,32'd4294967208,32'd4294967280,32'd162,32'd4,32'd19,32'd4294967269,32'd18,32'd4294967263,32'd139,32'd4294967213,32'd4294967288,32'd4294967276,32'd4294967292,32'd4294967265,32'd4294963456,32'd4294967062,32'd4294967217,32'd153,32'd46,32'd4294967294,32'd2,32'd4294967277,32'd20,32'd4294967219,32'd5,32'd34,32'd62,32'd4294967227,32'd4294967167,32'd4294967273,32'd4294967291,32'd40,32'd44,32'd4294967288,32'd19,32'd4294967273,32'd4294967245,32'd4294967277,32'd0,32'd4294967273,32'd4294967255,32'd149,32'd10,32'd1,32'd4294967252,32'd4294967291,32'd17,32'd58,32'd61,32'd4294967231,32'd18,32'd4294967256,32'd40,32'd4294967270,32'd4294967240,32'd24,32'd56,32'd4294967290,32'd4294967265,32'd63,32'd20,32'd4294967244,32'd152,32'd4294967079,32'd3,32'd4294967275,32'd25,32'd4294967214,32'd4294966817,32'd4294967198,32'd59,32'd4294967291,32'd30,32'd4,32'd4294967285,32'd66,32'd4294966834,32'd4294967225,32'd4294967252,32'd4294967276,32'd91,32'd20,32'd7,32'd4294967274,32'd17,32'd4294967270,32'd4294967183,32'd4294967266,32'd7,32'd4294967290,32'd4294967230,32'd54,32'd4294967271,32'd119,32'd142,32'd4294967205,32'd19,32'd4294967276,32'd17,32'd4294967197,32'd4294967271,32'd4294967164,32'd18,32'd9,32'd45,32'd4294967292,32'd119,32'd32,32'd4294967274,32'd4294967226,32'd4294967276,32'd65,32'd18,32'd4294967166,32'd102,32'd216,32'd89,32'd4294967236,32'd17,32'd4294967074,32'd14,32'd16,32'd4294967289,32'd74,32'd4294967234,32'd4294967211,32'd4294967222,32'd4294967159,32'd26,32'd4294967294,32'd4294967263,32'd75,32'd24,32'd102,32'd8,32'd4294967211,32'd4294967256,32'd116,32'd78,32'd31,32'd4294967288,32'd12,32'd25,32'd4294967181,32'd18,32'd66,32'd4294967177,32'd20,32'd108,32'd4294967261,32'd6,32'd2,32'd50,32'd4294967275,32'd4294967205,32'd4294967276,32'd9,32'd54,32'd4294967292,32'd4294967189,32'd22,32'd86,32'd26,32'd4294967292,32'd4294967262,32'd4294967248,32'd74,32'd4294967187,32'd58,32'd132,32'd29,32'd4294967204,32'd4294967207,32'd4294967256,32'd4294967085,32'd4294967150,32'd4294967218,32'd4294967145,32'd76,32'd4294967233,32'd4294967220,32'd4294967157,32'd17,32'd4294967271,32'd4294967106,32'd19,32'd29,32'd4294967275,32'd43,32'd4294967237,32'd4294967266,32'd5,32'd4294967272,32'd61,32'd91,32'd4294967267,32'd4294967273,32'd4294967247,32'd4294967248,32'd4294967181,32'd28,32'd117,32'd4294967274,32'd595,32'd4294967273,32'd21,32'd4294967288,32'd4294967090,32'd4294967289,32'd20,32'd4294967271,32'd93,32'd4294967260,32'd15,32'd4294967272,32'd77,32'd14,32'd4294967284,32'd131,32'd17,32'd4294967050,32'd4294967096,32'd51,32'd60,32'd4294967293,32'd17,32'd4294967056,32'd31,32'd4294967183,32'd97,32'd4294967276,32'd41,32'd4294967276,32'd4294967220,32'd4294967272,32'd4294967247,32'd4294967256,32'd63,32'd4294967150,32'd17,32'd4294967176,32'd22,32'd4294967293,32'd48,32'd4294966790,32'd165,32'd4294967268,32'd29,32'd4294967279,32'd122,32'd5,32'd4294967284,32'd7,32'd178,32'd223,32'd123,32'd4294967252,32'd18,32'd4294967268,32'd4294967228,32'd4294967292,32'd4294967224,32'd4294967291,32'd4294966840,32'd4294967224,32'd21,32'd4294967269,32'd60,32'd30,32'd6,32'd4294967170,32'd4294967257,32'd4294967259,32'd18,32'd19,32'd7,32'd4294967237,32'd22,32'd6,32'd23,32'd4294967232,32'd4294967293,32'd51,32'd27,32'd4294967238,32'd4294967202,32'd4294967293,32'd4294967278,32'd4294967193,32'd4294967060,32'd20,32'd21,32'd103,32'd16,32'd4294967273,32'd4294967123,32'd4294967291,32'd15,32'd107,32'd29,32'd4294967170,32'd4294967239,32'd10,32'd82,32'd37,32'd44,32'd4294967260,32'd282,32'd51,32'd5,32'd4294967239,32'd4294967260,32'd4294967277,32'd23,32'd4294967269,32'd66,32'd4294967269,32'd4294967235,32'd4294967164,32'd83,32'd162,32'd0,32'd4294967271,32'd19,32'd23,32'd3,32'd55,32'd31,32'd4294967277,32'd72,32'd44,32'd4294967223,32'd37,32'd56,32'd4294967031,32'd4294967285,32'd125,32'd4294967278,32'd4294967293,32'd74,32'd4294967273,32'd4294967240,32'd4294967175,32'd2,32'd4294967290,32'd128,32'd93,32'd0,32'd0,32'd120,32'd26,32'd21,32'd4294967273,32'd4294967282,32'd4294967289,32'd15,32'd25,32'd92,32'd4294967295,32'd4294967226,32'd4294967178,32'd109,32'd0,32'd49,32'd4294967260,32'd122,32'd9,32'd4294967280,32'd87,32'd4294967200,32'd9,32'd4294967205,32'd4294967173,32'd22,32'd3,32'd47,32'd59,32'd4294967237,32'd4294967214,32'd4294967255,32'd4294967193,32'd4294967268,32'd82,32'd4294967290,32'd18,32'd4294967125,32'd53,32'd4294967205,32'd147,32'd20,32'd4294967262,32'd40,32'd21,32'd4294967244,32'd17,32'd4294967262,32'd11,32'd4294967199,32'd25,32'd37,32'd32,32'd4294967267,32'd4294967257,32'd4294967280,32'd4294967237,32'd79,32'd28,32'd4294967273,32'd9,32'd4294967147,32'd165,32'd4294967287,32'd4294967268,32'd4294967274,32'd3,32'd4294967242,32'd4294967034,32'd4294967294,32'd4294967218,32'd4294967195,32'd14,32'd134,32'd4294967278,32'd4294967273,32'd22,32'd108,32'd17,32'd4294967271,32'd5,32'd57,32'd27,32'd86,32'd15,32'd10,32'd4294967164,32'd18,32'd113,32'd4294967109,32'd4294966902,32'd35,32'd9,32'd4294967276,32'd34,32'd4294967238,32'd4294967273,32'd4294967293,32'd4294967287,32'd4294967275,32'd19,32'd4294967276,32'd24,32'd4294967292,32'd4294967266,32'd4294967248,32'd19,32'd91,32'd8,32'd4294967294,32'd18,32'd120,32'd8,32'd4294966961,32'd32,32'd4294967224,32'd4294967288,32'd4294967278,32'd4294966900,32'd4294967247,32'd220,32'd4294967246,32'd20,32'd4294967267,32'd4294967045,32'd84,32'd37,32'd4294967157,32'd52,32'd4294967220,32'd17,32'd4,32'd4294967287,32'd4294967210,32'd4294967190,32'd34,32'd4294967290,32'd58,32'd43,32'd4294967210,32'd9,32'd84,32'd0,32'd4294967128,32'd15,32'd4294967092,32'd29,32'd98,32'd4294967288,32'd4294967126,32'd21,32'd109,32'd96,32'd4294967223,32'd26,32'd25,32'd4294967292,32'd4294967216,32'd4294967254,32'd4294967288,32'd24,32'd26,32'd2,32'd0,32'd4294967274,32'd4294967235,32'd101,32'd4294967293,32'd4294967263,32'd50,32'd4294967282,32'd4294967228,32'd23,32'd4294967294,32'd17,32'd18,32'd140,32'd4294967147,32'd112,32'd4294967246,32'd68,32'd51,32'd4294967241,32'd11,32'd4294967214,32'd4294967271,32'd10,32'd4294967101,32'd4294967289,32'd69,32'd4294967182,32'd49,32'd4294967281,32'd4294967254,32'd23,32'd4294967267,32'd84,32'd4294967185,32'd4294967153,32'd4294967257,32'd65,32'd4294967160,32'd4294967236,32'd4294967212,32'd4294967284,32'd0,32'd4294967224,32'd3,32'd81,32'd4294967169,32'd33,32'd4294967184,32'd4294967127,32'd4294967259,32'd45,32'd54,32'd83,32'd4294967155,32'd21,32'd53,32'd4294967233,32'd4294967261,32'd4294967238,32'd3,32'd4294967158,32'd23,32'd4294967201,32'd4294967221,32'd92,32'd4294967227,32'd34,32'd32,32'd40,32'd4294967186,32'd29,32'd33,32'd4294967136,32'd4294967269,32'd6,32'd169,32'd181,32'd4294967290,32'd24,32'd4294967271,32'd5,32'd4294967224,32'd111,32'd4294967198,32'd51,32'd64,32'd4294967042,32'd5,32'd73,32'd4294967203,32'd19,32'd4294967191,32'd103,32'd4294967290,32'd22,32'd4294967266,32'd24,32'd98,32'd41,32'd4294967286,32'd2,32'd221,32'd37,32'd4294967195,32'd26,32'd4294967289,32'd21,32'd4294967211,32'd17,32'd4294967141,32'd4294967258,32'd42,32'd4294967288,32'd24,32'd4294967171,32'd10,32'd4294967257,32'd4294967252,32'd4294967288,32'd4294967217,32'd4294967292,32'd47,32'd70,32'd4294967277,32'd4294967187,32'd4294967196,32'd4294967111,32'd160,32'd4294967203,32'd4294967267,32'd118,32'd4294967205,32'd20,32'd249,32'd4294967279,32'd4294967262,32'd4294967290,32'd4294967141,32'd37,32'd4294967236,32'd4294967285,32'd57,32'd83,32'd4294967209,32'd4294967277,32'd58,32'd4294967267,32'd4294967151,32'd22,32'd4294967290,32'd17,32'd4294967273,32'd1,32'd4294967264,32'd4294967287,32'd4294967269,32'd4294967234,32'd113,32'd4294967229,32'd4294967277,32'd23,32'd3,32'd4294967281,32'd4294967268,32'd18,32'd4294967266,32'd4294967294,32'd4294967110,32'd40,32'd4294967261,32'd308,32'd4294967007,32'd22,32'd1,32'd24,32'd4294967274,32'd4294967205,32'd4294967052,32'd32,32'd4294967269,32'd2,32'd23,32'd4294967270,32'd4294967232,32'd4294967269,32'd4294967244,32'd4294967287,32'd4294967231,32'd4294967271,32'd22,32'd83,32'd4294967229,32'd15,32'd4294967249,32'd4294967288,32'd4294967292,32'd4294967280,32'd4294967275,32'd4294967290,32'd25,32'd18,32'd4294967193,32'd35,32'd142,32'd14,32'd4294967197,32'd21,32'd4294967098,32'd6,32'd4294967276,32'd4294967157,32'd4294967268,32'd4294967277,32'd5,32'd4294967249,32'd3,32'd4294967221,32'd4294967229,32'd4294967295,32'd44,32'd4294967295,32'd3,32'd84,32'd4294967289,32'd4294967293,32'd125,32'd4,32'd4294967174,32'd39,32'd4294967295,32'd4294967273,32'd4294967268,32'd4294967068,32'd4294967291,32'd30,32'd4294967272,32'd4294967233,32'd4294967189,32'd34,32'd4294967291,32'd4294967113,32'd4294967249,32'd4294967295,32'd0,32'd26,32'd4294967244,32'd4294967283,32'd4294967195,32'd4294967284,32'd31,32'd4294967198,32'd4294967295,32'd4294967256,32'd2,32'd4294967226,32'd121,32'd4294967278,32'd14,32'd4294967255,32'd4294967254,32'd4294967232,32'd4294967227,32'd68,32'd4,32'd4294967163,32'd57,32'd4294967154,32'd43,32'd4294967219,32'd4294966921,32'd65,32'd4294966976,32'd43,32'd18,32'd4294967185,32'd25,32'd4294967295,32'd83,32'd4294967076,32'd14,32'd4294967269,32'd4294967270,32'd4294967161,32'd4294967281,32'd0,32'd20,32'd306,32'd69,32'd31,32'd22,32'd82,32'd111,32'd4294967255,32'd26,32'd4294967288,32'd23,32'd57,32'd3,32'd4294967225,32'd4,32'd4294967118,32'd4294967192,32'd206,32'd18,32'd4294967272,32'd4294967058,32'd4294967278,32'd10,32'd10,32'd4294967295,32'd4294967292,32'd31,32'd4294967268,32'd38,32'd135,32'd2,32'd4294967214,32'd45,32'd4294967272,32'd96,32'd19,32'd53,32'd4294967237,32'd4294967261,32'd4294967273,32'd30,32'd4294967238,32'd4294967270,32'd4294967292,32'd4294967079,32'd4294967270,32'd52,32'd4294967272,32'd4294967294,32'd3,32'd27,32'd4294967273,32'd4294967294,32'd2,32'd4294967227,32'd4294967262,32'd118,32'd4294967270,32'd4294967286,32'd15,32'd4294967235,32'd4294967210,32'd4294967147,32'd4294967182,32'd240,32'd63,32'd4294967245,32'd4294967147,32'd18,32'd4294967263,32'd4294967253,32'd169,32'd81,32'd4294967144,32'd92,32'd4294967157,32'd22,32'd4294967262,32'd50,32'd4294967266,32'd4294967265,32'd4294967292,32'd4294967273,32'd4294967288,32'd4294967188,32'd4294967217,32'd80,32'd67,32'd7,32'd4294967187,32'd43,32'd4294967275,32'd6,32'd4294967139,32'd41,32'd60,32'd4294967293,32'd50,32'd90,32'd4294967217,32'd0,32'd4294967295,32'd212,32'd4294967295,32'd23,32'd4294967239,32'd4294967259,32'd44,32'd4294967164,32'd4294967215,32'd23,32'd59,32'd4294967207,32'd4294967264,32'd4294967260,32'd4294967206,32'd4294967173,32'd4294967293,32'd4294967290,32'd6,32'd4294967198,32'd58,32'd4294967198,32'd4294967214,32'd4294967260,32'd80,32'd21,32'd4294967182,32'd4294967143,32'd4294967253,32'd69,32'd4294967191,32'd4294967294,32'd129,32'd4294967205,32'd6,32'd172,32'd4294967233,32'd4294967269,32'd4294967208,32'd4294967255,32'd4294967252,32'd4294967261,32'd4294967186,32'd4294967249,32'd91,32'd4294967270,32'd87,32'd9,32'd4294967294,32'd4294967227,32'd4294967271,32'd58,32'd3,32'd4,32'd4294967279,32'd4294967262,32'd44,32'd4294967289,32'd4294967294,32'd4294967288,32'd100,32'd4294967158,32'd4294967220,32'd4294967273,32'd19,32'd4294967295,32'd7,32'd4294967288,32'd4294967220,32'd4294967287,32'd132,32'd4,32'd5,32'd4294967290,32'd5,32'd4294967288,32'd16,32'd4294967174,32'd40,32'd28,32'd21,32'd4294967264,32'd4294966968,32'd4294967226,32'd4294967262,32'd248,32'd24,32'd4294967225,32'd4294967284,32'd25,32'd4294967269,32'd4294967180,32'd4294967294,32'd4294967295,32'd31,32'd182,32'd45,32'd4294967295,32'd4294967222,32'd61,32'd4294966944,32'd48,32'd4294967294,32'd0,32'd176,32'd4294967254,32'd2,32'd74,32'd26,32'd4294967295,32'd15,32'd4294967251,32'd4294967203,32'd4294967262,32'd12,32'd29,32'd54,32'd4294967219,32'd1,32'd4294967263,32'd72,32'd4294967186,32'd22,32'd4294967263,32'd26,32'd125,32'd31,32'd4294967292,32'd66,32'd4294967236,32'd16,32'd108,32'd25,32'd4294967115,32'd4294967198,32'd4294967270,32'd57,32'd4294967295,32'd4294967268,32'd0,32'd4294967269,32'd4,32'd3,32'd4294967144,32'd4294967232,32'd81,32'd4294967227,32'd164,32'd21,32'd25,32'd4294967267,32'd4294967199,32'd35,32'd4294967267,32'd21,32'd4294967294,32'd4294967146,32'd76,32'd76,32'd4294967292,32'd0,32'd46,32'd4294967288,32'd4294967187,32'd3,32'd38,32'd97,32'd4294967151,32'd17,32'd4294967292,32'd78,32'd4294967188,32'd4294967176,32'd8,32'd4294967285,32'd79,32'd4294967166,32'd115,32'd4294967163,32'd122,32'd4294967157,32'd5,32'd4294967234,32'd4294967169,32'd4294967281,32'd4294967253,32'd17,32'd185,32'd4294967275,32'd18,32'd4294967192,32'd4294967193,32'd4294967224,32'd4294967218,32'd4294967222,32'd30,32'd35,32'd42,32'd4294967175,32'd4294967236,32'd4294967270,32'd18,32'd4294967278,32'd18,32'd5,32'd4294967210,32'd4294967195,32'd4294967187,32'd51,32'd78,32'd63,32'd30,32'd232,32'd15,32'd4294967238,32'd4294967288,32'd124,32'd4294967271,32'd4294967288,32'd30,32'd4294967184,32'd44,32'd4294967207,32'd23,32'd4294967266,32'd81,32'd4294967268,32'd77,32'd4294967269,32'd4294967047,32'd6,32'd4294967175,32'd107,32'd104,32'd4294967248,32'd25,32'd4294967277,32'd17,32'd4294967292,32'd17,32'd4294967139,32'd9,32'd4294967204,32'd4294967001,32'd155,32'd4294967238,32'd4294967288,32'd4294967227,32'd19,32'd15,32'd37,32'd14,32'd4294967292,32'd4294967293,32'd54,32'd1,32'd4294967292,32'd4294967293,32'd4294967272,32'd4294967262,32'd59,32'd4294967211,32'd4294966997,32'd43,32'd58,32'd6,32'd23,32'd4294967216,32'd2,32'd4294967289,32'd0,32'd4294967196,32'd4294967229,32'd84,32'd4294967294,32'd4294967139,32'd4294967254,32'd4294967293,32'd4294967260,32'd60,32'd14,32'd4294967293,32'd4294967291,32'd4294967251,32'd4294967292,32'd33,32'd4294967209,32'd19,32'd49,32'd20,32'd86,32'd4294967283,32'd48,32'd4294967295,32'd4294967149,32'd4294967291,32'd78,32'd4294967191,32'd4294967266,32'd4294967288,32'd150,32'd64,32'd4294967273,32'd26,32'd4294967269,32'd4294967193,32'd4294967293,32'd19,32'd4294967290,32'd4294967282,32'd4294967261,32'd4294967267,32'd4294967245,32'd12,32'd4294967292,32'd22,32'd5,32'd4294967286,32'd4294967176,32'd31,32'd80,32'd23,32'd4294967227,32'd4294967261,32'd4294967147,32'd4294967290,32'd4294967256,32'd30,32'd4294967295,32'd15,32'd354,32'd22,32'd4294967203,32'd4294967205,32'd4294967192,32'd19,32'd103,32'd113,32'd4294966986,32'd37,32'd30,32'd4294967129,32'd4294967258,32'd4294967244,32'd4294967271,32'd4294967155,32'd4294967187,32'd4294967209,32'd152,32'd50,32'd2,32'd4294967230,32'd58,32'd4294967259,32'd4294967213,32'd4294967259,32'd28,32'd4294967247,32'd73,32'd73,32'd20,32'd4294967264,32'd21,32'd4294967216,32'd20,32'd4294967270,32'd41,32'd4294967269,32'd17,32'd58,32'd24,32'd4294967272,32'd19,32'd39,32'd86,32'd4294967210,32'd34,32'd4294967289,32'd4294967266,32'd4294967194,32'd4294967272,32'd4294967188,32'd23,32'd4294967290,32'd4294967217,32'd4294967273,32'd11,32'd4294967246,32'd3,32'd4294967264,32'd17,32'd17,32'd4294967238,32'd4294967186,32'd4294967293,32'd66,32'd19,32'd4294967294,32'd75,32'd4294967291,32'd70,32'd4294967075,32'd49,32'd4294967186,32'd4294967030,32'd109,32'd4294967295,32'd4294967292,32'd4294967213,32'd89,32'd4294967292,32'd4294967259,32'd4294967278,32'd4294967183,32'd45,32'd107,32'd4294967144,32'd4294967274,32'd67,32'd4294967250,32'd79,32'd2,32'd16,32'd4294967133,32'd4294967287,32'd4294967270,32'd22,32'd4294967288,32'd61,32'd4294967131,32'd4294967287,32'd4294967192,32'd15,32'd4294967183,32'd4294967196,32'd131,32'd4294967282,32'd4294967274,32'd4294967131,32'd4294967228,32'd4294967218,32'd4294967258,32'd79,32'd4294967192,32'd30,32'd4294967142,32'd4294967286,32'd30,32'd4294967219,32'd4294967233,32'd4294967233,32'd74,32'd4294967291,32'd4294967205,32'd4294967119,32'd4294967129,32'd22,32'd4294967097,32'd4294967094,32'd200,32'd1,32'd4294967224,32'd4294967120,32'd4294967257,32'd4294967217,32'd6,32'd4294967220,32'd4294967208,32'd32,32'd4294967204,32'd135,32'd4294967256,32'd4294967241,32'd65,32'd22,32'd4294967093,32'd77,32'd110,32'd114,32'd4294967247,32'd4294967284,32'd56,32'd56,32'd5,32'd20,32'd4294967149,32'd20,32'd4294967184,32'd4294967265,32'd4294967244,32'd49,32'd4294967115,32'd4294967195,32'd4294967224,32'd119,32'd4294967192,32'd20,32'd92,32'd311,32'd4294967144,32'd1,32'd18,32'd4294967202,32'd4294967177,32'd30,32'd4294967275,32'd27,32'd4294967171,32'd4294967081,32'd4294967246,32'd147,32'd4294967254,32'd4294967290,32'd279,32'd14,32'd4294967292,32'd4294967241,32'd105,32'd25,32'd4294967276,32'd4294967203,32'd4294967254,32'd4294967244,32'd4294967290,32'd15,32'd4294967274,32'd27,32'd4294967290,32'd49,32'd60,32'd4294967265,32'd4294967257,32'd0,32'd4294967289,32'd4294967254,32'd32,32'd29,32'd4294967264,32'd156,32'd4294967294,32'd15,32'd4294967268,32'd4294967231,32'd4294967265,32'd20,32'd4294967226,32'd69,32'd4294967178,32'd4294967289,32'd4294967213,32'd4294967274,32'd4294967112,32'd33,32'd39,32'd1,32'd84,32'd4294967192,32'd4294967130,32'd4294966935,32'd4294967185,32'd21,32'd29,32'd1,32'd122,32'd4294966591,32'd4294967163,32'd49,32'd4294967171,32'd4294967282,32'd4294967264,32'd19,32'd4294967253,32'd4294967213,32'd3,32'd4294967222,32'd4294967295,32'd4294967247,32'd4294967229,32'd4294967277,32'd4294967272,32'd23,32'd4294967262,32'd4294967286,32'd4294967294,32'd4294967237,32'd4294967295,32'd40,32'd4294967271,32'd14,32'd4294967295,32'd4294967259,32'd4294967264,32'd21,32'd81,32'd4294967164,32'd4294967261,32'd4294967176,32'd6,32'd4294967264,32'd4294967113,32'd53,32'd0,32'd36,32'd4294967245,32'd4294967277,32'd22,32'd20,32'd75,32'd4294967291,32'd4294967264,32'd146,32'd9,32'd69,32'd4294967110,32'd4294967152,32'd4294967264,32'd4294967286,32'd4294967185,32'd4294967289,32'd75,32'd4294967132,32'd4294967177,32'd4294967187,32'd58,32'd52,32'd4294967266,32'd65,32'd4294967235,32'd4294967242,32'd4294967232,32'd4294967180,32'd84,32'd4294967277,32'd11,32'd4294967165,32'd6,32'd4294967124,32'd8,32'd13,32'd4294967156,32'd4294967278,32'd4294967174,32'd4294967270,32'd27,32'd4294967289,32'd4294967066,32'd4294967256,32'd39,32'd4294967293,32'd22,32'd4294967036,32'd58,32'd4294967289,32'd4294967282,32'd4294967260,32'd38,32'd4294967210,32'd22,32'd7,32'd4294967223,32'd78,32'd4294967289,32'd4294967211,32'd4294967291,32'd4294967294,32'd4294967281,32'd264,32'd4294967271,32'd4294967292,32'd109,32'd4294967215,32'd4294967198,32'd4294967057,32'd283,32'd4294967145,32'd4294967112,32'd4294967251,32'd42,32'd4294967291,32'd4294967259,32'd4294967295,32'd33,32'd4294967268,32'd24,32'd137,32'd4294967283,32'd4294967294,32'd4294967207,32'd98,32'd4294967253,32'd176,32'd19,32'd4294967275,32'd4294967242,32'd4294967248,32'd0,32'd4294967179,32'd4294967243,32'd86,32'd162,32'd4294967274,32'd72,32'd5,32'd4294967293,32'd147,32'd4294967285,32'd4294967246,32'd4294966781,32'd4294967234,32'd78,32'd4294967274,32'd4294967252,32'd15,32'd17,32'd49,32'd77,32'd4294967262,32'd4294967290,32'd36,32'd4294967156,32'd4294967143,32'd22,32'd4294967293,32'd26,32'd4294967099,32'd45,32'd4294967148,32'd27,32'd53,32'd130,32'd4294967154,32'd61,32'd4294967270,32'd4294967295,32'd88,32'd26,32'd4294967267,32'd4,32'd4294967265,32'd4294967129,32'd20,32'd58,32'd1,32'd43,32'd5,32'd4294967274,32'd4294967107,32'd28,32'd20,32'd24,32'd4294967245,32'd29,32'd4294967180,32'd27,32'd4294967257,32'd158,32'd104,32'd4294967174,32'd86,32'd27,32'd4294967236,32'd4294967204,32'd4294967159,32'd4294967225,32'd46,32'd4294967224,32'd4294967181,32'd87,32'd70,32'd23,32'd51,32'd4294967292,32'd4294967222,32'd4294967169,32'd192,32'd4294967252,32'd4294967295,32'd4294967236,32'd0,32'd4294967295,32'd14,32'd17,32'd4294967276,32'd46,32'd8,32'd4294967120,32'd42,32'd4294967194,32'd118,32'd38,32'd4294967207,32'd70,32'd4294967273,32'd4294967263,32'd4294967290,32'd28,32'd4294967097,32'd50,32'd19,32'd1,32'd8,32'd4294967292,32'd23,32'd4294967207,32'd4294967264,32'd245,32'd4294967265,32'd4294967295,32'd10,32'd4294967090,32'd4294967257,32'd2,32'd2,32'd4294967262,32'd103,32'd4294967154,32'd15,32'd42,32'd24,32'd4294967261,32'd37,32'd18,32'd4294967102,32'd4294967162,32'd17,32'd4294967265,32'd19,32'd4294967160,32'd43,32'd4294967294,32'd87,32'd4294967239,32'd4294967272,32'd4294967291,32'd177,32'd4294967135,32'd42,32'd104,32'd4294967244,32'd95,32'd19,32'd4294967256,32'd4294967077,32'd4294967121,32'd21,32'd31,32'd4294967230,32'd117,32'd74,32'd4294967203,32'd4294967244,32'd4294967132,32'd4294967050,32'd4294967293,32'd4294967246,32'd9,32'd25,32'd4294967255,32'd73,32'd228,32'd1,32'd4294967180,32'd17,32'd105,32'd4294967295,32'd35,32'd4294967286,32'd75,32'd63,32'd4294967250,32'd4294967159,32'd4294967146,32'd15,32'd4294967140,32'd4294967191,32'd156,32'd175,32'd4294967259,32'd20,32'd36,32'd4294967212,32'd0,32'd4294967283,32'd30,32'd4294967284,32'd4294967169,32'd4294967231,32'd4294967162,32'd4294967231,32'd42,32'd4294967144,32'd4294967249,32'd4294967192,32'd4294967187,32'd4294967217,32'd21,32'd3,32'd20,32'd49,32'd7,32'd4294967261,32'd6,32'd9,32'd24,32'd3,32'd16,32'd36,32'd4294967289,32'd4294967291,32'd4294967283,32'd4294967275,32'd20,32'd100,32'd232,32'd4294967271,32'd25,32'd4294967271,32'd62,32'd4294967050,32'd4294967286,32'd5,32'd4294967292,32'd4294967160,32'd4294967293,32'd155,32'd4294967294,32'd48,32'd4294967194,32'd4294967269,32'd39,32'd223,32'd88,32'd8,32'd4294967268,32'd4294967226,32'd18,32'd151,32'd4294967265,32'd4294967073,32'd12,32'd25,32'd29,32'd4294967253,32'd81,32'd4294967079,32'd10,32'd5,32'd1,32'd4294967265,32'd4294967074,32'd4294967294,32'd4294967278,32'd4294967294,32'd19,32'd6,32'd4294967168,32'd4294967258,32'd48,32'd4294967007,32'd4294967112,32'd4294967258,32'd48,32'd4294967140,32'd4294967233,32'd0,32'd4294967117,32'd4294967271,32'd45,32'd4294967180,32'd4294967290,32'd4294967270,32'd103,32'd101,32'd3,32'd4294967240,32'd4294967179,32'd4294967261,32'd4294967226,32'd4294967145,32'd34,32'd4294967257,32'd4294967267,32'd4294967185,32'd4294967205,32'd118,32'd4294967228,32'd4294967176,32'd4294967252,32'd4294967180,32'd4294967201,32'd30,32'd44,32'd11,32'd42,32'd74,32'd4294967217,32'd4294967260,32'd34,32'd118,32'd4294967200,32'd4294967186,32'd151,32'd4294967247,32'd4294967222,32'd15,32'd4294967177,32'd4294967221,32'd4294967243,32'd4294967166,32'd78,32'd4294967283,32'd125,32'd4294967213,32'd4294967244,32'd89,32'd4294967291,32'd83,32'd1,32'd4294967283,32'd122,32'd0,32'd29,32'd4294966903,32'd123,32'd47,32'd4294967175,32'd24,32'd8,32'd4294967267,32'd4294967264,32'd53,32'd4294967230,32'd4294967262,32'd4294967294,32'd4294967290,32'd4294967131,32'd23,32'd4294967176,32'd6,32'd4294967219,32'd117,32'd124,32'd76,32'd4294967257,32'd4294967221,32'd4294967248,32'd4294967279,32'd7,32'd87,32'd4294967293,32'd104,32'd4294967158,32'd4294967152,32'd85,32'd4294967217,32'd77,32'd382,32'd207,32'd66,32'd4294967163,32'd32,32'd4294967266,32'd24,32'd4294967209,32'd4294967272,32'd125,32'd26,32'd4294967128,32'd4294967193,32'd33,32'd59,32'd4294967171,32'd21,32'd98,32'd4,32'd4294967100,32'd0,32'd4294967292,32'd128,32'd4294967292,32'd4294967272,32'd136,32'd4294967289,32'd25,32'd33,32'd4294967151,32'd22,32'd4294967229,32'd4294967173,32'd61,32'd126,32'd4294967171,32'd4294967275,32'd3,32'd20,32'd21,32'd4294967186,32'd4294967131,32'd37,32'd4294967162,32'd4294967108,32'd117,32'd59,32'd4294967242,32'd4294967181,32'd4294967257,32'd4294967195,32'd4294967180,32'd4294967171,32'd56,32'd4294967275,32'd89,32'd4294967186,32'd4294967265,32'd4294967260,32'd19,32'd4294967139,32'd4294967226,32'd4294967293,32'd4294967222,32'd145,32'd2,32'd106,32'd4294967181,32'd100,32'd4294967286,32'd4294967249,32'd16,32'd96,32'd4294967285,32'd33,32'd4294967276,32'd4294967143,32'd4294967093,32'd4294967267,32'd177,32'd37,32'd4294967104,32'd22,32'd99,32'd4294967034,32'd4294967129,32'd48,32'd4294967214,32'd4294967260,32'd126,32'd4294967151,32'd60,32'd7,32'd4294967250,32'd4294967203,32'd25,32'd108,32'd4294967213,32'd4294967122,32'd4294967293,32'd4294967271,32'd105,32'd4294967228,32'd1,32'd123,32'd23,32'd4294967260,32'd107,32'd4294967149,32'd27,32'd4294966902,32'd4294967081,32'd25,32'd47,32'd5,32'd4294967177,32'd24,32'd81,32'd4294967145,32'd17,32'd15,32'd4294967192,32'd4294967108,32'd129,32'd2,32'd27,32'd4294967182,32'd4294967240,32'd3,32'd76,32'd4294967255,32'd4294967041,32'd20,32'd34,32'd108,32'd4294967283,32'd4294967226,32'd4294967206,32'd4294967247,32'd4294967244,32'd4294967153,32'd4294967205,32'd4294967224,32'd91,32'd4294967219,32'd4294967263,32'd29,32'd4294967235,32'd76,32'd4294967292,32'd4294967259,32'd4294967267,32'd4294967263,32'd4294967008,32'd4294967195,32'd4294967292,32'd54,32'd63,32'd4294967127,32'd4294967269,32'd18,32'd4294967168,32'd48,32'd4294967292,32'd4294967219,32'd4294967258,32'd4294967233,32'd6,32'd4294967289,32'd4294967264,32'd51,32'd4294967038,32'd4294967174,32'd58,32'd4294967295,32'd2,32'd32,32'd87,32'd73,32'd4294967023,32'd4294967105,32'd99,32'd218,32'd4294967195,32'd4294967286,32'd4294967263,32'd47,32'd4294967127,32'd4294967292,32'd6,32'd4294967019,32'd4294967235,32'd22,32'd4294967150,32'd25,32'd17,32'd4294967177,32'd8,32'd4294967283,32'd4294967261,32'd27,32'd12,32'd4294967179,32'd6,32'd26,32'd4294967228,32'd4294967229,32'd4,32'd20,32'd4294967220,32'd4294967190,32'd96,32'd0,32'd51,32'd4294967282,32'd4294967255,32'd42,32'd4294967140,32'd30,32'd4294967076,32'd39,32'd4294967223,32'd4294967150,32'd4294967165,32'd130,32'd4294967216,32'd4294967041,32'd4294967244,32'd20,32'd3,32'd54,32'd4294967107,32'd4294967214,32'd4294967018,32'd125,32'd61,32'd44,32'd4294967158,32'd4294967282,32'd4294967272,32'd4294967215,32'd25,32'd4294967211,32'd4294967092,32'd4294967178,32'd54,32'd4294967156,32'd4294967162,32'd4294967148,32'd106,32'd4294967274,32'd4294967152,32'd4294967146,32'd27,32'd251,32'd4294967177,32'd24,32'd4294967268,32'd4294967262,32'd4294967156,32'd4294967155,32'd91,32'd60,32'd123,32'd4294967071,32'd9,32'd4294967281,32'd4294967197,32'd20,32'd4294967166,32'd19,32'd4294967055,32'd4294967157,32'd4,32'd50,32'd4294967004,32'd4294967195,32'd43,32'd4294967238,32'd4294967181,32'd18,32'd5,32'd4294967231,32'd32,32'd4294967208,32'd21,32'd4294967162,32'd40,32'd4294967263,32'd107,32'd4294967156,32'd4294967239,32'd71,32'd4294967204,32'd4294967246,32'd4294967199,32'd4294967138,32'd4294967163,32'd25,32'd4294967173,32'd102,32'd4294967083,32'd18,32'd134,32'd113,32'd4294967269,32'd4294967164,32'd4294967165,32'd27,32'd4294967247,32'd26,32'd4294967161,32'd4294967193,32'd4294967248,32'd4294967166,32'd1,32'd120,32'd56,32'd27,32'd4294967245,32'd37,32'd4294967263,32'd75,32'd81,32'd4294967100,32'd4294967244,32'd4294967187,32'd103,32'd72,32'd4294967177,32'd4294967192,32'd4294967136,32'd24,32'd45,32'd4294967188,32'd4294967238,32'd4294967234,32'd4294967059,32'd71,32'd11,32'd4294967246,32'd4,32'd20,32'd4294967194,32'd38,32'd4294967182,32'd46,32'd4294967243,32'd4294967237,32'd167,32'd73,32'd4294967161,32'd223,32'd4294967131,32'd4294967225,32'd4294967223,32'd33,32'd4294967167,32'd4294967153,32'd4294967182,32'd4294967259,32'd4294967011,32'd4294967244,32'd26,32'd4294967252,32'd2,32'd4294967155,32'd18,32'd10,32'd4294967100,32'd4294967261,32'd37,32'd4294967000,32'd4294967260,32'd42,32'd27,32'd4294967121,32'd31,32'd4294967141,32'd4294967266,32'd37,32'd4294967265,32'd4294967107,32'd4294967164,32'd4294967092,32'd28,32'd132,32'd4294967165,32'd7,32'd45,32'd4294967254,32'd159,32'd4294967176,32'd32,32'd4294967243,32'd4294967284,32'd52,32'd4294967138,32'd33,32'd39,32'd4294967156,32'd4294967261,32'd201,32'd141,32'd4294967252,32'd4294967265,32'd82,32'd4294967170,32'd4294967134,32'd4294967200,32'd4294967186,32'd4294967135,32'd4294967182,32'd25,32'd110,32'd89,32'd4294967253,32'd4294967221,32'd4294967251,32'd4294967227,32'd8,32'd4294967118,32'd111,32'd4294967134,32'd29,32'd97,32'd34,32'd48,32'd4294967149,32'd4294967286,32'd2,32'd4294967222,32'd4294967248,32'd185,32'd4294967168,32'd4294967291,32'd4294967120,32'd4294967161,32'd4294967128,32'd4294967130,32'd26,32'd26,32'd106,32'd4294967162,32'd4294967251,32'd4294967288,32'd4294967262,32'd95,32'd4294967090,32'd4294967271,32'd4294967074,32'd58,32'd4294967128,32'd34,32'd62,32'd36,32'd4294967220,32'd160,32'd39,32'd4294967272,32'd4294967240,32'd4294967142,32'd4294967158,32'd4294967234,32'd4294967140,32'd4294966870,32'd142,32'd54,32'd4294966999,32'd4294967249,32'd4294967199,32'd32,32'd19,32'd50,32'd9,32'd23,32'd4294967111,32'd4294967188,32'd4294966998,32'd4294967233,32'd184,32'd4294966966,32'd127,32'd4294967045,32'd23,32'd62,32'd22,32'd4294966983,32'd4294967173,32'd191,32'd4294967240,32'd4294967256,32'd4294967189,32'd4294967109,32'd4294967222,32'd4294967096,32'd148,32'd4294967062,32'd4294967289,32'd4294967176,32'd4294967072,32'd8,32'd4294967248,32'd114,32'd22,32'd4294967244,32'd4294967283,32'd4294967256,32'd226,32'd194,32'd4294967275,32'd4294967166,32'd36,32'd4294967088,32'd135,32'd4294967244,32'd4294967257,32'd47,32'd4294967231,32'd4294967117,32'd4294967212,32'd59,32'd4294967085,32'd4294967166,32'd50,32'd4294967218,32'd4294967251,32'd143,32'd187,32'd4294967242,32'd148,32'd119,32'd4294967251,32'd4294967157,32'd4294966954,32'd34,32'd4294967225,32'd4294967047,32'd4294967089,32'd159,32'd4294967186,32'd4294967107,32'd4294967080,32'd71,32'd4294967196,32'd4294967184,32'd4294967103,32'd4294967057,32'd267}
