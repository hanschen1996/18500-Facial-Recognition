`include "vj_weights.vh"

module vj_pipeline(
  input  logic clock, reset,
  input  logic [`WINDOW_SIZE-1:0][`WINDOW_SIZE-1:0][31:0] scan_win,
  input  logic [31:0] input_std_dev,
  input  logic [1:0][31:0] scan_win_index,
  output logic [1:0][31:0] top_left,
  output logic top_left_ready);

  logic [`WINDOW_SIZE-1:0][`WINDOW_SIZE-1:0][31:0] scan_win0, scan_win1,scan_win2,scan_win3,scan_win4,scan_win5,scan_win6,scan_win7,scan_win8,scan_win9,scan_win10,scan_win11,scan_win12,scan_win13,scan_win14,scan_win15,scan_win16,scan_win17,scan_win18,scan_win19,scan_win20,scan_win21,scan_win22,scan_win23,scan_win24,scan_win25,scan_win26,scan_win27,scan_win28,scan_win29,scan_win30,scan_win31,scan_win32,scan_win33,scan_win34,scan_win35,scan_win36,scan_win37,scan_win38,scan_win39,scan_win40,scan_win41,scan_win42,scan_win43,scan_win44,scan_win45,scan_win46,scan_win47,scan_win48,scan_win49,scan_win50,scan_win51,scan_win52,scan_win53,scan_win54,scan_win55,scan_win56,scan_win57,scan_win58,scan_win59,scan_win60,scan_win61,scan_win62,scan_win63,scan_win64,scan_win65,scan_win66,scan_win67,scan_win68,scan_win69,scan_win70,scan_win71,scan_win72,scan_win73,scan_win74,scan_win75,scan_win76,scan_win77,scan_win78,scan_win79,scan_win80,scan_win81,scan_win82,scan_win83,scan_win84,scan_win85,scan_win86,scan_win87,scan_win88,scan_win89,scan_win90,scan_win91,scan_win92,scan_win93,scan_win94,scan_win95,scan_win96,scan_win97,scan_win98,scan_win99,scan_win100,scan_win101,scan_win102,scan_win103,scan_win104,scan_win105,scan_win106,scan_win107,scan_win108,scan_win109,scan_win110,scan_win111,scan_win112,scan_win113,scan_win114,scan_win115,scan_win116,scan_win117,scan_win118,scan_win119,scan_win120,scan_win121,scan_win122,scan_win123,scan_win124,scan_win125,scan_win126,scan_win127,scan_win128,scan_win129,scan_win130,scan_win131,scan_win132,scan_win133,scan_win134,scan_win135,scan_win136,scan_win137,scan_win138,scan_win139,scan_win140,scan_win141,scan_win142,scan_win143,scan_win144,scan_win145,scan_win146,scan_win147,scan_win148,scan_win149,scan_win150,scan_win151,scan_win152,scan_win153,scan_win154,scan_win155,scan_win156,scan_win157,scan_win158,scan_win159,scan_win160,scan_win161,scan_win162,scan_win163,scan_win164,scan_win165,scan_win166,scan_win167,scan_win168,scan_win169,scan_win170,scan_win171,scan_win172,scan_win173,scan_win174,scan_win175,scan_win176,scan_win177,scan_win178,scan_win179,scan_win180,scan_win181,scan_win182,scan_win183,scan_win184,scan_win185,scan_win186,scan_win187,scan_win188,scan_win189,scan_win190,scan_win191,scan_win192,scan_win193,scan_win194,scan_win195,scan_win196,scan_win197,scan_win198,scan_win199,scan_win200,
  scan_win201,scan_win202,scan_win203,scan_win204,scan_win205,scan_win206,scan_win207,scan_win208,scan_win209,scan_win210,scan_win211,scan_win212,scan_win213,scan_win214,scan_win215,scan_win216,scan_win217,scan_win218,scan_win219,scan_win220,scan_win221,scan_win222,scan_win223,scan_win224,scan_win225,scan_win226,scan_win227,scan_win228,scan_win229,scan_win230,scan_win231,scan_win232,scan_win233,scan_win234,scan_win235,scan_win236,scan_win237,scan_win238,scan_win239,scan_win240,scan_win241,scan_win242,scan_win243,scan_win244,scan_win245,scan_win246,scan_win247,scan_win248,scan_win249,scan_win250,scan_win251,scan_win252,scan_win253,scan_win254,scan_win255,scan_win256,scan_win257,scan_win258,scan_win259,scan_win260,scan_win261,scan_win262,scan_win263,scan_win264,scan_win265,scan_win266,scan_win267,scan_win268,scan_win269,scan_win270,scan_win271,scan_win272,scan_win273,scan_win274,scan_win275,scan_win276,scan_win277,scan_win278,scan_win279,scan_win280,scan_win281,scan_win282,scan_win283,scan_win284,scan_win285,scan_win286,scan_win287,scan_win288,scan_win289,scan_win290,scan_win291,scan_win292,scan_win293,scan_win294,scan_win295,scan_win296,scan_win297,scan_win298,scan_win299,scan_win300,scan_win301,scan_win302,scan_win303,scan_win304,scan_win305,scan_win306,scan_win307,scan_win308,scan_win309,scan_win310,scan_win311,scan_win312,scan_win313,scan_win314,scan_win315,scan_win316,scan_win317,scan_win318,scan_win319,scan_win320,scan_win321,scan_win322,scan_win323,scan_win324,scan_win325,scan_win326,scan_win327,scan_win328,scan_win329,scan_win330,scan_win331,scan_win332,scan_win333,scan_win334,scan_win335,scan_win336,scan_win337,scan_win338,scan_win339,scan_win340,scan_win341,scan_win342,scan_win343,scan_win344,scan_win345,scan_win346,scan_win347,scan_win348,scan_win349,scan_win350,scan_win351,scan_win352,scan_win353,scan_win354,scan_win355,scan_win356,scan_win357,scan_win358,scan_win359,scan_win360,scan_win361,scan_win362,scan_win363,scan_win364,scan_win365,scan_win366,scan_win367,scan_win368,scan_win369,scan_win370,scan_win371,scan_win372,scan_win373,scan_win374,scan_win375,scan_win376,scan_win377,scan_win378,scan_win379,scan_win380,scan_win381,scan_win382,scan_win383,scan_win384,scan_win385,scan_win386,scan_win387,scan_win388,scan_win389,scan_win390,scan_win391,scan_win392,scan_win393,scan_win394,scan_win395,scan_win396,scan_win397,scan_win398,scan_win399,scan_win400,
  scan_win401,scan_win402,scan_win403,scan_win404,scan_win405,scan_win406,scan_win407,scan_win408,scan_win409,scan_win410,scan_win411,scan_win412,scan_win413,scan_win414,scan_win415,scan_win416,scan_win417,scan_win418,scan_win419,scan_win420,scan_win421,scan_win422,scan_win423,scan_win424,scan_win425,scan_win426,scan_win427,scan_win428,scan_win429,scan_win430,scan_win431,scan_win432,scan_win433,scan_win434,scan_win435,scan_win436,scan_win437,scan_win438,scan_win439,scan_win440,scan_win441,scan_win442,scan_win443,scan_win444,scan_win445,scan_win446,scan_win447,scan_win448,scan_win449,scan_win450,scan_win451,scan_win452,scan_win453,scan_win454,scan_win455,scan_win456,scan_win457,scan_win458,scan_win459,scan_win460,scan_win461,scan_win462,scan_win463,scan_win464,scan_win465,scan_win466,scan_win467,scan_win468,scan_win469,scan_win470,scan_win471,scan_win472,scan_win473,scan_win474,scan_win475,scan_win476,scan_win477,scan_win478,scan_win479,scan_win480,scan_win481,scan_win482,scan_win483,scan_win484,scan_win485,scan_win486,scan_win487,scan_win488,scan_win489,scan_win490,scan_win491,scan_win492,scan_win493,scan_win494,scan_win495,scan_win496,scan_win497,scan_win498,scan_win499,scan_win500,scan_win501,scan_win502,scan_win503,scan_win504,scan_win505,scan_win506,scan_win507,scan_win508,scan_win509,scan_win510,scan_win511,scan_win512,scan_win513,scan_win514,scan_win515,scan_win516,scan_win517,scan_win518,scan_win519,scan_win520,scan_win521,scan_win522,scan_win523,scan_win524,scan_win525,scan_win526,scan_win527,scan_win528,scan_win529,scan_win530,scan_win531,scan_win532,scan_win533,scan_win534,scan_win535,scan_win536,scan_win537,scan_win538,scan_win539,scan_win540,scan_win541,scan_win542,scan_win543,scan_win544,scan_win545,scan_win546,scan_win547,scan_win548,scan_win549,scan_win550,scan_win551,scan_win552,scan_win553,scan_win554,scan_win555,scan_win556,scan_win557,scan_win558,scan_win559,scan_win560,scan_win561,scan_win562,scan_win563,scan_win564,scan_win565,scan_win566,scan_win567,scan_win568,scan_win569,scan_win570,scan_win571,scan_win572,scan_win573,scan_win574,scan_win575,scan_win576,scan_win577,scan_win578,scan_win579,scan_win580,scan_win581,scan_win582,scan_win583,scan_win584,scan_win585,scan_win586,scan_win587,scan_win588,scan_win589,scan_win590,scan_win591,scan_win592,scan_win593,scan_win594,scan_win595,scan_win596,scan_win597,scan_win598,scan_win599,scan_win600,
  scan_win601,scan_win602,scan_win603,scan_win604,scan_win605,scan_win606,scan_win607,scan_win608,scan_win609,scan_win610,scan_win611,scan_win612,scan_win613,scan_win614,scan_win615,scan_win616,scan_win617,scan_win618,scan_win619,scan_win620,scan_win621,scan_win622,scan_win623,scan_win624,scan_win625,scan_win626,scan_win627,scan_win628,scan_win629,scan_win630,scan_win631,scan_win632,scan_win633,scan_win634,scan_win635,scan_win636,scan_win637,scan_win638,scan_win639,scan_win640,scan_win641,scan_win642,scan_win643,scan_win644,scan_win645,scan_win646,scan_win647,scan_win648,scan_win649,scan_win650,scan_win651,scan_win652,scan_win653,scan_win654,scan_win655,scan_win656,scan_win657,scan_win658,scan_win659,scan_win660,scan_win661,scan_win662,scan_win663,scan_win664,scan_win665,scan_win666,scan_win667,scan_win668,scan_win669,scan_win670,scan_win671,scan_win672,scan_win673,scan_win674,scan_win675,scan_win676,scan_win677,scan_win678,scan_win679,scan_win680,scan_win681,scan_win682,scan_win683,scan_win684,scan_win685,scan_win686,scan_win687,scan_win688,scan_win689,scan_win690,scan_win691,scan_win692,scan_win693,scan_win694,scan_win695,scan_win696,scan_win697,scan_win698,scan_win699,scan_win700,scan_win701,scan_win702,scan_win703,scan_win704,scan_win705,scan_win706,scan_win707,scan_win708,scan_win709,scan_win710,scan_win711,scan_win712,scan_win713,scan_win714,scan_win715,scan_win716,scan_win717,scan_win718,scan_win719,scan_win720,scan_win721,scan_win722,scan_win723,scan_win724,scan_win725,scan_win726,scan_win727,scan_win728,scan_win729,scan_win730,scan_win731,scan_win732,scan_win733,scan_win734,scan_win735,scan_win736,scan_win737,scan_win738,scan_win739,scan_win740,scan_win741,scan_win742,scan_win743,scan_win744,scan_win745,scan_win746,scan_win747,scan_win748,scan_win749,scan_win750,scan_win751,scan_win752,scan_win753,scan_win754,scan_win755,scan_win756,scan_win757,scan_win758,scan_win759,scan_win760,scan_win761,scan_win762,scan_win763,scan_win764,scan_win765,scan_win766,scan_win767,scan_win768,scan_win769,scan_win770,scan_win771,scan_win772,scan_win773,scan_win774,scan_win775,scan_win776,scan_win777,scan_win778,scan_win779,scan_win780,scan_win781,scan_win782,scan_win783,scan_win784,scan_win785,scan_win786,scan_win787,scan_win788,scan_win789,scan_win790,scan_win791,scan_win792,scan_win793,scan_win794,scan_win795,scan_win796,scan_win797,scan_win798,scan_win799,scan_win800,
  scan_win801,scan_win802,scan_win803,scan_win804,scan_win805,scan_win806,scan_win807,scan_win808,scan_win809,scan_win810,scan_win811,scan_win812,scan_win813,scan_win814,scan_win815,scan_win816,scan_win817,scan_win818,scan_win819,scan_win820,scan_win821,scan_win822,scan_win823,scan_win824,scan_win825,scan_win826,scan_win827,scan_win828,scan_win829,scan_win830,scan_win831,scan_win832,scan_win833,scan_win834,scan_win835,scan_win836,scan_win837,scan_win838,scan_win839,scan_win840,scan_win841,scan_win842,scan_win843,scan_win844,scan_win845,scan_win846,scan_win847,scan_win848,scan_win849,scan_win850,scan_win851,scan_win852,scan_win853,scan_win854,scan_win855,scan_win856,scan_win857,scan_win858,scan_win859,scan_win860,scan_win861,scan_win862,scan_win863,scan_win864,scan_win865,scan_win866,scan_win867,scan_win868,scan_win869,scan_win870,scan_win871,scan_win872,scan_win873,scan_win874,scan_win875,scan_win876,scan_win877,scan_win878,scan_win879,scan_win880,scan_win881,scan_win882,scan_win883,scan_win884,scan_win885,scan_win886,scan_win887,scan_win888,scan_win889,scan_win890,scan_win891,scan_win892,scan_win893,scan_win894,scan_win895,scan_win896,scan_win897,scan_win898,scan_win899,scan_win900,scan_win901,scan_win902,scan_win903,scan_win904,scan_win905,scan_win906,scan_win907,scan_win908,scan_win909,scan_win910,scan_win911,scan_win912,scan_win913,scan_win914,scan_win915,scan_win916,scan_win917,scan_win918,scan_win919,scan_win920,scan_win921,scan_win922,scan_win923,scan_win924,scan_win925,scan_win926,scan_win927,scan_win928,scan_win929,scan_win930,scan_win931,scan_win932,scan_win933,scan_win934,scan_win935,scan_win936,scan_win937,scan_win938,scan_win939,scan_win940,scan_win941,scan_win942,scan_win943,scan_win944,scan_win945,scan_win946,scan_win947,scan_win948,scan_win949,scan_win950,scan_win951,scan_win952,scan_win953,scan_win954,scan_win955,scan_win956,scan_win957,scan_win958,scan_win959,scan_win960,scan_win961,scan_win962,scan_win963,scan_win964,scan_win965,scan_win966,scan_win967,scan_win968,scan_win969,scan_win970,scan_win971,scan_win972,scan_win973,scan_win974,scan_win975,scan_win976,scan_win977,scan_win978,scan_win979,scan_win980,scan_win981,scan_win982,scan_win983,scan_win984,scan_win985,scan_win986,scan_win987,scan_win988,scan_win989,scan_win990,scan_win991,scan_win992,scan_win993,scan_win994,scan_win995,scan_win996,scan_win997,scan_win998,scan_win999,scan_win1000,
  scan_win1001,scan_win1002,scan_win1003,scan_win1004,scan_win1005,scan_win1006,scan_win1007,scan_win1008,scan_win1009,scan_win1010,scan_win1011,scan_win1012,scan_win1013,scan_win1014,scan_win1015,scan_win1016,scan_win1017,scan_win1018,scan_win1019,scan_win1020,scan_win1021,scan_win1022,scan_win1023,scan_win1024,scan_win1025,scan_win1026,scan_win1027,scan_win1028,scan_win1029,scan_win1030,scan_win1031,scan_win1032,scan_win1033,scan_win1034,scan_win1035,scan_win1036,scan_win1037,scan_win1038,scan_win1039,scan_win1040,scan_win1041,scan_win1042,scan_win1043,scan_win1044,scan_win1045,scan_win1046,scan_win1047,scan_win1048,scan_win1049,scan_win1050,scan_win1051,scan_win1052,scan_win1053,scan_win1054,scan_win1055,scan_win1056,scan_win1057,scan_win1058,scan_win1059,scan_win1060,scan_win1061,scan_win1062,scan_win1063,scan_win1064,scan_win1065,scan_win1066,scan_win1067,scan_win1068,scan_win1069,scan_win1070,scan_win1071,scan_win1072,scan_win1073,scan_win1074,scan_win1075,scan_win1076,scan_win1077,scan_win1078,scan_win1079,scan_win1080,scan_win1081,scan_win1082,scan_win1083,scan_win1084,scan_win1085,scan_win1086,scan_win1087,scan_win1088,scan_win1089,scan_win1090,scan_win1091,scan_win1092,scan_win1093,scan_win1094,scan_win1095,scan_win1096,scan_win1097,scan_win1098,scan_win1099,scan_win1100,scan_win1101,scan_win1102,scan_win1103,scan_win1104,scan_win1105,scan_win1106,scan_win1107,scan_win1108,scan_win1109,scan_win1110,scan_win1111,scan_win1112,scan_win1113,scan_win1114,scan_win1115,scan_win1116,scan_win1117,scan_win1118,scan_win1119,scan_win1120,scan_win1121,scan_win1122,scan_win1123,scan_win1124,scan_win1125,scan_win1126,scan_win1127,scan_win1128,scan_win1129,scan_win1130,scan_win1131,scan_win1132,scan_win1133,scan_win1134,scan_win1135,scan_win1136,scan_win1137,scan_win1138,scan_win1139,scan_win1140,scan_win1141,scan_win1142,scan_win1143,scan_win1144,scan_win1145,scan_win1146,scan_win1147,scan_win1148,scan_win1149,scan_win1150,scan_win1151,scan_win1152,scan_win1153,scan_win1154,scan_win1155,scan_win1156,scan_win1157,scan_win1158,scan_win1159,scan_win1160,scan_win1161,scan_win1162,scan_win1163,scan_win1164,scan_win1165,scan_win1166,scan_win1167,scan_win1168,scan_win1169,scan_win1170,scan_win1171,scan_win1172,scan_win1173,scan_win1174,scan_win1175,scan_win1176,scan_win1177,scan_win1178,scan_win1179,scan_win1180,scan_win1181,scan_win1182,scan_win1183,scan_win1184,scan_win1185,scan_win1186,scan_win1187,scan_win1188,scan_win1189,scan_win1190,scan_win1191,scan_win1192,scan_win1193,scan_win1194,scan_win1195,scan_win1196,scan_win1197,scan_win1198,scan_win1199,scan_win1200,
  scan_win1201,scan_win1202,scan_win1203,scan_win1204,scan_win1205,scan_win1206,scan_win1207,scan_win1208,scan_win1209,scan_win1210,scan_win1211,scan_win1212,scan_win1213,scan_win1214,scan_win1215,scan_win1216,scan_win1217,scan_win1218,scan_win1219,scan_win1220,scan_win1221,scan_win1222,scan_win1223,scan_win1224,scan_win1225,scan_win1226,scan_win1227,scan_win1228,scan_win1229,scan_win1230,scan_win1231,scan_win1232,scan_win1233,scan_win1234,scan_win1235,scan_win1236,scan_win1237,scan_win1238,scan_win1239,scan_win1240,scan_win1241,scan_win1242,scan_win1243,scan_win1244,scan_win1245,scan_win1246,scan_win1247,scan_win1248,scan_win1249,scan_win1250,scan_win1251,scan_win1252,scan_win1253,scan_win1254,scan_win1255,scan_win1256,scan_win1257,scan_win1258,scan_win1259,scan_win1260,scan_win1261,scan_win1262,scan_win1263,scan_win1264,scan_win1265,scan_win1266,scan_win1267,scan_win1268,scan_win1269,scan_win1270,scan_win1271,scan_win1272,scan_win1273,scan_win1274,scan_win1275,scan_win1276,scan_win1277,scan_win1278,scan_win1279,scan_win1280,scan_win1281,scan_win1282,scan_win1283,scan_win1284,scan_win1285,scan_win1286,scan_win1287,scan_win1288,scan_win1289,scan_win1290,scan_win1291,scan_win1292,scan_win1293,scan_win1294,scan_win1295,scan_win1296,scan_win1297,scan_win1298,scan_win1299,scan_win1300,scan_win1301,scan_win1302,scan_win1303,scan_win1304,scan_win1305,scan_win1306,scan_win1307,scan_win1308,scan_win1309,scan_win1310,scan_win1311,scan_win1312,scan_win1313,scan_win1314,scan_win1315,scan_win1316,scan_win1317,scan_win1318,scan_win1319,scan_win1320,scan_win1321,scan_win1322,scan_win1323,scan_win1324,scan_win1325,scan_win1326,scan_win1327,scan_win1328,scan_win1329,scan_win1330,scan_win1331,scan_win1332,scan_win1333,scan_win1334,scan_win1335,scan_win1336,scan_win1337,scan_win1338,scan_win1339,scan_win1340,scan_win1341,scan_win1342,scan_win1343,scan_win1344,scan_win1345,scan_win1346,scan_win1347,scan_win1348,scan_win1349,scan_win1350,scan_win1351,scan_win1352,scan_win1353,scan_win1354,scan_win1355,scan_win1356,scan_win1357,scan_win1358,scan_win1359,scan_win1360,scan_win1361,scan_win1362,scan_win1363,scan_win1364,scan_win1365,scan_win1366,scan_win1367,scan_win1368,scan_win1369,scan_win1370,scan_win1371,scan_win1372,scan_win1373,scan_win1374,scan_win1375,scan_win1376,scan_win1377,scan_win1378,scan_win1379,scan_win1380,scan_win1381,scan_win1382,scan_win1383,scan_win1384,scan_win1385,scan_win1386,scan_win1387,scan_win1388,scan_win1389,scan_win1390,scan_win1391,scan_win1392,scan_win1393,scan_win1394,scan_win1395,scan_win1396,scan_win1397,scan_win1398,scan_win1399,scan_win1400,
  scan_win1401,scan_win1402,scan_win1403,scan_win1404,scan_win1405,scan_win1406,scan_win1407,scan_win1408,scan_win1409,scan_win1410,scan_win1411,scan_win1412,scan_win1413,scan_win1414,scan_win1415,scan_win1416,scan_win1417,scan_win1418,scan_win1419,scan_win1420,scan_win1421,scan_win1422,scan_win1423,scan_win1424,scan_win1425,scan_win1426,scan_win1427,scan_win1428,scan_win1429,scan_win1430,scan_win1431,scan_win1432,scan_win1433,scan_win1434,scan_win1435,scan_win1436,scan_win1437,scan_win1438,scan_win1439,scan_win1440,scan_win1441,scan_win1442,scan_win1443,scan_win1444,scan_win1445,scan_win1446,scan_win1447,scan_win1448,scan_win1449,scan_win1450,scan_win1451,scan_win1452,scan_win1453,scan_win1454,scan_win1455,scan_win1456,scan_win1457,scan_win1458,scan_win1459,scan_win1460,scan_win1461,scan_win1462,scan_win1463,scan_win1464,scan_win1465,scan_win1466,scan_win1467,scan_win1468,scan_win1469,scan_win1470,scan_win1471,scan_win1472,scan_win1473,scan_win1474,scan_win1475,scan_win1476,scan_win1477,scan_win1478,scan_win1479,scan_win1480,scan_win1481,scan_win1482,scan_win1483,scan_win1484,scan_win1485,scan_win1486,scan_win1487,scan_win1488,scan_win1489,scan_win1490,scan_win1491,scan_win1492,scan_win1493,scan_win1494,scan_win1495,scan_win1496,scan_win1497,scan_win1498,scan_win1499,scan_win1500,scan_win1501,scan_win1502,scan_win1503,scan_win1504,scan_win1505,scan_win1506,scan_win1507,scan_win1508,scan_win1509,scan_win1510,scan_win1511,scan_win1512,scan_win1513,scan_win1514,scan_win1515,scan_win1516,scan_win1517,scan_win1518,scan_win1519,scan_win1520,scan_win1521,scan_win1522,scan_win1523,scan_win1524,scan_win1525,scan_win1526,scan_win1527,scan_win1528,scan_win1529,scan_win1530,scan_win1531,scan_win1532,scan_win1533,scan_win1534,scan_win1535,scan_win1536,scan_win1537,scan_win1538,scan_win1539,scan_win1540,scan_win1541,scan_win1542,scan_win1543,scan_win1544,scan_win1545,scan_win1546,scan_win1547,scan_win1548,scan_win1549,scan_win1550,scan_win1551,scan_win1552,scan_win1553,scan_win1554,scan_win1555,scan_win1556,scan_win1557,scan_win1558,scan_win1559,scan_win1560,scan_win1561,scan_win1562,scan_win1563,scan_win1564,scan_win1565,scan_win1566,scan_win1567,scan_win1568,scan_win1569,scan_win1570,scan_win1571,scan_win1572,scan_win1573,scan_win1574,scan_win1575,scan_win1576,scan_win1577,scan_win1578,scan_win1579,scan_win1580,scan_win1581,scan_win1582,scan_win1583,scan_win1584,scan_win1585,scan_win1586,scan_win1587,scan_win1588,scan_win1589,scan_win1590,scan_win1591,scan_win1592,scan_win1593,scan_win1594,scan_win1595,scan_win1596,scan_win1597,scan_win1598,scan_win1599,scan_win1600,
  scan_win1601,scan_win1602,scan_win1603,scan_win1604,scan_win1605,scan_win1606,scan_win1607,scan_win1608,scan_win1609,scan_win1610,scan_win1611,scan_win1612,scan_win1613,scan_win1614,scan_win1615,scan_win1616,scan_win1617,scan_win1618,scan_win1619,scan_win1620,scan_win1621,scan_win1622,scan_win1623,scan_win1624,scan_win1625,scan_win1626,scan_win1627,scan_win1628,scan_win1629,scan_win1630,scan_win1631,scan_win1632,scan_win1633,scan_win1634,scan_win1635,scan_win1636,scan_win1637,scan_win1638,scan_win1639,scan_win1640,scan_win1641,scan_win1642,scan_win1643,scan_win1644,scan_win1645,scan_win1646,scan_win1647,scan_win1648,scan_win1649,scan_win1650,scan_win1651,scan_win1652,scan_win1653,scan_win1654,scan_win1655,scan_win1656,scan_win1657,scan_win1658,scan_win1659,scan_win1660,scan_win1661,scan_win1662,scan_win1663,scan_win1664,scan_win1665,scan_win1666,scan_win1667,scan_win1668,scan_win1669,scan_win1670,scan_win1671,scan_win1672,scan_win1673,scan_win1674,scan_win1675,scan_win1676,scan_win1677,scan_win1678,scan_win1679,scan_win1680,scan_win1681,scan_win1682,scan_win1683,scan_win1684,scan_win1685,scan_win1686,scan_win1687,scan_win1688,scan_win1689,scan_win1690,scan_win1691,scan_win1692,scan_win1693,scan_win1694,scan_win1695,scan_win1696,scan_win1697,scan_win1698,scan_win1699,scan_win1700,scan_win1701,scan_win1702,scan_win1703,scan_win1704,scan_win1705,scan_win1706,scan_win1707,scan_win1708,scan_win1709,scan_win1710,scan_win1711,scan_win1712,scan_win1713,scan_win1714,scan_win1715,scan_win1716,scan_win1717,scan_win1718,scan_win1719,scan_win1720,scan_win1721,scan_win1722,scan_win1723,scan_win1724,scan_win1725,scan_win1726,scan_win1727,scan_win1728,scan_win1729,scan_win1730,scan_win1731,scan_win1732,scan_win1733,scan_win1734,scan_win1735,scan_win1736,scan_win1737,scan_win1738,scan_win1739,scan_win1740,scan_win1741,scan_win1742,scan_win1743,scan_win1744,scan_win1745,scan_win1746,scan_win1747,scan_win1748,scan_win1749,scan_win1750,scan_win1751,scan_win1752,scan_win1753,scan_win1754,scan_win1755,scan_win1756,scan_win1757,scan_win1758,scan_win1759,scan_win1760,scan_win1761,scan_win1762,scan_win1763,scan_win1764,scan_win1765,scan_win1766,scan_win1767,scan_win1768,scan_win1769,scan_win1770,scan_win1771,scan_win1772,scan_win1773,scan_win1774,scan_win1775,scan_win1776,scan_win1777,scan_win1778,scan_win1779,scan_win1780,scan_win1781,scan_win1782,scan_win1783,scan_win1784,scan_win1785,scan_win1786,scan_win1787,scan_win1788,scan_win1789,scan_win1790,scan_win1791,scan_win1792,scan_win1793,scan_win1794,scan_win1795,scan_win1796,scan_win1797,scan_win1798,scan_win1799,scan_win1800,
  scan_win1801,scan_win1802,scan_win1803,scan_win1804,scan_win1805,scan_win1806,scan_win1807,scan_win1808,scan_win1809,scan_win1810,scan_win1811,scan_win1812,scan_win1813,scan_win1814,scan_win1815,scan_win1816,scan_win1817,scan_win1818,scan_win1819,scan_win1820,scan_win1821,scan_win1822,scan_win1823,scan_win1824,scan_win1825,scan_win1826,scan_win1827,scan_win1828,scan_win1829,scan_win1830,scan_win1831,scan_win1832,scan_win1833,scan_win1834,scan_win1835,scan_win1836,scan_win1837,scan_win1838,scan_win1839,scan_win1840,scan_win1841,scan_win1842,scan_win1843,scan_win1844,scan_win1845,scan_win1846,scan_win1847,scan_win1848,scan_win1849,scan_win1850,scan_win1851,scan_win1852,scan_win1853,scan_win1854,scan_win1855,scan_win1856,scan_win1857,scan_win1858,scan_win1859,scan_win1860,scan_win1861,scan_win1862,scan_win1863,scan_win1864,scan_win1865,scan_win1866,scan_win1867,scan_win1868,scan_win1869,scan_win1870,scan_win1871,scan_win1872,scan_win1873,scan_win1874,scan_win1875,scan_win1876,scan_win1877,scan_win1878,scan_win1879,scan_win1880,scan_win1881,scan_win1882,scan_win1883,scan_win1884,scan_win1885,scan_win1886,scan_win1887,scan_win1888,scan_win1889,scan_win1890,scan_win1891,scan_win1892,scan_win1893,scan_win1894,scan_win1895,scan_win1896,scan_win1897,scan_win1898,scan_win1899,scan_win1900,scan_win1901,scan_win1902,scan_win1903,scan_win1904,scan_win1905,scan_win1906,scan_win1907,scan_win1908,scan_win1909,scan_win1910,scan_win1911,scan_win1912,scan_win1913,scan_win1914,scan_win1915,scan_win1916,scan_win1917,scan_win1918,scan_win1919,scan_win1920,scan_win1921,scan_win1922,scan_win1923,scan_win1924,scan_win1925,scan_win1926,scan_win1927,scan_win1928,scan_win1929,scan_win1930,scan_win1931,scan_win1932,scan_win1933,scan_win1934,scan_win1935,scan_win1936,scan_win1937,scan_win1938,scan_win1939,scan_win1940,scan_win1941,scan_win1942,scan_win1943,scan_win1944,scan_win1945,scan_win1946,scan_win1947,scan_win1948,scan_win1949,scan_win1950,scan_win1951,scan_win1952,scan_win1953,scan_win1954,scan_win1955,scan_win1956,scan_win1957,scan_win1958,scan_win1959,scan_win1960,scan_win1961,scan_win1962,scan_win1963,scan_win1964,scan_win1965,scan_win1966,scan_win1967,scan_win1968,scan_win1969,scan_win1970,scan_win1971,scan_win1972,scan_win1973,scan_win1974,scan_win1975,scan_win1976,scan_win1977,scan_win1978,scan_win1979,scan_win1980,scan_win1981,scan_win1982,scan_win1983,scan_win1984,scan_win1985,scan_win1986,scan_win1987,scan_win1988,scan_win1989,scan_win1990,scan_win1991,scan_win1992,scan_win1993,scan_win1994,scan_win1995,scan_win1996,scan_win1997,scan_win1998,scan_win1999,scan_win2000,
  scan_win2001,scan_win2002,scan_win2003,scan_win2004,scan_win2005,scan_win2006,scan_win2007,scan_win2008,scan_win2009,scan_win2010,scan_win2011,scan_win2012,scan_win2013,scan_win2014,scan_win2015,scan_win2016,scan_win2017,scan_win2018,scan_win2019,scan_win2020,scan_win2021,scan_win2022,scan_win2023,scan_win2024,scan_win2025,scan_win2026,scan_win2027,scan_win2028,scan_win2029,scan_win2030,scan_win2031,scan_win2032,scan_win2033,scan_win2034,scan_win2035,scan_win2036,scan_win2037,scan_win2038,scan_win2039,scan_win2040,scan_win2041,scan_win2042,scan_win2043,scan_win2044,scan_win2045,scan_win2046,scan_win2047,scan_win2048,scan_win2049,scan_win2050,scan_win2051,scan_win2052,scan_win2053,scan_win2054,scan_win2055,scan_win2056,scan_win2057,scan_win2058,scan_win2059,scan_win2060,scan_win2061,scan_win2062,scan_win2063,scan_win2064,scan_win2065,scan_win2066,scan_win2067,scan_win2068,scan_win2069,scan_win2070,scan_win2071,scan_win2072,scan_win2073,scan_win2074,scan_win2075,scan_win2076,scan_win2077,scan_win2078,scan_win2079,scan_win2080,scan_win2081,scan_win2082,scan_win2083,scan_win2084,scan_win2085,scan_win2086,scan_win2087,scan_win2088,scan_win2089,scan_win2090,scan_win2091,scan_win2092,scan_win2093,scan_win2094,scan_win2095,scan_win2096,scan_win2097,scan_win2098,scan_win2099,scan_win2100,scan_win2101,scan_win2102,scan_win2103,scan_win2104,scan_win2105,scan_win2106,scan_win2107,scan_win2108,scan_win2109,scan_win2110,scan_win2111,scan_win2112,scan_win2113,scan_win2114,scan_win2115,scan_win2116,scan_win2117,scan_win2118,scan_win2119,scan_win2120,scan_win2121,scan_win2122,scan_win2123,scan_win2124,scan_win2125,scan_win2126,scan_win2127,scan_win2128,scan_win2129,scan_win2130,scan_win2131,scan_win2132,scan_win2133,scan_win2134,scan_win2135,scan_win2136,scan_win2137,scan_win2138,scan_win2139,scan_win2140,scan_win2141,scan_win2142,scan_win2143,scan_win2144,scan_win2145,scan_win2146,scan_win2147,scan_win2148,scan_win2149,scan_win2150,scan_win2151,scan_win2152,scan_win2153,scan_win2154,scan_win2155,scan_win2156,scan_win2157,scan_win2158,scan_win2159,scan_win2160,scan_win2161,scan_win2162,scan_win2163,scan_win2164,scan_win2165,scan_win2166,scan_win2167,scan_win2168,scan_win2169,scan_win2170,scan_win2171,scan_win2172,scan_win2173,scan_win2174,scan_win2175,scan_win2176,scan_win2177,scan_win2178,scan_win2179,scan_win2180,scan_win2181,scan_win2182,scan_win2183,scan_win2184,scan_win2185,scan_win2186,scan_win2187,scan_win2188,scan_win2189,scan_win2190,scan_win2191,scan_win2192,scan_win2193,scan_win2194,scan_win2195,scan_win2196,scan_win2197,scan_win2198,scan_win2199,scan_win2200,
  scan_win2201,scan_win2202,scan_win2203,scan_win2204,scan_win2205,scan_win2206,scan_win2207,scan_win2208,scan_win2209,scan_win2210,scan_win2211,scan_win2212,scan_win2213,scan_win2214,scan_win2215,scan_win2216,scan_win2217,scan_win2218,scan_win2219,scan_win2220,scan_win2221,scan_win2222,scan_win2223,scan_win2224,scan_win2225,scan_win2226,scan_win2227,scan_win2228,scan_win2229,scan_win2230,scan_win2231,scan_win2232,scan_win2233,scan_win2234,scan_win2235,scan_win2236,scan_win2237,scan_win2238,scan_win2239,scan_win2240,scan_win2241,scan_win2242,scan_win2243,scan_win2244,scan_win2245,scan_win2246,scan_win2247,scan_win2248,scan_win2249,scan_win2250,scan_win2251,scan_win2252,scan_win2253,scan_win2254,scan_win2255,scan_win2256,scan_win2257,scan_win2258,scan_win2259,scan_win2260,scan_win2261,scan_win2262,scan_win2263,scan_win2264,scan_win2265,scan_win2266,scan_win2267,scan_win2268,scan_win2269,scan_win2270,scan_win2271,scan_win2272,scan_win2273,scan_win2274,scan_win2275,scan_win2276,scan_win2277,scan_win2278,scan_win2279,scan_win2280,scan_win2281,scan_win2282,scan_win2283,scan_win2284,scan_win2285,scan_win2286,scan_win2287,scan_win2288,scan_win2289,scan_win2290,scan_win2291,scan_win2292,scan_win2293,scan_win2294,scan_win2295,scan_win2296,scan_win2297,scan_win2298,scan_win2299,scan_win2300,scan_win2301,scan_win2302,scan_win2303,scan_win2304,scan_win2305,scan_win2306,scan_win2307,scan_win2308,scan_win2309,scan_win2310,scan_win2311,scan_win2312,scan_win2313,scan_win2314,scan_win2315,scan_win2316,scan_win2317,scan_win2318,scan_win2319,scan_win2320,scan_win2321,scan_win2322,scan_win2323,scan_win2324,scan_win2325,scan_win2326,scan_win2327,scan_win2328,scan_win2329,scan_win2330,scan_win2331,scan_win2332,scan_win2333,scan_win2334,scan_win2335,scan_win2336,scan_win2337,scan_win2338,scan_win2339,scan_win2340,scan_win2341,scan_win2342,scan_win2343,scan_win2344,scan_win2345,scan_win2346,scan_win2347,scan_win2348,scan_win2349,scan_win2350,scan_win2351,scan_win2352,scan_win2353,scan_win2354,scan_win2355,scan_win2356,scan_win2357,scan_win2358,scan_win2359,scan_win2360,scan_win2361,scan_win2362,scan_win2363,scan_win2364,scan_win2365,scan_win2366,scan_win2367,scan_win2368,scan_win2369,scan_win2370,scan_win2371,scan_win2372,scan_win2373,scan_win2374,scan_win2375,scan_win2376,scan_win2377,scan_win2378,scan_win2379,scan_win2380,scan_win2381,scan_win2382,scan_win2383,scan_win2384,scan_win2385,scan_win2386,scan_win2387,scan_win2388,scan_win2389,scan_win2390,scan_win2391,scan_win2392,scan_win2393,scan_win2394,scan_win2395,scan_win2396,scan_win2397,scan_win2398,scan_win2399,scan_win2400,
  scan_win2401,scan_win2402,scan_win2403,scan_win2404,scan_win2405,scan_win2406,scan_win2407,scan_win2408,scan_win2409,scan_win2410,scan_win2411,scan_win2412,scan_win2413,scan_win2414,scan_win2415,scan_win2416,scan_win2417,scan_win2418,scan_win2419,scan_win2420,scan_win2421,scan_win2422,scan_win2423,scan_win2424,scan_win2425,scan_win2426,scan_win2427,scan_win2428,scan_win2429,scan_win2430,scan_win2431,scan_win2432,scan_win2433,scan_win2434,scan_win2435,scan_win2436,scan_win2437,scan_win2438,scan_win2439,scan_win2440,scan_win2441,scan_win2442,scan_win2443,scan_win2444,scan_win2445,scan_win2446,scan_win2447,scan_win2448,scan_win2449,scan_win2450,scan_win2451,scan_win2452,scan_win2453,scan_win2454,scan_win2455,scan_win2456,scan_win2457,scan_win2458,scan_win2459,scan_win2460,scan_win2461,scan_win2462,scan_win2463,scan_win2464,scan_win2465,scan_win2466,scan_win2467,scan_win2468,scan_win2469,scan_win2470,scan_win2471,scan_win2472,scan_win2473,scan_win2474,scan_win2475,scan_win2476,scan_win2477,scan_win2478,scan_win2479,scan_win2480,scan_win2481,scan_win2482,scan_win2483,scan_win2484,scan_win2485,scan_win2486,scan_win2487,scan_win2488,scan_win2489,scan_win2490,scan_win2491,scan_win2492,scan_win2493,scan_win2494,scan_win2495,scan_win2496,scan_win2497,scan_win2498,scan_win2499,scan_win2500,scan_win2501,scan_win2502,scan_win2503,scan_win2504,scan_win2505,scan_win2506,scan_win2507,scan_win2508,scan_win2509,scan_win2510,scan_win2511,scan_win2512,scan_win2513,scan_win2514,scan_win2515,scan_win2516,scan_win2517,scan_win2518,scan_win2519,scan_win2520,scan_win2521,scan_win2522,scan_win2523,scan_win2524,scan_win2525,scan_win2526,scan_win2527,scan_win2528,scan_win2529,scan_win2530,scan_win2531,scan_win2532,scan_win2533,scan_win2534,scan_win2535,scan_win2536,scan_win2537,scan_win2538,scan_win2539,scan_win2540,scan_win2541,scan_win2542,scan_win2543,scan_win2544,scan_win2545,scan_win2546,scan_win2547,scan_win2548,scan_win2549,scan_win2550,scan_win2551,scan_win2552,scan_win2553,scan_win2554,scan_win2555,scan_win2556,scan_win2557,scan_win2558,scan_win2559,scan_win2560,scan_win2561,scan_win2562,scan_win2563,scan_win2564,scan_win2565,scan_win2566,scan_win2567,scan_win2568,scan_win2569,scan_win2570,scan_win2571,scan_win2572,scan_win2573,scan_win2574,scan_win2575,scan_win2576,scan_win2577,scan_win2578,scan_win2579,scan_win2580,scan_win2581,scan_win2582,scan_win2583,scan_win2584,scan_win2585,scan_win2586,scan_win2587,scan_win2588,scan_win2589,scan_win2590,scan_win2591,scan_win2592,scan_win2593,scan_win2594,scan_win2595,scan_win2596,scan_win2597,scan_win2598,scan_win2599,scan_win2600,
  scan_win2601,scan_win2602,scan_win2603,scan_win2604,scan_win2605,scan_win2606,scan_win2607,scan_win2608,scan_win2609,scan_win2610,scan_win2611,scan_win2612,scan_win2613,scan_win2614,scan_win2615,scan_win2616,scan_win2617,scan_win2618,scan_win2619,scan_win2620,scan_win2621,scan_win2622,scan_win2623,scan_win2624,scan_win2625,scan_win2626,scan_win2627,scan_win2628,scan_win2629,scan_win2630,scan_win2631,scan_win2632,scan_win2633,scan_win2634,scan_win2635,scan_win2636,scan_win2637,scan_win2638,scan_win2639,scan_win2640,scan_win2641,scan_win2642,scan_win2643,scan_win2644,scan_win2645,scan_win2646,scan_win2647,scan_win2648,scan_win2649,scan_win2650,scan_win2651,scan_win2652,scan_win2653,scan_win2654,scan_win2655,scan_win2656,scan_win2657,scan_win2658,scan_win2659,scan_win2660,scan_win2661,scan_win2662,scan_win2663,scan_win2664,scan_win2665,scan_win2666,scan_win2667,scan_win2668,scan_win2669,scan_win2670,scan_win2671,scan_win2672,scan_win2673,scan_win2674,scan_win2675,scan_win2676,scan_win2677,scan_win2678,scan_win2679,scan_win2680,scan_win2681,scan_win2682,scan_win2683,scan_win2684,scan_win2685,scan_win2686,scan_win2687,scan_win2688,scan_win2689,scan_win2690,scan_win2691,scan_win2692,scan_win2693,scan_win2694,scan_win2695,scan_win2696,scan_win2697,scan_win2698,scan_win2699,scan_win2700,scan_win2701,scan_win2702,scan_win2703,scan_win2704,scan_win2705,scan_win2706,scan_win2707,scan_win2708,scan_win2709,scan_win2710,scan_win2711,scan_win2712,scan_win2713,scan_win2714,scan_win2715,scan_win2716,scan_win2717,scan_win2718,scan_win2719,scan_win2720,scan_win2721,scan_win2722,scan_win2723,scan_win2724,scan_win2725,scan_win2726,scan_win2727,scan_win2728,scan_win2729,scan_win2730,scan_win2731,scan_win2732,scan_win2733,scan_win2734,scan_win2735,scan_win2736,scan_win2737,scan_win2738,scan_win2739,scan_win2740,scan_win2741,scan_win2742,scan_win2743,scan_win2744,scan_win2745,scan_win2746,scan_win2747,scan_win2748,scan_win2749,scan_win2750,scan_win2751,scan_win2752,scan_win2753,scan_win2754,scan_win2755,scan_win2756,scan_win2757,scan_win2758,scan_win2759,scan_win2760,scan_win2761,scan_win2762,scan_win2763,scan_win2764,scan_win2765,scan_win2766,scan_win2767,scan_win2768,scan_win2769,scan_win2770,scan_win2771,scan_win2772,scan_win2773,scan_win2774,scan_win2775,scan_win2776,scan_win2777,scan_win2778,scan_win2779,scan_win2780,scan_win2781,scan_win2782,scan_win2783,scan_win2784,scan_win2785,scan_win2786,scan_win2787,scan_win2788,scan_win2789,scan_win2790,scan_win2791,scan_win2792,scan_win2793,scan_win2794,scan_win2795,scan_win2796,scan_win2797,scan_win2798,scan_win2799,scan_win2800,
  scan_win2801,scan_win2802,scan_win2803,scan_win2804,scan_win2805,scan_win2806,scan_win2807,scan_win2808,scan_win2809,scan_win2810,scan_win2811,scan_win2812,scan_win2813,scan_win2814,scan_win2815,scan_win2816,scan_win2817,scan_win2818,scan_win2819,scan_win2820,scan_win2821,scan_win2822,scan_win2823,scan_win2824,scan_win2825,scan_win2826,scan_win2827,scan_win2828,scan_win2829,scan_win2830,scan_win2831,scan_win2832,scan_win2833,scan_win2834,scan_win2835,scan_win2836,scan_win2837,scan_win2838,scan_win2839,scan_win2840,scan_win2841,scan_win2842,scan_win2843,scan_win2844,scan_win2845,scan_win2846,scan_win2847,scan_win2848,scan_win2849,scan_win2850,scan_win2851,scan_win2852,scan_win2853,scan_win2854,scan_win2855,scan_win2856,scan_win2857,scan_win2858,scan_win2859,scan_win2860,scan_win2861,scan_win2862,scan_win2863,scan_win2864,scan_win2865,scan_win2866,scan_win2867,scan_win2868,scan_win2869,scan_win2870,scan_win2871,scan_win2872,scan_win2873,scan_win2874,scan_win2875,scan_win2876,scan_win2877,scan_win2878,scan_win2879,scan_win2880,scan_win2881,scan_win2882,scan_win2883,scan_win2884,scan_win2885,scan_win2886,scan_win2887,scan_win2888,scan_win2889,scan_win2890,scan_win2891,scan_win2892,scan_win2893,scan_win2894,scan_win2895,scan_win2896,scan_win2897,scan_win2898,scan_win2899,scan_win2900,scan_win2901,scan_win2902,scan_win2903,scan_win2904,scan_win2905,scan_win2906,scan_win2907,scan_win2908,scan_win2909,scan_win2910,scan_win2911,scan_win2912;
  logic [`NUM_FEATURE-1:0][1:0][31:0] scan_coords;
  logic [`NUM_FEATURE-1:0][31:0] scan_win_std_dev;

  localparam [`NUM_STAGE:0][31:0] stage_num_feature = `STAGE_NUM_FEATURE;
  logic [`NUM_STAGE-1:0][31:0] stage_threshold = `STAGE_THRESHOLD;
  logic [`NUM_FEATURE-1:0][31:0] rectangle1_xs = `RECTANGLE1_XS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle1_ys = `RECTANGLE1_YS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle1_widths = `RECTANGLE1_WIDTHS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle1_heights = `RECTANGLE1_HEIGHTS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle1_weights = `RECTANGLE1_WEIGHTS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle2_xs = `RECTANGLE2_XS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle2_ys = `RECTANGLE2_YS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle2_widths = `RECTANGLE2_WIDTHS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle2_heights = `RECTANGLE2_HEIGHTS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle2_weights = `RECTANGLE2_WEIGHTS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle3_xs = `RECTANGLE3_XS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle3_ys = `RECTANGLE3_YS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle3_widths = `RECTANGLE3_WIDTHS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle3_heights = `RECTANGLE3_HEIGHTS;
  logic [`NUM_FEATURE-1:0][31:0] rectangle3_weights = `RECTANGLE3_WEIGHTS;
  logic [`NUM_FEATURE-1:0][31:0] feature_threshold = `FEATURE_THRESHOLD;
  logic [`NUM_FEATURE-1:0][31:0] feature_aboves = `FEATURE_ABOVE;
  logic [`NUM_FEATURE-1:0][31:0] feature_belows = `FEATURE_BELOW;

  always_ff @(posedge clock, posedge reset) begin: set_scan_coords_and_scan_win_std_devs
    if (reset) begin: reset_scanning_windows
       scan_coords <= 'd0;
       scan_win_std_dev <= 'd0;
       top_left <= 'd0;
    end else begin: move_scan_coords_and_scan_win_std_devs
      scan_coords[0] <= scan_win_index;
      scan_win_std_dev[0] <= input_std_dev;
      for (int i = 0; i < `NUM_FEATURE-1; i++) begin
        scan_coords[i+1] <= scan_coords[i];
        scan_win_std_dev[i+1] <= scan_win_std_dev[i];
      end
      top_left <= scan_coords[`NUM_FEATURE-1];
    end
  end

  logic [`NUM_FEATURE-1:0][31:0] rectangle1_vals, rectangle2_vals, rectangle3_vals,
                                rectangle1_products, rectangle2_products, rectangle3_products,
                                feature_sums, feature_thresholds, feature_products,
                                feature_accums;
  logic [`NUM_FEATURE-1:0] feature_comparisons;

  logic [`NUM_FEATURE:0][31:0] stage_accums; // stage_accums[0] is wire to zero and stage_accums[2913] is reg to zero
  logic [`NUM_FEATURE:0] is_feature; // is_feature[0] is wire to one and is_feature[2913] is reg to face_coords_ready
  logic [`NUM_STAGE:1] stage_comparisons;
  assign top_left_ready = is_feature[`NUM_FEATURE];

  always_ff @(posedge clock, posedge reset) begin: set_accums_and_is_feature
    if (reset) begin
      for (int m = 1; m < `NUM_FEATURE; m++) begin
        stage_accums[m] <= 32'd0;
        is_feature[m] <= 1'd0;
      end
      stage_accums[0] <= 32'd0;
      is_feature[0] <= 1'd1;
    end else begin
      stage_accums[0] <= 32'd0;
      is_feature[0] <= 1'd1;
      for (int k = 1; k < 26; k++) begin
        for (int l = stage_num_feature[k-1]; l < stage_num_feature[k] - 1; l++) begin
          stage_accums[l+1] <= stage_accums[l] + feature_accums[l];
          is_feature[l+1] <= is_feature[l];
        end
        is_feature[stage_num_feature[k]] <= stage_comparisons[k] & is_feature[stage_num_feature[k] - 1];
        stage_accums[stage_num_feature[k]] <= 32'd0;
      end
    end
  end

  genvar m;
  generate
    for (m = 1; m < `NUM_STAGE+1; m=m+1) begin: stage_threshold_check
      signed_comparator stage_c(.gt(stage_comparisons[m]), .A(stage_accums[stage_num_feature[m] - 1] + feature_accums[stage_num_feature[m] - 1]), .B(stage_threshold[m-1]));
    end
  endgenerate

  always_ff @(posedge clock, posedge reset) begin : set_scan_wins
    if (reset) begin: reset_scan_wins
      scan_win0 <= 32'd0; 
      scan_win1 <= 32'd0; scan_win2 <= 32'd0; scan_win3 <= 32'd0; scan_win4 <= 32'd0; scan_win5 <= 32'd0; scan_win6 <= 32'd0; scan_win7 <= 32'd0; scan_win8 <= 32'd0; scan_win9 <= 32'd0; scan_win10 <= 32'd0; scan_win11 <= 32'd0; scan_win12 <= 32'd0; scan_win13 <= 32'd0; scan_win14 <= 32'd0; scan_win15 <= 32'd0; scan_win16 <= 32'd0; scan_win17 <= 32'd0; scan_win18 <= 32'd0; scan_win19 <= 32'd0; scan_win20 <= 32'd0; scan_win21 <= 32'd0; scan_win22 <= 32'd0; scan_win23 <= 32'd0; scan_win24 <= 32'd0; scan_win25 <= 32'd0; scan_win26 <= 32'd0; scan_win27 <= 32'd0; scan_win28 <= 32'd0; scan_win29 <= 32'd0; scan_win30 <= 32'd0; scan_win31 <= 32'd0; scan_win32 <= 32'd0; scan_win33 <= 32'd0; scan_win34 <= 32'd0; scan_win35 <= 32'd0; scan_win36 <= 32'd0; scan_win37 <= 32'd0; scan_win38 <= 32'd0; scan_win39 <= 32'd0; scan_win40 <= 32'd0; scan_win41 <= 32'd0; scan_win42 <= 32'd0; scan_win43 <= 32'd0; scan_win44 <= 32'd0; scan_win45 <= 32'd0; scan_win46 <= 32'd0; scan_win47 <= 32'd0; scan_win48 <= 32'd0; scan_win49 <= 32'd0; scan_win50 <= 32'd0; scan_win51 <= 32'd0; scan_win52 <= 32'd0; scan_win53 <= 32'd0; scan_win54 <= 32'd0; scan_win55 <= 32'd0; scan_win56 <= 32'd0; scan_win57 <= 32'd0; scan_win58 <= 32'd0; scan_win59 <= 32'd0; scan_win60 <= 32'd0; scan_win61 <= 32'd0; scan_win62 <= 32'd0; scan_win63 <= 32'd0; scan_win64 <= 32'd0; scan_win65 <= 32'd0; scan_win66 <= 32'd0; scan_win67 <= 32'd0; scan_win68 <= 32'd0; scan_win69 <= 32'd0; scan_win70 <= 32'd0; scan_win71 <= 32'd0; scan_win72 <= 32'd0; scan_win73 <= 32'd0; scan_win74 <= 32'd0; scan_win75 <= 32'd0; scan_win76 <= 32'd0; scan_win77 <= 32'd0; scan_win78 <= 32'd0; scan_win79 <= 32'd0; scan_win80 <= 32'd0; scan_win81 <= 32'd0; scan_win82 <= 32'd0; scan_win83 <= 32'd0; scan_win84 <= 32'd0; scan_win85 <= 32'd0; scan_win86 <= 32'd0; scan_win87 <= 32'd0; scan_win88 <= 32'd0; scan_win89 <= 32'd0; scan_win90 <= 32'd0; scan_win91 <= 32'd0; scan_win92 <= 32'd0; scan_win93 <= 32'd0; scan_win94 <= 32'd0; scan_win95 <= 32'd0; scan_win96 <= 32'd0; scan_win97 <= 32'd0; scan_win98 <= 32'd0; scan_win99 <= 32'd0; scan_win100 <= 32'd0; scan_win101 <= 32'd0; scan_win102 <= 32'd0; scan_win103 <= 32'd0; scan_win104 <= 32'd0; scan_win105 <= 32'd0; scan_win106 <= 32'd0; scan_win107 <= 32'd0; scan_win108 <= 32'd0; scan_win109 <= 32'd0; scan_win110 <= 32'd0; scan_win111 <= 32'd0; scan_win112 <= 32'd0; scan_win113 <= 32'd0; scan_win114 <= 32'd0; scan_win115 <= 32'd0; scan_win116 <= 32'd0; scan_win117 <= 32'd0; scan_win118 <= 32'd0; scan_win119 <= 32'd0; scan_win120 <= 32'd0; scan_win121 <= 32'd0; scan_win122 <= 32'd0; scan_win123 <= 32'd0; scan_win124 <= 32'd0; scan_win125 <= 32'd0; scan_win126 <= 32'd0; scan_win127 <= 32'd0; scan_win128 <= 32'd0; scan_win129 <= 32'd0; scan_win130 <= 32'd0; scan_win131 <= 32'd0; scan_win132 <= 32'd0; scan_win133 <= 32'd0; scan_win134 <= 32'd0; scan_win135 <= 32'd0; scan_win136 <= 32'd0; scan_win137 <= 32'd0; scan_win138 <= 32'd0; scan_win139 <= 32'd0; scan_win140 <= 32'd0; scan_win141 <= 32'd0; scan_win142 <= 32'd0; scan_win143 <= 32'd0; scan_win144 <= 32'd0; scan_win145 <= 32'd0; scan_win146 <= 32'd0; scan_win147 <= 32'd0; scan_win148 <= 32'd0; scan_win149 <= 32'd0; scan_win150 <= 32'd0; scan_win151 <= 32'd0; scan_win152 <= 32'd0; scan_win153 <= 32'd0; scan_win154 <= 32'd0; scan_win155 <= 32'd0; scan_win156 <= 32'd0; scan_win157 <= 32'd0; scan_win158 <= 32'd0; scan_win159 <= 32'd0; scan_win160 <= 32'd0; scan_win161 <= 32'd0; scan_win162 <= 32'd0; scan_win163 <= 32'd0; scan_win164 <= 32'd0; scan_win165 <= 32'd0; scan_win166 <= 32'd0; scan_win167 <= 32'd0; scan_win168 <= 32'd0; scan_win169 <= 32'd0; scan_win170 <= 32'd0; scan_win171 <= 32'd0; scan_win172 <= 32'd0; scan_win173 <= 32'd0; scan_win174 <= 32'd0; scan_win175 <= 32'd0; scan_win176 <= 32'd0; scan_win177 <= 32'd0; scan_win178 <= 32'd0; scan_win179 <= 32'd0; scan_win180 <= 32'd0; scan_win181 <= 32'd0; scan_win182 <= 32'd0; scan_win183 <= 32'd0; scan_win184 <= 32'd0; scan_win185 <= 32'd0; scan_win186 <= 32'd0; scan_win187 <= 32'd0; scan_win188 <= 32'd0; scan_win189 <= 32'd0; scan_win190 <= 32'd0; scan_win191 <= 32'd0; scan_win192 <= 32'd0; scan_win193 <= 32'd0; scan_win194 <= 32'd0; scan_win195 <= 32'd0; scan_win196 <= 32'd0; scan_win197 <= 32'd0; scan_win198 <= 32'd0; scan_win199 <= 32'd0; scan_win200 <= 32'd0; 
      scan_win201 <= 32'd0; scan_win202 <= 32'd0; scan_win203 <= 32'd0; scan_win204 <= 32'd0; scan_win205 <= 32'd0; scan_win206 <= 32'd0; scan_win207 <= 32'd0; scan_win208 <= 32'd0; scan_win209 <= 32'd0; scan_win210 <= 32'd0; scan_win211 <= 32'd0; scan_win212 <= 32'd0; scan_win213 <= 32'd0; scan_win214 <= 32'd0; scan_win215 <= 32'd0; scan_win216 <= 32'd0; scan_win217 <= 32'd0; scan_win218 <= 32'd0; scan_win219 <= 32'd0; scan_win220 <= 32'd0; scan_win221 <= 32'd0; scan_win222 <= 32'd0; scan_win223 <= 32'd0; scan_win224 <= 32'd0; scan_win225 <= 32'd0; scan_win226 <= 32'd0; scan_win227 <= 32'd0; scan_win228 <= 32'd0; scan_win229 <= 32'd0; scan_win230 <= 32'd0; scan_win231 <= 32'd0; scan_win232 <= 32'd0; scan_win233 <= 32'd0; scan_win234 <= 32'd0; scan_win235 <= 32'd0; scan_win236 <= 32'd0; scan_win237 <= 32'd0; scan_win238 <= 32'd0; scan_win239 <= 32'd0; scan_win240 <= 32'd0; scan_win241 <= 32'd0; scan_win242 <= 32'd0; scan_win243 <= 32'd0; scan_win244 <= 32'd0; scan_win245 <= 32'd0; scan_win246 <= 32'd0; scan_win247 <= 32'd0; scan_win248 <= 32'd0; scan_win249 <= 32'd0; scan_win250 <= 32'd0; scan_win251 <= 32'd0; scan_win252 <= 32'd0; scan_win253 <= 32'd0; scan_win254 <= 32'd0; scan_win255 <= 32'd0; scan_win256 <= 32'd0; scan_win257 <= 32'd0; scan_win258 <= 32'd0; scan_win259 <= 32'd0; scan_win260 <= 32'd0; scan_win261 <= 32'd0; scan_win262 <= 32'd0; scan_win263 <= 32'd0; scan_win264 <= 32'd0; scan_win265 <= 32'd0; scan_win266 <= 32'd0; scan_win267 <= 32'd0; scan_win268 <= 32'd0; scan_win269 <= 32'd0; scan_win270 <= 32'd0; scan_win271 <= 32'd0; scan_win272 <= 32'd0; scan_win273 <= 32'd0; scan_win274 <= 32'd0; scan_win275 <= 32'd0; scan_win276 <= 32'd0; scan_win277 <= 32'd0; scan_win278 <= 32'd0; scan_win279 <= 32'd0; scan_win280 <= 32'd0; scan_win281 <= 32'd0; scan_win282 <= 32'd0; scan_win283 <= 32'd0; scan_win284 <= 32'd0; scan_win285 <= 32'd0; scan_win286 <= 32'd0; scan_win287 <= 32'd0; scan_win288 <= 32'd0; scan_win289 <= 32'd0; scan_win290 <= 32'd0; scan_win291 <= 32'd0; scan_win292 <= 32'd0; scan_win293 <= 32'd0; scan_win294 <= 32'd0; scan_win295 <= 32'd0; scan_win296 <= 32'd0; scan_win297 <= 32'd0; scan_win298 <= 32'd0; scan_win299 <= 32'd0; scan_win300 <= 32'd0; scan_win301 <= 32'd0; scan_win302 <= 32'd0; scan_win303 <= 32'd0; scan_win304 <= 32'd0; scan_win305 <= 32'd0; scan_win306 <= 32'd0; scan_win307 <= 32'd0; scan_win308 <= 32'd0; scan_win309 <= 32'd0; scan_win310 <= 32'd0; scan_win311 <= 32'd0; scan_win312 <= 32'd0; scan_win313 <= 32'd0; scan_win314 <= 32'd0; scan_win315 <= 32'd0; scan_win316 <= 32'd0; scan_win317 <= 32'd0; scan_win318 <= 32'd0; scan_win319 <= 32'd0; scan_win320 <= 32'd0; scan_win321 <= 32'd0; scan_win322 <= 32'd0; scan_win323 <= 32'd0; scan_win324 <= 32'd0; scan_win325 <= 32'd0; scan_win326 <= 32'd0; scan_win327 <= 32'd0; scan_win328 <= 32'd0; scan_win329 <= 32'd0; scan_win330 <= 32'd0; scan_win331 <= 32'd0; scan_win332 <= 32'd0; scan_win333 <= 32'd0; scan_win334 <= 32'd0; scan_win335 <= 32'd0; scan_win336 <= 32'd0; scan_win337 <= 32'd0; scan_win338 <= 32'd0; scan_win339 <= 32'd0; scan_win340 <= 32'd0; scan_win341 <= 32'd0; scan_win342 <= 32'd0; scan_win343 <= 32'd0; scan_win344 <= 32'd0; scan_win345 <= 32'd0; scan_win346 <= 32'd0; scan_win347 <= 32'd0; scan_win348 <= 32'd0; scan_win349 <= 32'd0; scan_win350 <= 32'd0; scan_win351 <= 32'd0; scan_win352 <= 32'd0; scan_win353 <= 32'd0; scan_win354 <= 32'd0; scan_win355 <= 32'd0; scan_win356 <= 32'd0; scan_win357 <= 32'd0; scan_win358 <= 32'd0; scan_win359 <= 32'd0; scan_win360 <= 32'd0; scan_win361 <= 32'd0; scan_win362 <= 32'd0; scan_win363 <= 32'd0; scan_win364 <= 32'd0; scan_win365 <= 32'd0; scan_win366 <= 32'd0; scan_win367 <= 32'd0; scan_win368 <= 32'd0; scan_win369 <= 32'd0; scan_win370 <= 32'd0; scan_win371 <= 32'd0; scan_win372 <= 32'd0; scan_win373 <= 32'd0; scan_win374 <= 32'd0; scan_win375 <= 32'd0; scan_win376 <= 32'd0; scan_win377 <= 32'd0; scan_win378 <= 32'd0; scan_win379 <= 32'd0; scan_win380 <= 32'd0; scan_win381 <= 32'd0; scan_win382 <= 32'd0; scan_win383 <= 32'd0; scan_win384 <= 32'd0; scan_win385 <= 32'd0; scan_win386 <= 32'd0; scan_win387 <= 32'd0; scan_win388 <= 32'd0; scan_win389 <= 32'd0; scan_win390 <= 32'd0; scan_win391 <= 32'd0; scan_win392 <= 32'd0; scan_win393 <= 32'd0; scan_win394 <= 32'd0; scan_win395 <= 32'd0; scan_win396 <= 32'd0; scan_win397 <= 32'd0; scan_win398 <= 32'd0; scan_win399 <= 32'd0; scan_win400 <= 32'd0; 
      scan_win401 <= 32'd0; scan_win402 <= 32'd0; scan_win403 <= 32'd0; scan_win404 <= 32'd0; scan_win405 <= 32'd0; scan_win406 <= 32'd0; scan_win407 <= 32'd0; scan_win408 <= 32'd0; scan_win409 <= 32'd0; scan_win410 <= 32'd0; scan_win411 <= 32'd0; scan_win412 <= 32'd0; scan_win413 <= 32'd0; scan_win414 <= 32'd0; scan_win415 <= 32'd0; scan_win416 <= 32'd0; scan_win417 <= 32'd0; scan_win418 <= 32'd0; scan_win419 <= 32'd0; scan_win420 <= 32'd0; scan_win421 <= 32'd0; scan_win422 <= 32'd0; scan_win423 <= 32'd0; scan_win424 <= 32'd0; scan_win425 <= 32'd0; scan_win426 <= 32'd0; scan_win427 <= 32'd0; scan_win428 <= 32'd0; scan_win429 <= 32'd0; scan_win430 <= 32'd0; scan_win431 <= 32'd0; scan_win432 <= 32'd0; scan_win433 <= 32'd0; scan_win434 <= 32'd0; scan_win435 <= 32'd0; scan_win436 <= 32'd0; scan_win437 <= 32'd0; scan_win438 <= 32'd0; scan_win439 <= 32'd0; scan_win440 <= 32'd0; scan_win441 <= 32'd0; scan_win442 <= 32'd0; scan_win443 <= 32'd0; scan_win444 <= 32'd0; scan_win445 <= 32'd0; scan_win446 <= 32'd0; scan_win447 <= 32'd0; scan_win448 <= 32'd0; scan_win449 <= 32'd0; scan_win450 <= 32'd0; scan_win451 <= 32'd0; scan_win452 <= 32'd0; scan_win453 <= 32'd0; scan_win454 <= 32'd0; scan_win455 <= 32'd0; scan_win456 <= 32'd0; scan_win457 <= 32'd0; scan_win458 <= 32'd0; scan_win459 <= 32'd0; scan_win460 <= 32'd0; scan_win461 <= 32'd0; scan_win462 <= 32'd0; scan_win463 <= 32'd0; scan_win464 <= 32'd0; scan_win465 <= 32'd0; scan_win466 <= 32'd0; scan_win467 <= 32'd0; scan_win468 <= 32'd0; scan_win469 <= 32'd0; scan_win470 <= 32'd0; scan_win471 <= 32'd0; scan_win472 <= 32'd0; scan_win473 <= 32'd0; scan_win474 <= 32'd0; scan_win475 <= 32'd0; scan_win476 <= 32'd0; scan_win477 <= 32'd0; scan_win478 <= 32'd0; scan_win479 <= 32'd0; scan_win480 <= 32'd0; scan_win481 <= 32'd0; scan_win482 <= 32'd0; scan_win483 <= 32'd0; scan_win484 <= 32'd0; scan_win485 <= 32'd0; scan_win486 <= 32'd0; scan_win487 <= 32'd0; scan_win488 <= 32'd0; scan_win489 <= 32'd0; scan_win490 <= 32'd0; scan_win491 <= 32'd0; scan_win492 <= 32'd0; scan_win493 <= 32'd0; scan_win494 <= 32'd0; scan_win495 <= 32'd0; scan_win496 <= 32'd0; scan_win497 <= 32'd0; scan_win498 <= 32'd0; scan_win499 <= 32'd0; scan_win500 <= 32'd0; scan_win501 <= 32'd0; scan_win502 <= 32'd0; scan_win503 <= 32'd0; scan_win504 <= 32'd0; scan_win505 <= 32'd0; scan_win506 <= 32'd0; scan_win507 <= 32'd0; scan_win508 <= 32'd0; scan_win509 <= 32'd0; scan_win510 <= 32'd0; scan_win511 <= 32'd0; scan_win512 <= 32'd0; scan_win513 <= 32'd0; scan_win514 <= 32'd0; scan_win515 <= 32'd0; scan_win516 <= 32'd0; scan_win517 <= 32'd0; scan_win518 <= 32'd0; scan_win519 <= 32'd0; scan_win520 <= 32'd0; scan_win521 <= 32'd0; scan_win522 <= 32'd0; scan_win523 <= 32'd0; scan_win524 <= 32'd0; scan_win525 <= 32'd0; scan_win526 <= 32'd0; scan_win527 <= 32'd0; scan_win528 <= 32'd0; scan_win529 <= 32'd0; scan_win530 <= 32'd0; scan_win531 <= 32'd0; scan_win532 <= 32'd0; scan_win533 <= 32'd0; scan_win534 <= 32'd0; scan_win535 <= 32'd0; scan_win536 <= 32'd0; scan_win537 <= 32'd0; scan_win538 <= 32'd0; scan_win539 <= 32'd0; scan_win540 <= 32'd0; scan_win541 <= 32'd0; scan_win542 <= 32'd0; scan_win543 <= 32'd0; scan_win544 <= 32'd0; scan_win545 <= 32'd0; scan_win546 <= 32'd0; scan_win547 <= 32'd0; scan_win548 <= 32'd0; scan_win549 <= 32'd0; scan_win550 <= 32'd0; scan_win551 <= 32'd0; scan_win552 <= 32'd0; scan_win553 <= 32'd0; scan_win554 <= 32'd0; scan_win555 <= 32'd0; scan_win556 <= 32'd0; scan_win557 <= 32'd0; scan_win558 <= 32'd0; scan_win559 <= 32'd0; scan_win560 <= 32'd0; scan_win561 <= 32'd0; scan_win562 <= 32'd0; scan_win563 <= 32'd0; scan_win564 <= 32'd0; scan_win565 <= 32'd0; scan_win566 <= 32'd0; scan_win567 <= 32'd0; scan_win568 <= 32'd0; scan_win569 <= 32'd0; scan_win570 <= 32'd0; scan_win571 <= 32'd0; scan_win572 <= 32'd0; scan_win573 <= 32'd0; scan_win574 <= 32'd0; scan_win575 <= 32'd0; scan_win576 <= 32'd0; scan_win577 <= 32'd0; scan_win578 <= 32'd0; scan_win579 <= 32'd0; scan_win580 <= 32'd0; scan_win581 <= 32'd0; scan_win582 <= 32'd0; scan_win583 <= 32'd0; scan_win584 <= 32'd0; scan_win585 <= 32'd0; scan_win586 <= 32'd0; scan_win587 <= 32'd0; scan_win588 <= 32'd0; scan_win589 <= 32'd0; scan_win590 <= 32'd0; scan_win591 <= 32'd0; scan_win592 <= 32'd0; scan_win593 <= 32'd0; scan_win594 <= 32'd0; scan_win595 <= 32'd0; scan_win596 <= 32'd0; scan_win597 <= 32'd0; scan_win598 <= 32'd0; scan_win599 <= 32'd0; scan_win600 <= 32'd0; 
      scan_win601 <= 32'd0; scan_win602 <= 32'd0; scan_win603 <= 32'd0; scan_win604 <= 32'd0; scan_win605 <= 32'd0; scan_win606 <= 32'd0; scan_win607 <= 32'd0; scan_win608 <= 32'd0; scan_win609 <= 32'd0; scan_win610 <= 32'd0; scan_win611 <= 32'd0; scan_win612 <= 32'd0; scan_win613 <= 32'd0; scan_win614 <= 32'd0; scan_win615 <= 32'd0; scan_win616 <= 32'd0; scan_win617 <= 32'd0; scan_win618 <= 32'd0; scan_win619 <= 32'd0; scan_win620 <= 32'd0; scan_win621 <= 32'd0; scan_win622 <= 32'd0; scan_win623 <= 32'd0; scan_win624 <= 32'd0; scan_win625 <= 32'd0; scan_win626 <= 32'd0; scan_win627 <= 32'd0; scan_win628 <= 32'd0; scan_win629 <= 32'd0; scan_win630 <= 32'd0; scan_win631 <= 32'd0; scan_win632 <= 32'd0; scan_win633 <= 32'd0; scan_win634 <= 32'd0; scan_win635 <= 32'd0; scan_win636 <= 32'd0; scan_win637 <= 32'd0; scan_win638 <= 32'd0; scan_win639 <= 32'd0; scan_win640 <= 32'd0; scan_win641 <= 32'd0; scan_win642 <= 32'd0; scan_win643 <= 32'd0; scan_win644 <= 32'd0; scan_win645 <= 32'd0; scan_win646 <= 32'd0; scan_win647 <= 32'd0; scan_win648 <= 32'd0; scan_win649 <= 32'd0; scan_win650 <= 32'd0; scan_win651 <= 32'd0; scan_win652 <= 32'd0; scan_win653 <= 32'd0; scan_win654 <= 32'd0; scan_win655 <= 32'd0; scan_win656 <= 32'd0; scan_win657 <= 32'd0; scan_win658 <= 32'd0; scan_win659 <= 32'd0; scan_win660 <= 32'd0; scan_win661 <= 32'd0; scan_win662 <= 32'd0; scan_win663 <= 32'd0; scan_win664 <= 32'd0; scan_win665 <= 32'd0; scan_win666 <= 32'd0; scan_win667 <= 32'd0; scan_win668 <= 32'd0; scan_win669 <= 32'd0; scan_win670 <= 32'd0; scan_win671 <= 32'd0; scan_win672 <= 32'd0; scan_win673 <= 32'd0; scan_win674 <= 32'd0; scan_win675 <= 32'd0; scan_win676 <= 32'd0; scan_win677 <= 32'd0; scan_win678 <= 32'd0; scan_win679 <= 32'd0; scan_win680 <= 32'd0; scan_win681 <= 32'd0; scan_win682 <= 32'd0; scan_win683 <= 32'd0; scan_win684 <= 32'd0; scan_win685 <= 32'd0; scan_win686 <= 32'd0; scan_win687 <= 32'd0; scan_win688 <= 32'd0; scan_win689 <= 32'd0; scan_win690 <= 32'd0; scan_win691 <= 32'd0; scan_win692 <= 32'd0; scan_win693 <= 32'd0; scan_win694 <= 32'd0; scan_win695 <= 32'd0; scan_win696 <= 32'd0; scan_win697 <= 32'd0; scan_win698 <= 32'd0; scan_win699 <= 32'd0; scan_win700 <= 32'd0; scan_win701 <= 32'd0; scan_win702 <= 32'd0; scan_win703 <= 32'd0; scan_win704 <= 32'd0; scan_win705 <= 32'd0; scan_win706 <= 32'd0; scan_win707 <= 32'd0; scan_win708 <= 32'd0; scan_win709 <= 32'd0; scan_win710 <= 32'd0; scan_win711 <= 32'd0; scan_win712 <= 32'd0; scan_win713 <= 32'd0; scan_win714 <= 32'd0; scan_win715 <= 32'd0; scan_win716 <= 32'd0; scan_win717 <= 32'd0; scan_win718 <= 32'd0; scan_win719 <= 32'd0; scan_win720 <= 32'd0; scan_win721 <= 32'd0; scan_win722 <= 32'd0; scan_win723 <= 32'd0; scan_win724 <= 32'd0; scan_win725 <= 32'd0; scan_win726 <= 32'd0; scan_win727 <= 32'd0; scan_win728 <= 32'd0; scan_win729 <= 32'd0; scan_win730 <= 32'd0; scan_win731 <= 32'd0; scan_win732 <= 32'd0; scan_win733 <= 32'd0; scan_win734 <= 32'd0; scan_win735 <= 32'd0; scan_win736 <= 32'd0; scan_win737 <= 32'd0; scan_win738 <= 32'd0; scan_win739 <= 32'd0; scan_win740 <= 32'd0; scan_win741 <= 32'd0; scan_win742 <= 32'd0; scan_win743 <= 32'd0; scan_win744 <= 32'd0; scan_win745 <= 32'd0; scan_win746 <= 32'd0; scan_win747 <= 32'd0; scan_win748 <= 32'd0; scan_win749 <= 32'd0; scan_win750 <= 32'd0; scan_win751 <= 32'd0; scan_win752 <= 32'd0; scan_win753 <= 32'd0; scan_win754 <= 32'd0; scan_win755 <= 32'd0; scan_win756 <= 32'd0; scan_win757 <= 32'd0; scan_win758 <= 32'd0; scan_win759 <= 32'd0; scan_win760 <= 32'd0; scan_win761 <= 32'd0; scan_win762 <= 32'd0; scan_win763 <= 32'd0; scan_win764 <= 32'd0; scan_win765 <= 32'd0; scan_win766 <= 32'd0; scan_win767 <= 32'd0; scan_win768 <= 32'd0; scan_win769 <= 32'd0; scan_win770 <= 32'd0; scan_win771 <= 32'd0; scan_win772 <= 32'd0; scan_win773 <= 32'd0; scan_win774 <= 32'd0; scan_win775 <= 32'd0; scan_win776 <= 32'd0; scan_win777 <= 32'd0; scan_win778 <= 32'd0; scan_win779 <= 32'd0; scan_win780 <= 32'd0; scan_win781 <= 32'd0; scan_win782 <= 32'd0; scan_win783 <= 32'd0; scan_win784 <= 32'd0; scan_win785 <= 32'd0; scan_win786 <= 32'd0; scan_win787 <= 32'd0; scan_win788 <= 32'd0; scan_win789 <= 32'd0; scan_win790 <= 32'd0; scan_win791 <= 32'd0; scan_win792 <= 32'd0; scan_win793 <= 32'd0; scan_win794 <= 32'd0; scan_win795 <= 32'd0; scan_win796 <= 32'd0; scan_win797 <= 32'd0; scan_win798 <= 32'd0; scan_win799 <= 32'd0; scan_win800 <= 32'd0; 
      scan_win801 <= 32'd0; scan_win802 <= 32'd0; scan_win803 <= 32'd0; scan_win804 <= 32'd0; scan_win805 <= 32'd0; scan_win806 <= 32'd0; scan_win807 <= 32'd0; scan_win808 <= 32'd0; scan_win809 <= 32'd0; scan_win810 <= 32'd0; scan_win811 <= 32'd0; scan_win812 <= 32'd0; scan_win813 <= 32'd0; scan_win814 <= 32'd0; scan_win815 <= 32'd0; scan_win816 <= 32'd0; scan_win817 <= 32'd0; scan_win818 <= 32'd0; scan_win819 <= 32'd0; scan_win820 <= 32'd0; scan_win821 <= 32'd0; scan_win822 <= 32'd0; scan_win823 <= 32'd0; scan_win824 <= 32'd0; scan_win825 <= 32'd0; scan_win826 <= 32'd0; scan_win827 <= 32'd0; scan_win828 <= 32'd0; scan_win829 <= 32'd0; scan_win830 <= 32'd0; scan_win831 <= 32'd0; scan_win832 <= 32'd0; scan_win833 <= 32'd0; scan_win834 <= 32'd0; scan_win835 <= 32'd0; scan_win836 <= 32'd0; scan_win837 <= 32'd0; scan_win838 <= 32'd0; scan_win839 <= 32'd0; scan_win840 <= 32'd0; scan_win841 <= 32'd0; scan_win842 <= 32'd0; scan_win843 <= 32'd0; scan_win844 <= 32'd0; scan_win845 <= 32'd0; scan_win846 <= 32'd0; scan_win847 <= 32'd0; scan_win848 <= 32'd0; scan_win849 <= 32'd0; scan_win850 <= 32'd0; scan_win851 <= 32'd0; scan_win852 <= 32'd0; scan_win853 <= 32'd0; scan_win854 <= 32'd0; scan_win855 <= 32'd0; scan_win856 <= 32'd0; scan_win857 <= 32'd0; scan_win858 <= 32'd0; scan_win859 <= 32'd0; scan_win860 <= 32'd0; scan_win861 <= 32'd0; scan_win862 <= 32'd0; scan_win863 <= 32'd0; scan_win864 <= 32'd0; scan_win865 <= 32'd0; scan_win866 <= 32'd0; scan_win867 <= 32'd0; scan_win868 <= 32'd0; scan_win869 <= 32'd0; scan_win870 <= 32'd0; scan_win871 <= 32'd0; scan_win872 <= 32'd0; scan_win873 <= 32'd0; scan_win874 <= 32'd0; scan_win875 <= 32'd0; scan_win876 <= 32'd0; scan_win877 <= 32'd0; scan_win878 <= 32'd0; scan_win879 <= 32'd0; scan_win880 <= 32'd0; scan_win881 <= 32'd0; scan_win882 <= 32'd0; scan_win883 <= 32'd0; scan_win884 <= 32'd0; scan_win885 <= 32'd0; scan_win886 <= 32'd0; scan_win887 <= 32'd0; scan_win888 <= 32'd0; scan_win889 <= 32'd0; scan_win890 <= 32'd0; scan_win891 <= 32'd0; scan_win892 <= 32'd0; scan_win893 <= 32'd0; scan_win894 <= 32'd0; scan_win895 <= 32'd0; scan_win896 <= 32'd0; scan_win897 <= 32'd0; scan_win898 <= 32'd0; scan_win899 <= 32'd0; scan_win900 <= 32'd0; scan_win901 <= 32'd0; scan_win902 <= 32'd0; scan_win903 <= 32'd0; scan_win904 <= 32'd0; scan_win905 <= 32'd0; scan_win906 <= 32'd0; scan_win907 <= 32'd0; scan_win908 <= 32'd0; scan_win909 <= 32'd0; scan_win910 <= 32'd0; scan_win911 <= 32'd0; scan_win912 <= 32'd0; scan_win913 <= 32'd0; scan_win914 <= 32'd0; scan_win915 <= 32'd0; scan_win916 <= 32'd0; scan_win917 <= 32'd0; scan_win918 <= 32'd0; scan_win919 <= 32'd0; scan_win920 <= 32'd0; scan_win921 <= 32'd0; scan_win922 <= 32'd0; scan_win923 <= 32'd0; scan_win924 <= 32'd0; scan_win925 <= 32'd0; scan_win926 <= 32'd0; scan_win927 <= 32'd0; scan_win928 <= 32'd0; scan_win929 <= 32'd0; scan_win930 <= 32'd0; scan_win931 <= 32'd0; scan_win932 <= 32'd0; scan_win933 <= 32'd0; scan_win934 <= 32'd0; scan_win935 <= 32'd0; scan_win936 <= 32'd0; scan_win937 <= 32'd0; scan_win938 <= 32'd0; scan_win939 <= 32'd0; scan_win940 <= 32'd0; scan_win941 <= 32'd0; scan_win942 <= 32'd0; scan_win943 <= 32'd0; scan_win944 <= 32'd0; scan_win945 <= 32'd0; scan_win946 <= 32'd0; scan_win947 <= 32'd0; scan_win948 <= 32'd0; scan_win949 <= 32'd0; scan_win950 <= 32'd0; scan_win951 <= 32'd0; scan_win952 <= 32'd0; scan_win953 <= 32'd0; scan_win954 <= 32'd0; scan_win955 <= 32'd0; scan_win956 <= 32'd0; scan_win957 <= 32'd0; scan_win958 <= 32'd0; scan_win959 <= 32'd0; scan_win960 <= 32'd0; scan_win961 <= 32'd0; scan_win962 <= 32'd0; scan_win963 <= 32'd0; scan_win964 <= 32'd0; scan_win965 <= 32'd0; scan_win966 <= 32'd0; scan_win967 <= 32'd0; scan_win968 <= 32'd0; scan_win969 <= 32'd0; scan_win970 <= 32'd0; scan_win971 <= 32'd0; scan_win972 <= 32'd0; scan_win973 <= 32'd0; scan_win974 <= 32'd0; scan_win975 <= 32'd0; scan_win976 <= 32'd0; scan_win977 <= 32'd0; scan_win978 <= 32'd0; scan_win979 <= 32'd0; scan_win980 <= 32'd0; scan_win981 <= 32'd0; scan_win982 <= 32'd0; scan_win983 <= 32'd0; scan_win984 <= 32'd0; scan_win985 <= 32'd0; scan_win986 <= 32'd0; scan_win987 <= 32'd0; scan_win988 <= 32'd0; scan_win989 <= 32'd0; scan_win990 <= 32'd0; scan_win991 <= 32'd0; scan_win992 <= 32'd0; scan_win993 <= 32'd0; scan_win994 <= 32'd0; scan_win995 <= 32'd0; scan_win996 <= 32'd0; scan_win997 <= 32'd0; scan_win998 <= 32'd0; scan_win999 <= 32'd0; scan_win1000 <= 32'd0; 
      scan_win1001 <= 32'd0; scan_win1002 <= 32'd0; scan_win1003 <= 32'd0; scan_win1004 <= 32'd0; scan_win1005 <= 32'd0; scan_win1006 <= 32'd0; scan_win1007 <= 32'd0; scan_win1008 <= 32'd0; scan_win1009 <= 32'd0; scan_win1010 <= 32'd0; scan_win1011 <= 32'd0; scan_win1012 <= 32'd0; scan_win1013 <= 32'd0; scan_win1014 <= 32'd0; scan_win1015 <= 32'd0; scan_win1016 <= 32'd0; scan_win1017 <= 32'd0; scan_win1018 <= 32'd0; scan_win1019 <= 32'd0; scan_win1020 <= 32'd0; scan_win1021 <= 32'd0; scan_win1022 <= 32'd0; scan_win1023 <= 32'd0; scan_win1024 <= 32'd0; scan_win1025 <= 32'd0; scan_win1026 <= 32'd0; scan_win1027 <= 32'd0; scan_win1028 <= 32'd0; scan_win1029 <= 32'd0; scan_win1030 <= 32'd0; scan_win1031 <= 32'd0; scan_win1032 <= 32'd0; scan_win1033 <= 32'd0; scan_win1034 <= 32'd0; scan_win1035 <= 32'd0; scan_win1036 <= 32'd0; scan_win1037 <= 32'd0; scan_win1038 <= 32'd0; scan_win1039 <= 32'd0; scan_win1040 <= 32'd0; scan_win1041 <= 32'd0; scan_win1042 <= 32'd0; scan_win1043 <= 32'd0; scan_win1044 <= 32'd0; scan_win1045 <= 32'd0; scan_win1046 <= 32'd0; scan_win1047 <= 32'd0; scan_win1048 <= 32'd0; scan_win1049 <= 32'd0; scan_win1050 <= 32'd0; scan_win1051 <= 32'd0; scan_win1052 <= 32'd0; scan_win1053 <= 32'd0; scan_win1054 <= 32'd0; scan_win1055 <= 32'd0; scan_win1056 <= 32'd0; scan_win1057 <= 32'd0; scan_win1058 <= 32'd0; scan_win1059 <= 32'd0; scan_win1060 <= 32'd0; scan_win1061 <= 32'd0; scan_win1062 <= 32'd0; scan_win1063 <= 32'd0; scan_win1064 <= 32'd0; scan_win1065 <= 32'd0; scan_win1066 <= 32'd0; scan_win1067 <= 32'd0; scan_win1068 <= 32'd0; scan_win1069 <= 32'd0; scan_win1070 <= 32'd0; scan_win1071 <= 32'd0; scan_win1072 <= 32'd0; scan_win1073 <= 32'd0; scan_win1074 <= 32'd0; scan_win1075 <= 32'd0; scan_win1076 <= 32'd0; scan_win1077 <= 32'd0; scan_win1078 <= 32'd0; scan_win1079 <= 32'd0; scan_win1080 <= 32'd0; scan_win1081 <= 32'd0; scan_win1082 <= 32'd0; scan_win1083 <= 32'd0; scan_win1084 <= 32'd0; scan_win1085 <= 32'd0; scan_win1086 <= 32'd0; scan_win1087 <= 32'd0; scan_win1088 <= 32'd0; scan_win1089 <= 32'd0; scan_win1090 <= 32'd0; scan_win1091 <= 32'd0; scan_win1092 <= 32'd0; scan_win1093 <= 32'd0; scan_win1094 <= 32'd0; scan_win1095 <= 32'd0; scan_win1096 <= 32'd0; scan_win1097 <= 32'd0; scan_win1098 <= 32'd0; scan_win1099 <= 32'd0; scan_win1100 <= 32'd0; scan_win1101 <= 32'd0; scan_win1102 <= 32'd0; scan_win1103 <= 32'd0; scan_win1104 <= 32'd0; scan_win1105 <= 32'd0; scan_win1106 <= 32'd0; scan_win1107 <= 32'd0; scan_win1108 <= 32'd0; scan_win1109 <= 32'd0; scan_win1110 <= 32'd0; scan_win1111 <= 32'd0; scan_win1112 <= 32'd0; scan_win1113 <= 32'd0; scan_win1114 <= 32'd0; scan_win1115 <= 32'd0; scan_win1116 <= 32'd0; scan_win1117 <= 32'd0; scan_win1118 <= 32'd0; scan_win1119 <= 32'd0; scan_win1120 <= 32'd0; scan_win1121 <= 32'd0; scan_win1122 <= 32'd0; scan_win1123 <= 32'd0; scan_win1124 <= 32'd0; scan_win1125 <= 32'd0; scan_win1126 <= 32'd0; scan_win1127 <= 32'd0; scan_win1128 <= 32'd0; scan_win1129 <= 32'd0; scan_win1130 <= 32'd0; scan_win1131 <= 32'd0; scan_win1132 <= 32'd0; scan_win1133 <= 32'd0; scan_win1134 <= 32'd0; scan_win1135 <= 32'd0; scan_win1136 <= 32'd0; scan_win1137 <= 32'd0; scan_win1138 <= 32'd0; scan_win1139 <= 32'd0; scan_win1140 <= 32'd0; scan_win1141 <= 32'd0; scan_win1142 <= 32'd0; scan_win1143 <= 32'd0; scan_win1144 <= 32'd0; scan_win1145 <= 32'd0; scan_win1146 <= 32'd0; scan_win1147 <= 32'd0; scan_win1148 <= 32'd0; scan_win1149 <= 32'd0; scan_win1150 <= 32'd0; scan_win1151 <= 32'd0; scan_win1152 <= 32'd0; scan_win1153 <= 32'd0; scan_win1154 <= 32'd0; scan_win1155 <= 32'd0; scan_win1156 <= 32'd0; scan_win1157 <= 32'd0; scan_win1158 <= 32'd0; scan_win1159 <= 32'd0; scan_win1160 <= 32'd0; scan_win1161 <= 32'd0; scan_win1162 <= 32'd0; scan_win1163 <= 32'd0; scan_win1164 <= 32'd0; scan_win1165 <= 32'd0; scan_win1166 <= 32'd0; scan_win1167 <= 32'd0; scan_win1168 <= 32'd0; scan_win1169 <= 32'd0; scan_win1170 <= 32'd0; scan_win1171 <= 32'd0; scan_win1172 <= 32'd0; scan_win1173 <= 32'd0; scan_win1174 <= 32'd0; scan_win1175 <= 32'd0; scan_win1176 <= 32'd0; scan_win1177 <= 32'd0; scan_win1178 <= 32'd0; scan_win1179 <= 32'd0; scan_win1180 <= 32'd0; scan_win1181 <= 32'd0; scan_win1182 <= 32'd0; scan_win1183 <= 32'd0; scan_win1184 <= 32'd0; scan_win1185 <= 32'd0; scan_win1186 <= 32'd0; scan_win1187 <= 32'd0; scan_win1188 <= 32'd0; scan_win1189 <= 32'd0; scan_win1190 <= 32'd0; scan_win1191 <= 32'd0; scan_win1192 <= 32'd0; scan_win1193 <= 32'd0; scan_win1194 <= 32'd0; scan_win1195 <= 32'd0; scan_win1196 <= 32'd0; scan_win1197 <= 32'd0; scan_win1198 <= 32'd0; scan_win1199 <= 32'd0; scan_win1200 <= 32'd0; 
      scan_win1201 <= 32'd0; scan_win1202 <= 32'd0; scan_win1203 <= 32'd0; scan_win1204 <= 32'd0; scan_win1205 <= 32'd0; scan_win1206 <= 32'd0; scan_win1207 <= 32'd0; scan_win1208 <= 32'd0; scan_win1209 <= 32'd0; scan_win1210 <= 32'd0; scan_win1211 <= 32'd0; scan_win1212 <= 32'd0; scan_win1213 <= 32'd0; scan_win1214 <= 32'd0; scan_win1215 <= 32'd0; scan_win1216 <= 32'd0; scan_win1217 <= 32'd0; scan_win1218 <= 32'd0; scan_win1219 <= 32'd0; scan_win1220 <= 32'd0; scan_win1221 <= 32'd0; scan_win1222 <= 32'd0; scan_win1223 <= 32'd0; scan_win1224 <= 32'd0; scan_win1225 <= 32'd0; scan_win1226 <= 32'd0; scan_win1227 <= 32'd0; scan_win1228 <= 32'd0; scan_win1229 <= 32'd0; scan_win1230 <= 32'd0; scan_win1231 <= 32'd0; scan_win1232 <= 32'd0; scan_win1233 <= 32'd0; scan_win1234 <= 32'd0; scan_win1235 <= 32'd0; scan_win1236 <= 32'd0; scan_win1237 <= 32'd0; scan_win1238 <= 32'd0; scan_win1239 <= 32'd0; scan_win1240 <= 32'd0; scan_win1241 <= 32'd0; scan_win1242 <= 32'd0; scan_win1243 <= 32'd0; scan_win1244 <= 32'd0; scan_win1245 <= 32'd0; scan_win1246 <= 32'd0; scan_win1247 <= 32'd0; scan_win1248 <= 32'd0; scan_win1249 <= 32'd0; scan_win1250 <= 32'd0; scan_win1251 <= 32'd0; scan_win1252 <= 32'd0; scan_win1253 <= 32'd0; scan_win1254 <= 32'd0; scan_win1255 <= 32'd0; scan_win1256 <= 32'd0; scan_win1257 <= 32'd0; scan_win1258 <= 32'd0; scan_win1259 <= 32'd0; scan_win1260 <= 32'd0; scan_win1261 <= 32'd0; scan_win1262 <= 32'd0; scan_win1263 <= 32'd0; scan_win1264 <= 32'd0; scan_win1265 <= 32'd0; scan_win1266 <= 32'd0; scan_win1267 <= 32'd0; scan_win1268 <= 32'd0; scan_win1269 <= 32'd0; scan_win1270 <= 32'd0; scan_win1271 <= 32'd0; scan_win1272 <= 32'd0; scan_win1273 <= 32'd0; scan_win1274 <= 32'd0; scan_win1275 <= 32'd0; scan_win1276 <= 32'd0; scan_win1277 <= 32'd0; scan_win1278 <= 32'd0; scan_win1279 <= 32'd0; scan_win1280 <= 32'd0; scan_win1281 <= 32'd0; scan_win1282 <= 32'd0; scan_win1283 <= 32'd0; scan_win1284 <= 32'd0; scan_win1285 <= 32'd0; scan_win1286 <= 32'd0; scan_win1287 <= 32'd0; scan_win1288 <= 32'd0; scan_win1289 <= 32'd0; scan_win1290 <= 32'd0; scan_win1291 <= 32'd0; scan_win1292 <= 32'd0; scan_win1293 <= 32'd0; scan_win1294 <= 32'd0; scan_win1295 <= 32'd0; scan_win1296 <= 32'd0; scan_win1297 <= 32'd0; scan_win1298 <= 32'd0; scan_win1299 <= 32'd0; scan_win1300 <= 32'd0; scan_win1301 <= 32'd0; scan_win1302 <= 32'd0; scan_win1303 <= 32'd0; scan_win1304 <= 32'd0; scan_win1305 <= 32'd0; scan_win1306 <= 32'd0; scan_win1307 <= 32'd0; scan_win1308 <= 32'd0; scan_win1309 <= 32'd0; scan_win1310 <= 32'd0; scan_win1311 <= 32'd0; scan_win1312 <= 32'd0; scan_win1313 <= 32'd0; scan_win1314 <= 32'd0; scan_win1315 <= 32'd0; scan_win1316 <= 32'd0; scan_win1317 <= 32'd0; scan_win1318 <= 32'd0; scan_win1319 <= 32'd0; scan_win1320 <= 32'd0; scan_win1321 <= 32'd0; scan_win1322 <= 32'd0; scan_win1323 <= 32'd0; scan_win1324 <= 32'd0; scan_win1325 <= 32'd0; scan_win1326 <= 32'd0; scan_win1327 <= 32'd0; scan_win1328 <= 32'd0; scan_win1329 <= 32'd0; scan_win1330 <= 32'd0; scan_win1331 <= 32'd0; scan_win1332 <= 32'd0; scan_win1333 <= 32'd0; scan_win1334 <= 32'd0; scan_win1335 <= 32'd0; scan_win1336 <= 32'd0; scan_win1337 <= 32'd0; scan_win1338 <= 32'd0; scan_win1339 <= 32'd0; scan_win1340 <= 32'd0; scan_win1341 <= 32'd0; scan_win1342 <= 32'd0; scan_win1343 <= 32'd0; scan_win1344 <= 32'd0; scan_win1345 <= 32'd0; scan_win1346 <= 32'd0; scan_win1347 <= 32'd0; scan_win1348 <= 32'd0; scan_win1349 <= 32'd0; scan_win1350 <= 32'd0; scan_win1351 <= 32'd0; scan_win1352 <= 32'd0; scan_win1353 <= 32'd0; scan_win1354 <= 32'd0; scan_win1355 <= 32'd0; scan_win1356 <= 32'd0; scan_win1357 <= 32'd0; scan_win1358 <= 32'd0; scan_win1359 <= 32'd0; scan_win1360 <= 32'd0; scan_win1361 <= 32'd0; scan_win1362 <= 32'd0; scan_win1363 <= 32'd0; scan_win1364 <= 32'd0; scan_win1365 <= 32'd0; scan_win1366 <= 32'd0; scan_win1367 <= 32'd0; scan_win1368 <= 32'd0; scan_win1369 <= 32'd0; scan_win1370 <= 32'd0; scan_win1371 <= 32'd0; scan_win1372 <= 32'd0; scan_win1373 <= 32'd0; scan_win1374 <= 32'd0; scan_win1375 <= 32'd0; scan_win1376 <= 32'd0; scan_win1377 <= 32'd0; scan_win1378 <= 32'd0; scan_win1379 <= 32'd0; scan_win1380 <= 32'd0; scan_win1381 <= 32'd0; scan_win1382 <= 32'd0; scan_win1383 <= 32'd0; scan_win1384 <= 32'd0; scan_win1385 <= 32'd0; scan_win1386 <= 32'd0; scan_win1387 <= 32'd0; scan_win1388 <= 32'd0; scan_win1389 <= 32'd0; scan_win1390 <= 32'd0; scan_win1391 <= 32'd0; scan_win1392 <= 32'd0; scan_win1393 <= 32'd0; scan_win1394 <= 32'd0; scan_win1395 <= 32'd0; scan_win1396 <= 32'd0; scan_win1397 <= 32'd0; scan_win1398 <= 32'd0; scan_win1399 <= 32'd0; scan_win1400 <= 32'd0; 
      scan_win1401 <= 32'd0; scan_win1402 <= 32'd0; scan_win1403 <= 32'd0; scan_win1404 <= 32'd0; scan_win1405 <= 32'd0; scan_win1406 <= 32'd0; scan_win1407 <= 32'd0; scan_win1408 <= 32'd0; scan_win1409 <= 32'd0; scan_win1410 <= 32'd0; scan_win1411 <= 32'd0; scan_win1412 <= 32'd0; scan_win1413 <= 32'd0; scan_win1414 <= 32'd0; scan_win1415 <= 32'd0; scan_win1416 <= 32'd0; scan_win1417 <= 32'd0; scan_win1418 <= 32'd0; scan_win1419 <= 32'd0; scan_win1420 <= 32'd0; scan_win1421 <= 32'd0; scan_win1422 <= 32'd0; scan_win1423 <= 32'd0; scan_win1424 <= 32'd0; scan_win1425 <= 32'd0; scan_win1426 <= 32'd0; scan_win1427 <= 32'd0; scan_win1428 <= 32'd0; scan_win1429 <= 32'd0; scan_win1430 <= 32'd0; scan_win1431 <= 32'd0; scan_win1432 <= 32'd0; scan_win1433 <= 32'd0; scan_win1434 <= 32'd0; scan_win1435 <= 32'd0; scan_win1436 <= 32'd0; scan_win1437 <= 32'd0; scan_win1438 <= 32'd0; scan_win1439 <= 32'd0; scan_win1440 <= 32'd0; scan_win1441 <= 32'd0; scan_win1442 <= 32'd0; scan_win1443 <= 32'd0; scan_win1444 <= 32'd0; scan_win1445 <= 32'd0; scan_win1446 <= 32'd0; scan_win1447 <= 32'd0; scan_win1448 <= 32'd0; scan_win1449 <= 32'd0; scan_win1450 <= 32'd0; scan_win1451 <= 32'd0; scan_win1452 <= 32'd0; scan_win1453 <= 32'd0; scan_win1454 <= 32'd0; scan_win1455 <= 32'd0; scan_win1456 <= 32'd0; scan_win1457 <= 32'd0; scan_win1458 <= 32'd0; scan_win1459 <= 32'd0; scan_win1460 <= 32'd0; scan_win1461 <= 32'd0; scan_win1462 <= 32'd0; scan_win1463 <= 32'd0; scan_win1464 <= 32'd0; scan_win1465 <= 32'd0; scan_win1466 <= 32'd0; scan_win1467 <= 32'd0; scan_win1468 <= 32'd0; scan_win1469 <= 32'd0; scan_win1470 <= 32'd0; scan_win1471 <= 32'd0; scan_win1472 <= 32'd0; scan_win1473 <= 32'd0; scan_win1474 <= 32'd0; scan_win1475 <= 32'd0; scan_win1476 <= 32'd0; scan_win1477 <= 32'd0; scan_win1478 <= 32'd0; scan_win1479 <= 32'd0; scan_win1480 <= 32'd0; scan_win1481 <= 32'd0; scan_win1482 <= 32'd0; scan_win1483 <= 32'd0; scan_win1484 <= 32'd0; scan_win1485 <= 32'd0; scan_win1486 <= 32'd0; scan_win1487 <= 32'd0; scan_win1488 <= 32'd0; scan_win1489 <= 32'd0; scan_win1490 <= 32'd0; scan_win1491 <= 32'd0; scan_win1492 <= 32'd0; scan_win1493 <= 32'd0; scan_win1494 <= 32'd0; scan_win1495 <= 32'd0; scan_win1496 <= 32'd0; scan_win1497 <= 32'd0; scan_win1498 <= 32'd0; scan_win1499 <= 32'd0; scan_win1500 <= 32'd0; scan_win1501 <= 32'd0; scan_win1502 <= 32'd0; scan_win1503 <= 32'd0; scan_win1504 <= 32'd0; scan_win1505 <= 32'd0; scan_win1506 <= 32'd0; scan_win1507 <= 32'd0; scan_win1508 <= 32'd0; scan_win1509 <= 32'd0; scan_win1510 <= 32'd0; scan_win1511 <= 32'd0; scan_win1512 <= 32'd0; scan_win1513 <= 32'd0; scan_win1514 <= 32'd0; scan_win1515 <= 32'd0; scan_win1516 <= 32'd0; scan_win1517 <= 32'd0; scan_win1518 <= 32'd0; scan_win1519 <= 32'd0; scan_win1520 <= 32'd0; scan_win1521 <= 32'd0; scan_win1522 <= 32'd0; scan_win1523 <= 32'd0; scan_win1524 <= 32'd0; scan_win1525 <= 32'd0; scan_win1526 <= 32'd0; scan_win1527 <= 32'd0; scan_win1528 <= 32'd0; scan_win1529 <= 32'd0; scan_win1530 <= 32'd0; scan_win1531 <= 32'd0; scan_win1532 <= 32'd0; scan_win1533 <= 32'd0; scan_win1534 <= 32'd0; scan_win1535 <= 32'd0; scan_win1536 <= 32'd0; scan_win1537 <= 32'd0; scan_win1538 <= 32'd0; scan_win1539 <= 32'd0; scan_win1540 <= 32'd0; scan_win1541 <= 32'd0; scan_win1542 <= 32'd0; scan_win1543 <= 32'd0; scan_win1544 <= 32'd0; scan_win1545 <= 32'd0; scan_win1546 <= 32'd0; scan_win1547 <= 32'd0; scan_win1548 <= 32'd0; scan_win1549 <= 32'd0; scan_win1550 <= 32'd0; scan_win1551 <= 32'd0; scan_win1552 <= 32'd0; scan_win1553 <= 32'd0; scan_win1554 <= 32'd0; scan_win1555 <= 32'd0; scan_win1556 <= 32'd0; scan_win1557 <= 32'd0; scan_win1558 <= 32'd0; scan_win1559 <= 32'd0; scan_win1560 <= 32'd0; scan_win1561 <= 32'd0; scan_win1562 <= 32'd0; scan_win1563 <= 32'd0; scan_win1564 <= 32'd0; scan_win1565 <= 32'd0; scan_win1566 <= 32'd0; scan_win1567 <= 32'd0; scan_win1568 <= 32'd0; scan_win1569 <= 32'd0; scan_win1570 <= 32'd0; scan_win1571 <= 32'd0; scan_win1572 <= 32'd0; scan_win1573 <= 32'd0; scan_win1574 <= 32'd0; scan_win1575 <= 32'd0; scan_win1576 <= 32'd0; scan_win1577 <= 32'd0; scan_win1578 <= 32'd0; scan_win1579 <= 32'd0; scan_win1580 <= 32'd0; scan_win1581 <= 32'd0; scan_win1582 <= 32'd0; scan_win1583 <= 32'd0; scan_win1584 <= 32'd0; scan_win1585 <= 32'd0; scan_win1586 <= 32'd0; scan_win1587 <= 32'd0; scan_win1588 <= 32'd0; scan_win1589 <= 32'd0; scan_win1590 <= 32'd0; scan_win1591 <= 32'd0; scan_win1592 <= 32'd0; scan_win1593 <= 32'd0; scan_win1594 <= 32'd0; scan_win1595 <= 32'd0; scan_win1596 <= 32'd0; scan_win1597 <= 32'd0; scan_win1598 <= 32'd0; scan_win1599 <= 32'd0; scan_win1600 <= 32'd0; 
      scan_win1601 <= 32'd0; scan_win1602 <= 32'd0; scan_win1603 <= 32'd0; scan_win1604 <= 32'd0; scan_win1605 <= 32'd0; scan_win1606 <= 32'd0; scan_win1607 <= 32'd0; scan_win1608 <= 32'd0; scan_win1609 <= 32'd0; scan_win1610 <= 32'd0; scan_win1611 <= 32'd0; scan_win1612 <= 32'd0; scan_win1613 <= 32'd0; scan_win1614 <= 32'd0; scan_win1615 <= 32'd0; scan_win1616 <= 32'd0; scan_win1617 <= 32'd0; scan_win1618 <= 32'd0; scan_win1619 <= 32'd0; scan_win1620 <= 32'd0; scan_win1621 <= 32'd0; scan_win1622 <= 32'd0; scan_win1623 <= 32'd0; scan_win1624 <= 32'd0; scan_win1625 <= 32'd0; scan_win1626 <= 32'd0; scan_win1627 <= 32'd0; scan_win1628 <= 32'd0; scan_win1629 <= 32'd0; scan_win1630 <= 32'd0; scan_win1631 <= 32'd0; scan_win1632 <= 32'd0; scan_win1633 <= 32'd0; scan_win1634 <= 32'd0; scan_win1635 <= 32'd0; scan_win1636 <= 32'd0; scan_win1637 <= 32'd0; scan_win1638 <= 32'd0; scan_win1639 <= 32'd0; scan_win1640 <= 32'd0; scan_win1641 <= 32'd0; scan_win1642 <= 32'd0; scan_win1643 <= 32'd0; scan_win1644 <= 32'd0; scan_win1645 <= 32'd0; scan_win1646 <= 32'd0; scan_win1647 <= 32'd0; scan_win1648 <= 32'd0; scan_win1649 <= 32'd0; scan_win1650 <= 32'd0; scan_win1651 <= 32'd0; scan_win1652 <= 32'd0; scan_win1653 <= 32'd0; scan_win1654 <= 32'd0; scan_win1655 <= 32'd0; scan_win1656 <= 32'd0; scan_win1657 <= 32'd0; scan_win1658 <= 32'd0; scan_win1659 <= 32'd0; scan_win1660 <= 32'd0; scan_win1661 <= 32'd0; scan_win1662 <= 32'd0; scan_win1663 <= 32'd0; scan_win1664 <= 32'd0; scan_win1665 <= 32'd0; scan_win1666 <= 32'd0; scan_win1667 <= 32'd0; scan_win1668 <= 32'd0; scan_win1669 <= 32'd0; scan_win1670 <= 32'd0; scan_win1671 <= 32'd0; scan_win1672 <= 32'd0; scan_win1673 <= 32'd0; scan_win1674 <= 32'd0; scan_win1675 <= 32'd0; scan_win1676 <= 32'd0; scan_win1677 <= 32'd0; scan_win1678 <= 32'd0; scan_win1679 <= 32'd0; scan_win1680 <= 32'd0; scan_win1681 <= 32'd0; scan_win1682 <= 32'd0; scan_win1683 <= 32'd0; scan_win1684 <= 32'd0; scan_win1685 <= 32'd0; scan_win1686 <= 32'd0; scan_win1687 <= 32'd0; scan_win1688 <= 32'd0; scan_win1689 <= 32'd0; scan_win1690 <= 32'd0; scan_win1691 <= 32'd0; scan_win1692 <= 32'd0; scan_win1693 <= 32'd0; scan_win1694 <= 32'd0; scan_win1695 <= 32'd0; scan_win1696 <= 32'd0; scan_win1697 <= 32'd0; scan_win1698 <= 32'd0; scan_win1699 <= 32'd0; scan_win1700 <= 32'd0; scan_win1701 <= 32'd0; scan_win1702 <= 32'd0; scan_win1703 <= 32'd0; scan_win1704 <= 32'd0; scan_win1705 <= 32'd0; scan_win1706 <= 32'd0; scan_win1707 <= 32'd0; scan_win1708 <= 32'd0; scan_win1709 <= 32'd0; scan_win1710 <= 32'd0; scan_win1711 <= 32'd0; scan_win1712 <= 32'd0; scan_win1713 <= 32'd0; scan_win1714 <= 32'd0; scan_win1715 <= 32'd0; scan_win1716 <= 32'd0; scan_win1717 <= 32'd0; scan_win1718 <= 32'd0; scan_win1719 <= 32'd0; scan_win1720 <= 32'd0; scan_win1721 <= 32'd0; scan_win1722 <= 32'd0; scan_win1723 <= 32'd0; scan_win1724 <= 32'd0; scan_win1725 <= 32'd0; scan_win1726 <= 32'd0; scan_win1727 <= 32'd0; scan_win1728 <= 32'd0; scan_win1729 <= 32'd0; scan_win1730 <= 32'd0; scan_win1731 <= 32'd0; scan_win1732 <= 32'd0; scan_win1733 <= 32'd0; scan_win1734 <= 32'd0; scan_win1735 <= 32'd0; scan_win1736 <= 32'd0; scan_win1737 <= 32'd0; scan_win1738 <= 32'd0; scan_win1739 <= 32'd0; scan_win1740 <= 32'd0; scan_win1741 <= 32'd0; scan_win1742 <= 32'd0; scan_win1743 <= 32'd0; scan_win1744 <= 32'd0; scan_win1745 <= 32'd0; scan_win1746 <= 32'd0; scan_win1747 <= 32'd0; scan_win1748 <= 32'd0; scan_win1749 <= 32'd0; scan_win1750 <= 32'd0; scan_win1751 <= 32'd0; scan_win1752 <= 32'd0; scan_win1753 <= 32'd0; scan_win1754 <= 32'd0; scan_win1755 <= 32'd0; scan_win1756 <= 32'd0; scan_win1757 <= 32'd0; scan_win1758 <= 32'd0; scan_win1759 <= 32'd0; scan_win1760 <= 32'd0; scan_win1761 <= 32'd0; scan_win1762 <= 32'd0; scan_win1763 <= 32'd0; scan_win1764 <= 32'd0; scan_win1765 <= 32'd0; scan_win1766 <= 32'd0; scan_win1767 <= 32'd0; scan_win1768 <= 32'd0; scan_win1769 <= 32'd0; scan_win1770 <= 32'd0; scan_win1771 <= 32'd0; scan_win1772 <= 32'd0; scan_win1773 <= 32'd0; scan_win1774 <= 32'd0; scan_win1775 <= 32'd0; scan_win1776 <= 32'd0; scan_win1777 <= 32'd0; scan_win1778 <= 32'd0; scan_win1779 <= 32'd0; scan_win1780 <= 32'd0; scan_win1781 <= 32'd0; scan_win1782 <= 32'd0; scan_win1783 <= 32'd0; scan_win1784 <= 32'd0; scan_win1785 <= 32'd0; scan_win1786 <= 32'd0; scan_win1787 <= 32'd0; scan_win1788 <= 32'd0; scan_win1789 <= 32'd0; scan_win1790 <= 32'd0; scan_win1791 <= 32'd0; scan_win1792 <= 32'd0; scan_win1793 <= 32'd0; scan_win1794 <= 32'd0; scan_win1795 <= 32'd0; scan_win1796 <= 32'd0; scan_win1797 <= 32'd0; scan_win1798 <= 32'd0; scan_win1799 <= 32'd0; scan_win1800 <= 32'd0; 
      scan_win1801 <= 32'd0; scan_win1802 <= 32'd0; scan_win1803 <= 32'd0; scan_win1804 <= 32'd0; scan_win1805 <= 32'd0; scan_win1806 <= 32'd0; scan_win1807 <= 32'd0; scan_win1808 <= 32'd0; scan_win1809 <= 32'd0; scan_win1810 <= 32'd0; scan_win1811 <= 32'd0; scan_win1812 <= 32'd0; scan_win1813 <= 32'd0; scan_win1814 <= 32'd0; scan_win1815 <= 32'd0; scan_win1816 <= 32'd0; scan_win1817 <= 32'd0; scan_win1818 <= 32'd0; scan_win1819 <= 32'd0; scan_win1820 <= 32'd0; scan_win1821 <= 32'd0; scan_win1822 <= 32'd0; scan_win1823 <= 32'd0; scan_win1824 <= 32'd0; scan_win1825 <= 32'd0; scan_win1826 <= 32'd0; scan_win1827 <= 32'd0; scan_win1828 <= 32'd0; scan_win1829 <= 32'd0; scan_win1830 <= 32'd0; scan_win1831 <= 32'd0; scan_win1832 <= 32'd0; scan_win1833 <= 32'd0; scan_win1834 <= 32'd0; scan_win1835 <= 32'd0; scan_win1836 <= 32'd0; scan_win1837 <= 32'd0; scan_win1838 <= 32'd0; scan_win1839 <= 32'd0; scan_win1840 <= 32'd0; scan_win1841 <= 32'd0; scan_win1842 <= 32'd0; scan_win1843 <= 32'd0; scan_win1844 <= 32'd0; scan_win1845 <= 32'd0; scan_win1846 <= 32'd0; scan_win1847 <= 32'd0; scan_win1848 <= 32'd0; scan_win1849 <= 32'd0; scan_win1850 <= 32'd0; scan_win1851 <= 32'd0; scan_win1852 <= 32'd0; scan_win1853 <= 32'd0; scan_win1854 <= 32'd0; scan_win1855 <= 32'd0; scan_win1856 <= 32'd0; scan_win1857 <= 32'd0; scan_win1858 <= 32'd0; scan_win1859 <= 32'd0; scan_win1860 <= 32'd0; scan_win1861 <= 32'd0; scan_win1862 <= 32'd0; scan_win1863 <= 32'd0; scan_win1864 <= 32'd0; scan_win1865 <= 32'd0; scan_win1866 <= 32'd0; scan_win1867 <= 32'd0; scan_win1868 <= 32'd0; scan_win1869 <= 32'd0; scan_win1870 <= 32'd0; scan_win1871 <= 32'd0; scan_win1872 <= 32'd0; scan_win1873 <= 32'd0; scan_win1874 <= 32'd0; scan_win1875 <= 32'd0; scan_win1876 <= 32'd0; scan_win1877 <= 32'd0; scan_win1878 <= 32'd0; scan_win1879 <= 32'd0; scan_win1880 <= 32'd0; scan_win1881 <= 32'd0; scan_win1882 <= 32'd0; scan_win1883 <= 32'd0; scan_win1884 <= 32'd0; scan_win1885 <= 32'd0; scan_win1886 <= 32'd0; scan_win1887 <= 32'd0; scan_win1888 <= 32'd0; scan_win1889 <= 32'd0; scan_win1890 <= 32'd0; scan_win1891 <= 32'd0; scan_win1892 <= 32'd0; scan_win1893 <= 32'd0; scan_win1894 <= 32'd0; scan_win1895 <= 32'd0; scan_win1896 <= 32'd0; scan_win1897 <= 32'd0; scan_win1898 <= 32'd0; scan_win1899 <= 32'd0; scan_win1900 <= 32'd0; scan_win1901 <= 32'd0; scan_win1902 <= 32'd0; scan_win1903 <= 32'd0; scan_win1904 <= 32'd0; scan_win1905 <= 32'd0; scan_win1906 <= 32'd0; scan_win1907 <= 32'd0; scan_win1908 <= 32'd0; scan_win1909 <= 32'd0; scan_win1910 <= 32'd0; scan_win1911 <= 32'd0; scan_win1912 <= 32'd0; scan_win1913 <= 32'd0; scan_win1914 <= 32'd0; scan_win1915 <= 32'd0; scan_win1916 <= 32'd0; scan_win1917 <= 32'd0; scan_win1918 <= 32'd0; scan_win1919 <= 32'd0; scan_win1920 <= 32'd0; scan_win1921 <= 32'd0; scan_win1922 <= 32'd0; scan_win1923 <= 32'd0; scan_win1924 <= 32'd0; scan_win1925 <= 32'd0; scan_win1926 <= 32'd0; scan_win1927 <= 32'd0; scan_win1928 <= 32'd0; scan_win1929 <= 32'd0; scan_win1930 <= 32'd0; scan_win1931 <= 32'd0; scan_win1932 <= 32'd0; scan_win1933 <= 32'd0; scan_win1934 <= 32'd0; scan_win1935 <= 32'd0; scan_win1936 <= 32'd0; scan_win1937 <= 32'd0; scan_win1938 <= 32'd0; scan_win1939 <= 32'd0; scan_win1940 <= 32'd0; scan_win1941 <= 32'd0; scan_win1942 <= 32'd0; scan_win1943 <= 32'd0; scan_win1944 <= 32'd0; scan_win1945 <= 32'd0; scan_win1946 <= 32'd0; scan_win1947 <= 32'd0; scan_win1948 <= 32'd0; scan_win1949 <= 32'd0; scan_win1950 <= 32'd0; scan_win1951 <= 32'd0; scan_win1952 <= 32'd0; scan_win1953 <= 32'd0; scan_win1954 <= 32'd0; scan_win1955 <= 32'd0; scan_win1956 <= 32'd0; scan_win1957 <= 32'd0; scan_win1958 <= 32'd0; scan_win1959 <= 32'd0; scan_win1960 <= 32'd0; scan_win1961 <= 32'd0; scan_win1962 <= 32'd0; scan_win1963 <= 32'd0; scan_win1964 <= 32'd0; scan_win1965 <= 32'd0; scan_win1966 <= 32'd0; scan_win1967 <= 32'd0; scan_win1968 <= 32'd0; scan_win1969 <= 32'd0; scan_win1970 <= 32'd0; scan_win1971 <= 32'd0; scan_win1972 <= 32'd0; scan_win1973 <= 32'd0; scan_win1974 <= 32'd0; scan_win1975 <= 32'd0; scan_win1976 <= 32'd0; scan_win1977 <= 32'd0; scan_win1978 <= 32'd0; scan_win1979 <= 32'd0; scan_win1980 <= 32'd0; scan_win1981 <= 32'd0; scan_win1982 <= 32'd0; scan_win1983 <= 32'd0; scan_win1984 <= 32'd0; scan_win1985 <= 32'd0; scan_win1986 <= 32'd0; scan_win1987 <= 32'd0; scan_win1988 <= 32'd0; scan_win1989 <= 32'd0; scan_win1990 <= 32'd0; scan_win1991 <= 32'd0; scan_win1992 <= 32'd0; scan_win1993 <= 32'd0; scan_win1994 <= 32'd0; scan_win1995 <= 32'd0; scan_win1996 <= 32'd0; scan_win1997 <= 32'd0; scan_win1998 <= 32'd0; scan_win1999 <= 32'd0; scan_win2000 <= 32'd0; 
      scan_win2001 <= 32'd0; scan_win2002 <= 32'd0; scan_win2003 <= 32'd0; scan_win2004 <= 32'd0; scan_win2005 <= 32'd0; scan_win2006 <= 32'd0; scan_win2007 <= 32'd0; scan_win2008 <= 32'd0; scan_win2009 <= 32'd0; scan_win2010 <= 32'd0; scan_win2011 <= 32'd0; scan_win2012 <= 32'd0; scan_win2013 <= 32'd0; scan_win2014 <= 32'd0; scan_win2015 <= 32'd0; scan_win2016 <= 32'd0; scan_win2017 <= 32'd0; scan_win2018 <= 32'd0; scan_win2019 <= 32'd0; scan_win2020 <= 32'd0; scan_win2021 <= 32'd0; scan_win2022 <= 32'd0; scan_win2023 <= 32'd0; scan_win2024 <= 32'd0; scan_win2025 <= 32'd0; scan_win2026 <= 32'd0; scan_win2027 <= 32'd0; scan_win2028 <= 32'd0; scan_win2029 <= 32'd0; scan_win2030 <= 32'd0; scan_win2031 <= 32'd0; scan_win2032 <= 32'd0; scan_win2033 <= 32'd0; scan_win2034 <= 32'd0; scan_win2035 <= 32'd0; scan_win2036 <= 32'd0; scan_win2037 <= 32'd0; scan_win2038 <= 32'd0; scan_win2039 <= 32'd0; scan_win2040 <= 32'd0; scan_win2041 <= 32'd0; scan_win2042 <= 32'd0; scan_win2043 <= 32'd0; scan_win2044 <= 32'd0; scan_win2045 <= 32'd0; scan_win2046 <= 32'd0; scan_win2047 <= 32'd0; scan_win2048 <= 32'd0; scan_win2049 <= 32'd0; scan_win2050 <= 32'd0; scan_win2051 <= 32'd0; scan_win2052 <= 32'd0; scan_win2053 <= 32'd0; scan_win2054 <= 32'd0; scan_win2055 <= 32'd0; scan_win2056 <= 32'd0; scan_win2057 <= 32'd0; scan_win2058 <= 32'd0; scan_win2059 <= 32'd0; scan_win2060 <= 32'd0; scan_win2061 <= 32'd0; scan_win2062 <= 32'd0; scan_win2063 <= 32'd0; scan_win2064 <= 32'd0; scan_win2065 <= 32'd0; scan_win2066 <= 32'd0; scan_win2067 <= 32'd0; scan_win2068 <= 32'd0; scan_win2069 <= 32'd0; scan_win2070 <= 32'd0; scan_win2071 <= 32'd0; scan_win2072 <= 32'd0; scan_win2073 <= 32'd0; scan_win2074 <= 32'd0; scan_win2075 <= 32'd0; scan_win2076 <= 32'd0; scan_win2077 <= 32'd0; scan_win2078 <= 32'd0; scan_win2079 <= 32'd0; scan_win2080 <= 32'd0; scan_win2081 <= 32'd0; scan_win2082 <= 32'd0; scan_win2083 <= 32'd0; scan_win2084 <= 32'd0; scan_win2085 <= 32'd0; scan_win2086 <= 32'd0; scan_win2087 <= 32'd0; scan_win2088 <= 32'd0; scan_win2089 <= 32'd0; scan_win2090 <= 32'd0; scan_win2091 <= 32'd0; scan_win2092 <= 32'd0; scan_win2093 <= 32'd0; scan_win2094 <= 32'd0; scan_win2095 <= 32'd0; scan_win2096 <= 32'd0; scan_win2097 <= 32'd0; scan_win2098 <= 32'd0; scan_win2099 <= 32'd0; scan_win2100 <= 32'd0; scan_win2101 <= 32'd0; scan_win2102 <= 32'd0; scan_win2103 <= 32'd0; scan_win2104 <= 32'd0; scan_win2105 <= 32'd0; scan_win2106 <= 32'd0; scan_win2107 <= 32'd0; scan_win2108 <= 32'd0; scan_win2109 <= 32'd0; scan_win2110 <= 32'd0; scan_win2111 <= 32'd0; scan_win2112 <= 32'd0; scan_win2113 <= 32'd0; scan_win2114 <= 32'd0; scan_win2115 <= 32'd0; scan_win2116 <= 32'd0; scan_win2117 <= 32'd0; scan_win2118 <= 32'd0; scan_win2119 <= 32'd0; scan_win2120 <= 32'd0; scan_win2121 <= 32'd0; scan_win2122 <= 32'd0; scan_win2123 <= 32'd0; scan_win2124 <= 32'd0; scan_win2125 <= 32'd0; scan_win2126 <= 32'd0; scan_win2127 <= 32'd0; scan_win2128 <= 32'd0; scan_win2129 <= 32'd0; scan_win2130 <= 32'd0; scan_win2131 <= 32'd0; scan_win2132 <= 32'd0; scan_win2133 <= 32'd0; scan_win2134 <= 32'd0; scan_win2135 <= 32'd0; scan_win2136 <= 32'd0; scan_win2137 <= 32'd0; scan_win2138 <= 32'd0; scan_win2139 <= 32'd0; scan_win2140 <= 32'd0; scan_win2141 <= 32'd0; scan_win2142 <= 32'd0; scan_win2143 <= 32'd0; scan_win2144 <= 32'd0; scan_win2145 <= 32'd0; scan_win2146 <= 32'd0; scan_win2147 <= 32'd0; scan_win2148 <= 32'd0; scan_win2149 <= 32'd0; scan_win2150 <= 32'd0; scan_win2151 <= 32'd0; scan_win2152 <= 32'd0; scan_win2153 <= 32'd0; scan_win2154 <= 32'd0; scan_win2155 <= 32'd0; scan_win2156 <= 32'd0; scan_win2157 <= 32'd0; scan_win2158 <= 32'd0; scan_win2159 <= 32'd0; scan_win2160 <= 32'd0; scan_win2161 <= 32'd0; scan_win2162 <= 32'd0; scan_win2163 <= 32'd0; scan_win2164 <= 32'd0; scan_win2165 <= 32'd0; scan_win2166 <= 32'd0; scan_win2167 <= 32'd0; scan_win2168 <= 32'd0; scan_win2169 <= 32'd0; scan_win2170 <= 32'd0; scan_win2171 <= 32'd0; scan_win2172 <= 32'd0; scan_win2173 <= 32'd0; scan_win2174 <= 32'd0; scan_win2175 <= 32'd0; scan_win2176 <= 32'd0; scan_win2177 <= 32'd0; scan_win2178 <= 32'd0; scan_win2179 <= 32'd0; scan_win2180 <= 32'd0; scan_win2181 <= 32'd0; scan_win2182 <= 32'd0; scan_win2183 <= 32'd0; scan_win2184 <= 32'd0; scan_win2185 <= 32'd0; scan_win2186 <= 32'd0; scan_win2187 <= 32'd0; scan_win2188 <= 32'd0; scan_win2189 <= 32'd0; scan_win2190 <= 32'd0; scan_win2191 <= 32'd0; scan_win2192 <= 32'd0; scan_win2193 <= 32'd0; scan_win2194 <= 32'd0; scan_win2195 <= 32'd0; scan_win2196 <= 32'd0; scan_win2197 <= 32'd0; scan_win2198 <= 32'd0; scan_win2199 <= 32'd0; scan_win2200 <= 32'd0; 
      scan_win2201 <= 32'd0; scan_win2202 <= 32'd0; scan_win2203 <= 32'd0; scan_win2204 <= 32'd0; scan_win2205 <= 32'd0; scan_win2206 <= 32'd0; scan_win2207 <= 32'd0; scan_win2208 <= 32'd0; scan_win2209 <= 32'd0; scan_win2210 <= 32'd0; scan_win2211 <= 32'd0; scan_win2212 <= 32'd0; scan_win2213 <= 32'd0; scan_win2214 <= 32'd0; scan_win2215 <= 32'd0; scan_win2216 <= 32'd0; scan_win2217 <= 32'd0; scan_win2218 <= 32'd0; scan_win2219 <= 32'd0; scan_win2220 <= 32'd0; scan_win2221 <= 32'd0; scan_win2222 <= 32'd0; scan_win2223 <= 32'd0; scan_win2224 <= 32'd0; scan_win2225 <= 32'd0; scan_win2226 <= 32'd0; scan_win2227 <= 32'd0; scan_win2228 <= 32'd0; scan_win2229 <= 32'd0; scan_win2230 <= 32'd0; scan_win2231 <= 32'd0; scan_win2232 <= 32'd0; scan_win2233 <= 32'd0; scan_win2234 <= 32'd0; scan_win2235 <= 32'd0; scan_win2236 <= 32'd0; scan_win2237 <= 32'd0; scan_win2238 <= 32'd0; scan_win2239 <= 32'd0; scan_win2240 <= 32'd0; scan_win2241 <= 32'd0; scan_win2242 <= 32'd0; scan_win2243 <= 32'd0; scan_win2244 <= 32'd0; scan_win2245 <= 32'd0; scan_win2246 <= 32'd0; scan_win2247 <= 32'd0; scan_win2248 <= 32'd0; scan_win2249 <= 32'd0; scan_win2250 <= 32'd0; scan_win2251 <= 32'd0; scan_win2252 <= 32'd0; scan_win2253 <= 32'd0; scan_win2254 <= 32'd0; scan_win2255 <= 32'd0; scan_win2256 <= 32'd0; scan_win2257 <= 32'd0; scan_win2258 <= 32'd0; scan_win2259 <= 32'd0; scan_win2260 <= 32'd0; scan_win2261 <= 32'd0; scan_win2262 <= 32'd0; scan_win2263 <= 32'd0; scan_win2264 <= 32'd0; scan_win2265 <= 32'd0; scan_win2266 <= 32'd0; scan_win2267 <= 32'd0; scan_win2268 <= 32'd0; scan_win2269 <= 32'd0; scan_win2270 <= 32'd0; scan_win2271 <= 32'd0; scan_win2272 <= 32'd0; scan_win2273 <= 32'd0; scan_win2274 <= 32'd0; scan_win2275 <= 32'd0; scan_win2276 <= 32'd0; scan_win2277 <= 32'd0; scan_win2278 <= 32'd0; scan_win2279 <= 32'd0; scan_win2280 <= 32'd0; scan_win2281 <= 32'd0; scan_win2282 <= 32'd0; scan_win2283 <= 32'd0; scan_win2284 <= 32'd0; scan_win2285 <= 32'd0; scan_win2286 <= 32'd0; scan_win2287 <= 32'd0; scan_win2288 <= 32'd0; scan_win2289 <= 32'd0; scan_win2290 <= 32'd0; scan_win2291 <= 32'd0; scan_win2292 <= 32'd0; scan_win2293 <= 32'd0; scan_win2294 <= 32'd0; scan_win2295 <= 32'd0; scan_win2296 <= 32'd0; scan_win2297 <= 32'd0; scan_win2298 <= 32'd0; scan_win2299 <= 32'd0; scan_win2300 <= 32'd0; scan_win2301 <= 32'd0; scan_win2302 <= 32'd0; scan_win2303 <= 32'd0; scan_win2304 <= 32'd0; scan_win2305 <= 32'd0; scan_win2306 <= 32'd0; scan_win2307 <= 32'd0; scan_win2308 <= 32'd0; scan_win2309 <= 32'd0; scan_win2310 <= 32'd0; scan_win2311 <= 32'd0; scan_win2312 <= 32'd0; scan_win2313 <= 32'd0; scan_win2314 <= 32'd0; scan_win2315 <= 32'd0; scan_win2316 <= 32'd0; scan_win2317 <= 32'd0; scan_win2318 <= 32'd0; scan_win2319 <= 32'd0; scan_win2320 <= 32'd0; scan_win2321 <= 32'd0; scan_win2322 <= 32'd0; scan_win2323 <= 32'd0; scan_win2324 <= 32'd0; scan_win2325 <= 32'd0; scan_win2326 <= 32'd0; scan_win2327 <= 32'd0; scan_win2328 <= 32'd0; scan_win2329 <= 32'd0; scan_win2330 <= 32'd0; scan_win2331 <= 32'd0; scan_win2332 <= 32'd0; scan_win2333 <= 32'd0; scan_win2334 <= 32'd0; scan_win2335 <= 32'd0; scan_win2336 <= 32'd0; scan_win2337 <= 32'd0; scan_win2338 <= 32'd0; scan_win2339 <= 32'd0; scan_win2340 <= 32'd0; scan_win2341 <= 32'd0; scan_win2342 <= 32'd0; scan_win2343 <= 32'd0; scan_win2344 <= 32'd0; scan_win2345 <= 32'd0; scan_win2346 <= 32'd0; scan_win2347 <= 32'd0; scan_win2348 <= 32'd0; scan_win2349 <= 32'd0; scan_win2350 <= 32'd0; scan_win2351 <= 32'd0; scan_win2352 <= 32'd0; scan_win2353 <= 32'd0; scan_win2354 <= 32'd0; scan_win2355 <= 32'd0; scan_win2356 <= 32'd0; scan_win2357 <= 32'd0; scan_win2358 <= 32'd0; scan_win2359 <= 32'd0; scan_win2360 <= 32'd0; scan_win2361 <= 32'd0; scan_win2362 <= 32'd0; scan_win2363 <= 32'd0; scan_win2364 <= 32'd0; scan_win2365 <= 32'd0; scan_win2366 <= 32'd0; scan_win2367 <= 32'd0; scan_win2368 <= 32'd0; scan_win2369 <= 32'd0; scan_win2370 <= 32'd0; scan_win2371 <= 32'd0; scan_win2372 <= 32'd0; scan_win2373 <= 32'd0; scan_win2374 <= 32'd0; scan_win2375 <= 32'd0; scan_win2376 <= 32'd0; scan_win2377 <= 32'd0; scan_win2378 <= 32'd0; scan_win2379 <= 32'd0; scan_win2380 <= 32'd0; scan_win2381 <= 32'd0; scan_win2382 <= 32'd0; scan_win2383 <= 32'd0; scan_win2384 <= 32'd0; scan_win2385 <= 32'd0; scan_win2386 <= 32'd0; scan_win2387 <= 32'd0; scan_win2388 <= 32'd0; scan_win2389 <= 32'd0; scan_win2390 <= 32'd0; scan_win2391 <= 32'd0; scan_win2392 <= 32'd0; scan_win2393 <= 32'd0; scan_win2394 <= 32'd0; scan_win2395 <= 32'd0; scan_win2396 <= 32'd0; scan_win2397 <= 32'd0; scan_win2398 <= 32'd0; scan_win2399 <= 32'd0; scan_win2400 <= 32'd0; 
      scan_win2401 <= 32'd0; scan_win2402 <= 32'd0; scan_win2403 <= 32'd0; scan_win2404 <= 32'd0; scan_win2405 <= 32'd0; scan_win2406 <= 32'd0; scan_win2407 <= 32'd0; scan_win2408 <= 32'd0; scan_win2409 <= 32'd0; scan_win2410 <= 32'd0; scan_win2411 <= 32'd0; scan_win2412 <= 32'd0; scan_win2413 <= 32'd0; scan_win2414 <= 32'd0; scan_win2415 <= 32'd0; scan_win2416 <= 32'd0; scan_win2417 <= 32'd0; scan_win2418 <= 32'd0; scan_win2419 <= 32'd0; scan_win2420 <= 32'd0; scan_win2421 <= 32'd0; scan_win2422 <= 32'd0; scan_win2423 <= 32'd0; scan_win2424 <= 32'd0; scan_win2425 <= 32'd0; scan_win2426 <= 32'd0; scan_win2427 <= 32'd0; scan_win2428 <= 32'd0; scan_win2429 <= 32'd0; scan_win2430 <= 32'd0; scan_win2431 <= 32'd0; scan_win2432 <= 32'd0; scan_win2433 <= 32'd0; scan_win2434 <= 32'd0; scan_win2435 <= 32'd0; scan_win2436 <= 32'd0; scan_win2437 <= 32'd0; scan_win2438 <= 32'd0; scan_win2439 <= 32'd0; scan_win2440 <= 32'd0; scan_win2441 <= 32'd0; scan_win2442 <= 32'd0; scan_win2443 <= 32'd0; scan_win2444 <= 32'd0; scan_win2445 <= 32'd0; scan_win2446 <= 32'd0; scan_win2447 <= 32'd0; scan_win2448 <= 32'd0; scan_win2449 <= 32'd0; scan_win2450 <= 32'd0; scan_win2451 <= 32'd0; scan_win2452 <= 32'd0; scan_win2453 <= 32'd0; scan_win2454 <= 32'd0; scan_win2455 <= 32'd0; scan_win2456 <= 32'd0; scan_win2457 <= 32'd0; scan_win2458 <= 32'd0; scan_win2459 <= 32'd0; scan_win2460 <= 32'd0; scan_win2461 <= 32'd0; scan_win2462 <= 32'd0; scan_win2463 <= 32'd0; scan_win2464 <= 32'd0; scan_win2465 <= 32'd0; scan_win2466 <= 32'd0; scan_win2467 <= 32'd0; scan_win2468 <= 32'd0; scan_win2469 <= 32'd0; scan_win2470 <= 32'd0; scan_win2471 <= 32'd0; scan_win2472 <= 32'd0; scan_win2473 <= 32'd0; scan_win2474 <= 32'd0; scan_win2475 <= 32'd0; scan_win2476 <= 32'd0; scan_win2477 <= 32'd0; scan_win2478 <= 32'd0; scan_win2479 <= 32'd0; scan_win2480 <= 32'd0; scan_win2481 <= 32'd0; scan_win2482 <= 32'd0; scan_win2483 <= 32'd0; scan_win2484 <= 32'd0; scan_win2485 <= 32'd0; scan_win2486 <= 32'd0; scan_win2487 <= 32'd0; scan_win2488 <= 32'd0; scan_win2489 <= 32'd0; scan_win2490 <= 32'd0; scan_win2491 <= 32'd0; scan_win2492 <= 32'd0; scan_win2493 <= 32'd0; scan_win2494 <= 32'd0; scan_win2495 <= 32'd0; scan_win2496 <= 32'd0; scan_win2497 <= 32'd0; scan_win2498 <= 32'd0; scan_win2499 <= 32'd0; scan_win2500 <= 32'd0; scan_win2501 <= 32'd0; scan_win2502 <= 32'd0; scan_win2503 <= 32'd0; scan_win2504 <= 32'd0; scan_win2505 <= 32'd0; scan_win2506 <= 32'd0; scan_win2507 <= 32'd0; scan_win2508 <= 32'd0; scan_win2509 <= 32'd0; scan_win2510 <= 32'd0; scan_win2511 <= 32'd0; scan_win2512 <= 32'd0; scan_win2513 <= 32'd0; scan_win2514 <= 32'd0; scan_win2515 <= 32'd0; scan_win2516 <= 32'd0; scan_win2517 <= 32'd0; scan_win2518 <= 32'd0; scan_win2519 <= 32'd0; scan_win2520 <= 32'd0; scan_win2521 <= 32'd0; scan_win2522 <= 32'd0; scan_win2523 <= 32'd0; scan_win2524 <= 32'd0; scan_win2525 <= 32'd0; scan_win2526 <= 32'd0; scan_win2527 <= 32'd0; scan_win2528 <= 32'd0; scan_win2529 <= 32'd0; scan_win2530 <= 32'd0; scan_win2531 <= 32'd0; scan_win2532 <= 32'd0; scan_win2533 <= 32'd0; scan_win2534 <= 32'd0; scan_win2535 <= 32'd0; scan_win2536 <= 32'd0; scan_win2537 <= 32'd0; scan_win2538 <= 32'd0; scan_win2539 <= 32'd0; scan_win2540 <= 32'd0; scan_win2541 <= 32'd0; scan_win2542 <= 32'd0; scan_win2543 <= 32'd0; scan_win2544 <= 32'd0; scan_win2545 <= 32'd0; scan_win2546 <= 32'd0; scan_win2547 <= 32'd0; scan_win2548 <= 32'd0; scan_win2549 <= 32'd0; scan_win2550 <= 32'd0; scan_win2551 <= 32'd0; scan_win2552 <= 32'd0; scan_win2553 <= 32'd0; scan_win2554 <= 32'd0; scan_win2555 <= 32'd0; scan_win2556 <= 32'd0; scan_win2557 <= 32'd0; scan_win2558 <= 32'd0; scan_win2559 <= 32'd0; scan_win2560 <= 32'd0; scan_win2561 <= 32'd0; scan_win2562 <= 32'd0; scan_win2563 <= 32'd0; scan_win2564 <= 32'd0; scan_win2565 <= 32'd0; scan_win2566 <= 32'd0; scan_win2567 <= 32'd0; scan_win2568 <= 32'd0; scan_win2569 <= 32'd0; scan_win2570 <= 32'd0; scan_win2571 <= 32'd0; scan_win2572 <= 32'd0; scan_win2573 <= 32'd0; scan_win2574 <= 32'd0; scan_win2575 <= 32'd0; scan_win2576 <= 32'd0; scan_win2577 <= 32'd0; scan_win2578 <= 32'd0; scan_win2579 <= 32'd0; scan_win2580 <= 32'd0; scan_win2581 <= 32'd0; scan_win2582 <= 32'd0; scan_win2583 <= 32'd0; scan_win2584 <= 32'd0; scan_win2585 <= 32'd0; scan_win2586 <= 32'd0; scan_win2587 <= 32'd0; scan_win2588 <= 32'd0; scan_win2589 <= 32'd0; scan_win2590 <= 32'd0; scan_win2591 <= 32'd0; scan_win2592 <= 32'd0; scan_win2593 <= 32'd0; scan_win2594 <= 32'd0; scan_win2595 <= 32'd0; scan_win2596 <= 32'd0; scan_win2597 <= 32'd0; scan_win2598 <= 32'd0; scan_win2599 <= 32'd0; scan_win2600 <= 32'd0; 
      scan_win2601 <= 32'd0; scan_win2602 <= 32'd0; scan_win2603 <= 32'd0; scan_win2604 <= 32'd0; scan_win2605 <= 32'd0; scan_win2606 <= 32'd0; scan_win2607 <= 32'd0; scan_win2608 <= 32'd0; scan_win2609 <= 32'd0; scan_win2610 <= 32'd0; scan_win2611 <= 32'd0; scan_win2612 <= 32'd0; scan_win2613 <= 32'd0; scan_win2614 <= 32'd0; scan_win2615 <= 32'd0; scan_win2616 <= 32'd0; scan_win2617 <= 32'd0; scan_win2618 <= 32'd0; scan_win2619 <= 32'd0; scan_win2620 <= 32'd0; scan_win2621 <= 32'd0; scan_win2622 <= 32'd0; scan_win2623 <= 32'd0; scan_win2624 <= 32'd0; scan_win2625 <= 32'd0; scan_win2626 <= 32'd0; scan_win2627 <= 32'd0; scan_win2628 <= 32'd0; scan_win2629 <= 32'd0; scan_win2630 <= 32'd0; scan_win2631 <= 32'd0; scan_win2632 <= 32'd0; scan_win2633 <= 32'd0; scan_win2634 <= 32'd0; scan_win2635 <= 32'd0; scan_win2636 <= 32'd0; scan_win2637 <= 32'd0; scan_win2638 <= 32'd0; scan_win2639 <= 32'd0; scan_win2640 <= 32'd0; scan_win2641 <= 32'd0; scan_win2642 <= 32'd0; scan_win2643 <= 32'd0; scan_win2644 <= 32'd0; scan_win2645 <= 32'd0; scan_win2646 <= 32'd0; scan_win2647 <= 32'd0; scan_win2648 <= 32'd0; scan_win2649 <= 32'd0; scan_win2650 <= 32'd0; scan_win2651 <= 32'd0; scan_win2652 <= 32'd0; scan_win2653 <= 32'd0; scan_win2654 <= 32'd0; scan_win2655 <= 32'd0; scan_win2656 <= 32'd0; scan_win2657 <= 32'd0; scan_win2658 <= 32'd0; scan_win2659 <= 32'd0; scan_win2660 <= 32'd0; scan_win2661 <= 32'd0; scan_win2662 <= 32'd0; scan_win2663 <= 32'd0; scan_win2664 <= 32'd0; scan_win2665 <= 32'd0; scan_win2666 <= 32'd0; scan_win2667 <= 32'd0; scan_win2668 <= 32'd0; scan_win2669 <= 32'd0; scan_win2670 <= 32'd0; scan_win2671 <= 32'd0; scan_win2672 <= 32'd0; scan_win2673 <= 32'd0; scan_win2674 <= 32'd0; scan_win2675 <= 32'd0; scan_win2676 <= 32'd0; scan_win2677 <= 32'd0; scan_win2678 <= 32'd0; scan_win2679 <= 32'd0; scan_win2680 <= 32'd0; scan_win2681 <= 32'd0; scan_win2682 <= 32'd0; scan_win2683 <= 32'd0; scan_win2684 <= 32'd0; scan_win2685 <= 32'd0; scan_win2686 <= 32'd0; scan_win2687 <= 32'd0; scan_win2688 <= 32'd0; scan_win2689 <= 32'd0; scan_win2690 <= 32'd0; scan_win2691 <= 32'd0; scan_win2692 <= 32'd0; scan_win2693 <= 32'd0; scan_win2694 <= 32'd0; scan_win2695 <= 32'd0; scan_win2696 <= 32'd0; scan_win2697 <= 32'd0; scan_win2698 <= 32'd0; scan_win2699 <= 32'd0; scan_win2700 <= 32'd0; scan_win2701 <= 32'd0; scan_win2702 <= 32'd0; scan_win2703 <= 32'd0; scan_win2704 <= 32'd0; scan_win2705 <= 32'd0; scan_win2706 <= 32'd0; scan_win2707 <= 32'd0; scan_win2708 <= 32'd0; scan_win2709 <= 32'd0; scan_win2710 <= 32'd0; scan_win2711 <= 32'd0; scan_win2712 <= 32'd0; scan_win2713 <= 32'd0; scan_win2714 <= 32'd0; scan_win2715 <= 32'd0; scan_win2716 <= 32'd0; scan_win2717 <= 32'd0; scan_win2718 <= 32'd0; scan_win2719 <= 32'd0; scan_win2720 <= 32'd0; scan_win2721 <= 32'd0; scan_win2722 <= 32'd0; scan_win2723 <= 32'd0; scan_win2724 <= 32'd0; scan_win2725 <= 32'd0; scan_win2726 <= 32'd0; scan_win2727 <= 32'd0; scan_win2728 <= 32'd0; scan_win2729 <= 32'd0; scan_win2730 <= 32'd0; scan_win2731 <= 32'd0; scan_win2732 <= 32'd0; scan_win2733 <= 32'd0; scan_win2734 <= 32'd0; scan_win2735 <= 32'd0; scan_win2736 <= 32'd0; scan_win2737 <= 32'd0; scan_win2738 <= 32'd0; scan_win2739 <= 32'd0; scan_win2740 <= 32'd0; scan_win2741 <= 32'd0; scan_win2742 <= 32'd0; scan_win2743 <= 32'd0; scan_win2744 <= 32'd0; scan_win2745 <= 32'd0; scan_win2746 <= 32'd0; scan_win2747 <= 32'd0; scan_win2748 <= 32'd0; scan_win2749 <= 32'd0; scan_win2750 <= 32'd0; scan_win2751 <= 32'd0; scan_win2752 <= 32'd0; scan_win2753 <= 32'd0; scan_win2754 <= 32'd0; scan_win2755 <= 32'd0; scan_win2756 <= 32'd0; scan_win2757 <= 32'd0; scan_win2758 <= 32'd0; scan_win2759 <= 32'd0; scan_win2760 <= 32'd0; scan_win2761 <= 32'd0; scan_win2762 <= 32'd0; scan_win2763 <= 32'd0; scan_win2764 <= 32'd0; scan_win2765 <= 32'd0; scan_win2766 <= 32'd0; scan_win2767 <= 32'd0; scan_win2768 <= 32'd0; scan_win2769 <= 32'd0; scan_win2770 <= 32'd0; scan_win2771 <= 32'd0; scan_win2772 <= 32'd0; scan_win2773 <= 32'd0; scan_win2774 <= 32'd0; scan_win2775 <= 32'd0; scan_win2776 <= 32'd0; scan_win2777 <= 32'd0; scan_win2778 <= 32'd0; scan_win2779 <= 32'd0; scan_win2780 <= 32'd0; scan_win2781 <= 32'd0; scan_win2782 <= 32'd0; scan_win2783 <= 32'd0; scan_win2784 <= 32'd0; scan_win2785 <= 32'd0; scan_win2786 <= 32'd0; scan_win2787 <= 32'd0; scan_win2788 <= 32'd0; scan_win2789 <= 32'd0; scan_win2790 <= 32'd0; scan_win2791 <= 32'd0; scan_win2792 <= 32'd0; scan_win2793 <= 32'd0; scan_win2794 <= 32'd0; scan_win2795 <= 32'd0; scan_win2796 <= 32'd0; scan_win2797 <= 32'd0; scan_win2798 <= 32'd0; scan_win2799 <= 32'd0; scan_win2800 <= 32'd0; 
      scan_win2801 <= 32'd0; scan_win2802 <= 32'd0; scan_win2803 <= 32'd0; scan_win2804 <= 32'd0; scan_win2805 <= 32'd0; scan_win2806 <= 32'd0; scan_win2807 <= 32'd0; scan_win2808 <= 32'd0; scan_win2809 <= 32'd0; scan_win2810 <= 32'd0; scan_win2811 <= 32'd0; scan_win2812 <= 32'd0; scan_win2813 <= 32'd0; scan_win2814 <= 32'd0; scan_win2815 <= 32'd0; scan_win2816 <= 32'd0; scan_win2817 <= 32'd0; scan_win2818 <= 32'd0; scan_win2819 <= 32'd0; scan_win2820 <= 32'd0; scan_win2821 <= 32'd0; scan_win2822 <= 32'd0; scan_win2823 <= 32'd0; scan_win2824 <= 32'd0; scan_win2825 <= 32'd0; scan_win2826 <= 32'd0; scan_win2827 <= 32'd0; scan_win2828 <= 32'd0; scan_win2829 <= 32'd0; scan_win2830 <= 32'd0; scan_win2831 <= 32'd0; scan_win2832 <= 32'd0; scan_win2833 <= 32'd0; scan_win2834 <= 32'd0; scan_win2835 <= 32'd0; scan_win2836 <= 32'd0; scan_win2837 <= 32'd0; scan_win2838 <= 32'd0; scan_win2839 <= 32'd0; scan_win2840 <= 32'd0; scan_win2841 <= 32'd0; scan_win2842 <= 32'd0; scan_win2843 <= 32'd0; scan_win2844 <= 32'd0; scan_win2845 <= 32'd0; scan_win2846 <= 32'd0; scan_win2847 <= 32'd0; scan_win2848 <= 32'd0; scan_win2849 <= 32'd0; scan_win2850 <= 32'd0; scan_win2851 <= 32'd0; scan_win2852 <= 32'd0; scan_win2853 <= 32'd0; scan_win2854 <= 32'd0; scan_win2855 <= 32'd0; scan_win2856 <= 32'd0; scan_win2857 <= 32'd0; scan_win2858 <= 32'd0; scan_win2859 <= 32'd0; scan_win2860 <= 32'd0; scan_win2861 <= 32'd0; scan_win2862 <= 32'd0; scan_win2863 <= 32'd0; scan_win2864 <= 32'd0; scan_win2865 <= 32'd0; scan_win2866 <= 32'd0; scan_win2867 <= 32'd0; scan_win2868 <= 32'd0; scan_win2869 <= 32'd0; scan_win2870 <= 32'd0; scan_win2871 <= 32'd0; scan_win2872 <= 32'd0; scan_win2873 <= 32'd0; scan_win2874 <= 32'd0; scan_win2875 <= 32'd0; scan_win2876 <= 32'd0; scan_win2877 <= 32'd0; scan_win2878 <= 32'd0; scan_win2879 <= 32'd0; scan_win2880 <= 32'd0; scan_win2881 <= 32'd0; scan_win2882 <= 32'd0; scan_win2883 <= 32'd0; scan_win2884 <= 32'd0; scan_win2885 <= 32'd0; scan_win2886 <= 32'd0; scan_win2887 <= 32'd0; scan_win2888 <= 32'd0; scan_win2889 <= 32'd0; scan_win2890 <= 32'd0; scan_win2891 <= 32'd0; scan_win2892 <= 32'd0; scan_win2893 <= 32'd0; scan_win2894 <= 32'd0; scan_win2895 <= 32'd0; scan_win2896 <= 32'd0; scan_win2897 <= 32'd0; scan_win2898 <= 32'd0; scan_win2899 <= 32'd0; scan_win2900 <= 32'd0; scan_win2901 <= 32'd0; scan_win2902 <= 32'd0; scan_win2903 <= 32'd0; scan_win2904 <= 32'd0; scan_win2905 <= 32'd0; scan_win2906 <= 32'd0; scan_win2907 <= 32'd0; scan_win2908 <= 32'd0; scan_win2909 <= 32'd0; scan_win2910 <= 32'd0; scan_win2911 <= 32'd0; scan_win2912 <= 32'd0;
    end else begin: move_scan_wins
      scan_win0 <= scan_win;
      scan_win1 <= scan_win0; scan_win2 <= scan_win1; scan_win3 <= scan_win2; scan_win4 <= scan_win3; scan_win5 <= scan_win4; scan_win6 <= scan_win5; scan_win7 <= scan_win6; scan_win8 <= scan_win7; scan_win9 <= scan_win8; scan_win10 <= scan_win9; scan_win11 <= scan_win10; scan_win12 <= scan_win11; scan_win13 <= scan_win12; scan_win14 <= scan_win13; scan_win15 <= scan_win14; scan_win16 <= scan_win15; scan_win17 <= scan_win16; scan_win18 <= scan_win17; scan_win19 <= scan_win18; scan_win20 <= scan_win19; scan_win21 <= scan_win20; scan_win22 <= scan_win21; scan_win23 <= scan_win22; scan_win24 <= scan_win23; scan_win25 <= scan_win24; scan_win26 <= scan_win25; scan_win27 <= scan_win26; scan_win28 <= scan_win27; scan_win29 <= scan_win28; scan_win30 <= scan_win29; scan_win31 <= scan_win30; scan_win32 <= scan_win31; scan_win33 <= scan_win32; scan_win34 <= scan_win33; scan_win35 <= scan_win34; scan_win36 <= scan_win35; scan_win37 <= scan_win36; scan_win38 <= scan_win37; scan_win39 <= scan_win38; scan_win40 <= scan_win39; scan_win41 <= scan_win40; scan_win42 <= scan_win41; scan_win43 <= scan_win42; scan_win44 <= scan_win43; scan_win45 <= scan_win44; scan_win46 <= scan_win45; scan_win47 <= scan_win46; scan_win48 <= scan_win47; scan_win49 <= scan_win48; scan_win50 <= scan_win49; scan_win51 <= scan_win50; scan_win52 <= scan_win51; scan_win53 <= scan_win52; scan_win54 <= scan_win53; scan_win55 <= scan_win54; scan_win56 <= scan_win55; scan_win57 <= scan_win56; scan_win58 <= scan_win57; scan_win59 <= scan_win58; scan_win60 <= scan_win59; scan_win61 <= scan_win60; scan_win62 <= scan_win61; scan_win63 <= scan_win62; scan_win64 <= scan_win63; scan_win65 <= scan_win64; scan_win66 <= scan_win65; scan_win67 <= scan_win66; scan_win68 <= scan_win67; scan_win69 <= scan_win68; scan_win70 <= scan_win69; scan_win71 <= scan_win70; scan_win72 <= scan_win71; scan_win73 <= scan_win72; scan_win74 <= scan_win73; scan_win75 <= scan_win74; scan_win76 <= scan_win75; scan_win77 <= scan_win76; scan_win78 <= scan_win77; scan_win79 <= scan_win78; scan_win80 <= scan_win79; scan_win81 <= scan_win80; scan_win82 <= scan_win81; scan_win83 <= scan_win82; scan_win84 <= scan_win83; scan_win85 <= scan_win84; scan_win86 <= scan_win85; scan_win87 <= scan_win86; scan_win88 <= scan_win87; scan_win89 <= scan_win88; scan_win90 <= scan_win89; scan_win91 <= scan_win90; scan_win92 <= scan_win91; scan_win93 <= scan_win92; scan_win94 <= scan_win93; scan_win95 <= scan_win94; scan_win96 <= scan_win95; scan_win97 <= scan_win96; scan_win98 <= scan_win97; scan_win99 <= scan_win98; scan_win100 <= scan_win99; scan_win101 <= scan_win100; scan_win102 <= scan_win101; scan_win103 <= scan_win102; scan_win104 <= scan_win103; scan_win105 <= scan_win104; scan_win106 <= scan_win105; scan_win107 <= scan_win106; scan_win108 <= scan_win107; scan_win109 <= scan_win108; scan_win110 <= scan_win109; scan_win111 <= scan_win110; scan_win112 <= scan_win111; scan_win113 <= scan_win112; scan_win114 <= scan_win113; scan_win115 <= scan_win114; scan_win116 <= scan_win115; scan_win117 <= scan_win116; scan_win118 <= scan_win117; scan_win119 <= scan_win118; scan_win120 <= scan_win119; scan_win121 <= scan_win120; scan_win122 <= scan_win121; scan_win123 <= scan_win122; scan_win124 <= scan_win123; scan_win125 <= scan_win124; scan_win126 <= scan_win125; scan_win127 <= scan_win126; scan_win128 <= scan_win127; scan_win129 <= scan_win128; scan_win130 <= scan_win129; scan_win131 <= scan_win130; scan_win132 <= scan_win131; scan_win133 <= scan_win132; scan_win134 <= scan_win133; scan_win135 <= scan_win134; scan_win136 <= scan_win135; scan_win137 <= scan_win136; scan_win138 <= scan_win137; scan_win139 <= scan_win138; scan_win140 <= scan_win139; scan_win141 <= scan_win140; scan_win142 <= scan_win141; scan_win143 <= scan_win142; scan_win144 <= scan_win143; scan_win145 <= scan_win144; scan_win146 <= scan_win145; scan_win147 <= scan_win146; scan_win148 <= scan_win147; scan_win149 <= scan_win148; scan_win150 <= scan_win149; scan_win151 <= scan_win150; scan_win152 <= scan_win151; scan_win153 <= scan_win152; scan_win154 <= scan_win153; scan_win155 <= scan_win154; scan_win156 <= scan_win155; scan_win157 <= scan_win156; scan_win158 <= scan_win157; scan_win159 <= scan_win158; scan_win160 <= scan_win159; scan_win161 <= scan_win160; scan_win162 <= scan_win161; scan_win163 <= scan_win162; scan_win164 <= scan_win163; scan_win165 <= scan_win164; scan_win166 <= scan_win165; scan_win167 <= scan_win166; scan_win168 <= scan_win167; scan_win169 <= scan_win168; scan_win170 <= scan_win169; scan_win171 <= scan_win170; scan_win172 <= scan_win171; scan_win173 <= scan_win172; scan_win174 <= scan_win173; scan_win175 <= scan_win174; scan_win176 <= scan_win175; scan_win177 <= scan_win176; scan_win178 <= scan_win177; scan_win179 <= scan_win178; scan_win180 <= scan_win179; scan_win181 <= scan_win180; scan_win182 <= scan_win181; scan_win183 <= scan_win182; scan_win184 <= scan_win183; scan_win185 <= scan_win184; scan_win186 <= scan_win185; scan_win187 <= scan_win186; scan_win188 <= scan_win187; scan_win189 <= scan_win188; scan_win190 <= scan_win189; scan_win191 <= scan_win190; scan_win192 <= scan_win191; scan_win193 <= scan_win192; scan_win194 <= scan_win193; scan_win195 <= scan_win194; scan_win196 <= scan_win195; scan_win197 <= scan_win196; scan_win198 <= scan_win197; scan_win199 <= scan_win198; scan_win200 <= scan_win199; 
      scan_win201 <= scan_win200; scan_win202 <= scan_win201; scan_win203 <= scan_win202; scan_win204 <= scan_win203; scan_win205 <= scan_win204; scan_win206 <= scan_win205; scan_win207 <= scan_win206; scan_win208 <= scan_win207; scan_win209 <= scan_win208; scan_win210 <= scan_win209; scan_win211 <= scan_win210; scan_win212 <= scan_win211; scan_win213 <= scan_win212; scan_win214 <= scan_win213; scan_win215 <= scan_win214; scan_win216 <= scan_win215; scan_win217 <= scan_win216; scan_win218 <= scan_win217; scan_win219 <= scan_win218; scan_win220 <= scan_win219; scan_win221 <= scan_win220; scan_win222 <= scan_win221; scan_win223 <= scan_win222; scan_win224 <= scan_win223; scan_win225 <= scan_win224; scan_win226 <= scan_win225; scan_win227 <= scan_win226; scan_win228 <= scan_win227; scan_win229 <= scan_win228; scan_win230 <= scan_win229; scan_win231 <= scan_win230; scan_win232 <= scan_win231; scan_win233 <= scan_win232; scan_win234 <= scan_win233; scan_win235 <= scan_win234; scan_win236 <= scan_win235; scan_win237 <= scan_win236; scan_win238 <= scan_win237; scan_win239 <= scan_win238; scan_win240 <= scan_win239; scan_win241 <= scan_win240; scan_win242 <= scan_win241; scan_win243 <= scan_win242; scan_win244 <= scan_win243; scan_win245 <= scan_win244; scan_win246 <= scan_win245; scan_win247 <= scan_win246; scan_win248 <= scan_win247; scan_win249 <= scan_win248; scan_win250 <= scan_win249; scan_win251 <= scan_win250; scan_win252 <= scan_win251; scan_win253 <= scan_win252; scan_win254 <= scan_win253; scan_win255 <= scan_win254; scan_win256 <= scan_win255; scan_win257 <= scan_win256; scan_win258 <= scan_win257; scan_win259 <= scan_win258; scan_win260 <= scan_win259; scan_win261 <= scan_win260; scan_win262 <= scan_win261; scan_win263 <= scan_win262; scan_win264 <= scan_win263; scan_win265 <= scan_win264; scan_win266 <= scan_win265; scan_win267 <= scan_win266; scan_win268 <= scan_win267; scan_win269 <= scan_win268; scan_win270 <= scan_win269; scan_win271 <= scan_win270; scan_win272 <= scan_win271; scan_win273 <= scan_win272; scan_win274 <= scan_win273; scan_win275 <= scan_win274; scan_win276 <= scan_win275; scan_win277 <= scan_win276; scan_win278 <= scan_win277; scan_win279 <= scan_win278; scan_win280 <= scan_win279; scan_win281 <= scan_win280; scan_win282 <= scan_win281; scan_win283 <= scan_win282; scan_win284 <= scan_win283; scan_win285 <= scan_win284; scan_win286 <= scan_win285; scan_win287 <= scan_win286; scan_win288 <= scan_win287; scan_win289 <= scan_win288; scan_win290 <= scan_win289; scan_win291 <= scan_win290; scan_win292 <= scan_win291; scan_win293 <= scan_win292; scan_win294 <= scan_win293; scan_win295 <= scan_win294; scan_win296 <= scan_win295; scan_win297 <= scan_win296; scan_win298 <= scan_win297; scan_win299 <= scan_win298; scan_win300 <= scan_win299; scan_win301 <= scan_win300; scan_win302 <= scan_win301; scan_win303 <= scan_win302; scan_win304 <= scan_win303; scan_win305 <= scan_win304; scan_win306 <= scan_win305; scan_win307 <= scan_win306; scan_win308 <= scan_win307; scan_win309 <= scan_win308; scan_win310 <= scan_win309; scan_win311 <= scan_win310; scan_win312 <= scan_win311; scan_win313 <= scan_win312; scan_win314 <= scan_win313; scan_win315 <= scan_win314; scan_win316 <= scan_win315; scan_win317 <= scan_win316; scan_win318 <= scan_win317; scan_win319 <= scan_win318; scan_win320 <= scan_win319; scan_win321 <= scan_win320; scan_win322 <= scan_win321; scan_win323 <= scan_win322; scan_win324 <= scan_win323; scan_win325 <= scan_win324; scan_win326 <= scan_win325; scan_win327 <= scan_win326; scan_win328 <= scan_win327; scan_win329 <= scan_win328; scan_win330 <= scan_win329; scan_win331 <= scan_win330; scan_win332 <= scan_win331; scan_win333 <= scan_win332; scan_win334 <= scan_win333; scan_win335 <= scan_win334; scan_win336 <= scan_win335; scan_win337 <= scan_win336; scan_win338 <= scan_win337; scan_win339 <= scan_win338; scan_win340 <= scan_win339; scan_win341 <= scan_win340; scan_win342 <= scan_win341; scan_win343 <= scan_win342; scan_win344 <= scan_win343; scan_win345 <= scan_win344; scan_win346 <= scan_win345; scan_win347 <= scan_win346; scan_win348 <= scan_win347; scan_win349 <= scan_win348; scan_win350 <= scan_win349; scan_win351 <= scan_win350; scan_win352 <= scan_win351; scan_win353 <= scan_win352; scan_win354 <= scan_win353; scan_win355 <= scan_win354; scan_win356 <= scan_win355; scan_win357 <= scan_win356; scan_win358 <= scan_win357; scan_win359 <= scan_win358; scan_win360 <= scan_win359; scan_win361 <= scan_win360; scan_win362 <= scan_win361; scan_win363 <= scan_win362; scan_win364 <= scan_win363; scan_win365 <= scan_win364; scan_win366 <= scan_win365; scan_win367 <= scan_win366; scan_win368 <= scan_win367; scan_win369 <= scan_win368; scan_win370 <= scan_win369; scan_win371 <= scan_win370; scan_win372 <= scan_win371; scan_win373 <= scan_win372; scan_win374 <= scan_win373; scan_win375 <= scan_win374; scan_win376 <= scan_win375; scan_win377 <= scan_win376; scan_win378 <= scan_win377; scan_win379 <= scan_win378; scan_win380 <= scan_win379; scan_win381 <= scan_win380; scan_win382 <= scan_win381; scan_win383 <= scan_win382; scan_win384 <= scan_win383; scan_win385 <= scan_win384; scan_win386 <= scan_win385; scan_win387 <= scan_win386; scan_win388 <= scan_win387; scan_win389 <= scan_win388; scan_win390 <= scan_win389; scan_win391 <= scan_win390; scan_win392 <= scan_win391; scan_win393 <= scan_win392; scan_win394 <= scan_win393; scan_win395 <= scan_win394; scan_win396 <= scan_win395; scan_win397 <= scan_win396; scan_win398 <= scan_win397; scan_win399 <= scan_win398; scan_win400 <= scan_win399; 
      scan_win401 <= scan_win400; scan_win402 <= scan_win401; scan_win403 <= scan_win402; scan_win404 <= scan_win403; scan_win405 <= scan_win404; scan_win406 <= scan_win405; scan_win407 <= scan_win406; scan_win408 <= scan_win407; scan_win409 <= scan_win408; scan_win410 <= scan_win409; scan_win411 <= scan_win410; scan_win412 <= scan_win411; scan_win413 <= scan_win412; scan_win414 <= scan_win413; scan_win415 <= scan_win414; scan_win416 <= scan_win415; scan_win417 <= scan_win416; scan_win418 <= scan_win417; scan_win419 <= scan_win418; scan_win420 <= scan_win419; scan_win421 <= scan_win420; scan_win422 <= scan_win421; scan_win423 <= scan_win422; scan_win424 <= scan_win423; scan_win425 <= scan_win424; scan_win426 <= scan_win425; scan_win427 <= scan_win426; scan_win428 <= scan_win427; scan_win429 <= scan_win428; scan_win430 <= scan_win429; scan_win431 <= scan_win430; scan_win432 <= scan_win431; scan_win433 <= scan_win432; scan_win434 <= scan_win433; scan_win435 <= scan_win434; scan_win436 <= scan_win435; scan_win437 <= scan_win436; scan_win438 <= scan_win437; scan_win439 <= scan_win438; scan_win440 <= scan_win439; scan_win441 <= scan_win440; scan_win442 <= scan_win441; scan_win443 <= scan_win442; scan_win444 <= scan_win443; scan_win445 <= scan_win444; scan_win446 <= scan_win445; scan_win447 <= scan_win446; scan_win448 <= scan_win447; scan_win449 <= scan_win448; scan_win450 <= scan_win449; scan_win451 <= scan_win450; scan_win452 <= scan_win451; scan_win453 <= scan_win452; scan_win454 <= scan_win453; scan_win455 <= scan_win454; scan_win456 <= scan_win455; scan_win457 <= scan_win456; scan_win458 <= scan_win457; scan_win459 <= scan_win458; scan_win460 <= scan_win459; scan_win461 <= scan_win460; scan_win462 <= scan_win461; scan_win463 <= scan_win462; scan_win464 <= scan_win463; scan_win465 <= scan_win464; scan_win466 <= scan_win465; scan_win467 <= scan_win466; scan_win468 <= scan_win467; scan_win469 <= scan_win468; scan_win470 <= scan_win469; scan_win471 <= scan_win470; scan_win472 <= scan_win471; scan_win473 <= scan_win472; scan_win474 <= scan_win473; scan_win475 <= scan_win474; scan_win476 <= scan_win475; scan_win477 <= scan_win476; scan_win478 <= scan_win477; scan_win479 <= scan_win478; scan_win480 <= scan_win479; scan_win481 <= scan_win480; scan_win482 <= scan_win481; scan_win483 <= scan_win482; scan_win484 <= scan_win483; scan_win485 <= scan_win484; scan_win486 <= scan_win485; scan_win487 <= scan_win486; scan_win488 <= scan_win487; scan_win489 <= scan_win488; scan_win490 <= scan_win489; scan_win491 <= scan_win490; scan_win492 <= scan_win491; scan_win493 <= scan_win492; scan_win494 <= scan_win493; scan_win495 <= scan_win494; scan_win496 <= scan_win495; scan_win497 <= scan_win496; scan_win498 <= scan_win497; scan_win499 <= scan_win498; scan_win500 <= scan_win499; scan_win501 <= scan_win500; scan_win502 <= scan_win501; scan_win503 <= scan_win502; scan_win504 <= scan_win503; scan_win505 <= scan_win504; scan_win506 <= scan_win505; scan_win507 <= scan_win506; scan_win508 <= scan_win507; scan_win509 <= scan_win508; scan_win510 <= scan_win509; scan_win511 <= scan_win510; scan_win512 <= scan_win511; scan_win513 <= scan_win512; scan_win514 <= scan_win513; scan_win515 <= scan_win514; scan_win516 <= scan_win515; scan_win517 <= scan_win516; scan_win518 <= scan_win517; scan_win519 <= scan_win518; scan_win520 <= scan_win519; scan_win521 <= scan_win520; scan_win522 <= scan_win521; scan_win523 <= scan_win522; scan_win524 <= scan_win523; scan_win525 <= scan_win524; scan_win526 <= scan_win525; scan_win527 <= scan_win526; scan_win528 <= scan_win527; scan_win529 <= scan_win528; scan_win530 <= scan_win529; scan_win531 <= scan_win530; scan_win532 <= scan_win531; scan_win533 <= scan_win532; scan_win534 <= scan_win533; scan_win535 <= scan_win534; scan_win536 <= scan_win535; scan_win537 <= scan_win536; scan_win538 <= scan_win537; scan_win539 <= scan_win538; scan_win540 <= scan_win539; scan_win541 <= scan_win540; scan_win542 <= scan_win541; scan_win543 <= scan_win542; scan_win544 <= scan_win543; scan_win545 <= scan_win544; scan_win546 <= scan_win545; scan_win547 <= scan_win546; scan_win548 <= scan_win547; scan_win549 <= scan_win548; scan_win550 <= scan_win549; scan_win551 <= scan_win550; scan_win552 <= scan_win551; scan_win553 <= scan_win552; scan_win554 <= scan_win553; scan_win555 <= scan_win554; scan_win556 <= scan_win555; scan_win557 <= scan_win556; scan_win558 <= scan_win557; scan_win559 <= scan_win558; scan_win560 <= scan_win559; scan_win561 <= scan_win560; scan_win562 <= scan_win561; scan_win563 <= scan_win562; scan_win564 <= scan_win563; scan_win565 <= scan_win564; scan_win566 <= scan_win565; scan_win567 <= scan_win566; scan_win568 <= scan_win567; scan_win569 <= scan_win568; scan_win570 <= scan_win569; scan_win571 <= scan_win570; scan_win572 <= scan_win571; scan_win573 <= scan_win572; scan_win574 <= scan_win573; scan_win575 <= scan_win574; scan_win576 <= scan_win575; scan_win577 <= scan_win576; scan_win578 <= scan_win577; scan_win579 <= scan_win578; scan_win580 <= scan_win579; scan_win581 <= scan_win580; scan_win582 <= scan_win581; scan_win583 <= scan_win582; scan_win584 <= scan_win583; scan_win585 <= scan_win584; scan_win586 <= scan_win585; scan_win587 <= scan_win586; scan_win588 <= scan_win587; scan_win589 <= scan_win588; scan_win590 <= scan_win589; scan_win591 <= scan_win590; scan_win592 <= scan_win591; scan_win593 <= scan_win592; scan_win594 <= scan_win593; scan_win595 <= scan_win594; scan_win596 <= scan_win595; scan_win597 <= scan_win596; scan_win598 <= scan_win597; scan_win599 <= scan_win598; scan_win600 <= scan_win599; 
      scan_win601 <= scan_win600; scan_win602 <= scan_win601; scan_win603 <= scan_win602; scan_win604 <= scan_win603; scan_win605 <= scan_win604; scan_win606 <= scan_win605; scan_win607 <= scan_win606; scan_win608 <= scan_win607; scan_win609 <= scan_win608; scan_win610 <= scan_win609; scan_win611 <= scan_win610; scan_win612 <= scan_win611; scan_win613 <= scan_win612; scan_win614 <= scan_win613; scan_win615 <= scan_win614; scan_win616 <= scan_win615; scan_win617 <= scan_win616; scan_win618 <= scan_win617; scan_win619 <= scan_win618; scan_win620 <= scan_win619; scan_win621 <= scan_win620; scan_win622 <= scan_win621; scan_win623 <= scan_win622; scan_win624 <= scan_win623; scan_win625 <= scan_win624; scan_win626 <= scan_win625; scan_win627 <= scan_win626; scan_win628 <= scan_win627; scan_win629 <= scan_win628; scan_win630 <= scan_win629; scan_win631 <= scan_win630; scan_win632 <= scan_win631; scan_win633 <= scan_win632; scan_win634 <= scan_win633; scan_win635 <= scan_win634; scan_win636 <= scan_win635; scan_win637 <= scan_win636; scan_win638 <= scan_win637; scan_win639 <= scan_win638; scan_win640 <= scan_win639; scan_win641 <= scan_win640; scan_win642 <= scan_win641; scan_win643 <= scan_win642; scan_win644 <= scan_win643; scan_win645 <= scan_win644; scan_win646 <= scan_win645; scan_win647 <= scan_win646; scan_win648 <= scan_win647; scan_win649 <= scan_win648; scan_win650 <= scan_win649; scan_win651 <= scan_win650; scan_win652 <= scan_win651; scan_win653 <= scan_win652; scan_win654 <= scan_win653; scan_win655 <= scan_win654; scan_win656 <= scan_win655; scan_win657 <= scan_win656; scan_win658 <= scan_win657; scan_win659 <= scan_win658; scan_win660 <= scan_win659; scan_win661 <= scan_win660; scan_win662 <= scan_win661; scan_win663 <= scan_win662; scan_win664 <= scan_win663; scan_win665 <= scan_win664; scan_win666 <= scan_win665; scan_win667 <= scan_win666; scan_win668 <= scan_win667; scan_win669 <= scan_win668; scan_win670 <= scan_win669; scan_win671 <= scan_win670; scan_win672 <= scan_win671; scan_win673 <= scan_win672; scan_win674 <= scan_win673; scan_win675 <= scan_win674; scan_win676 <= scan_win675; scan_win677 <= scan_win676; scan_win678 <= scan_win677; scan_win679 <= scan_win678; scan_win680 <= scan_win679; scan_win681 <= scan_win680; scan_win682 <= scan_win681; scan_win683 <= scan_win682; scan_win684 <= scan_win683; scan_win685 <= scan_win684; scan_win686 <= scan_win685; scan_win687 <= scan_win686; scan_win688 <= scan_win687; scan_win689 <= scan_win688; scan_win690 <= scan_win689; scan_win691 <= scan_win690; scan_win692 <= scan_win691; scan_win693 <= scan_win692; scan_win694 <= scan_win693; scan_win695 <= scan_win694; scan_win696 <= scan_win695; scan_win697 <= scan_win696; scan_win698 <= scan_win697; scan_win699 <= scan_win698; scan_win700 <= scan_win699; scan_win701 <= scan_win700; scan_win702 <= scan_win701; scan_win703 <= scan_win702; scan_win704 <= scan_win703; scan_win705 <= scan_win704; scan_win706 <= scan_win705; scan_win707 <= scan_win706; scan_win708 <= scan_win707; scan_win709 <= scan_win708; scan_win710 <= scan_win709; scan_win711 <= scan_win710; scan_win712 <= scan_win711; scan_win713 <= scan_win712; scan_win714 <= scan_win713; scan_win715 <= scan_win714; scan_win716 <= scan_win715; scan_win717 <= scan_win716; scan_win718 <= scan_win717; scan_win719 <= scan_win718; scan_win720 <= scan_win719; scan_win721 <= scan_win720; scan_win722 <= scan_win721; scan_win723 <= scan_win722; scan_win724 <= scan_win723; scan_win725 <= scan_win724; scan_win726 <= scan_win725; scan_win727 <= scan_win726; scan_win728 <= scan_win727; scan_win729 <= scan_win728; scan_win730 <= scan_win729; scan_win731 <= scan_win730; scan_win732 <= scan_win731; scan_win733 <= scan_win732; scan_win734 <= scan_win733; scan_win735 <= scan_win734; scan_win736 <= scan_win735; scan_win737 <= scan_win736; scan_win738 <= scan_win737; scan_win739 <= scan_win738; scan_win740 <= scan_win739; scan_win741 <= scan_win740; scan_win742 <= scan_win741; scan_win743 <= scan_win742; scan_win744 <= scan_win743; scan_win745 <= scan_win744; scan_win746 <= scan_win745; scan_win747 <= scan_win746; scan_win748 <= scan_win747; scan_win749 <= scan_win748; scan_win750 <= scan_win749; scan_win751 <= scan_win750; scan_win752 <= scan_win751; scan_win753 <= scan_win752; scan_win754 <= scan_win753; scan_win755 <= scan_win754; scan_win756 <= scan_win755; scan_win757 <= scan_win756; scan_win758 <= scan_win757; scan_win759 <= scan_win758; scan_win760 <= scan_win759; scan_win761 <= scan_win760; scan_win762 <= scan_win761; scan_win763 <= scan_win762; scan_win764 <= scan_win763; scan_win765 <= scan_win764; scan_win766 <= scan_win765; scan_win767 <= scan_win766; scan_win768 <= scan_win767; scan_win769 <= scan_win768; scan_win770 <= scan_win769; scan_win771 <= scan_win770; scan_win772 <= scan_win771; scan_win773 <= scan_win772; scan_win774 <= scan_win773; scan_win775 <= scan_win774; scan_win776 <= scan_win775; scan_win777 <= scan_win776; scan_win778 <= scan_win777; scan_win779 <= scan_win778; scan_win780 <= scan_win779; scan_win781 <= scan_win780; scan_win782 <= scan_win781; scan_win783 <= scan_win782; scan_win784 <= scan_win783; scan_win785 <= scan_win784; scan_win786 <= scan_win785; scan_win787 <= scan_win786; scan_win788 <= scan_win787; scan_win789 <= scan_win788; scan_win790 <= scan_win789; scan_win791 <= scan_win790; scan_win792 <= scan_win791; scan_win793 <= scan_win792; scan_win794 <= scan_win793; scan_win795 <= scan_win794; scan_win796 <= scan_win795; scan_win797 <= scan_win796; scan_win798 <= scan_win797; scan_win799 <= scan_win798; scan_win800 <= scan_win799; 
      scan_win801 <= scan_win800; scan_win802 <= scan_win801; scan_win803 <= scan_win802; scan_win804 <= scan_win803; scan_win805 <= scan_win804; scan_win806 <= scan_win805; scan_win807 <= scan_win806; scan_win808 <= scan_win807; scan_win809 <= scan_win808; scan_win810 <= scan_win809; scan_win811 <= scan_win810; scan_win812 <= scan_win811; scan_win813 <= scan_win812; scan_win814 <= scan_win813; scan_win815 <= scan_win814; scan_win816 <= scan_win815; scan_win817 <= scan_win816; scan_win818 <= scan_win817; scan_win819 <= scan_win818; scan_win820 <= scan_win819; scan_win821 <= scan_win820; scan_win822 <= scan_win821; scan_win823 <= scan_win822; scan_win824 <= scan_win823; scan_win825 <= scan_win824; scan_win826 <= scan_win825; scan_win827 <= scan_win826; scan_win828 <= scan_win827; scan_win829 <= scan_win828; scan_win830 <= scan_win829; scan_win831 <= scan_win830; scan_win832 <= scan_win831; scan_win833 <= scan_win832; scan_win834 <= scan_win833; scan_win835 <= scan_win834; scan_win836 <= scan_win835; scan_win837 <= scan_win836; scan_win838 <= scan_win837; scan_win839 <= scan_win838; scan_win840 <= scan_win839; scan_win841 <= scan_win840; scan_win842 <= scan_win841; scan_win843 <= scan_win842; scan_win844 <= scan_win843; scan_win845 <= scan_win844; scan_win846 <= scan_win845; scan_win847 <= scan_win846; scan_win848 <= scan_win847; scan_win849 <= scan_win848; scan_win850 <= scan_win849; scan_win851 <= scan_win850; scan_win852 <= scan_win851; scan_win853 <= scan_win852; scan_win854 <= scan_win853; scan_win855 <= scan_win854; scan_win856 <= scan_win855; scan_win857 <= scan_win856; scan_win858 <= scan_win857; scan_win859 <= scan_win858; scan_win860 <= scan_win859; scan_win861 <= scan_win860; scan_win862 <= scan_win861; scan_win863 <= scan_win862; scan_win864 <= scan_win863; scan_win865 <= scan_win864; scan_win866 <= scan_win865; scan_win867 <= scan_win866; scan_win868 <= scan_win867; scan_win869 <= scan_win868; scan_win870 <= scan_win869; scan_win871 <= scan_win870; scan_win872 <= scan_win871; scan_win873 <= scan_win872; scan_win874 <= scan_win873; scan_win875 <= scan_win874; scan_win876 <= scan_win875; scan_win877 <= scan_win876; scan_win878 <= scan_win877; scan_win879 <= scan_win878; scan_win880 <= scan_win879; scan_win881 <= scan_win880; scan_win882 <= scan_win881; scan_win883 <= scan_win882; scan_win884 <= scan_win883; scan_win885 <= scan_win884; scan_win886 <= scan_win885; scan_win887 <= scan_win886; scan_win888 <= scan_win887; scan_win889 <= scan_win888; scan_win890 <= scan_win889; scan_win891 <= scan_win890; scan_win892 <= scan_win891; scan_win893 <= scan_win892; scan_win894 <= scan_win893; scan_win895 <= scan_win894; scan_win896 <= scan_win895; scan_win897 <= scan_win896; scan_win898 <= scan_win897; scan_win899 <= scan_win898; scan_win900 <= scan_win899; scan_win901 <= scan_win900; scan_win902 <= scan_win901; scan_win903 <= scan_win902; scan_win904 <= scan_win903; scan_win905 <= scan_win904; scan_win906 <= scan_win905; scan_win907 <= scan_win906; scan_win908 <= scan_win907; scan_win909 <= scan_win908; scan_win910 <= scan_win909; scan_win911 <= scan_win910; scan_win912 <= scan_win911; scan_win913 <= scan_win912; scan_win914 <= scan_win913; scan_win915 <= scan_win914; scan_win916 <= scan_win915; scan_win917 <= scan_win916; scan_win918 <= scan_win917; scan_win919 <= scan_win918; scan_win920 <= scan_win919; scan_win921 <= scan_win920; scan_win922 <= scan_win921; scan_win923 <= scan_win922; scan_win924 <= scan_win923; scan_win925 <= scan_win924; scan_win926 <= scan_win925; scan_win927 <= scan_win926; scan_win928 <= scan_win927; scan_win929 <= scan_win928; scan_win930 <= scan_win929; scan_win931 <= scan_win930; scan_win932 <= scan_win931; scan_win933 <= scan_win932; scan_win934 <= scan_win933; scan_win935 <= scan_win934; scan_win936 <= scan_win935; scan_win937 <= scan_win936; scan_win938 <= scan_win937; scan_win939 <= scan_win938; scan_win940 <= scan_win939; scan_win941 <= scan_win940; scan_win942 <= scan_win941; scan_win943 <= scan_win942; scan_win944 <= scan_win943; scan_win945 <= scan_win944; scan_win946 <= scan_win945; scan_win947 <= scan_win946; scan_win948 <= scan_win947; scan_win949 <= scan_win948; scan_win950 <= scan_win949; scan_win951 <= scan_win950; scan_win952 <= scan_win951; scan_win953 <= scan_win952; scan_win954 <= scan_win953; scan_win955 <= scan_win954; scan_win956 <= scan_win955; scan_win957 <= scan_win956; scan_win958 <= scan_win957; scan_win959 <= scan_win958; scan_win960 <= scan_win959; scan_win961 <= scan_win960; scan_win962 <= scan_win961; scan_win963 <= scan_win962; scan_win964 <= scan_win963; scan_win965 <= scan_win964; scan_win966 <= scan_win965; scan_win967 <= scan_win966; scan_win968 <= scan_win967; scan_win969 <= scan_win968; scan_win970 <= scan_win969; scan_win971 <= scan_win970; scan_win972 <= scan_win971; scan_win973 <= scan_win972; scan_win974 <= scan_win973; scan_win975 <= scan_win974; scan_win976 <= scan_win975; scan_win977 <= scan_win976; scan_win978 <= scan_win977; scan_win979 <= scan_win978; scan_win980 <= scan_win979; scan_win981 <= scan_win980; scan_win982 <= scan_win981; scan_win983 <= scan_win982; scan_win984 <= scan_win983; scan_win985 <= scan_win984; scan_win986 <= scan_win985; scan_win987 <= scan_win986; scan_win988 <= scan_win987; scan_win989 <= scan_win988; scan_win990 <= scan_win989; scan_win991 <= scan_win990; scan_win992 <= scan_win991; scan_win993 <= scan_win992; scan_win994 <= scan_win993; scan_win995 <= scan_win994; scan_win996 <= scan_win995; scan_win997 <= scan_win996; scan_win998 <= scan_win997; scan_win999 <= scan_win998; scan_win1000 <= scan_win999; 
      scan_win1001 <= scan_win1000; scan_win1002 <= scan_win1001; scan_win1003 <= scan_win1002; scan_win1004 <= scan_win1003; scan_win1005 <= scan_win1004; scan_win1006 <= scan_win1005; scan_win1007 <= scan_win1006; scan_win1008 <= scan_win1007; scan_win1009 <= scan_win1008; scan_win1010 <= scan_win1009; scan_win1011 <= scan_win1010; scan_win1012 <= scan_win1011; scan_win1013 <= scan_win1012; scan_win1014 <= scan_win1013; scan_win1015 <= scan_win1014; scan_win1016 <= scan_win1015; scan_win1017 <= scan_win1016; scan_win1018 <= scan_win1017; scan_win1019 <= scan_win1018; scan_win1020 <= scan_win1019; scan_win1021 <= scan_win1020; scan_win1022 <= scan_win1021; scan_win1023 <= scan_win1022; scan_win1024 <= scan_win1023; scan_win1025 <= scan_win1024; scan_win1026 <= scan_win1025; scan_win1027 <= scan_win1026; scan_win1028 <= scan_win1027; scan_win1029 <= scan_win1028; scan_win1030 <= scan_win1029; scan_win1031 <= scan_win1030; scan_win1032 <= scan_win1031; scan_win1033 <= scan_win1032; scan_win1034 <= scan_win1033; scan_win1035 <= scan_win1034; scan_win1036 <= scan_win1035; scan_win1037 <= scan_win1036; scan_win1038 <= scan_win1037; scan_win1039 <= scan_win1038; scan_win1040 <= scan_win1039; scan_win1041 <= scan_win1040; scan_win1042 <= scan_win1041; scan_win1043 <= scan_win1042; scan_win1044 <= scan_win1043; scan_win1045 <= scan_win1044; scan_win1046 <= scan_win1045; scan_win1047 <= scan_win1046; scan_win1048 <= scan_win1047; scan_win1049 <= scan_win1048; scan_win1050 <= scan_win1049; scan_win1051 <= scan_win1050; scan_win1052 <= scan_win1051; scan_win1053 <= scan_win1052; scan_win1054 <= scan_win1053; scan_win1055 <= scan_win1054; scan_win1056 <= scan_win1055; scan_win1057 <= scan_win1056; scan_win1058 <= scan_win1057; scan_win1059 <= scan_win1058; scan_win1060 <= scan_win1059; scan_win1061 <= scan_win1060; scan_win1062 <= scan_win1061; scan_win1063 <= scan_win1062; scan_win1064 <= scan_win1063; scan_win1065 <= scan_win1064; scan_win1066 <= scan_win1065; scan_win1067 <= scan_win1066; scan_win1068 <= scan_win1067; scan_win1069 <= scan_win1068; scan_win1070 <= scan_win1069; scan_win1071 <= scan_win1070; scan_win1072 <= scan_win1071; scan_win1073 <= scan_win1072; scan_win1074 <= scan_win1073; scan_win1075 <= scan_win1074; scan_win1076 <= scan_win1075; scan_win1077 <= scan_win1076; scan_win1078 <= scan_win1077; scan_win1079 <= scan_win1078; scan_win1080 <= scan_win1079; scan_win1081 <= scan_win1080; scan_win1082 <= scan_win1081; scan_win1083 <= scan_win1082; scan_win1084 <= scan_win1083; scan_win1085 <= scan_win1084; scan_win1086 <= scan_win1085; scan_win1087 <= scan_win1086; scan_win1088 <= scan_win1087; scan_win1089 <= scan_win1088; scan_win1090 <= scan_win1089; scan_win1091 <= scan_win1090; scan_win1092 <= scan_win1091; scan_win1093 <= scan_win1092; scan_win1094 <= scan_win1093; scan_win1095 <= scan_win1094; scan_win1096 <= scan_win1095; scan_win1097 <= scan_win1096; scan_win1098 <= scan_win1097; scan_win1099 <= scan_win1098; scan_win1100 <= scan_win1099; scan_win1101 <= scan_win1100; scan_win1102 <= scan_win1101; scan_win1103 <= scan_win1102; scan_win1104 <= scan_win1103; scan_win1105 <= scan_win1104; scan_win1106 <= scan_win1105; scan_win1107 <= scan_win1106; scan_win1108 <= scan_win1107; scan_win1109 <= scan_win1108; scan_win1110 <= scan_win1109; scan_win1111 <= scan_win1110; scan_win1112 <= scan_win1111; scan_win1113 <= scan_win1112; scan_win1114 <= scan_win1113; scan_win1115 <= scan_win1114; scan_win1116 <= scan_win1115; scan_win1117 <= scan_win1116; scan_win1118 <= scan_win1117; scan_win1119 <= scan_win1118; scan_win1120 <= scan_win1119; scan_win1121 <= scan_win1120; scan_win1122 <= scan_win1121; scan_win1123 <= scan_win1122; scan_win1124 <= scan_win1123; scan_win1125 <= scan_win1124; scan_win1126 <= scan_win1125; scan_win1127 <= scan_win1126; scan_win1128 <= scan_win1127; scan_win1129 <= scan_win1128; scan_win1130 <= scan_win1129; scan_win1131 <= scan_win1130; scan_win1132 <= scan_win1131; scan_win1133 <= scan_win1132; scan_win1134 <= scan_win1133; scan_win1135 <= scan_win1134; scan_win1136 <= scan_win1135; scan_win1137 <= scan_win1136; scan_win1138 <= scan_win1137; scan_win1139 <= scan_win1138; scan_win1140 <= scan_win1139; scan_win1141 <= scan_win1140; scan_win1142 <= scan_win1141; scan_win1143 <= scan_win1142; scan_win1144 <= scan_win1143; scan_win1145 <= scan_win1144; scan_win1146 <= scan_win1145; scan_win1147 <= scan_win1146; scan_win1148 <= scan_win1147; scan_win1149 <= scan_win1148; scan_win1150 <= scan_win1149; scan_win1151 <= scan_win1150; scan_win1152 <= scan_win1151; scan_win1153 <= scan_win1152; scan_win1154 <= scan_win1153; scan_win1155 <= scan_win1154; scan_win1156 <= scan_win1155; scan_win1157 <= scan_win1156; scan_win1158 <= scan_win1157; scan_win1159 <= scan_win1158; scan_win1160 <= scan_win1159; scan_win1161 <= scan_win1160; scan_win1162 <= scan_win1161; scan_win1163 <= scan_win1162; scan_win1164 <= scan_win1163; scan_win1165 <= scan_win1164; scan_win1166 <= scan_win1165; scan_win1167 <= scan_win1166; scan_win1168 <= scan_win1167; scan_win1169 <= scan_win1168; scan_win1170 <= scan_win1169; scan_win1171 <= scan_win1170; scan_win1172 <= scan_win1171; scan_win1173 <= scan_win1172; scan_win1174 <= scan_win1173; scan_win1175 <= scan_win1174; scan_win1176 <= scan_win1175; scan_win1177 <= scan_win1176; scan_win1178 <= scan_win1177; scan_win1179 <= scan_win1178; scan_win1180 <= scan_win1179; scan_win1181 <= scan_win1180; scan_win1182 <= scan_win1181; scan_win1183 <= scan_win1182; scan_win1184 <= scan_win1183; scan_win1185 <= scan_win1184; scan_win1186 <= scan_win1185; scan_win1187 <= scan_win1186; scan_win1188 <= scan_win1187; scan_win1189 <= scan_win1188; scan_win1190 <= scan_win1189; scan_win1191 <= scan_win1190; scan_win1192 <= scan_win1191; scan_win1193 <= scan_win1192; scan_win1194 <= scan_win1193; scan_win1195 <= scan_win1194; scan_win1196 <= scan_win1195; scan_win1197 <= scan_win1196; scan_win1198 <= scan_win1197; scan_win1199 <= scan_win1198; scan_win1200 <= scan_win1199; 
      scan_win1201 <= scan_win1200; scan_win1202 <= scan_win1201; scan_win1203 <= scan_win1202; scan_win1204 <= scan_win1203; scan_win1205 <= scan_win1204; scan_win1206 <= scan_win1205; scan_win1207 <= scan_win1206; scan_win1208 <= scan_win1207; scan_win1209 <= scan_win1208; scan_win1210 <= scan_win1209; scan_win1211 <= scan_win1210; scan_win1212 <= scan_win1211; scan_win1213 <= scan_win1212; scan_win1214 <= scan_win1213; scan_win1215 <= scan_win1214; scan_win1216 <= scan_win1215; scan_win1217 <= scan_win1216; scan_win1218 <= scan_win1217; scan_win1219 <= scan_win1218; scan_win1220 <= scan_win1219; scan_win1221 <= scan_win1220; scan_win1222 <= scan_win1221; scan_win1223 <= scan_win1222; scan_win1224 <= scan_win1223; scan_win1225 <= scan_win1224; scan_win1226 <= scan_win1225; scan_win1227 <= scan_win1226; scan_win1228 <= scan_win1227; scan_win1229 <= scan_win1228; scan_win1230 <= scan_win1229; scan_win1231 <= scan_win1230; scan_win1232 <= scan_win1231; scan_win1233 <= scan_win1232; scan_win1234 <= scan_win1233; scan_win1235 <= scan_win1234; scan_win1236 <= scan_win1235; scan_win1237 <= scan_win1236; scan_win1238 <= scan_win1237; scan_win1239 <= scan_win1238; scan_win1240 <= scan_win1239; scan_win1241 <= scan_win1240; scan_win1242 <= scan_win1241; scan_win1243 <= scan_win1242; scan_win1244 <= scan_win1243; scan_win1245 <= scan_win1244; scan_win1246 <= scan_win1245; scan_win1247 <= scan_win1246; scan_win1248 <= scan_win1247; scan_win1249 <= scan_win1248; scan_win1250 <= scan_win1249; scan_win1251 <= scan_win1250; scan_win1252 <= scan_win1251; scan_win1253 <= scan_win1252; scan_win1254 <= scan_win1253; scan_win1255 <= scan_win1254; scan_win1256 <= scan_win1255; scan_win1257 <= scan_win1256; scan_win1258 <= scan_win1257; scan_win1259 <= scan_win1258; scan_win1260 <= scan_win1259; scan_win1261 <= scan_win1260; scan_win1262 <= scan_win1261; scan_win1263 <= scan_win1262; scan_win1264 <= scan_win1263; scan_win1265 <= scan_win1264; scan_win1266 <= scan_win1265; scan_win1267 <= scan_win1266; scan_win1268 <= scan_win1267; scan_win1269 <= scan_win1268; scan_win1270 <= scan_win1269; scan_win1271 <= scan_win1270; scan_win1272 <= scan_win1271; scan_win1273 <= scan_win1272; scan_win1274 <= scan_win1273; scan_win1275 <= scan_win1274; scan_win1276 <= scan_win1275; scan_win1277 <= scan_win1276; scan_win1278 <= scan_win1277; scan_win1279 <= scan_win1278; scan_win1280 <= scan_win1279; scan_win1281 <= scan_win1280; scan_win1282 <= scan_win1281; scan_win1283 <= scan_win1282; scan_win1284 <= scan_win1283; scan_win1285 <= scan_win1284; scan_win1286 <= scan_win1285; scan_win1287 <= scan_win1286; scan_win1288 <= scan_win1287; scan_win1289 <= scan_win1288; scan_win1290 <= scan_win1289; scan_win1291 <= scan_win1290; scan_win1292 <= scan_win1291; scan_win1293 <= scan_win1292; scan_win1294 <= scan_win1293; scan_win1295 <= scan_win1294; scan_win1296 <= scan_win1295; scan_win1297 <= scan_win1296; scan_win1298 <= scan_win1297; scan_win1299 <= scan_win1298; scan_win1300 <= scan_win1299; scan_win1301 <= scan_win1300; scan_win1302 <= scan_win1301; scan_win1303 <= scan_win1302; scan_win1304 <= scan_win1303; scan_win1305 <= scan_win1304; scan_win1306 <= scan_win1305; scan_win1307 <= scan_win1306; scan_win1308 <= scan_win1307; scan_win1309 <= scan_win1308; scan_win1310 <= scan_win1309; scan_win1311 <= scan_win1310; scan_win1312 <= scan_win1311; scan_win1313 <= scan_win1312; scan_win1314 <= scan_win1313; scan_win1315 <= scan_win1314; scan_win1316 <= scan_win1315; scan_win1317 <= scan_win1316; scan_win1318 <= scan_win1317; scan_win1319 <= scan_win1318; scan_win1320 <= scan_win1319; scan_win1321 <= scan_win1320; scan_win1322 <= scan_win1321; scan_win1323 <= scan_win1322; scan_win1324 <= scan_win1323; scan_win1325 <= scan_win1324; scan_win1326 <= scan_win1325; scan_win1327 <= scan_win1326; scan_win1328 <= scan_win1327; scan_win1329 <= scan_win1328; scan_win1330 <= scan_win1329; scan_win1331 <= scan_win1330; scan_win1332 <= scan_win1331; scan_win1333 <= scan_win1332; scan_win1334 <= scan_win1333; scan_win1335 <= scan_win1334; scan_win1336 <= scan_win1335; scan_win1337 <= scan_win1336; scan_win1338 <= scan_win1337; scan_win1339 <= scan_win1338; scan_win1340 <= scan_win1339; scan_win1341 <= scan_win1340; scan_win1342 <= scan_win1341; scan_win1343 <= scan_win1342; scan_win1344 <= scan_win1343; scan_win1345 <= scan_win1344; scan_win1346 <= scan_win1345; scan_win1347 <= scan_win1346; scan_win1348 <= scan_win1347; scan_win1349 <= scan_win1348; scan_win1350 <= scan_win1349; scan_win1351 <= scan_win1350; scan_win1352 <= scan_win1351; scan_win1353 <= scan_win1352; scan_win1354 <= scan_win1353; scan_win1355 <= scan_win1354; scan_win1356 <= scan_win1355; scan_win1357 <= scan_win1356; scan_win1358 <= scan_win1357; scan_win1359 <= scan_win1358; scan_win1360 <= scan_win1359; scan_win1361 <= scan_win1360; scan_win1362 <= scan_win1361; scan_win1363 <= scan_win1362; scan_win1364 <= scan_win1363; scan_win1365 <= scan_win1364; scan_win1366 <= scan_win1365; scan_win1367 <= scan_win1366; scan_win1368 <= scan_win1367; scan_win1369 <= scan_win1368; scan_win1370 <= scan_win1369; scan_win1371 <= scan_win1370; scan_win1372 <= scan_win1371; scan_win1373 <= scan_win1372; scan_win1374 <= scan_win1373; scan_win1375 <= scan_win1374; scan_win1376 <= scan_win1375; scan_win1377 <= scan_win1376; scan_win1378 <= scan_win1377; scan_win1379 <= scan_win1378; scan_win1380 <= scan_win1379; scan_win1381 <= scan_win1380; scan_win1382 <= scan_win1381; scan_win1383 <= scan_win1382; scan_win1384 <= scan_win1383; scan_win1385 <= scan_win1384; scan_win1386 <= scan_win1385; scan_win1387 <= scan_win1386; scan_win1388 <= scan_win1387; scan_win1389 <= scan_win1388; scan_win1390 <= scan_win1389; scan_win1391 <= scan_win1390; scan_win1392 <= scan_win1391; scan_win1393 <= scan_win1392; scan_win1394 <= scan_win1393; scan_win1395 <= scan_win1394; scan_win1396 <= scan_win1395; scan_win1397 <= scan_win1396; scan_win1398 <= scan_win1397; scan_win1399 <= scan_win1398; scan_win1400 <= scan_win1399; 
      scan_win1401 <= scan_win1400; scan_win1402 <= scan_win1401; scan_win1403 <= scan_win1402; scan_win1404 <= scan_win1403; scan_win1405 <= scan_win1404; scan_win1406 <= scan_win1405; scan_win1407 <= scan_win1406; scan_win1408 <= scan_win1407; scan_win1409 <= scan_win1408; scan_win1410 <= scan_win1409; scan_win1411 <= scan_win1410; scan_win1412 <= scan_win1411; scan_win1413 <= scan_win1412; scan_win1414 <= scan_win1413; scan_win1415 <= scan_win1414; scan_win1416 <= scan_win1415; scan_win1417 <= scan_win1416; scan_win1418 <= scan_win1417; scan_win1419 <= scan_win1418; scan_win1420 <= scan_win1419; scan_win1421 <= scan_win1420; scan_win1422 <= scan_win1421; scan_win1423 <= scan_win1422; scan_win1424 <= scan_win1423; scan_win1425 <= scan_win1424; scan_win1426 <= scan_win1425; scan_win1427 <= scan_win1426; scan_win1428 <= scan_win1427; scan_win1429 <= scan_win1428; scan_win1430 <= scan_win1429; scan_win1431 <= scan_win1430; scan_win1432 <= scan_win1431; scan_win1433 <= scan_win1432; scan_win1434 <= scan_win1433; scan_win1435 <= scan_win1434; scan_win1436 <= scan_win1435; scan_win1437 <= scan_win1436; scan_win1438 <= scan_win1437; scan_win1439 <= scan_win1438; scan_win1440 <= scan_win1439; scan_win1441 <= scan_win1440; scan_win1442 <= scan_win1441; scan_win1443 <= scan_win1442; scan_win1444 <= scan_win1443; scan_win1445 <= scan_win1444; scan_win1446 <= scan_win1445; scan_win1447 <= scan_win1446; scan_win1448 <= scan_win1447; scan_win1449 <= scan_win1448; scan_win1450 <= scan_win1449; scan_win1451 <= scan_win1450; scan_win1452 <= scan_win1451; scan_win1453 <= scan_win1452; scan_win1454 <= scan_win1453; scan_win1455 <= scan_win1454; scan_win1456 <= scan_win1455; scan_win1457 <= scan_win1456; scan_win1458 <= scan_win1457; scan_win1459 <= scan_win1458; scan_win1460 <= scan_win1459; scan_win1461 <= scan_win1460; scan_win1462 <= scan_win1461; scan_win1463 <= scan_win1462; scan_win1464 <= scan_win1463; scan_win1465 <= scan_win1464; scan_win1466 <= scan_win1465; scan_win1467 <= scan_win1466; scan_win1468 <= scan_win1467; scan_win1469 <= scan_win1468; scan_win1470 <= scan_win1469; scan_win1471 <= scan_win1470; scan_win1472 <= scan_win1471; scan_win1473 <= scan_win1472; scan_win1474 <= scan_win1473; scan_win1475 <= scan_win1474; scan_win1476 <= scan_win1475; scan_win1477 <= scan_win1476; scan_win1478 <= scan_win1477; scan_win1479 <= scan_win1478; scan_win1480 <= scan_win1479; scan_win1481 <= scan_win1480; scan_win1482 <= scan_win1481; scan_win1483 <= scan_win1482; scan_win1484 <= scan_win1483; scan_win1485 <= scan_win1484; scan_win1486 <= scan_win1485; scan_win1487 <= scan_win1486; scan_win1488 <= scan_win1487; scan_win1489 <= scan_win1488; scan_win1490 <= scan_win1489; scan_win1491 <= scan_win1490; scan_win1492 <= scan_win1491; scan_win1493 <= scan_win1492; scan_win1494 <= scan_win1493; scan_win1495 <= scan_win1494; scan_win1496 <= scan_win1495; scan_win1497 <= scan_win1496; scan_win1498 <= scan_win1497; scan_win1499 <= scan_win1498; scan_win1500 <= scan_win1499; scan_win1501 <= scan_win1500; scan_win1502 <= scan_win1501; scan_win1503 <= scan_win1502; scan_win1504 <= scan_win1503; scan_win1505 <= scan_win1504; scan_win1506 <= scan_win1505; scan_win1507 <= scan_win1506; scan_win1508 <= scan_win1507; scan_win1509 <= scan_win1508; scan_win1510 <= scan_win1509; scan_win1511 <= scan_win1510; scan_win1512 <= scan_win1511; scan_win1513 <= scan_win1512; scan_win1514 <= scan_win1513; scan_win1515 <= scan_win1514; scan_win1516 <= scan_win1515; scan_win1517 <= scan_win1516; scan_win1518 <= scan_win1517; scan_win1519 <= scan_win1518; scan_win1520 <= scan_win1519; scan_win1521 <= scan_win1520; scan_win1522 <= scan_win1521; scan_win1523 <= scan_win1522; scan_win1524 <= scan_win1523; scan_win1525 <= scan_win1524; scan_win1526 <= scan_win1525; scan_win1527 <= scan_win1526; scan_win1528 <= scan_win1527; scan_win1529 <= scan_win1528; scan_win1530 <= scan_win1529; scan_win1531 <= scan_win1530; scan_win1532 <= scan_win1531; scan_win1533 <= scan_win1532; scan_win1534 <= scan_win1533; scan_win1535 <= scan_win1534; scan_win1536 <= scan_win1535; scan_win1537 <= scan_win1536; scan_win1538 <= scan_win1537; scan_win1539 <= scan_win1538; scan_win1540 <= scan_win1539; scan_win1541 <= scan_win1540; scan_win1542 <= scan_win1541; scan_win1543 <= scan_win1542; scan_win1544 <= scan_win1543; scan_win1545 <= scan_win1544; scan_win1546 <= scan_win1545; scan_win1547 <= scan_win1546; scan_win1548 <= scan_win1547; scan_win1549 <= scan_win1548; scan_win1550 <= scan_win1549; scan_win1551 <= scan_win1550; scan_win1552 <= scan_win1551; scan_win1553 <= scan_win1552; scan_win1554 <= scan_win1553; scan_win1555 <= scan_win1554; scan_win1556 <= scan_win1555; scan_win1557 <= scan_win1556; scan_win1558 <= scan_win1557; scan_win1559 <= scan_win1558; scan_win1560 <= scan_win1559; scan_win1561 <= scan_win1560; scan_win1562 <= scan_win1561; scan_win1563 <= scan_win1562; scan_win1564 <= scan_win1563; scan_win1565 <= scan_win1564; scan_win1566 <= scan_win1565; scan_win1567 <= scan_win1566; scan_win1568 <= scan_win1567; scan_win1569 <= scan_win1568; scan_win1570 <= scan_win1569; scan_win1571 <= scan_win1570; scan_win1572 <= scan_win1571; scan_win1573 <= scan_win1572; scan_win1574 <= scan_win1573; scan_win1575 <= scan_win1574; scan_win1576 <= scan_win1575; scan_win1577 <= scan_win1576; scan_win1578 <= scan_win1577; scan_win1579 <= scan_win1578; scan_win1580 <= scan_win1579; scan_win1581 <= scan_win1580; scan_win1582 <= scan_win1581; scan_win1583 <= scan_win1582; scan_win1584 <= scan_win1583; scan_win1585 <= scan_win1584; scan_win1586 <= scan_win1585; scan_win1587 <= scan_win1586; scan_win1588 <= scan_win1587; scan_win1589 <= scan_win1588; scan_win1590 <= scan_win1589; scan_win1591 <= scan_win1590; scan_win1592 <= scan_win1591; scan_win1593 <= scan_win1592; scan_win1594 <= scan_win1593; scan_win1595 <= scan_win1594; scan_win1596 <= scan_win1595; scan_win1597 <= scan_win1596; scan_win1598 <= scan_win1597; scan_win1599 <= scan_win1598; scan_win1600 <= scan_win1599; 
      scan_win1601 <= scan_win1600; scan_win1602 <= scan_win1601; scan_win1603 <= scan_win1602; scan_win1604 <= scan_win1603; scan_win1605 <= scan_win1604; scan_win1606 <= scan_win1605; scan_win1607 <= scan_win1606; scan_win1608 <= scan_win1607; scan_win1609 <= scan_win1608; scan_win1610 <= scan_win1609; scan_win1611 <= scan_win1610; scan_win1612 <= scan_win1611; scan_win1613 <= scan_win1612; scan_win1614 <= scan_win1613; scan_win1615 <= scan_win1614; scan_win1616 <= scan_win1615; scan_win1617 <= scan_win1616; scan_win1618 <= scan_win1617; scan_win1619 <= scan_win1618; scan_win1620 <= scan_win1619; scan_win1621 <= scan_win1620; scan_win1622 <= scan_win1621; scan_win1623 <= scan_win1622; scan_win1624 <= scan_win1623; scan_win1625 <= scan_win1624; scan_win1626 <= scan_win1625; scan_win1627 <= scan_win1626; scan_win1628 <= scan_win1627; scan_win1629 <= scan_win1628; scan_win1630 <= scan_win1629; scan_win1631 <= scan_win1630; scan_win1632 <= scan_win1631; scan_win1633 <= scan_win1632; scan_win1634 <= scan_win1633; scan_win1635 <= scan_win1634; scan_win1636 <= scan_win1635; scan_win1637 <= scan_win1636; scan_win1638 <= scan_win1637; scan_win1639 <= scan_win1638; scan_win1640 <= scan_win1639; scan_win1641 <= scan_win1640; scan_win1642 <= scan_win1641; scan_win1643 <= scan_win1642; scan_win1644 <= scan_win1643; scan_win1645 <= scan_win1644; scan_win1646 <= scan_win1645; scan_win1647 <= scan_win1646; scan_win1648 <= scan_win1647; scan_win1649 <= scan_win1648; scan_win1650 <= scan_win1649; scan_win1651 <= scan_win1650; scan_win1652 <= scan_win1651; scan_win1653 <= scan_win1652; scan_win1654 <= scan_win1653; scan_win1655 <= scan_win1654; scan_win1656 <= scan_win1655; scan_win1657 <= scan_win1656; scan_win1658 <= scan_win1657; scan_win1659 <= scan_win1658; scan_win1660 <= scan_win1659; scan_win1661 <= scan_win1660; scan_win1662 <= scan_win1661; scan_win1663 <= scan_win1662; scan_win1664 <= scan_win1663; scan_win1665 <= scan_win1664; scan_win1666 <= scan_win1665; scan_win1667 <= scan_win1666; scan_win1668 <= scan_win1667; scan_win1669 <= scan_win1668; scan_win1670 <= scan_win1669; scan_win1671 <= scan_win1670; scan_win1672 <= scan_win1671; scan_win1673 <= scan_win1672; scan_win1674 <= scan_win1673; scan_win1675 <= scan_win1674; scan_win1676 <= scan_win1675; scan_win1677 <= scan_win1676; scan_win1678 <= scan_win1677; scan_win1679 <= scan_win1678; scan_win1680 <= scan_win1679; scan_win1681 <= scan_win1680; scan_win1682 <= scan_win1681; scan_win1683 <= scan_win1682; scan_win1684 <= scan_win1683; scan_win1685 <= scan_win1684; scan_win1686 <= scan_win1685; scan_win1687 <= scan_win1686; scan_win1688 <= scan_win1687; scan_win1689 <= scan_win1688; scan_win1690 <= scan_win1689; scan_win1691 <= scan_win1690; scan_win1692 <= scan_win1691; scan_win1693 <= scan_win1692; scan_win1694 <= scan_win1693; scan_win1695 <= scan_win1694; scan_win1696 <= scan_win1695; scan_win1697 <= scan_win1696; scan_win1698 <= scan_win1697; scan_win1699 <= scan_win1698; scan_win1700 <= scan_win1699; scan_win1701 <= scan_win1700; scan_win1702 <= scan_win1701; scan_win1703 <= scan_win1702; scan_win1704 <= scan_win1703; scan_win1705 <= scan_win1704; scan_win1706 <= scan_win1705; scan_win1707 <= scan_win1706; scan_win1708 <= scan_win1707; scan_win1709 <= scan_win1708; scan_win1710 <= scan_win1709; scan_win1711 <= scan_win1710; scan_win1712 <= scan_win1711; scan_win1713 <= scan_win1712; scan_win1714 <= scan_win1713; scan_win1715 <= scan_win1714; scan_win1716 <= scan_win1715; scan_win1717 <= scan_win1716; scan_win1718 <= scan_win1717; scan_win1719 <= scan_win1718; scan_win1720 <= scan_win1719; scan_win1721 <= scan_win1720; scan_win1722 <= scan_win1721; scan_win1723 <= scan_win1722; scan_win1724 <= scan_win1723; scan_win1725 <= scan_win1724; scan_win1726 <= scan_win1725; scan_win1727 <= scan_win1726; scan_win1728 <= scan_win1727; scan_win1729 <= scan_win1728; scan_win1730 <= scan_win1729; scan_win1731 <= scan_win1730; scan_win1732 <= scan_win1731; scan_win1733 <= scan_win1732; scan_win1734 <= scan_win1733; scan_win1735 <= scan_win1734; scan_win1736 <= scan_win1735; scan_win1737 <= scan_win1736; scan_win1738 <= scan_win1737; scan_win1739 <= scan_win1738; scan_win1740 <= scan_win1739; scan_win1741 <= scan_win1740; scan_win1742 <= scan_win1741; scan_win1743 <= scan_win1742; scan_win1744 <= scan_win1743; scan_win1745 <= scan_win1744; scan_win1746 <= scan_win1745; scan_win1747 <= scan_win1746; scan_win1748 <= scan_win1747; scan_win1749 <= scan_win1748; scan_win1750 <= scan_win1749; scan_win1751 <= scan_win1750; scan_win1752 <= scan_win1751; scan_win1753 <= scan_win1752; scan_win1754 <= scan_win1753; scan_win1755 <= scan_win1754; scan_win1756 <= scan_win1755; scan_win1757 <= scan_win1756; scan_win1758 <= scan_win1757; scan_win1759 <= scan_win1758; scan_win1760 <= scan_win1759; scan_win1761 <= scan_win1760; scan_win1762 <= scan_win1761; scan_win1763 <= scan_win1762; scan_win1764 <= scan_win1763; scan_win1765 <= scan_win1764; scan_win1766 <= scan_win1765; scan_win1767 <= scan_win1766; scan_win1768 <= scan_win1767; scan_win1769 <= scan_win1768; scan_win1770 <= scan_win1769; scan_win1771 <= scan_win1770; scan_win1772 <= scan_win1771; scan_win1773 <= scan_win1772; scan_win1774 <= scan_win1773; scan_win1775 <= scan_win1774; scan_win1776 <= scan_win1775; scan_win1777 <= scan_win1776; scan_win1778 <= scan_win1777; scan_win1779 <= scan_win1778; scan_win1780 <= scan_win1779; scan_win1781 <= scan_win1780; scan_win1782 <= scan_win1781; scan_win1783 <= scan_win1782; scan_win1784 <= scan_win1783; scan_win1785 <= scan_win1784; scan_win1786 <= scan_win1785; scan_win1787 <= scan_win1786; scan_win1788 <= scan_win1787; scan_win1789 <= scan_win1788; scan_win1790 <= scan_win1789; scan_win1791 <= scan_win1790; scan_win1792 <= scan_win1791; scan_win1793 <= scan_win1792; scan_win1794 <= scan_win1793; scan_win1795 <= scan_win1794; scan_win1796 <= scan_win1795; scan_win1797 <= scan_win1796; scan_win1798 <= scan_win1797; scan_win1799 <= scan_win1798; scan_win1800 <= scan_win1799; 
      scan_win1801 <= scan_win1800; scan_win1802 <= scan_win1801; scan_win1803 <= scan_win1802; scan_win1804 <= scan_win1803; scan_win1805 <= scan_win1804; scan_win1806 <= scan_win1805; scan_win1807 <= scan_win1806; scan_win1808 <= scan_win1807; scan_win1809 <= scan_win1808; scan_win1810 <= scan_win1809; scan_win1811 <= scan_win1810; scan_win1812 <= scan_win1811; scan_win1813 <= scan_win1812; scan_win1814 <= scan_win1813; scan_win1815 <= scan_win1814; scan_win1816 <= scan_win1815; scan_win1817 <= scan_win1816; scan_win1818 <= scan_win1817; scan_win1819 <= scan_win1818; scan_win1820 <= scan_win1819; scan_win1821 <= scan_win1820; scan_win1822 <= scan_win1821; scan_win1823 <= scan_win1822; scan_win1824 <= scan_win1823; scan_win1825 <= scan_win1824; scan_win1826 <= scan_win1825; scan_win1827 <= scan_win1826; scan_win1828 <= scan_win1827; scan_win1829 <= scan_win1828; scan_win1830 <= scan_win1829; scan_win1831 <= scan_win1830; scan_win1832 <= scan_win1831; scan_win1833 <= scan_win1832; scan_win1834 <= scan_win1833; scan_win1835 <= scan_win1834; scan_win1836 <= scan_win1835; scan_win1837 <= scan_win1836; scan_win1838 <= scan_win1837; scan_win1839 <= scan_win1838; scan_win1840 <= scan_win1839; scan_win1841 <= scan_win1840; scan_win1842 <= scan_win1841; scan_win1843 <= scan_win1842; scan_win1844 <= scan_win1843; scan_win1845 <= scan_win1844; scan_win1846 <= scan_win1845; scan_win1847 <= scan_win1846; scan_win1848 <= scan_win1847; scan_win1849 <= scan_win1848; scan_win1850 <= scan_win1849; scan_win1851 <= scan_win1850; scan_win1852 <= scan_win1851; scan_win1853 <= scan_win1852; scan_win1854 <= scan_win1853; scan_win1855 <= scan_win1854; scan_win1856 <= scan_win1855; scan_win1857 <= scan_win1856; scan_win1858 <= scan_win1857; scan_win1859 <= scan_win1858; scan_win1860 <= scan_win1859; scan_win1861 <= scan_win1860; scan_win1862 <= scan_win1861; scan_win1863 <= scan_win1862; scan_win1864 <= scan_win1863; scan_win1865 <= scan_win1864; scan_win1866 <= scan_win1865; scan_win1867 <= scan_win1866; scan_win1868 <= scan_win1867; scan_win1869 <= scan_win1868; scan_win1870 <= scan_win1869; scan_win1871 <= scan_win1870; scan_win1872 <= scan_win1871; scan_win1873 <= scan_win1872; scan_win1874 <= scan_win1873; scan_win1875 <= scan_win1874; scan_win1876 <= scan_win1875; scan_win1877 <= scan_win1876; scan_win1878 <= scan_win1877; scan_win1879 <= scan_win1878; scan_win1880 <= scan_win1879; scan_win1881 <= scan_win1880; scan_win1882 <= scan_win1881; scan_win1883 <= scan_win1882; scan_win1884 <= scan_win1883; scan_win1885 <= scan_win1884; scan_win1886 <= scan_win1885; scan_win1887 <= scan_win1886; scan_win1888 <= scan_win1887; scan_win1889 <= scan_win1888; scan_win1890 <= scan_win1889; scan_win1891 <= scan_win1890; scan_win1892 <= scan_win1891; scan_win1893 <= scan_win1892; scan_win1894 <= scan_win1893; scan_win1895 <= scan_win1894; scan_win1896 <= scan_win1895; scan_win1897 <= scan_win1896; scan_win1898 <= scan_win1897; scan_win1899 <= scan_win1898; scan_win1900 <= scan_win1899; scan_win1901 <= scan_win1900; scan_win1902 <= scan_win1901; scan_win1903 <= scan_win1902; scan_win1904 <= scan_win1903; scan_win1905 <= scan_win1904; scan_win1906 <= scan_win1905; scan_win1907 <= scan_win1906; scan_win1908 <= scan_win1907; scan_win1909 <= scan_win1908; scan_win1910 <= scan_win1909; scan_win1911 <= scan_win1910; scan_win1912 <= scan_win1911; scan_win1913 <= scan_win1912; scan_win1914 <= scan_win1913; scan_win1915 <= scan_win1914; scan_win1916 <= scan_win1915; scan_win1917 <= scan_win1916; scan_win1918 <= scan_win1917; scan_win1919 <= scan_win1918; scan_win1920 <= scan_win1919; scan_win1921 <= scan_win1920; scan_win1922 <= scan_win1921; scan_win1923 <= scan_win1922; scan_win1924 <= scan_win1923; scan_win1925 <= scan_win1924; scan_win1926 <= scan_win1925; scan_win1927 <= scan_win1926; scan_win1928 <= scan_win1927; scan_win1929 <= scan_win1928; scan_win1930 <= scan_win1929; scan_win1931 <= scan_win1930; scan_win1932 <= scan_win1931; scan_win1933 <= scan_win1932; scan_win1934 <= scan_win1933; scan_win1935 <= scan_win1934; scan_win1936 <= scan_win1935; scan_win1937 <= scan_win1936; scan_win1938 <= scan_win1937; scan_win1939 <= scan_win1938; scan_win1940 <= scan_win1939; scan_win1941 <= scan_win1940; scan_win1942 <= scan_win1941; scan_win1943 <= scan_win1942; scan_win1944 <= scan_win1943; scan_win1945 <= scan_win1944; scan_win1946 <= scan_win1945; scan_win1947 <= scan_win1946; scan_win1948 <= scan_win1947; scan_win1949 <= scan_win1948; scan_win1950 <= scan_win1949; scan_win1951 <= scan_win1950; scan_win1952 <= scan_win1951; scan_win1953 <= scan_win1952; scan_win1954 <= scan_win1953; scan_win1955 <= scan_win1954; scan_win1956 <= scan_win1955; scan_win1957 <= scan_win1956; scan_win1958 <= scan_win1957; scan_win1959 <= scan_win1958; scan_win1960 <= scan_win1959; scan_win1961 <= scan_win1960; scan_win1962 <= scan_win1961; scan_win1963 <= scan_win1962; scan_win1964 <= scan_win1963; scan_win1965 <= scan_win1964; scan_win1966 <= scan_win1965; scan_win1967 <= scan_win1966; scan_win1968 <= scan_win1967; scan_win1969 <= scan_win1968; scan_win1970 <= scan_win1969; scan_win1971 <= scan_win1970; scan_win1972 <= scan_win1971; scan_win1973 <= scan_win1972; scan_win1974 <= scan_win1973; scan_win1975 <= scan_win1974; scan_win1976 <= scan_win1975; scan_win1977 <= scan_win1976; scan_win1978 <= scan_win1977; scan_win1979 <= scan_win1978; scan_win1980 <= scan_win1979; scan_win1981 <= scan_win1980; scan_win1982 <= scan_win1981; scan_win1983 <= scan_win1982; scan_win1984 <= scan_win1983; scan_win1985 <= scan_win1984; scan_win1986 <= scan_win1985; scan_win1987 <= scan_win1986; scan_win1988 <= scan_win1987; scan_win1989 <= scan_win1988; scan_win1990 <= scan_win1989; scan_win1991 <= scan_win1990; scan_win1992 <= scan_win1991; scan_win1993 <= scan_win1992; scan_win1994 <= scan_win1993; scan_win1995 <= scan_win1994; scan_win1996 <= scan_win1995; scan_win1997 <= scan_win1996; scan_win1998 <= scan_win1997; scan_win1999 <= scan_win1998; scan_win2000 <= scan_win1999; 
      scan_win2001 <= scan_win2000; scan_win2002 <= scan_win2001; scan_win2003 <= scan_win2002; scan_win2004 <= scan_win2003; scan_win2005 <= scan_win2004; scan_win2006 <= scan_win2005; scan_win2007 <= scan_win2006; scan_win2008 <= scan_win2007; scan_win2009 <= scan_win2008; scan_win2010 <= scan_win2009; scan_win2011 <= scan_win2010; scan_win2012 <= scan_win2011; scan_win2013 <= scan_win2012; scan_win2014 <= scan_win2013; scan_win2015 <= scan_win2014; scan_win2016 <= scan_win2015; scan_win2017 <= scan_win2016; scan_win2018 <= scan_win2017; scan_win2019 <= scan_win2018; scan_win2020 <= scan_win2019; scan_win2021 <= scan_win2020; scan_win2022 <= scan_win2021; scan_win2023 <= scan_win2022; scan_win2024 <= scan_win2023; scan_win2025 <= scan_win2024; scan_win2026 <= scan_win2025; scan_win2027 <= scan_win2026; scan_win2028 <= scan_win2027; scan_win2029 <= scan_win2028; scan_win2030 <= scan_win2029; scan_win2031 <= scan_win2030; scan_win2032 <= scan_win2031; scan_win2033 <= scan_win2032; scan_win2034 <= scan_win2033; scan_win2035 <= scan_win2034; scan_win2036 <= scan_win2035; scan_win2037 <= scan_win2036; scan_win2038 <= scan_win2037; scan_win2039 <= scan_win2038; scan_win2040 <= scan_win2039; scan_win2041 <= scan_win2040; scan_win2042 <= scan_win2041; scan_win2043 <= scan_win2042; scan_win2044 <= scan_win2043; scan_win2045 <= scan_win2044; scan_win2046 <= scan_win2045; scan_win2047 <= scan_win2046; scan_win2048 <= scan_win2047; scan_win2049 <= scan_win2048; scan_win2050 <= scan_win2049; scan_win2051 <= scan_win2050; scan_win2052 <= scan_win2051; scan_win2053 <= scan_win2052; scan_win2054 <= scan_win2053; scan_win2055 <= scan_win2054; scan_win2056 <= scan_win2055; scan_win2057 <= scan_win2056; scan_win2058 <= scan_win2057; scan_win2059 <= scan_win2058; scan_win2060 <= scan_win2059; scan_win2061 <= scan_win2060; scan_win2062 <= scan_win2061; scan_win2063 <= scan_win2062; scan_win2064 <= scan_win2063; scan_win2065 <= scan_win2064; scan_win2066 <= scan_win2065; scan_win2067 <= scan_win2066; scan_win2068 <= scan_win2067; scan_win2069 <= scan_win2068; scan_win2070 <= scan_win2069; scan_win2071 <= scan_win2070; scan_win2072 <= scan_win2071; scan_win2073 <= scan_win2072; scan_win2074 <= scan_win2073; scan_win2075 <= scan_win2074; scan_win2076 <= scan_win2075; scan_win2077 <= scan_win2076; scan_win2078 <= scan_win2077; scan_win2079 <= scan_win2078; scan_win2080 <= scan_win2079; scan_win2081 <= scan_win2080; scan_win2082 <= scan_win2081; scan_win2083 <= scan_win2082; scan_win2084 <= scan_win2083; scan_win2085 <= scan_win2084; scan_win2086 <= scan_win2085; scan_win2087 <= scan_win2086; scan_win2088 <= scan_win2087; scan_win2089 <= scan_win2088; scan_win2090 <= scan_win2089; scan_win2091 <= scan_win2090; scan_win2092 <= scan_win2091; scan_win2093 <= scan_win2092; scan_win2094 <= scan_win2093; scan_win2095 <= scan_win2094; scan_win2096 <= scan_win2095; scan_win2097 <= scan_win2096; scan_win2098 <= scan_win2097; scan_win2099 <= scan_win2098; scan_win2100 <= scan_win2099; scan_win2101 <= scan_win2100; scan_win2102 <= scan_win2101; scan_win2103 <= scan_win2102; scan_win2104 <= scan_win2103; scan_win2105 <= scan_win2104; scan_win2106 <= scan_win2105; scan_win2107 <= scan_win2106; scan_win2108 <= scan_win2107; scan_win2109 <= scan_win2108; scan_win2110 <= scan_win2109; scan_win2111 <= scan_win2110; scan_win2112 <= scan_win2111; scan_win2113 <= scan_win2112; scan_win2114 <= scan_win2113; scan_win2115 <= scan_win2114; scan_win2116 <= scan_win2115; scan_win2117 <= scan_win2116; scan_win2118 <= scan_win2117; scan_win2119 <= scan_win2118; scan_win2120 <= scan_win2119; scan_win2121 <= scan_win2120; scan_win2122 <= scan_win2121; scan_win2123 <= scan_win2122; scan_win2124 <= scan_win2123; scan_win2125 <= scan_win2124; scan_win2126 <= scan_win2125; scan_win2127 <= scan_win2126; scan_win2128 <= scan_win2127; scan_win2129 <= scan_win2128; scan_win2130 <= scan_win2129; scan_win2131 <= scan_win2130; scan_win2132 <= scan_win2131; scan_win2133 <= scan_win2132; scan_win2134 <= scan_win2133; scan_win2135 <= scan_win2134; scan_win2136 <= scan_win2135; scan_win2137 <= scan_win2136; scan_win2138 <= scan_win2137; scan_win2139 <= scan_win2138; scan_win2140 <= scan_win2139; scan_win2141 <= scan_win2140; scan_win2142 <= scan_win2141; scan_win2143 <= scan_win2142; scan_win2144 <= scan_win2143; scan_win2145 <= scan_win2144; scan_win2146 <= scan_win2145; scan_win2147 <= scan_win2146; scan_win2148 <= scan_win2147; scan_win2149 <= scan_win2148; scan_win2150 <= scan_win2149; scan_win2151 <= scan_win2150; scan_win2152 <= scan_win2151; scan_win2153 <= scan_win2152; scan_win2154 <= scan_win2153; scan_win2155 <= scan_win2154; scan_win2156 <= scan_win2155; scan_win2157 <= scan_win2156; scan_win2158 <= scan_win2157; scan_win2159 <= scan_win2158; scan_win2160 <= scan_win2159; scan_win2161 <= scan_win2160; scan_win2162 <= scan_win2161; scan_win2163 <= scan_win2162; scan_win2164 <= scan_win2163; scan_win2165 <= scan_win2164; scan_win2166 <= scan_win2165; scan_win2167 <= scan_win2166; scan_win2168 <= scan_win2167; scan_win2169 <= scan_win2168; scan_win2170 <= scan_win2169; scan_win2171 <= scan_win2170; scan_win2172 <= scan_win2171; scan_win2173 <= scan_win2172; scan_win2174 <= scan_win2173; scan_win2175 <= scan_win2174; scan_win2176 <= scan_win2175; scan_win2177 <= scan_win2176; scan_win2178 <= scan_win2177; scan_win2179 <= scan_win2178; scan_win2180 <= scan_win2179; scan_win2181 <= scan_win2180; scan_win2182 <= scan_win2181; scan_win2183 <= scan_win2182; scan_win2184 <= scan_win2183; scan_win2185 <= scan_win2184; scan_win2186 <= scan_win2185; scan_win2187 <= scan_win2186; scan_win2188 <= scan_win2187; scan_win2189 <= scan_win2188; scan_win2190 <= scan_win2189; scan_win2191 <= scan_win2190; scan_win2192 <= scan_win2191; scan_win2193 <= scan_win2192; scan_win2194 <= scan_win2193; scan_win2195 <= scan_win2194; scan_win2196 <= scan_win2195; scan_win2197 <= scan_win2196; scan_win2198 <= scan_win2197; scan_win2199 <= scan_win2198; scan_win2200 <= scan_win2199; 
      scan_win2201 <= scan_win2200; scan_win2202 <= scan_win2201; scan_win2203 <= scan_win2202; scan_win2204 <= scan_win2203; scan_win2205 <= scan_win2204; scan_win2206 <= scan_win2205; scan_win2207 <= scan_win2206; scan_win2208 <= scan_win2207; scan_win2209 <= scan_win2208; scan_win2210 <= scan_win2209; scan_win2211 <= scan_win2210; scan_win2212 <= scan_win2211; scan_win2213 <= scan_win2212; scan_win2214 <= scan_win2213; scan_win2215 <= scan_win2214; scan_win2216 <= scan_win2215; scan_win2217 <= scan_win2216; scan_win2218 <= scan_win2217; scan_win2219 <= scan_win2218; scan_win2220 <= scan_win2219; scan_win2221 <= scan_win2220; scan_win2222 <= scan_win2221; scan_win2223 <= scan_win2222; scan_win2224 <= scan_win2223; scan_win2225 <= scan_win2224; scan_win2226 <= scan_win2225; scan_win2227 <= scan_win2226; scan_win2228 <= scan_win2227; scan_win2229 <= scan_win2228; scan_win2230 <= scan_win2229; scan_win2231 <= scan_win2230; scan_win2232 <= scan_win2231; scan_win2233 <= scan_win2232; scan_win2234 <= scan_win2233; scan_win2235 <= scan_win2234; scan_win2236 <= scan_win2235; scan_win2237 <= scan_win2236; scan_win2238 <= scan_win2237; scan_win2239 <= scan_win2238; scan_win2240 <= scan_win2239; scan_win2241 <= scan_win2240; scan_win2242 <= scan_win2241; scan_win2243 <= scan_win2242; scan_win2244 <= scan_win2243; scan_win2245 <= scan_win2244; scan_win2246 <= scan_win2245; scan_win2247 <= scan_win2246; scan_win2248 <= scan_win2247; scan_win2249 <= scan_win2248; scan_win2250 <= scan_win2249; scan_win2251 <= scan_win2250; scan_win2252 <= scan_win2251; scan_win2253 <= scan_win2252; scan_win2254 <= scan_win2253; scan_win2255 <= scan_win2254; scan_win2256 <= scan_win2255; scan_win2257 <= scan_win2256; scan_win2258 <= scan_win2257; scan_win2259 <= scan_win2258; scan_win2260 <= scan_win2259; scan_win2261 <= scan_win2260; scan_win2262 <= scan_win2261; scan_win2263 <= scan_win2262; scan_win2264 <= scan_win2263; scan_win2265 <= scan_win2264; scan_win2266 <= scan_win2265; scan_win2267 <= scan_win2266; scan_win2268 <= scan_win2267; scan_win2269 <= scan_win2268; scan_win2270 <= scan_win2269; scan_win2271 <= scan_win2270; scan_win2272 <= scan_win2271; scan_win2273 <= scan_win2272; scan_win2274 <= scan_win2273; scan_win2275 <= scan_win2274; scan_win2276 <= scan_win2275; scan_win2277 <= scan_win2276; scan_win2278 <= scan_win2277; scan_win2279 <= scan_win2278; scan_win2280 <= scan_win2279; scan_win2281 <= scan_win2280; scan_win2282 <= scan_win2281; scan_win2283 <= scan_win2282; scan_win2284 <= scan_win2283; scan_win2285 <= scan_win2284; scan_win2286 <= scan_win2285; scan_win2287 <= scan_win2286; scan_win2288 <= scan_win2287; scan_win2289 <= scan_win2288; scan_win2290 <= scan_win2289; scan_win2291 <= scan_win2290; scan_win2292 <= scan_win2291; scan_win2293 <= scan_win2292; scan_win2294 <= scan_win2293; scan_win2295 <= scan_win2294; scan_win2296 <= scan_win2295; scan_win2297 <= scan_win2296; scan_win2298 <= scan_win2297; scan_win2299 <= scan_win2298; scan_win2300 <= scan_win2299; scan_win2301 <= scan_win2300; scan_win2302 <= scan_win2301; scan_win2303 <= scan_win2302; scan_win2304 <= scan_win2303; scan_win2305 <= scan_win2304; scan_win2306 <= scan_win2305; scan_win2307 <= scan_win2306; scan_win2308 <= scan_win2307; scan_win2309 <= scan_win2308; scan_win2310 <= scan_win2309; scan_win2311 <= scan_win2310; scan_win2312 <= scan_win2311; scan_win2313 <= scan_win2312; scan_win2314 <= scan_win2313; scan_win2315 <= scan_win2314; scan_win2316 <= scan_win2315; scan_win2317 <= scan_win2316; scan_win2318 <= scan_win2317; scan_win2319 <= scan_win2318; scan_win2320 <= scan_win2319; scan_win2321 <= scan_win2320; scan_win2322 <= scan_win2321; scan_win2323 <= scan_win2322; scan_win2324 <= scan_win2323; scan_win2325 <= scan_win2324; scan_win2326 <= scan_win2325; scan_win2327 <= scan_win2326; scan_win2328 <= scan_win2327; scan_win2329 <= scan_win2328; scan_win2330 <= scan_win2329; scan_win2331 <= scan_win2330; scan_win2332 <= scan_win2331; scan_win2333 <= scan_win2332; scan_win2334 <= scan_win2333; scan_win2335 <= scan_win2334; scan_win2336 <= scan_win2335; scan_win2337 <= scan_win2336; scan_win2338 <= scan_win2337; scan_win2339 <= scan_win2338; scan_win2340 <= scan_win2339; scan_win2341 <= scan_win2340; scan_win2342 <= scan_win2341; scan_win2343 <= scan_win2342; scan_win2344 <= scan_win2343; scan_win2345 <= scan_win2344; scan_win2346 <= scan_win2345; scan_win2347 <= scan_win2346; scan_win2348 <= scan_win2347; scan_win2349 <= scan_win2348; scan_win2350 <= scan_win2349; scan_win2351 <= scan_win2350; scan_win2352 <= scan_win2351; scan_win2353 <= scan_win2352; scan_win2354 <= scan_win2353; scan_win2355 <= scan_win2354; scan_win2356 <= scan_win2355; scan_win2357 <= scan_win2356; scan_win2358 <= scan_win2357; scan_win2359 <= scan_win2358; scan_win2360 <= scan_win2359; scan_win2361 <= scan_win2360; scan_win2362 <= scan_win2361; scan_win2363 <= scan_win2362; scan_win2364 <= scan_win2363; scan_win2365 <= scan_win2364; scan_win2366 <= scan_win2365; scan_win2367 <= scan_win2366; scan_win2368 <= scan_win2367; scan_win2369 <= scan_win2368; scan_win2370 <= scan_win2369; scan_win2371 <= scan_win2370; scan_win2372 <= scan_win2371; scan_win2373 <= scan_win2372; scan_win2374 <= scan_win2373; scan_win2375 <= scan_win2374; scan_win2376 <= scan_win2375; scan_win2377 <= scan_win2376; scan_win2378 <= scan_win2377; scan_win2379 <= scan_win2378; scan_win2380 <= scan_win2379; scan_win2381 <= scan_win2380; scan_win2382 <= scan_win2381; scan_win2383 <= scan_win2382; scan_win2384 <= scan_win2383; scan_win2385 <= scan_win2384; scan_win2386 <= scan_win2385; scan_win2387 <= scan_win2386; scan_win2388 <= scan_win2387; scan_win2389 <= scan_win2388; scan_win2390 <= scan_win2389; scan_win2391 <= scan_win2390; scan_win2392 <= scan_win2391; scan_win2393 <= scan_win2392; scan_win2394 <= scan_win2393; scan_win2395 <= scan_win2394; scan_win2396 <= scan_win2395; scan_win2397 <= scan_win2396; scan_win2398 <= scan_win2397; scan_win2399 <= scan_win2398; scan_win2400 <= scan_win2399; 
      scan_win2401 <= scan_win2400; scan_win2402 <= scan_win2401; scan_win2403 <= scan_win2402; scan_win2404 <= scan_win2403; scan_win2405 <= scan_win2404; scan_win2406 <= scan_win2405; scan_win2407 <= scan_win2406; scan_win2408 <= scan_win2407; scan_win2409 <= scan_win2408; scan_win2410 <= scan_win2409; scan_win2411 <= scan_win2410; scan_win2412 <= scan_win2411; scan_win2413 <= scan_win2412; scan_win2414 <= scan_win2413; scan_win2415 <= scan_win2414; scan_win2416 <= scan_win2415; scan_win2417 <= scan_win2416; scan_win2418 <= scan_win2417; scan_win2419 <= scan_win2418; scan_win2420 <= scan_win2419; scan_win2421 <= scan_win2420; scan_win2422 <= scan_win2421; scan_win2423 <= scan_win2422; scan_win2424 <= scan_win2423; scan_win2425 <= scan_win2424; scan_win2426 <= scan_win2425; scan_win2427 <= scan_win2426; scan_win2428 <= scan_win2427; scan_win2429 <= scan_win2428; scan_win2430 <= scan_win2429; scan_win2431 <= scan_win2430; scan_win2432 <= scan_win2431; scan_win2433 <= scan_win2432; scan_win2434 <= scan_win2433; scan_win2435 <= scan_win2434; scan_win2436 <= scan_win2435; scan_win2437 <= scan_win2436; scan_win2438 <= scan_win2437; scan_win2439 <= scan_win2438; scan_win2440 <= scan_win2439; scan_win2441 <= scan_win2440; scan_win2442 <= scan_win2441; scan_win2443 <= scan_win2442; scan_win2444 <= scan_win2443; scan_win2445 <= scan_win2444; scan_win2446 <= scan_win2445; scan_win2447 <= scan_win2446; scan_win2448 <= scan_win2447; scan_win2449 <= scan_win2448; scan_win2450 <= scan_win2449; scan_win2451 <= scan_win2450; scan_win2452 <= scan_win2451; scan_win2453 <= scan_win2452; scan_win2454 <= scan_win2453; scan_win2455 <= scan_win2454; scan_win2456 <= scan_win2455; scan_win2457 <= scan_win2456; scan_win2458 <= scan_win2457; scan_win2459 <= scan_win2458; scan_win2460 <= scan_win2459; scan_win2461 <= scan_win2460; scan_win2462 <= scan_win2461; scan_win2463 <= scan_win2462; scan_win2464 <= scan_win2463; scan_win2465 <= scan_win2464; scan_win2466 <= scan_win2465; scan_win2467 <= scan_win2466; scan_win2468 <= scan_win2467; scan_win2469 <= scan_win2468; scan_win2470 <= scan_win2469; scan_win2471 <= scan_win2470; scan_win2472 <= scan_win2471; scan_win2473 <= scan_win2472; scan_win2474 <= scan_win2473; scan_win2475 <= scan_win2474; scan_win2476 <= scan_win2475; scan_win2477 <= scan_win2476; scan_win2478 <= scan_win2477; scan_win2479 <= scan_win2478; scan_win2480 <= scan_win2479; scan_win2481 <= scan_win2480; scan_win2482 <= scan_win2481; scan_win2483 <= scan_win2482; scan_win2484 <= scan_win2483; scan_win2485 <= scan_win2484; scan_win2486 <= scan_win2485; scan_win2487 <= scan_win2486; scan_win2488 <= scan_win2487; scan_win2489 <= scan_win2488; scan_win2490 <= scan_win2489; scan_win2491 <= scan_win2490; scan_win2492 <= scan_win2491; scan_win2493 <= scan_win2492; scan_win2494 <= scan_win2493; scan_win2495 <= scan_win2494; scan_win2496 <= scan_win2495; scan_win2497 <= scan_win2496; scan_win2498 <= scan_win2497; scan_win2499 <= scan_win2498; scan_win2500 <= scan_win2499; scan_win2501 <= scan_win2500; scan_win2502 <= scan_win2501; scan_win2503 <= scan_win2502; scan_win2504 <= scan_win2503; scan_win2505 <= scan_win2504; scan_win2506 <= scan_win2505; scan_win2507 <= scan_win2506; scan_win2508 <= scan_win2507; scan_win2509 <= scan_win2508; scan_win2510 <= scan_win2509; scan_win2511 <= scan_win2510; scan_win2512 <= scan_win2511; scan_win2513 <= scan_win2512; scan_win2514 <= scan_win2513; scan_win2515 <= scan_win2514; scan_win2516 <= scan_win2515; scan_win2517 <= scan_win2516; scan_win2518 <= scan_win2517; scan_win2519 <= scan_win2518; scan_win2520 <= scan_win2519; scan_win2521 <= scan_win2520; scan_win2522 <= scan_win2521; scan_win2523 <= scan_win2522; scan_win2524 <= scan_win2523; scan_win2525 <= scan_win2524; scan_win2526 <= scan_win2525; scan_win2527 <= scan_win2526; scan_win2528 <= scan_win2527; scan_win2529 <= scan_win2528; scan_win2530 <= scan_win2529; scan_win2531 <= scan_win2530; scan_win2532 <= scan_win2531; scan_win2533 <= scan_win2532; scan_win2534 <= scan_win2533; scan_win2535 <= scan_win2534; scan_win2536 <= scan_win2535; scan_win2537 <= scan_win2536; scan_win2538 <= scan_win2537; scan_win2539 <= scan_win2538; scan_win2540 <= scan_win2539; scan_win2541 <= scan_win2540; scan_win2542 <= scan_win2541; scan_win2543 <= scan_win2542; scan_win2544 <= scan_win2543; scan_win2545 <= scan_win2544; scan_win2546 <= scan_win2545; scan_win2547 <= scan_win2546; scan_win2548 <= scan_win2547; scan_win2549 <= scan_win2548; scan_win2550 <= scan_win2549; scan_win2551 <= scan_win2550; scan_win2552 <= scan_win2551; scan_win2553 <= scan_win2552; scan_win2554 <= scan_win2553; scan_win2555 <= scan_win2554; scan_win2556 <= scan_win2555; scan_win2557 <= scan_win2556; scan_win2558 <= scan_win2557; scan_win2559 <= scan_win2558; scan_win2560 <= scan_win2559; scan_win2561 <= scan_win2560; scan_win2562 <= scan_win2561; scan_win2563 <= scan_win2562; scan_win2564 <= scan_win2563; scan_win2565 <= scan_win2564; scan_win2566 <= scan_win2565; scan_win2567 <= scan_win2566; scan_win2568 <= scan_win2567; scan_win2569 <= scan_win2568; scan_win2570 <= scan_win2569; scan_win2571 <= scan_win2570; scan_win2572 <= scan_win2571; scan_win2573 <= scan_win2572; scan_win2574 <= scan_win2573; scan_win2575 <= scan_win2574; scan_win2576 <= scan_win2575; scan_win2577 <= scan_win2576; scan_win2578 <= scan_win2577; scan_win2579 <= scan_win2578; scan_win2580 <= scan_win2579; scan_win2581 <= scan_win2580; scan_win2582 <= scan_win2581; scan_win2583 <= scan_win2582; scan_win2584 <= scan_win2583; scan_win2585 <= scan_win2584; scan_win2586 <= scan_win2585; scan_win2587 <= scan_win2586; scan_win2588 <= scan_win2587; scan_win2589 <= scan_win2588; scan_win2590 <= scan_win2589; scan_win2591 <= scan_win2590; scan_win2592 <= scan_win2591; scan_win2593 <= scan_win2592; scan_win2594 <= scan_win2593; scan_win2595 <= scan_win2594; scan_win2596 <= scan_win2595; scan_win2597 <= scan_win2596; scan_win2598 <= scan_win2597; scan_win2599 <= scan_win2598; scan_win2600 <= scan_win2599; 
      scan_win2601 <= scan_win2600; scan_win2602 <= scan_win2601; scan_win2603 <= scan_win2602; scan_win2604 <= scan_win2603; scan_win2605 <= scan_win2604; scan_win2606 <= scan_win2605; scan_win2607 <= scan_win2606; scan_win2608 <= scan_win2607; scan_win2609 <= scan_win2608; scan_win2610 <= scan_win2609; scan_win2611 <= scan_win2610; scan_win2612 <= scan_win2611; scan_win2613 <= scan_win2612; scan_win2614 <= scan_win2613; scan_win2615 <= scan_win2614; scan_win2616 <= scan_win2615; scan_win2617 <= scan_win2616; scan_win2618 <= scan_win2617; scan_win2619 <= scan_win2618; scan_win2620 <= scan_win2619; scan_win2621 <= scan_win2620; scan_win2622 <= scan_win2621; scan_win2623 <= scan_win2622; scan_win2624 <= scan_win2623; scan_win2625 <= scan_win2624; scan_win2626 <= scan_win2625; scan_win2627 <= scan_win2626; scan_win2628 <= scan_win2627; scan_win2629 <= scan_win2628; scan_win2630 <= scan_win2629; scan_win2631 <= scan_win2630; scan_win2632 <= scan_win2631; scan_win2633 <= scan_win2632; scan_win2634 <= scan_win2633; scan_win2635 <= scan_win2634; scan_win2636 <= scan_win2635; scan_win2637 <= scan_win2636; scan_win2638 <= scan_win2637; scan_win2639 <= scan_win2638; scan_win2640 <= scan_win2639; scan_win2641 <= scan_win2640; scan_win2642 <= scan_win2641; scan_win2643 <= scan_win2642; scan_win2644 <= scan_win2643; scan_win2645 <= scan_win2644; scan_win2646 <= scan_win2645; scan_win2647 <= scan_win2646; scan_win2648 <= scan_win2647; scan_win2649 <= scan_win2648; scan_win2650 <= scan_win2649; scan_win2651 <= scan_win2650; scan_win2652 <= scan_win2651; scan_win2653 <= scan_win2652; scan_win2654 <= scan_win2653; scan_win2655 <= scan_win2654; scan_win2656 <= scan_win2655; scan_win2657 <= scan_win2656; scan_win2658 <= scan_win2657; scan_win2659 <= scan_win2658; scan_win2660 <= scan_win2659; scan_win2661 <= scan_win2660; scan_win2662 <= scan_win2661; scan_win2663 <= scan_win2662; scan_win2664 <= scan_win2663; scan_win2665 <= scan_win2664; scan_win2666 <= scan_win2665; scan_win2667 <= scan_win2666; scan_win2668 <= scan_win2667; scan_win2669 <= scan_win2668; scan_win2670 <= scan_win2669; scan_win2671 <= scan_win2670; scan_win2672 <= scan_win2671; scan_win2673 <= scan_win2672; scan_win2674 <= scan_win2673; scan_win2675 <= scan_win2674; scan_win2676 <= scan_win2675; scan_win2677 <= scan_win2676; scan_win2678 <= scan_win2677; scan_win2679 <= scan_win2678; scan_win2680 <= scan_win2679; scan_win2681 <= scan_win2680; scan_win2682 <= scan_win2681; scan_win2683 <= scan_win2682; scan_win2684 <= scan_win2683; scan_win2685 <= scan_win2684; scan_win2686 <= scan_win2685; scan_win2687 <= scan_win2686; scan_win2688 <= scan_win2687; scan_win2689 <= scan_win2688; scan_win2690 <= scan_win2689; scan_win2691 <= scan_win2690; scan_win2692 <= scan_win2691; scan_win2693 <= scan_win2692; scan_win2694 <= scan_win2693; scan_win2695 <= scan_win2694; scan_win2696 <= scan_win2695; scan_win2697 <= scan_win2696; scan_win2698 <= scan_win2697; scan_win2699 <= scan_win2698; scan_win2700 <= scan_win2699; scan_win2701 <= scan_win2700; scan_win2702 <= scan_win2701; scan_win2703 <= scan_win2702; scan_win2704 <= scan_win2703; scan_win2705 <= scan_win2704; scan_win2706 <= scan_win2705; scan_win2707 <= scan_win2706; scan_win2708 <= scan_win2707; scan_win2709 <= scan_win2708; scan_win2710 <= scan_win2709; scan_win2711 <= scan_win2710; scan_win2712 <= scan_win2711; scan_win2713 <= scan_win2712; scan_win2714 <= scan_win2713; scan_win2715 <= scan_win2714; scan_win2716 <= scan_win2715; scan_win2717 <= scan_win2716; scan_win2718 <= scan_win2717; scan_win2719 <= scan_win2718; scan_win2720 <= scan_win2719; scan_win2721 <= scan_win2720; scan_win2722 <= scan_win2721; scan_win2723 <= scan_win2722; scan_win2724 <= scan_win2723; scan_win2725 <= scan_win2724; scan_win2726 <= scan_win2725; scan_win2727 <= scan_win2726; scan_win2728 <= scan_win2727; scan_win2729 <= scan_win2728; scan_win2730 <= scan_win2729; scan_win2731 <= scan_win2730; scan_win2732 <= scan_win2731; scan_win2733 <= scan_win2732; scan_win2734 <= scan_win2733; scan_win2735 <= scan_win2734; scan_win2736 <= scan_win2735; scan_win2737 <= scan_win2736; scan_win2738 <= scan_win2737; scan_win2739 <= scan_win2738; scan_win2740 <= scan_win2739; scan_win2741 <= scan_win2740; scan_win2742 <= scan_win2741; scan_win2743 <= scan_win2742; scan_win2744 <= scan_win2743; scan_win2745 <= scan_win2744; scan_win2746 <= scan_win2745; scan_win2747 <= scan_win2746; scan_win2748 <= scan_win2747; scan_win2749 <= scan_win2748; scan_win2750 <= scan_win2749; scan_win2751 <= scan_win2750; scan_win2752 <= scan_win2751; scan_win2753 <= scan_win2752; scan_win2754 <= scan_win2753; scan_win2755 <= scan_win2754; scan_win2756 <= scan_win2755; scan_win2757 <= scan_win2756; scan_win2758 <= scan_win2757; scan_win2759 <= scan_win2758; scan_win2760 <= scan_win2759; scan_win2761 <= scan_win2760; scan_win2762 <= scan_win2761; scan_win2763 <= scan_win2762; scan_win2764 <= scan_win2763; scan_win2765 <= scan_win2764; scan_win2766 <= scan_win2765; scan_win2767 <= scan_win2766; scan_win2768 <= scan_win2767; scan_win2769 <= scan_win2768; scan_win2770 <= scan_win2769; scan_win2771 <= scan_win2770; scan_win2772 <= scan_win2771; scan_win2773 <= scan_win2772; scan_win2774 <= scan_win2773; scan_win2775 <= scan_win2774; scan_win2776 <= scan_win2775; scan_win2777 <= scan_win2776; scan_win2778 <= scan_win2777; scan_win2779 <= scan_win2778; scan_win2780 <= scan_win2779; scan_win2781 <= scan_win2780; scan_win2782 <= scan_win2781; scan_win2783 <= scan_win2782; scan_win2784 <= scan_win2783; scan_win2785 <= scan_win2784; scan_win2786 <= scan_win2785; scan_win2787 <= scan_win2786; scan_win2788 <= scan_win2787; scan_win2789 <= scan_win2788; scan_win2790 <= scan_win2789; scan_win2791 <= scan_win2790; scan_win2792 <= scan_win2791; scan_win2793 <= scan_win2792; scan_win2794 <= scan_win2793; scan_win2795 <= scan_win2794; scan_win2796 <= scan_win2795; scan_win2797 <= scan_win2796; scan_win2798 <= scan_win2797; scan_win2799 <= scan_win2798; scan_win2800 <= scan_win2799; 
      scan_win2801 <= scan_win2800; scan_win2802 <= scan_win2801; scan_win2803 <= scan_win2802; scan_win2804 <= scan_win2803; scan_win2805 <= scan_win2804; scan_win2806 <= scan_win2805; scan_win2807 <= scan_win2806; scan_win2808 <= scan_win2807; scan_win2809 <= scan_win2808; scan_win2810 <= scan_win2809; scan_win2811 <= scan_win2810; scan_win2812 <= scan_win2811; scan_win2813 <= scan_win2812; scan_win2814 <= scan_win2813; scan_win2815 <= scan_win2814; scan_win2816 <= scan_win2815; scan_win2817 <= scan_win2816; scan_win2818 <= scan_win2817; scan_win2819 <= scan_win2818; scan_win2820 <= scan_win2819; scan_win2821 <= scan_win2820; scan_win2822 <= scan_win2821; scan_win2823 <= scan_win2822; scan_win2824 <= scan_win2823; scan_win2825 <= scan_win2824; scan_win2826 <= scan_win2825; scan_win2827 <= scan_win2826; scan_win2828 <= scan_win2827; scan_win2829 <= scan_win2828; scan_win2830 <= scan_win2829; scan_win2831 <= scan_win2830; scan_win2832 <= scan_win2831; scan_win2833 <= scan_win2832; scan_win2834 <= scan_win2833; scan_win2835 <= scan_win2834; scan_win2836 <= scan_win2835; scan_win2837 <= scan_win2836; scan_win2838 <= scan_win2837; scan_win2839 <= scan_win2838; scan_win2840 <= scan_win2839; scan_win2841 <= scan_win2840; scan_win2842 <= scan_win2841; scan_win2843 <= scan_win2842; scan_win2844 <= scan_win2843; scan_win2845 <= scan_win2844; scan_win2846 <= scan_win2845; scan_win2847 <= scan_win2846; scan_win2848 <= scan_win2847; scan_win2849 <= scan_win2848; scan_win2850 <= scan_win2849; scan_win2851 <= scan_win2850; scan_win2852 <= scan_win2851; scan_win2853 <= scan_win2852; scan_win2854 <= scan_win2853; scan_win2855 <= scan_win2854; scan_win2856 <= scan_win2855; scan_win2857 <= scan_win2856; scan_win2858 <= scan_win2857; scan_win2859 <= scan_win2858; scan_win2860 <= scan_win2859; scan_win2861 <= scan_win2860; scan_win2862 <= scan_win2861; scan_win2863 <= scan_win2862; scan_win2864 <= scan_win2863; scan_win2865 <= scan_win2864; scan_win2866 <= scan_win2865; scan_win2867 <= scan_win2866; scan_win2868 <= scan_win2867; scan_win2869 <= scan_win2868; scan_win2870 <= scan_win2869; scan_win2871 <= scan_win2870; scan_win2872 <= scan_win2871; scan_win2873 <= scan_win2872; scan_win2874 <= scan_win2873; scan_win2875 <= scan_win2874; scan_win2876 <= scan_win2875; scan_win2877 <= scan_win2876; scan_win2878 <= scan_win2877; scan_win2879 <= scan_win2878; scan_win2880 <= scan_win2879; scan_win2881 <= scan_win2880; scan_win2882 <= scan_win2881; scan_win2883 <= scan_win2882; scan_win2884 <= scan_win2883; scan_win2885 <= scan_win2884; scan_win2886 <= scan_win2885; scan_win2887 <= scan_win2886; scan_win2888 <= scan_win2887; scan_win2889 <= scan_win2888; scan_win2890 <= scan_win2889; scan_win2891 <= scan_win2890; scan_win2892 <= scan_win2891; scan_win2893 <= scan_win2892; scan_win2894 <= scan_win2893; scan_win2895 <= scan_win2894; scan_win2896 <= scan_win2895; scan_win2897 <= scan_win2896; scan_win2898 <= scan_win2897; scan_win2899 <= scan_win2898; scan_win2900 <= scan_win2899; scan_win2901 <= scan_win2900; scan_win2902 <= scan_win2901; scan_win2903 <= scan_win2902; scan_win2904 <= scan_win2903; scan_win2905 <= scan_win2904; scan_win2906 <= scan_win2905; scan_win2907 <= scan_win2906; scan_win2908 <= scan_win2907; scan_win2909 <= scan_win2908; scan_win2910 <= scan_win2909; scan_win2911 <= scan_win2910; scan_win2912 <= scan_win2911; 
    end
  end

  accum_calculator ac0(.scan_win(scan_win0), .rectangle1_x(rectangle1_xs[0]), .rectangle1_y(rectangle1_ys[0]), .rectangle1_width(rectangle1_widths[0]), .rectangle1_height(rectangle1_heights[0]), .rectangle1_weight(rectangle1_weights[0]), .rectangle2_x(rectangle2_xs[0]), .rectangle2_y(rectangle2_ys[0]), .rectangle2_width(rectangle2_widths[0]), .rectangle2_height(rectangle2_heights[0]), .rectangle2_weight(rectangle2_weights[0]), .rectangle3_x(rectangle3_xs[0]), .rectangle3_y(rectangle3_ys[0]), .rectangle3_width(rectangle3_widths[0]), .rectangle3_height(rectangle3_heights[0]), .rectangle3_weight(rectangle3_weights[0]), .feature_threshold(feature_thresholds[0]), .feature_above(feature_aboves[0]), .feature_below(feature_belows[0]), .scan_win_std_dev(scan_win_std_dev[0]), .feature_accum(feature_accums[0]));
  accum_calculator ac1(.scan_win(scan_win1), .rectangle1_x(rectangle1_xs[1]), .rectangle1_y(rectangle1_ys[1]), .rectangle1_width(rectangle1_widths[1]), .rectangle1_height(rectangle1_heights[1]), .rectangle1_weight(rectangle1_weights[1]), .rectangle2_x(rectangle2_xs[1]), .rectangle2_y(rectangle2_ys[1]), .rectangle2_width(rectangle2_widths[1]), .rectangle2_height(rectangle2_heights[1]), .rectangle2_weight(rectangle2_weights[1]), .rectangle3_x(rectangle3_xs[1]), .rectangle3_y(rectangle3_ys[1]), .rectangle3_width(rectangle3_widths[1]), .rectangle3_height(rectangle3_heights[1]), .rectangle3_weight(rectangle3_weights[1]), .feature_threshold(feature_thresholds[1]), .feature_above(feature_aboves[1]), .feature_below(feature_belows[1]), .scan_win_std_dev(scan_win_std_dev[1]), .feature_accum(feature_accums[1]));
  accum_calculator ac2(.scan_win(scan_win2), .rectangle1_x(rectangle1_xs[2]), .rectangle1_y(rectangle1_ys[2]), .rectangle1_width(rectangle1_widths[2]), .rectangle1_height(rectangle1_heights[2]), .rectangle1_weight(rectangle1_weights[2]), .rectangle2_x(rectangle2_xs[2]), .rectangle2_y(rectangle2_ys[2]), .rectangle2_width(rectangle2_widths[2]), .rectangle2_height(rectangle2_heights[2]), .rectangle2_weight(rectangle2_weights[2]), .rectangle3_x(rectangle3_xs[2]), .rectangle3_y(rectangle3_ys[2]), .rectangle3_width(rectangle3_widths[2]), .rectangle3_height(rectangle3_heights[2]), .rectangle3_weight(rectangle3_weights[2]), .feature_threshold(feature_thresholds[2]), .feature_above(feature_aboves[2]), .feature_below(feature_belows[2]), .scan_win_std_dev(scan_win_std_dev[2]), .feature_accum(feature_accums[2]));
  accum_calculator ac3(.scan_win(scan_win3), .rectangle1_x(rectangle1_xs[3]), .rectangle1_y(rectangle1_ys[3]), .rectangle1_width(rectangle1_widths[3]), .rectangle1_height(rectangle1_heights[3]), .rectangle1_weight(rectangle1_weights[3]), .rectangle2_x(rectangle2_xs[3]), .rectangle2_y(rectangle2_ys[3]), .rectangle2_width(rectangle2_widths[3]), .rectangle2_height(rectangle2_heights[3]), .rectangle2_weight(rectangle2_weights[3]), .rectangle3_x(rectangle3_xs[3]), .rectangle3_y(rectangle3_ys[3]), .rectangle3_width(rectangle3_widths[3]), .rectangle3_height(rectangle3_heights[3]), .rectangle3_weight(rectangle3_weights[3]), .feature_threshold(feature_thresholds[3]), .feature_above(feature_aboves[3]), .feature_below(feature_belows[3]), .scan_win_std_dev(scan_win_std_dev[3]), .feature_accum(feature_accums[3]));
  accum_calculator ac4(.scan_win(scan_win4), .rectangle1_x(rectangle1_xs[4]), .rectangle1_y(rectangle1_ys[4]), .rectangle1_width(rectangle1_widths[4]), .rectangle1_height(rectangle1_heights[4]), .rectangle1_weight(rectangle1_weights[4]), .rectangle2_x(rectangle2_xs[4]), .rectangle2_y(rectangle2_ys[4]), .rectangle2_width(rectangle2_widths[4]), .rectangle2_height(rectangle2_heights[4]), .rectangle2_weight(rectangle2_weights[4]), .rectangle3_x(rectangle3_xs[4]), .rectangle3_y(rectangle3_ys[4]), .rectangle3_width(rectangle3_widths[4]), .rectangle3_height(rectangle3_heights[4]), .rectangle3_weight(rectangle3_weights[4]), .feature_threshold(feature_thresholds[4]), .feature_above(feature_aboves[4]), .feature_below(feature_belows[4]), .scan_win_std_dev(scan_win_std_dev[4]), .feature_accum(feature_accums[4]));
  accum_calculator ac5(.scan_win(scan_win5), .rectangle1_x(rectangle1_xs[5]), .rectangle1_y(rectangle1_ys[5]), .rectangle1_width(rectangle1_widths[5]), .rectangle1_height(rectangle1_heights[5]), .rectangle1_weight(rectangle1_weights[5]), .rectangle2_x(rectangle2_xs[5]), .rectangle2_y(rectangle2_ys[5]), .rectangle2_width(rectangle2_widths[5]), .rectangle2_height(rectangle2_heights[5]), .rectangle2_weight(rectangle2_weights[5]), .rectangle3_x(rectangle3_xs[5]), .rectangle3_y(rectangle3_ys[5]), .rectangle3_width(rectangle3_widths[5]), .rectangle3_height(rectangle3_heights[5]), .rectangle3_weight(rectangle3_weights[5]), .feature_threshold(feature_thresholds[5]), .feature_above(feature_aboves[5]), .feature_below(feature_belows[5]), .scan_win_std_dev(scan_win_std_dev[5]), .feature_accum(feature_accums[5]));
  accum_calculator ac6(.scan_win(scan_win6), .rectangle1_x(rectangle1_xs[6]), .rectangle1_y(rectangle1_ys[6]), .rectangle1_width(rectangle1_widths[6]), .rectangle1_height(rectangle1_heights[6]), .rectangle1_weight(rectangle1_weights[6]), .rectangle2_x(rectangle2_xs[6]), .rectangle2_y(rectangle2_ys[6]), .rectangle2_width(rectangle2_widths[6]), .rectangle2_height(rectangle2_heights[6]), .rectangle2_weight(rectangle2_weights[6]), .rectangle3_x(rectangle3_xs[6]), .rectangle3_y(rectangle3_ys[6]), .rectangle3_width(rectangle3_widths[6]), .rectangle3_height(rectangle3_heights[6]), .rectangle3_weight(rectangle3_weights[6]), .feature_threshold(feature_thresholds[6]), .feature_above(feature_aboves[6]), .feature_below(feature_belows[6]), .scan_win_std_dev(scan_win_std_dev[6]), .feature_accum(feature_accums[6]));
  accum_calculator ac7(.scan_win(scan_win7), .rectangle1_x(rectangle1_xs[7]), .rectangle1_y(rectangle1_ys[7]), .rectangle1_width(rectangle1_widths[7]), .rectangle1_height(rectangle1_heights[7]), .rectangle1_weight(rectangle1_weights[7]), .rectangle2_x(rectangle2_xs[7]), .rectangle2_y(rectangle2_ys[7]), .rectangle2_width(rectangle2_widths[7]), .rectangle2_height(rectangle2_heights[7]), .rectangle2_weight(rectangle2_weights[7]), .rectangle3_x(rectangle3_xs[7]), .rectangle3_y(rectangle3_ys[7]), .rectangle3_width(rectangle3_widths[7]), .rectangle3_height(rectangle3_heights[7]), .rectangle3_weight(rectangle3_weights[7]), .feature_threshold(feature_thresholds[7]), .feature_above(feature_aboves[7]), .feature_below(feature_belows[7]), .scan_win_std_dev(scan_win_std_dev[7]), .feature_accum(feature_accums[7]));
  accum_calculator ac8(.scan_win(scan_win8), .rectangle1_x(rectangle1_xs[8]), .rectangle1_y(rectangle1_ys[8]), .rectangle1_width(rectangle1_widths[8]), .rectangle1_height(rectangle1_heights[8]), .rectangle1_weight(rectangle1_weights[8]), .rectangle2_x(rectangle2_xs[8]), .rectangle2_y(rectangle2_ys[8]), .rectangle2_width(rectangle2_widths[8]), .rectangle2_height(rectangle2_heights[8]), .rectangle2_weight(rectangle2_weights[8]), .rectangle3_x(rectangle3_xs[8]), .rectangle3_y(rectangle3_ys[8]), .rectangle3_width(rectangle3_widths[8]), .rectangle3_height(rectangle3_heights[8]), .rectangle3_weight(rectangle3_weights[8]), .feature_threshold(feature_thresholds[8]), .feature_above(feature_aboves[8]), .feature_below(feature_belows[8]), .scan_win_std_dev(scan_win_std_dev[8]), .feature_accum(feature_accums[8]));
  accum_calculator ac9(.scan_win(scan_win9), .rectangle1_x(rectangle1_xs[9]), .rectangle1_y(rectangle1_ys[9]), .rectangle1_width(rectangle1_widths[9]), .rectangle1_height(rectangle1_heights[9]), .rectangle1_weight(rectangle1_weights[9]), .rectangle2_x(rectangle2_xs[9]), .rectangle2_y(rectangle2_ys[9]), .rectangle2_width(rectangle2_widths[9]), .rectangle2_height(rectangle2_heights[9]), .rectangle2_weight(rectangle2_weights[9]), .rectangle3_x(rectangle3_xs[9]), .rectangle3_y(rectangle3_ys[9]), .rectangle3_width(rectangle3_widths[9]), .rectangle3_height(rectangle3_heights[9]), .rectangle3_weight(rectangle3_weights[9]), .feature_threshold(feature_thresholds[9]), .feature_above(feature_aboves[9]), .feature_below(feature_belows[9]), .scan_win_std_dev(scan_win_std_dev[9]), .feature_accum(feature_accums[9]));
  accum_calculator ac10(.scan_win(scan_win10), .rectangle1_x(rectangle1_xs[10]), .rectangle1_y(rectangle1_ys[10]), .rectangle1_width(rectangle1_widths[10]), .rectangle1_height(rectangle1_heights[10]), .rectangle1_weight(rectangle1_weights[10]), .rectangle2_x(rectangle2_xs[10]), .rectangle2_y(rectangle2_ys[10]), .rectangle2_width(rectangle2_widths[10]), .rectangle2_height(rectangle2_heights[10]), .rectangle2_weight(rectangle2_weights[10]), .rectangle3_x(rectangle3_xs[10]), .rectangle3_y(rectangle3_ys[10]), .rectangle3_width(rectangle3_widths[10]), .rectangle3_height(rectangle3_heights[10]), .rectangle3_weight(rectangle3_weights[10]), .feature_threshold(feature_thresholds[10]), .feature_above(feature_aboves[10]), .feature_below(feature_belows[10]), .scan_win_std_dev(scan_win_std_dev[10]), .feature_accum(feature_accums[10]));
  accum_calculator ac11(.scan_win(scan_win11), .rectangle1_x(rectangle1_xs[11]), .rectangle1_y(rectangle1_ys[11]), .rectangle1_width(rectangle1_widths[11]), .rectangle1_height(rectangle1_heights[11]), .rectangle1_weight(rectangle1_weights[11]), .rectangle2_x(rectangle2_xs[11]), .rectangle2_y(rectangle2_ys[11]), .rectangle2_width(rectangle2_widths[11]), .rectangle2_height(rectangle2_heights[11]), .rectangle2_weight(rectangle2_weights[11]), .rectangle3_x(rectangle3_xs[11]), .rectangle3_y(rectangle3_ys[11]), .rectangle3_width(rectangle3_widths[11]), .rectangle3_height(rectangle3_heights[11]), .rectangle3_weight(rectangle3_weights[11]), .feature_threshold(feature_thresholds[11]), .feature_above(feature_aboves[11]), .feature_below(feature_belows[11]), .scan_win_std_dev(scan_win_std_dev[11]), .feature_accum(feature_accums[11]));
  accum_calculator ac12(.scan_win(scan_win12), .rectangle1_x(rectangle1_xs[12]), .rectangle1_y(rectangle1_ys[12]), .rectangle1_width(rectangle1_widths[12]), .rectangle1_height(rectangle1_heights[12]), .rectangle1_weight(rectangle1_weights[12]), .rectangle2_x(rectangle2_xs[12]), .rectangle2_y(rectangle2_ys[12]), .rectangle2_width(rectangle2_widths[12]), .rectangle2_height(rectangle2_heights[12]), .rectangle2_weight(rectangle2_weights[12]), .rectangle3_x(rectangle3_xs[12]), .rectangle3_y(rectangle3_ys[12]), .rectangle3_width(rectangle3_widths[12]), .rectangle3_height(rectangle3_heights[12]), .rectangle3_weight(rectangle3_weights[12]), .feature_threshold(feature_thresholds[12]), .feature_above(feature_aboves[12]), .feature_below(feature_belows[12]), .scan_win_std_dev(scan_win_std_dev[12]), .feature_accum(feature_accums[12]));
  accum_calculator ac13(.scan_win(scan_win13), .rectangle1_x(rectangle1_xs[13]), .rectangle1_y(rectangle1_ys[13]), .rectangle1_width(rectangle1_widths[13]), .rectangle1_height(rectangle1_heights[13]), .rectangle1_weight(rectangle1_weights[13]), .rectangle2_x(rectangle2_xs[13]), .rectangle2_y(rectangle2_ys[13]), .rectangle2_width(rectangle2_widths[13]), .rectangle2_height(rectangle2_heights[13]), .rectangle2_weight(rectangle2_weights[13]), .rectangle3_x(rectangle3_xs[13]), .rectangle3_y(rectangle3_ys[13]), .rectangle3_width(rectangle3_widths[13]), .rectangle3_height(rectangle3_heights[13]), .rectangle3_weight(rectangle3_weights[13]), .feature_threshold(feature_thresholds[13]), .feature_above(feature_aboves[13]), .feature_below(feature_belows[13]), .scan_win_std_dev(scan_win_std_dev[13]), .feature_accum(feature_accums[13]));
  accum_calculator ac14(.scan_win(scan_win14), .rectangle1_x(rectangle1_xs[14]), .rectangle1_y(rectangle1_ys[14]), .rectangle1_width(rectangle1_widths[14]), .rectangle1_height(rectangle1_heights[14]), .rectangle1_weight(rectangle1_weights[14]), .rectangle2_x(rectangle2_xs[14]), .rectangle2_y(rectangle2_ys[14]), .rectangle2_width(rectangle2_widths[14]), .rectangle2_height(rectangle2_heights[14]), .rectangle2_weight(rectangle2_weights[14]), .rectangle3_x(rectangle3_xs[14]), .rectangle3_y(rectangle3_ys[14]), .rectangle3_width(rectangle3_widths[14]), .rectangle3_height(rectangle3_heights[14]), .rectangle3_weight(rectangle3_weights[14]), .feature_threshold(feature_thresholds[14]), .feature_above(feature_aboves[14]), .feature_below(feature_belows[14]), .scan_win_std_dev(scan_win_std_dev[14]), .feature_accum(feature_accums[14]));
  accum_calculator ac15(.scan_win(scan_win15), .rectangle1_x(rectangle1_xs[15]), .rectangle1_y(rectangle1_ys[15]), .rectangle1_width(rectangle1_widths[15]), .rectangle1_height(rectangle1_heights[15]), .rectangle1_weight(rectangle1_weights[15]), .rectangle2_x(rectangle2_xs[15]), .rectangle2_y(rectangle2_ys[15]), .rectangle2_width(rectangle2_widths[15]), .rectangle2_height(rectangle2_heights[15]), .rectangle2_weight(rectangle2_weights[15]), .rectangle3_x(rectangle3_xs[15]), .rectangle3_y(rectangle3_ys[15]), .rectangle3_width(rectangle3_widths[15]), .rectangle3_height(rectangle3_heights[15]), .rectangle3_weight(rectangle3_weights[15]), .feature_threshold(feature_thresholds[15]), .feature_above(feature_aboves[15]), .feature_below(feature_belows[15]), .scan_win_std_dev(scan_win_std_dev[15]), .feature_accum(feature_accums[15]));
  accum_calculator ac16(.scan_win(scan_win16), .rectangle1_x(rectangle1_xs[16]), .rectangle1_y(rectangle1_ys[16]), .rectangle1_width(rectangle1_widths[16]), .rectangle1_height(rectangle1_heights[16]), .rectangle1_weight(rectangle1_weights[16]), .rectangle2_x(rectangle2_xs[16]), .rectangle2_y(rectangle2_ys[16]), .rectangle2_width(rectangle2_widths[16]), .rectangle2_height(rectangle2_heights[16]), .rectangle2_weight(rectangle2_weights[16]), .rectangle3_x(rectangle3_xs[16]), .rectangle3_y(rectangle3_ys[16]), .rectangle3_width(rectangle3_widths[16]), .rectangle3_height(rectangle3_heights[16]), .rectangle3_weight(rectangle3_weights[16]), .feature_threshold(feature_thresholds[16]), .feature_above(feature_aboves[16]), .feature_below(feature_belows[16]), .scan_win_std_dev(scan_win_std_dev[16]), .feature_accum(feature_accums[16]));
  accum_calculator ac17(.scan_win(scan_win17), .rectangle1_x(rectangle1_xs[17]), .rectangle1_y(rectangle1_ys[17]), .rectangle1_width(rectangle1_widths[17]), .rectangle1_height(rectangle1_heights[17]), .rectangle1_weight(rectangle1_weights[17]), .rectangle2_x(rectangle2_xs[17]), .rectangle2_y(rectangle2_ys[17]), .rectangle2_width(rectangle2_widths[17]), .rectangle2_height(rectangle2_heights[17]), .rectangle2_weight(rectangle2_weights[17]), .rectangle3_x(rectangle3_xs[17]), .rectangle3_y(rectangle3_ys[17]), .rectangle3_width(rectangle3_widths[17]), .rectangle3_height(rectangle3_heights[17]), .rectangle3_weight(rectangle3_weights[17]), .feature_threshold(feature_thresholds[17]), .feature_above(feature_aboves[17]), .feature_below(feature_belows[17]), .scan_win_std_dev(scan_win_std_dev[17]), .feature_accum(feature_accums[17]));
  accum_calculator ac18(.scan_win(scan_win18), .rectangle1_x(rectangle1_xs[18]), .rectangle1_y(rectangle1_ys[18]), .rectangle1_width(rectangle1_widths[18]), .rectangle1_height(rectangle1_heights[18]), .rectangle1_weight(rectangle1_weights[18]), .rectangle2_x(rectangle2_xs[18]), .rectangle2_y(rectangle2_ys[18]), .rectangle2_width(rectangle2_widths[18]), .rectangle2_height(rectangle2_heights[18]), .rectangle2_weight(rectangle2_weights[18]), .rectangle3_x(rectangle3_xs[18]), .rectangle3_y(rectangle3_ys[18]), .rectangle3_width(rectangle3_widths[18]), .rectangle3_height(rectangle3_heights[18]), .rectangle3_weight(rectangle3_weights[18]), .feature_threshold(feature_thresholds[18]), .feature_above(feature_aboves[18]), .feature_below(feature_belows[18]), .scan_win_std_dev(scan_win_std_dev[18]), .feature_accum(feature_accums[18]));
  accum_calculator ac19(.scan_win(scan_win19), .rectangle1_x(rectangle1_xs[19]), .rectangle1_y(rectangle1_ys[19]), .rectangle1_width(rectangle1_widths[19]), .rectangle1_height(rectangle1_heights[19]), .rectangle1_weight(rectangle1_weights[19]), .rectangle2_x(rectangle2_xs[19]), .rectangle2_y(rectangle2_ys[19]), .rectangle2_width(rectangle2_widths[19]), .rectangle2_height(rectangle2_heights[19]), .rectangle2_weight(rectangle2_weights[19]), .rectangle3_x(rectangle3_xs[19]), .rectangle3_y(rectangle3_ys[19]), .rectangle3_width(rectangle3_widths[19]), .rectangle3_height(rectangle3_heights[19]), .rectangle3_weight(rectangle3_weights[19]), .feature_threshold(feature_thresholds[19]), .feature_above(feature_aboves[19]), .feature_below(feature_belows[19]), .scan_win_std_dev(scan_win_std_dev[19]), .feature_accum(feature_accums[19]));
  accum_calculator ac20(.scan_win(scan_win20), .rectangle1_x(rectangle1_xs[20]), .rectangle1_y(rectangle1_ys[20]), .rectangle1_width(rectangle1_widths[20]), .rectangle1_height(rectangle1_heights[20]), .rectangle1_weight(rectangle1_weights[20]), .rectangle2_x(rectangle2_xs[20]), .rectangle2_y(rectangle2_ys[20]), .rectangle2_width(rectangle2_widths[20]), .rectangle2_height(rectangle2_heights[20]), .rectangle2_weight(rectangle2_weights[20]), .rectangle3_x(rectangle3_xs[20]), .rectangle3_y(rectangle3_ys[20]), .rectangle3_width(rectangle3_widths[20]), .rectangle3_height(rectangle3_heights[20]), .rectangle3_weight(rectangle3_weights[20]), .feature_threshold(feature_thresholds[20]), .feature_above(feature_aboves[20]), .feature_below(feature_belows[20]), .scan_win_std_dev(scan_win_std_dev[20]), .feature_accum(feature_accums[20]));
  accum_calculator ac21(.scan_win(scan_win21), .rectangle1_x(rectangle1_xs[21]), .rectangle1_y(rectangle1_ys[21]), .rectangle1_width(rectangle1_widths[21]), .rectangle1_height(rectangle1_heights[21]), .rectangle1_weight(rectangle1_weights[21]), .rectangle2_x(rectangle2_xs[21]), .rectangle2_y(rectangle2_ys[21]), .rectangle2_width(rectangle2_widths[21]), .rectangle2_height(rectangle2_heights[21]), .rectangle2_weight(rectangle2_weights[21]), .rectangle3_x(rectangle3_xs[21]), .rectangle3_y(rectangle3_ys[21]), .rectangle3_width(rectangle3_widths[21]), .rectangle3_height(rectangle3_heights[21]), .rectangle3_weight(rectangle3_weights[21]), .feature_threshold(feature_thresholds[21]), .feature_above(feature_aboves[21]), .feature_below(feature_belows[21]), .scan_win_std_dev(scan_win_std_dev[21]), .feature_accum(feature_accums[21]));
  accum_calculator ac22(.scan_win(scan_win22), .rectangle1_x(rectangle1_xs[22]), .rectangle1_y(rectangle1_ys[22]), .rectangle1_width(rectangle1_widths[22]), .rectangle1_height(rectangle1_heights[22]), .rectangle1_weight(rectangle1_weights[22]), .rectangle2_x(rectangle2_xs[22]), .rectangle2_y(rectangle2_ys[22]), .rectangle2_width(rectangle2_widths[22]), .rectangle2_height(rectangle2_heights[22]), .rectangle2_weight(rectangle2_weights[22]), .rectangle3_x(rectangle3_xs[22]), .rectangle3_y(rectangle3_ys[22]), .rectangle3_width(rectangle3_widths[22]), .rectangle3_height(rectangle3_heights[22]), .rectangle3_weight(rectangle3_weights[22]), .feature_threshold(feature_thresholds[22]), .feature_above(feature_aboves[22]), .feature_below(feature_belows[22]), .scan_win_std_dev(scan_win_std_dev[22]), .feature_accum(feature_accums[22]));
  accum_calculator ac23(.scan_win(scan_win23), .rectangle1_x(rectangle1_xs[23]), .rectangle1_y(rectangle1_ys[23]), .rectangle1_width(rectangle1_widths[23]), .rectangle1_height(rectangle1_heights[23]), .rectangle1_weight(rectangle1_weights[23]), .rectangle2_x(rectangle2_xs[23]), .rectangle2_y(rectangle2_ys[23]), .rectangle2_width(rectangle2_widths[23]), .rectangle2_height(rectangle2_heights[23]), .rectangle2_weight(rectangle2_weights[23]), .rectangle3_x(rectangle3_xs[23]), .rectangle3_y(rectangle3_ys[23]), .rectangle3_width(rectangle3_widths[23]), .rectangle3_height(rectangle3_heights[23]), .rectangle3_weight(rectangle3_weights[23]), .feature_threshold(feature_thresholds[23]), .feature_above(feature_aboves[23]), .feature_below(feature_belows[23]), .scan_win_std_dev(scan_win_std_dev[23]), .feature_accum(feature_accums[23]));
  accum_calculator ac24(.scan_win(scan_win24), .rectangle1_x(rectangle1_xs[24]), .rectangle1_y(rectangle1_ys[24]), .rectangle1_width(rectangle1_widths[24]), .rectangle1_height(rectangle1_heights[24]), .rectangle1_weight(rectangle1_weights[24]), .rectangle2_x(rectangle2_xs[24]), .rectangle2_y(rectangle2_ys[24]), .rectangle2_width(rectangle2_widths[24]), .rectangle2_height(rectangle2_heights[24]), .rectangle2_weight(rectangle2_weights[24]), .rectangle3_x(rectangle3_xs[24]), .rectangle3_y(rectangle3_ys[24]), .rectangle3_width(rectangle3_widths[24]), .rectangle3_height(rectangle3_heights[24]), .rectangle3_weight(rectangle3_weights[24]), .feature_threshold(feature_thresholds[24]), .feature_above(feature_aboves[24]), .feature_below(feature_belows[24]), .scan_win_std_dev(scan_win_std_dev[24]), .feature_accum(feature_accums[24]));
  accum_calculator ac25(.scan_win(scan_win25), .rectangle1_x(rectangle1_xs[25]), .rectangle1_y(rectangle1_ys[25]), .rectangle1_width(rectangle1_widths[25]), .rectangle1_height(rectangle1_heights[25]), .rectangle1_weight(rectangle1_weights[25]), .rectangle2_x(rectangle2_xs[25]), .rectangle2_y(rectangle2_ys[25]), .rectangle2_width(rectangle2_widths[25]), .rectangle2_height(rectangle2_heights[25]), .rectangle2_weight(rectangle2_weights[25]), .rectangle3_x(rectangle3_xs[25]), .rectangle3_y(rectangle3_ys[25]), .rectangle3_width(rectangle3_widths[25]), .rectangle3_height(rectangle3_heights[25]), .rectangle3_weight(rectangle3_weights[25]), .feature_threshold(feature_thresholds[25]), .feature_above(feature_aboves[25]), .feature_below(feature_belows[25]), .scan_win_std_dev(scan_win_std_dev[25]), .feature_accum(feature_accums[25]));
  accum_calculator ac26(.scan_win(scan_win26), .rectangle1_x(rectangle1_xs[26]), .rectangle1_y(rectangle1_ys[26]), .rectangle1_width(rectangle1_widths[26]), .rectangle1_height(rectangle1_heights[26]), .rectangle1_weight(rectangle1_weights[26]), .rectangle2_x(rectangle2_xs[26]), .rectangle2_y(rectangle2_ys[26]), .rectangle2_width(rectangle2_widths[26]), .rectangle2_height(rectangle2_heights[26]), .rectangle2_weight(rectangle2_weights[26]), .rectangle3_x(rectangle3_xs[26]), .rectangle3_y(rectangle3_ys[26]), .rectangle3_width(rectangle3_widths[26]), .rectangle3_height(rectangle3_heights[26]), .rectangle3_weight(rectangle3_weights[26]), .feature_threshold(feature_thresholds[26]), .feature_above(feature_aboves[26]), .feature_below(feature_belows[26]), .scan_win_std_dev(scan_win_std_dev[26]), .feature_accum(feature_accums[26]));
  accum_calculator ac27(.scan_win(scan_win27), .rectangle1_x(rectangle1_xs[27]), .rectangle1_y(rectangle1_ys[27]), .rectangle1_width(rectangle1_widths[27]), .rectangle1_height(rectangle1_heights[27]), .rectangle1_weight(rectangle1_weights[27]), .rectangle2_x(rectangle2_xs[27]), .rectangle2_y(rectangle2_ys[27]), .rectangle2_width(rectangle2_widths[27]), .rectangle2_height(rectangle2_heights[27]), .rectangle2_weight(rectangle2_weights[27]), .rectangle3_x(rectangle3_xs[27]), .rectangle3_y(rectangle3_ys[27]), .rectangle3_width(rectangle3_widths[27]), .rectangle3_height(rectangle3_heights[27]), .rectangle3_weight(rectangle3_weights[27]), .feature_threshold(feature_thresholds[27]), .feature_above(feature_aboves[27]), .feature_below(feature_belows[27]), .scan_win_std_dev(scan_win_std_dev[27]), .feature_accum(feature_accums[27]));
  accum_calculator ac28(.scan_win(scan_win28), .rectangle1_x(rectangle1_xs[28]), .rectangle1_y(rectangle1_ys[28]), .rectangle1_width(rectangle1_widths[28]), .rectangle1_height(rectangle1_heights[28]), .rectangle1_weight(rectangle1_weights[28]), .rectangle2_x(rectangle2_xs[28]), .rectangle2_y(rectangle2_ys[28]), .rectangle2_width(rectangle2_widths[28]), .rectangle2_height(rectangle2_heights[28]), .rectangle2_weight(rectangle2_weights[28]), .rectangle3_x(rectangle3_xs[28]), .rectangle3_y(rectangle3_ys[28]), .rectangle3_width(rectangle3_widths[28]), .rectangle3_height(rectangle3_heights[28]), .rectangle3_weight(rectangle3_weights[28]), .feature_threshold(feature_thresholds[28]), .feature_above(feature_aboves[28]), .feature_below(feature_belows[28]), .scan_win_std_dev(scan_win_std_dev[28]), .feature_accum(feature_accums[28]));
  accum_calculator ac29(.scan_win(scan_win29), .rectangle1_x(rectangle1_xs[29]), .rectangle1_y(rectangle1_ys[29]), .rectangle1_width(rectangle1_widths[29]), .rectangle1_height(rectangle1_heights[29]), .rectangle1_weight(rectangle1_weights[29]), .rectangle2_x(rectangle2_xs[29]), .rectangle2_y(rectangle2_ys[29]), .rectangle2_width(rectangle2_widths[29]), .rectangle2_height(rectangle2_heights[29]), .rectangle2_weight(rectangle2_weights[29]), .rectangle3_x(rectangle3_xs[29]), .rectangle3_y(rectangle3_ys[29]), .rectangle3_width(rectangle3_widths[29]), .rectangle3_height(rectangle3_heights[29]), .rectangle3_weight(rectangle3_weights[29]), .feature_threshold(feature_thresholds[29]), .feature_above(feature_aboves[29]), .feature_below(feature_belows[29]), .scan_win_std_dev(scan_win_std_dev[29]), .feature_accum(feature_accums[29]));
  accum_calculator ac30(.scan_win(scan_win30), .rectangle1_x(rectangle1_xs[30]), .rectangle1_y(rectangle1_ys[30]), .rectangle1_width(rectangle1_widths[30]), .rectangle1_height(rectangle1_heights[30]), .rectangle1_weight(rectangle1_weights[30]), .rectangle2_x(rectangle2_xs[30]), .rectangle2_y(rectangle2_ys[30]), .rectangle2_width(rectangle2_widths[30]), .rectangle2_height(rectangle2_heights[30]), .rectangle2_weight(rectangle2_weights[30]), .rectangle3_x(rectangle3_xs[30]), .rectangle3_y(rectangle3_ys[30]), .rectangle3_width(rectangle3_widths[30]), .rectangle3_height(rectangle3_heights[30]), .rectangle3_weight(rectangle3_weights[30]), .feature_threshold(feature_thresholds[30]), .feature_above(feature_aboves[30]), .feature_below(feature_belows[30]), .scan_win_std_dev(scan_win_std_dev[30]), .feature_accum(feature_accums[30]));
  accum_calculator ac31(.scan_win(scan_win31), .rectangle1_x(rectangle1_xs[31]), .rectangle1_y(rectangle1_ys[31]), .rectangle1_width(rectangle1_widths[31]), .rectangle1_height(rectangle1_heights[31]), .rectangle1_weight(rectangle1_weights[31]), .rectangle2_x(rectangle2_xs[31]), .rectangle2_y(rectangle2_ys[31]), .rectangle2_width(rectangle2_widths[31]), .rectangle2_height(rectangle2_heights[31]), .rectangle2_weight(rectangle2_weights[31]), .rectangle3_x(rectangle3_xs[31]), .rectangle3_y(rectangle3_ys[31]), .rectangle3_width(rectangle3_widths[31]), .rectangle3_height(rectangle3_heights[31]), .rectangle3_weight(rectangle3_weights[31]), .feature_threshold(feature_thresholds[31]), .feature_above(feature_aboves[31]), .feature_below(feature_belows[31]), .scan_win_std_dev(scan_win_std_dev[31]), .feature_accum(feature_accums[31]));
  accum_calculator ac32(.scan_win(scan_win32), .rectangle1_x(rectangle1_xs[32]), .rectangle1_y(rectangle1_ys[32]), .rectangle1_width(rectangle1_widths[32]), .rectangle1_height(rectangle1_heights[32]), .rectangle1_weight(rectangle1_weights[32]), .rectangle2_x(rectangle2_xs[32]), .rectangle2_y(rectangle2_ys[32]), .rectangle2_width(rectangle2_widths[32]), .rectangle2_height(rectangle2_heights[32]), .rectangle2_weight(rectangle2_weights[32]), .rectangle3_x(rectangle3_xs[32]), .rectangle3_y(rectangle3_ys[32]), .rectangle3_width(rectangle3_widths[32]), .rectangle3_height(rectangle3_heights[32]), .rectangle3_weight(rectangle3_weights[32]), .feature_threshold(feature_thresholds[32]), .feature_above(feature_aboves[32]), .feature_below(feature_belows[32]), .scan_win_std_dev(scan_win_std_dev[32]), .feature_accum(feature_accums[32]));
  accum_calculator ac33(.scan_win(scan_win33), .rectangle1_x(rectangle1_xs[33]), .rectangle1_y(rectangle1_ys[33]), .rectangle1_width(rectangle1_widths[33]), .rectangle1_height(rectangle1_heights[33]), .rectangle1_weight(rectangle1_weights[33]), .rectangle2_x(rectangle2_xs[33]), .rectangle2_y(rectangle2_ys[33]), .rectangle2_width(rectangle2_widths[33]), .rectangle2_height(rectangle2_heights[33]), .rectangle2_weight(rectangle2_weights[33]), .rectangle3_x(rectangle3_xs[33]), .rectangle3_y(rectangle3_ys[33]), .rectangle3_width(rectangle3_widths[33]), .rectangle3_height(rectangle3_heights[33]), .rectangle3_weight(rectangle3_weights[33]), .feature_threshold(feature_thresholds[33]), .feature_above(feature_aboves[33]), .feature_below(feature_belows[33]), .scan_win_std_dev(scan_win_std_dev[33]), .feature_accum(feature_accums[33]));
  accum_calculator ac34(.scan_win(scan_win34), .rectangle1_x(rectangle1_xs[34]), .rectangle1_y(rectangle1_ys[34]), .rectangle1_width(rectangle1_widths[34]), .rectangle1_height(rectangle1_heights[34]), .rectangle1_weight(rectangle1_weights[34]), .rectangle2_x(rectangle2_xs[34]), .rectangle2_y(rectangle2_ys[34]), .rectangle2_width(rectangle2_widths[34]), .rectangle2_height(rectangle2_heights[34]), .rectangle2_weight(rectangle2_weights[34]), .rectangle3_x(rectangle3_xs[34]), .rectangle3_y(rectangle3_ys[34]), .rectangle3_width(rectangle3_widths[34]), .rectangle3_height(rectangle3_heights[34]), .rectangle3_weight(rectangle3_weights[34]), .feature_threshold(feature_thresholds[34]), .feature_above(feature_aboves[34]), .feature_below(feature_belows[34]), .scan_win_std_dev(scan_win_std_dev[34]), .feature_accum(feature_accums[34]));
  accum_calculator ac35(.scan_win(scan_win35), .rectangle1_x(rectangle1_xs[35]), .rectangle1_y(rectangle1_ys[35]), .rectangle1_width(rectangle1_widths[35]), .rectangle1_height(rectangle1_heights[35]), .rectangle1_weight(rectangle1_weights[35]), .rectangle2_x(rectangle2_xs[35]), .rectangle2_y(rectangle2_ys[35]), .rectangle2_width(rectangle2_widths[35]), .rectangle2_height(rectangle2_heights[35]), .rectangle2_weight(rectangle2_weights[35]), .rectangle3_x(rectangle3_xs[35]), .rectangle3_y(rectangle3_ys[35]), .rectangle3_width(rectangle3_widths[35]), .rectangle3_height(rectangle3_heights[35]), .rectangle3_weight(rectangle3_weights[35]), .feature_threshold(feature_thresholds[35]), .feature_above(feature_aboves[35]), .feature_below(feature_belows[35]), .scan_win_std_dev(scan_win_std_dev[35]), .feature_accum(feature_accums[35]));
  accum_calculator ac36(.scan_win(scan_win36), .rectangle1_x(rectangle1_xs[36]), .rectangle1_y(rectangle1_ys[36]), .rectangle1_width(rectangle1_widths[36]), .rectangle1_height(rectangle1_heights[36]), .rectangle1_weight(rectangle1_weights[36]), .rectangle2_x(rectangle2_xs[36]), .rectangle2_y(rectangle2_ys[36]), .rectangle2_width(rectangle2_widths[36]), .rectangle2_height(rectangle2_heights[36]), .rectangle2_weight(rectangle2_weights[36]), .rectangle3_x(rectangle3_xs[36]), .rectangle3_y(rectangle3_ys[36]), .rectangle3_width(rectangle3_widths[36]), .rectangle3_height(rectangle3_heights[36]), .rectangle3_weight(rectangle3_weights[36]), .feature_threshold(feature_thresholds[36]), .feature_above(feature_aboves[36]), .feature_below(feature_belows[36]), .scan_win_std_dev(scan_win_std_dev[36]), .feature_accum(feature_accums[36]));
  accum_calculator ac37(.scan_win(scan_win37), .rectangle1_x(rectangle1_xs[37]), .rectangle1_y(rectangle1_ys[37]), .rectangle1_width(rectangle1_widths[37]), .rectangle1_height(rectangle1_heights[37]), .rectangle1_weight(rectangle1_weights[37]), .rectangle2_x(rectangle2_xs[37]), .rectangle2_y(rectangle2_ys[37]), .rectangle2_width(rectangle2_widths[37]), .rectangle2_height(rectangle2_heights[37]), .rectangle2_weight(rectangle2_weights[37]), .rectangle3_x(rectangle3_xs[37]), .rectangle3_y(rectangle3_ys[37]), .rectangle3_width(rectangle3_widths[37]), .rectangle3_height(rectangle3_heights[37]), .rectangle3_weight(rectangle3_weights[37]), .feature_threshold(feature_thresholds[37]), .feature_above(feature_aboves[37]), .feature_below(feature_belows[37]), .scan_win_std_dev(scan_win_std_dev[37]), .feature_accum(feature_accums[37]));
  accum_calculator ac38(.scan_win(scan_win38), .rectangle1_x(rectangle1_xs[38]), .rectangle1_y(rectangle1_ys[38]), .rectangle1_width(rectangle1_widths[38]), .rectangle1_height(rectangle1_heights[38]), .rectangle1_weight(rectangle1_weights[38]), .rectangle2_x(rectangle2_xs[38]), .rectangle2_y(rectangle2_ys[38]), .rectangle2_width(rectangle2_widths[38]), .rectangle2_height(rectangle2_heights[38]), .rectangle2_weight(rectangle2_weights[38]), .rectangle3_x(rectangle3_xs[38]), .rectangle3_y(rectangle3_ys[38]), .rectangle3_width(rectangle3_widths[38]), .rectangle3_height(rectangle3_heights[38]), .rectangle3_weight(rectangle3_weights[38]), .feature_threshold(feature_thresholds[38]), .feature_above(feature_aboves[38]), .feature_below(feature_belows[38]), .scan_win_std_dev(scan_win_std_dev[38]), .feature_accum(feature_accums[38]));
  accum_calculator ac39(.scan_win(scan_win39), .rectangle1_x(rectangle1_xs[39]), .rectangle1_y(rectangle1_ys[39]), .rectangle1_width(rectangle1_widths[39]), .rectangle1_height(rectangle1_heights[39]), .rectangle1_weight(rectangle1_weights[39]), .rectangle2_x(rectangle2_xs[39]), .rectangle2_y(rectangle2_ys[39]), .rectangle2_width(rectangle2_widths[39]), .rectangle2_height(rectangle2_heights[39]), .rectangle2_weight(rectangle2_weights[39]), .rectangle3_x(rectangle3_xs[39]), .rectangle3_y(rectangle3_ys[39]), .rectangle3_width(rectangle3_widths[39]), .rectangle3_height(rectangle3_heights[39]), .rectangle3_weight(rectangle3_weights[39]), .feature_threshold(feature_thresholds[39]), .feature_above(feature_aboves[39]), .feature_below(feature_belows[39]), .scan_win_std_dev(scan_win_std_dev[39]), .feature_accum(feature_accums[39]));
  accum_calculator ac40(.scan_win(scan_win40), .rectangle1_x(rectangle1_xs[40]), .rectangle1_y(rectangle1_ys[40]), .rectangle1_width(rectangle1_widths[40]), .rectangle1_height(rectangle1_heights[40]), .rectangle1_weight(rectangle1_weights[40]), .rectangle2_x(rectangle2_xs[40]), .rectangle2_y(rectangle2_ys[40]), .rectangle2_width(rectangle2_widths[40]), .rectangle2_height(rectangle2_heights[40]), .rectangle2_weight(rectangle2_weights[40]), .rectangle3_x(rectangle3_xs[40]), .rectangle3_y(rectangle3_ys[40]), .rectangle3_width(rectangle3_widths[40]), .rectangle3_height(rectangle3_heights[40]), .rectangle3_weight(rectangle3_weights[40]), .feature_threshold(feature_thresholds[40]), .feature_above(feature_aboves[40]), .feature_below(feature_belows[40]), .scan_win_std_dev(scan_win_std_dev[40]), .feature_accum(feature_accums[40]));
  accum_calculator ac41(.scan_win(scan_win41), .rectangle1_x(rectangle1_xs[41]), .rectangle1_y(rectangle1_ys[41]), .rectangle1_width(rectangle1_widths[41]), .rectangle1_height(rectangle1_heights[41]), .rectangle1_weight(rectangle1_weights[41]), .rectangle2_x(rectangle2_xs[41]), .rectangle2_y(rectangle2_ys[41]), .rectangle2_width(rectangle2_widths[41]), .rectangle2_height(rectangle2_heights[41]), .rectangle2_weight(rectangle2_weights[41]), .rectangle3_x(rectangle3_xs[41]), .rectangle3_y(rectangle3_ys[41]), .rectangle3_width(rectangle3_widths[41]), .rectangle3_height(rectangle3_heights[41]), .rectangle3_weight(rectangle3_weights[41]), .feature_threshold(feature_thresholds[41]), .feature_above(feature_aboves[41]), .feature_below(feature_belows[41]), .scan_win_std_dev(scan_win_std_dev[41]), .feature_accum(feature_accums[41]));
  accum_calculator ac42(.scan_win(scan_win42), .rectangle1_x(rectangle1_xs[42]), .rectangle1_y(rectangle1_ys[42]), .rectangle1_width(rectangle1_widths[42]), .rectangle1_height(rectangle1_heights[42]), .rectangle1_weight(rectangle1_weights[42]), .rectangle2_x(rectangle2_xs[42]), .rectangle2_y(rectangle2_ys[42]), .rectangle2_width(rectangle2_widths[42]), .rectangle2_height(rectangle2_heights[42]), .rectangle2_weight(rectangle2_weights[42]), .rectangle3_x(rectangle3_xs[42]), .rectangle3_y(rectangle3_ys[42]), .rectangle3_width(rectangle3_widths[42]), .rectangle3_height(rectangle3_heights[42]), .rectangle3_weight(rectangle3_weights[42]), .feature_threshold(feature_thresholds[42]), .feature_above(feature_aboves[42]), .feature_below(feature_belows[42]), .scan_win_std_dev(scan_win_std_dev[42]), .feature_accum(feature_accums[42]));
  accum_calculator ac43(.scan_win(scan_win43), .rectangle1_x(rectangle1_xs[43]), .rectangle1_y(rectangle1_ys[43]), .rectangle1_width(rectangle1_widths[43]), .rectangle1_height(rectangle1_heights[43]), .rectangle1_weight(rectangle1_weights[43]), .rectangle2_x(rectangle2_xs[43]), .rectangle2_y(rectangle2_ys[43]), .rectangle2_width(rectangle2_widths[43]), .rectangle2_height(rectangle2_heights[43]), .rectangle2_weight(rectangle2_weights[43]), .rectangle3_x(rectangle3_xs[43]), .rectangle3_y(rectangle3_ys[43]), .rectangle3_width(rectangle3_widths[43]), .rectangle3_height(rectangle3_heights[43]), .rectangle3_weight(rectangle3_weights[43]), .feature_threshold(feature_thresholds[43]), .feature_above(feature_aboves[43]), .feature_below(feature_belows[43]), .scan_win_std_dev(scan_win_std_dev[43]), .feature_accum(feature_accums[43]));
  accum_calculator ac44(.scan_win(scan_win44), .rectangle1_x(rectangle1_xs[44]), .rectangle1_y(rectangle1_ys[44]), .rectangle1_width(rectangle1_widths[44]), .rectangle1_height(rectangle1_heights[44]), .rectangle1_weight(rectangle1_weights[44]), .rectangle2_x(rectangle2_xs[44]), .rectangle2_y(rectangle2_ys[44]), .rectangle2_width(rectangle2_widths[44]), .rectangle2_height(rectangle2_heights[44]), .rectangle2_weight(rectangle2_weights[44]), .rectangle3_x(rectangle3_xs[44]), .rectangle3_y(rectangle3_ys[44]), .rectangle3_width(rectangle3_widths[44]), .rectangle3_height(rectangle3_heights[44]), .rectangle3_weight(rectangle3_weights[44]), .feature_threshold(feature_thresholds[44]), .feature_above(feature_aboves[44]), .feature_below(feature_belows[44]), .scan_win_std_dev(scan_win_std_dev[44]), .feature_accum(feature_accums[44]));
  accum_calculator ac45(.scan_win(scan_win45), .rectangle1_x(rectangle1_xs[45]), .rectangle1_y(rectangle1_ys[45]), .rectangle1_width(rectangle1_widths[45]), .rectangle1_height(rectangle1_heights[45]), .rectangle1_weight(rectangle1_weights[45]), .rectangle2_x(rectangle2_xs[45]), .rectangle2_y(rectangle2_ys[45]), .rectangle2_width(rectangle2_widths[45]), .rectangle2_height(rectangle2_heights[45]), .rectangle2_weight(rectangle2_weights[45]), .rectangle3_x(rectangle3_xs[45]), .rectangle3_y(rectangle3_ys[45]), .rectangle3_width(rectangle3_widths[45]), .rectangle3_height(rectangle3_heights[45]), .rectangle3_weight(rectangle3_weights[45]), .feature_threshold(feature_thresholds[45]), .feature_above(feature_aboves[45]), .feature_below(feature_belows[45]), .scan_win_std_dev(scan_win_std_dev[45]), .feature_accum(feature_accums[45]));
  accum_calculator ac46(.scan_win(scan_win46), .rectangle1_x(rectangle1_xs[46]), .rectangle1_y(rectangle1_ys[46]), .rectangle1_width(rectangle1_widths[46]), .rectangle1_height(rectangle1_heights[46]), .rectangle1_weight(rectangle1_weights[46]), .rectangle2_x(rectangle2_xs[46]), .rectangle2_y(rectangle2_ys[46]), .rectangle2_width(rectangle2_widths[46]), .rectangle2_height(rectangle2_heights[46]), .rectangle2_weight(rectangle2_weights[46]), .rectangle3_x(rectangle3_xs[46]), .rectangle3_y(rectangle3_ys[46]), .rectangle3_width(rectangle3_widths[46]), .rectangle3_height(rectangle3_heights[46]), .rectangle3_weight(rectangle3_weights[46]), .feature_threshold(feature_thresholds[46]), .feature_above(feature_aboves[46]), .feature_below(feature_belows[46]), .scan_win_std_dev(scan_win_std_dev[46]), .feature_accum(feature_accums[46]));
  accum_calculator ac47(.scan_win(scan_win47), .rectangle1_x(rectangle1_xs[47]), .rectangle1_y(rectangle1_ys[47]), .rectangle1_width(rectangle1_widths[47]), .rectangle1_height(rectangle1_heights[47]), .rectangle1_weight(rectangle1_weights[47]), .rectangle2_x(rectangle2_xs[47]), .rectangle2_y(rectangle2_ys[47]), .rectangle2_width(rectangle2_widths[47]), .rectangle2_height(rectangle2_heights[47]), .rectangle2_weight(rectangle2_weights[47]), .rectangle3_x(rectangle3_xs[47]), .rectangle3_y(rectangle3_ys[47]), .rectangle3_width(rectangle3_widths[47]), .rectangle3_height(rectangle3_heights[47]), .rectangle3_weight(rectangle3_weights[47]), .feature_threshold(feature_thresholds[47]), .feature_above(feature_aboves[47]), .feature_below(feature_belows[47]), .scan_win_std_dev(scan_win_std_dev[47]), .feature_accum(feature_accums[47]));
  accum_calculator ac48(.scan_win(scan_win48), .rectangle1_x(rectangle1_xs[48]), .rectangle1_y(rectangle1_ys[48]), .rectangle1_width(rectangle1_widths[48]), .rectangle1_height(rectangle1_heights[48]), .rectangle1_weight(rectangle1_weights[48]), .rectangle2_x(rectangle2_xs[48]), .rectangle2_y(rectangle2_ys[48]), .rectangle2_width(rectangle2_widths[48]), .rectangle2_height(rectangle2_heights[48]), .rectangle2_weight(rectangle2_weights[48]), .rectangle3_x(rectangle3_xs[48]), .rectangle3_y(rectangle3_ys[48]), .rectangle3_width(rectangle3_widths[48]), .rectangle3_height(rectangle3_heights[48]), .rectangle3_weight(rectangle3_weights[48]), .feature_threshold(feature_thresholds[48]), .feature_above(feature_aboves[48]), .feature_below(feature_belows[48]), .scan_win_std_dev(scan_win_std_dev[48]), .feature_accum(feature_accums[48]));
  accum_calculator ac49(.scan_win(scan_win49), .rectangle1_x(rectangle1_xs[49]), .rectangle1_y(rectangle1_ys[49]), .rectangle1_width(rectangle1_widths[49]), .rectangle1_height(rectangle1_heights[49]), .rectangle1_weight(rectangle1_weights[49]), .rectangle2_x(rectangle2_xs[49]), .rectangle2_y(rectangle2_ys[49]), .rectangle2_width(rectangle2_widths[49]), .rectangle2_height(rectangle2_heights[49]), .rectangle2_weight(rectangle2_weights[49]), .rectangle3_x(rectangle3_xs[49]), .rectangle3_y(rectangle3_ys[49]), .rectangle3_width(rectangle3_widths[49]), .rectangle3_height(rectangle3_heights[49]), .rectangle3_weight(rectangle3_weights[49]), .feature_threshold(feature_thresholds[49]), .feature_above(feature_aboves[49]), .feature_below(feature_belows[49]), .scan_win_std_dev(scan_win_std_dev[49]), .feature_accum(feature_accums[49]));
  accum_calculator ac50(.scan_win(scan_win50), .rectangle1_x(rectangle1_xs[50]), .rectangle1_y(rectangle1_ys[50]), .rectangle1_width(rectangle1_widths[50]), .rectangle1_height(rectangle1_heights[50]), .rectangle1_weight(rectangle1_weights[50]), .rectangle2_x(rectangle2_xs[50]), .rectangle2_y(rectangle2_ys[50]), .rectangle2_width(rectangle2_widths[50]), .rectangle2_height(rectangle2_heights[50]), .rectangle2_weight(rectangle2_weights[50]), .rectangle3_x(rectangle3_xs[50]), .rectangle3_y(rectangle3_ys[50]), .rectangle3_width(rectangle3_widths[50]), .rectangle3_height(rectangle3_heights[50]), .rectangle3_weight(rectangle3_weights[50]), .feature_threshold(feature_thresholds[50]), .feature_above(feature_aboves[50]), .feature_below(feature_belows[50]), .scan_win_std_dev(scan_win_std_dev[50]), .feature_accum(feature_accums[50]));
  accum_calculator ac51(.scan_win(scan_win51), .rectangle1_x(rectangle1_xs[51]), .rectangle1_y(rectangle1_ys[51]), .rectangle1_width(rectangle1_widths[51]), .rectangle1_height(rectangle1_heights[51]), .rectangle1_weight(rectangle1_weights[51]), .rectangle2_x(rectangle2_xs[51]), .rectangle2_y(rectangle2_ys[51]), .rectangle2_width(rectangle2_widths[51]), .rectangle2_height(rectangle2_heights[51]), .rectangle2_weight(rectangle2_weights[51]), .rectangle3_x(rectangle3_xs[51]), .rectangle3_y(rectangle3_ys[51]), .rectangle3_width(rectangle3_widths[51]), .rectangle3_height(rectangle3_heights[51]), .rectangle3_weight(rectangle3_weights[51]), .feature_threshold(feature_thresholds[51]), .feature_above(feature_aboves[51]), .feature_below(feature_belows[51]), .scan_win_std_dev(scan_win_std_dev[51]), .feature_accum(feature_accums[51]));
  accum_calculator ac52(.scan_win(scan_win52), .rectangle1_x(rectangle1_xs[52]), .rectangle1_y(rectangle1_ys[52]), .rectangle1_width(rectangle1_widths[52]), .rectangle1_height(rectangle1_heights[52]), .rectangle1_weight(rectangle1_weights[52]), .rectangle2_x(rectangle2_xs[52]), .rectangle2_y(rectangle2_ys[52]), .rectangle2_width(rectangle2_widths[52]), .rectangle2_height(rectangle2_heights[52]), .rectangle2_weight(rectangle2_weights[52]), .rectangle3_x(rectangle3_xs[52]), .rectangle3_y(rectangle3_ys[52]), .rectangle3_width(rectangle3_widths[52]), .rectangle3_height(rectangle3_heights[52]), .rectangle3_weight(rectangle3_weights[52]), .feature_threshold(feature_thresholds[52]), .feature_above(feature_aboves[52]), .feature_below(feature_belows[52]), .scan_win_std_dev(scan_win_std_dev[52]), .feature_accum(feature_accums[52]));
  accum_calculator ac53(.scan_win(scan_win53), .rectangle1_x(rectangle1_xs[53]), .rectangle1_y(rectangle1_ys[53]), .rectangle1_width(rectangle1_widths[53]), .rectangle1_height(rectangle1_heights[53]), .rectangle1_weight(rectangle1_weights[53]), .rectangle2_x(rectangle2_xs[53]), .rectangle2_y(rectangle2_ys[53]), .rectangle2_width(rectangle2_widths[53]), .rectangle2_height(rectangle2_heights[53]), .rectangle2_weight(rectangle2_weights[53]), .rectangle3_x(rectangle3_xs[53]), .rectangle3_y(rectangle3_ys[53]), .rectangle3_width(rectangle3_widths[53]), .rectangle3_height(rectangle3_heights[53]), .rectangle3_weight(rectangle3_weights[53]), .feature_threshold(feature_thresholds[53]), .feature_above(feature_aboves[53]), .feature_below(feature_belows[53]), .scan_win_std_dev(scan_win_std_dev[53]), .feature_accum(feature_accums[53]));
  accum_calculator ac54(.scan_win(scan_win54), .rectangle1_x(rectangle1_xs[54]), .rectangle1_y(rectangle1_ys[54]), .rectangle1_width(rectangle1_widths[54]), .rectangle1_height(rectangle1_heights[54]), .rectangle1_weight(rectangle1_weights[54]), .rectangle2_x(rectangle2_xs[54]), .rectangle2_y(rectangle2_ys[54]), .rectangle2_width(rectangle2_widths[54]), .rectangle2_height(rectangle2_heights[54]), .rectangle2_weight(rectangle2_weights[54]), .rectangle3_x(rectangle3_xs[54]), .rectangle3_y(rectangle3_ys[54]), .rectangle3_width(rectangle3_widths[54]), .rectangle3_height(rectangle3_heights[54]), .rectangle3_weight(rectangle3_weights[54]), .feature_threshold(feature_thresholds[54]), .feature_above(feature_aboves[54]), .feature_below(feature_belows[54]), .scan_win_std_dev(scan_win_std_dev[54]), .feature_accum(feature_accums[54]));
  accum_calculator ac55(.scan_win(scan_win55), .rectangle1_x(rectangle1_xs[55]), .rectangle1_y(rectangle1_ys[55]), .rectangle1_width(rectangle1_widths[55]), .rectangle1_height(rectangle1_heights[55]), .rectangle1_weight(rectangle1_weights[55]), .rectangle2_x(rectangle2_xs[55]), .rectangle2_y(rectangle2_ys[55]), .rectangle2_width(rectangle2_widths[55]), .rectangle2_height(rectangle2_heights[55]), .rectangle2_weight(rectangle2_weights[55]), .rectangle3_x(rectangle3_xs[55]), .rectangle3_y(rectangle3_ys[55]), .rectangle3_width(rectangle3_widths[55]), .rectangle3_height(rectangle3_heights[55]), .rectangle3_weight(rectangle3_weights[55]), .feature_threshold(feature_thresholds[55]), .feature_above(feature_aboves[55]), .feature_below(feature_belows[55]), .scan_win_std_dev(scan_win_std_dev[55]), .feature_accum(feature_accums[55]));
  accum_calculator ac56(.scan_win(scan_win56), .rectangle1_x(rectangle1_xs[56]), .rectangle1_y(rectangle1_ys[56]), .rectangle1_width(rectangle1_widths[56]), .rectangle1_height(rectangle1_heights[56]), .rectangle1_weight(rectangle1_weights[56]), .rectangle2_x(rectangle2_xs[56]), .rectangle2_y(rectangle2_ys[56]), .rectangle2_width(rectangle2_widths[56]), .rectangle2_height(rectangle2_heights[56]), .rectangle2_weight(rectangle2_weights[56]), .rectangle3_x(rectangle3_xs[56]), .rectangle3_y(rectangle3_ys[56]), .rectangle3_width(rectangle3_widths[56]), .rectangle3_height(rectangle3_heights[56]), .rectangle3_weight(rectangle3_weights[56]), .feature_threshold(feature_thresholds[56]), .feature_above(feature_aboves[56]), .feature_below(feature_belows[56]), .scan_win_std_dev(scan_win_std_dev[56]), .feature_accum(feature_accums[56]));
  accum_calculator ac57(.scan_win(scan_win57), .rectangle1_x(rectangle1_xs[57]), .rectangle1_y(rectangle1_ys[57]), .rectangle1_width(rectangle1_widths[57]), .rectangle1_height(rectangle1_heights[57]), .rectangle1_weight(rectangle1_weights[57]), .rectangle2_x(rectangle2_xs[57]), .rectangle2_y(rectangle2_ys[57]), .rectangle2_width(rectangle2_widths[57]), .rectangle2_height(rectangle2_heights[57]), .rectangle2_weight(rectangle2_weights[57]), .rectangle3_x(rectangle3_xs[57]), .rectangle3_y(rectangle3_ys[57]), .rectangle3_width(rectangle3_widths[57]), .rectangle3_height(rectangle3_heights[57]), .rectangle3_weight(rectangle3_weights[57]), .feature_threshold(feature_thresholds[57]), .feature_above(feature_aboves[57]), .feature_below(feature_belows[57]), .scan_win_std_dev(scan_win_std_dev[57]), .feature_accum(feature_accums[57]));
  accum_calculator ac58(.scan_win(scan_win58), .rectangle1_x(rectangle1_xs[58]), .rectangle1_y(rectangle1_ys[58]), .rectangle1_width(rectangle1_widths[58]), .rectangle1_height(rectangle1_heights[58]), .rectangle1_weight(rectangle1_weights[58]), .rectangle2_x(rectangle2_xs[58]), .rectangle2_y(rectangle2_ys[58]), .rectangle2_width(rectangle2_widths[58]), .rectangle2_height(rectangle2_heights[58]), .rectangle2_weight(rectangle2_weights[58]), .rectangle3_x(rectangle3_xs[58]), .rectangle3_y(rectangle3_ys[58]), .rectangle3_width(rectangle3_widths[58]), .rectangle3_height(rectangle3_heights[58]), .rectangle3_weight(rectangle3_weights[58]), .feature_threshold(feature_thresholds[58]), .feature_above(feature_aboves[58]), .feature_below(feature_belows[58]), .scan_win_std_dev(scan_win_std_dev[58]), .feature_accum(feature_accums[58]));
  accum_calculator ac59(.scan_win(scan_win59), .rectangle1_x(rectangle1_xs[59]), .rectangle1_y(rectangle1_ys[59]), .rectangle1_width(rectangle1_widths[59]), .rectangle1_height(rectangle1_heights[59]), .rectangle1_weight(rectangle1_weights[59]), .rectangle2_x(rectangle2_xs[59]), .rectangle2_y(rectangle2_ys[59]), .rectangle2_width(rectangle2_widths[59]), .rectangle2_height(rectangle2_heights[59]), .rectangle2_weight(rectangle2_weights[59]), .rectangle3_x(rectangle3_xs[59]), .rectangle3_y(rectangle3_ys[59]), .rectangle3_width(rectangle3_widths[59]), .rectangle3_height(rectangle3_heights[59]), .rectangle3_weight(rectangle3_weights[59]), .feature_threshold(feature_thresholds[59]), .feature_above(feature_aboves[59]), .feature_below(feature_belows[59]), .scan_win_std_dev(scan_win_std_dev[59]), .feature_accum(feature_accums[59]));
  accum_calculator ac60(.scan_win(scan_win60), .rectangle1_x(rectangle1_xs[60]), .rectangle1_y(rectangle1_ys[60]), .rectangle1_width(rectangle1_widths[60]), .rectangle1_height(rectangle1_heights[60]), .rectangle1_weight(rectangle1_weights[60]), .rectangle2_x(rectangle2_xs[60]), .rectangle2_y(rectangle2_ys[60]), .rectangle2_width(rectangle2_widths[60]), .rectangle2_height(rectangle2_heights[60]), .rectangle2_weight(rectangle2_weights[60]), .rectangle3_x(rectangle3_xs[60]), .rectangle3_y(rectangle3_ys[60]), .rectangle3_width(rectangle3_widths[60]), .rectangle3_height(rectangle3_heights[60]), .rectangle3_weight(rectangle3_weights[60]), .feature_threshold(feature_thresholds[60]), .feature_above(feature_aboves[60]), .feature_below(feature_belows[60]), .scan_win_std_dev(scan_win_std_dev[60]), .feature_accum(feature_accums[60]));
  accum_calculator ac61(.scan_win(scan_win61), .rectangle1_x(rectangle1_xs[61]), .rectangle1_y(rectangle1_ys[61]), .rectangle1_width(rectangle1_widths[61]), .rectangle1_height(rectangle1_heights[61]), .rectangle1_weight(rectangle1_weights[61]), .rectangle2_x(rectangle2_xs[61]), .rectangle2_y(rectangle2_ys[61]), .rectangle2_width(rectangle2_widths[61]), .rectangle2_height(rectangle2_heights[61]), .rectangle2_weight(rectangle2_weights[61]), .rectangle3_x(rectangle3_xs[61]), .rectangle3_y(rectangle3_ys[61]), .rectangle3_width(rectangle3_widths[61]), .rectangle3_height(rectangle3_heights[61]), .rectangle3_weight(rectangle3_weights[61]), .feature_threshold(feature_thresholds[61]), .feature_above(feature_aboves[61]), .feature_below(feature_belows[61]), .scan_win_std_dev(scan_win_std_dev[61]), .feature_accum(feature_accums[61]));
  accum_calculator ac62(.scan_win(scan_win62), .rectangle1_x(rectangle1_xs[62]), .rectangle1_y(rectangle1_ys[62]), .rectangle1_width(rectangle1_widths[62]), .rectangle1_height(rectangle1_heights[62]), .rectangle1_weight(rectangle1_weights[62]), .rectangle2_x(rectangle2_xs[62]), .rectangle2_y(rectangle2_ys[62]), .rectangle2_width(rectangle2_widths[62]), .rectangle2_height(rectangle2_heights[62]), .rectangle2_weight(rectangle2_weights[62]), .rectangle3_x(rectangle3_xs[62]), .rectangle3_y(rectangle3_ys[62]), .rectangle3_width(rectangle3_widths[62]), .rectangle3_height(rectangle3_heights[62]), .rectangle3_weight(rectangle3_weights[62]), .feature_threshold(feature_thresholds[62]), .feature_above(feature_aboves[62]), .feature_below(feature_belows[62]), .scan_win_std_dev(scan_win_std_dev[62]), .feature_accum(feature_accums[62]));
  accum_calculator ac63(.scan_win(scan_win63), .rectangle1_x(rectangle1_xs[63]), .rectangle1_y(rectangle1_ys[63]), .rectangle1_width(rectangle1_widths[63]), .rectangle1_height(rectangle1_heights[63]), .rectangle1_weight(rectangle1_weights[63]), .rectangle2_x(rectangle2_xs[63]), .rectangle2_y(rectangle2_ys[63]), .rectangle2_width(rectangle2_widths[63]), .rectangle2_height(rectangle2_heights[63]), .rectangle2_weight(rectangle2_weights[63]), .rectangle3_x(rectangle3_xs[63]), .rectangle3_y(rectangle3_ys[63]), .rectangle3_width(rectangle3_widths[63]), .rectangle3_height(rectangle3_heights[63]), .rectangle3_weight(rectangle3_weights[63]), .feature_threshold(feature_thresholds[63]), .feature_above(feature_aboves[63]), .feature_below(feature_belows[63]), .scan_win_std_dev(scan_win_std_dev[63]), .feature_accum(feature_accums[63]));
  accum_calculator ac64(.scan_win(scan_win64), .rectangle1_x(rectangle1_xs[64]), .rectangle1_y(rectangle1_ys[64]), .rectangle1_width(rectangle1_widths[64]), .rectangle1_height(rectangle1_heights[64]), .rectangle1_weight(rectangle1_weights[64]), .rectangle2_x(rectangle2_xs[64]), .rectangle2_y(rectangle2_ys[64]), .rectangle2_width(rectangle2_widths[64]), .rectangle2_height(rectangle2_heights[64]), .rectangle2_weight(rectangle2_weights[64]), .rectangle3_x(rectangle3_xs[64]), .rectangle3_y(rectangle3_ys[64]), .rectangle3_width(rectangle3_widths[64]), .rectangle3_height(rectangle3_heights[64]), .rectangle3_weight(rectangle3_weights[64]), .feature_threshold(feature_thresholds[64]), .feature_above(feature_aboves[64]), .feature_below(feature_belows[64]), .scan_win_std_dev(scan_win_std_dev[64]), .feature_accum(feature_accums[64]));
  accum_calculator ac65(.scan_win(scan_win65), .rectangle1_x(rectangle1_xs[65]), .rectangle1_y(rectangle1_ys[65]), .rectangle1_width(rectangle1_widths[65]), .rectangle1_height(rectangle1_heights[65]), .rectangle1_weight(rectangle1_weights[65]), .rectangle2_x(rectangle2_xs[65]), .rectangle2_y(rectangle2_ys[65]), .rectangle2_width(rectangle2_widths[65]), .rectangle2_height(rectangle2_heights[65]), .rectangle2_weight(rectangle2_weights[65]), .rectangle3_x(rectangle3_xs[65]), .rectangle3_y(rectangle3_ys[65]), .rectangle3_width(rectangle3_widths[65]), .rectangle3_height(rectangle3_heights[65]), .rectangle3_weight(rectangle3_weights[65]), .feature_threshold(feature_thresholds[65]), .feature_above(feature_aboves[65]), .feature_below(feature_belows[65]), .scan_win_std_dev(scan_win_std_dev[65]), .feature_accum(feature_accums[65]));
  accum_calculator ac66(.scan_win(scan_win66), .rectangle1_x(rectangle1_xs[66]), .rectangle1_y(rectangle1_ys[66]), .rectangle1_width(rectangle1_widths[66]), .rectangle1_height(rectangle1_heights[66]), .rectangle1_weight(rectangle1_weights[66]), .rectangle2_x(rectangle2_xs[66]), .rectangle2_y(rectangle2_ys[66]), .rectangle2_width(rectangle2_widths[66]), .rectangle2_height(rectangle2_heights[66]), .rectangle2_weight(rectangle2_weights[66]), .rectangle3_x(rectangle3_xs[66]), .rectangle3_y(rectangle3_ys[66]), .rectangle3_width(rectangle3_widths[66]), .rectangle3_height(rectangle3_heights[66]), .rectangle3_weight(rectangle3_weights[66]), .feature_threshold(feature_thresholds[66]), .feature_above(feature_aboves[66]), .feature_below(feature_belows[66]), .scan_win_std_dev(scan_win_std_dev[66]), .feature_accum(feature_accums[66]));
  accum_calculator ac67(.scan_win(scan_win67), .rectangle1_x(rectangle1_xs[67]), .rectangle1_y(rectangle1_ys[67]), .rectangle1_width(rectangle1_widths[67]), .rectangle1_height(rectangle1_heights[67]), .rectangle1_weight(rectangle1_weights[67]), .rectangle2_x(rectangle2_xs[67]), .rectangle2_y(rectangle2_ys[67]), .rectangle2_width(rectangle2_widths[67]), .rectangle2_height(rectangle2_heights[67]), .rectangle2_weight(rectangle2_weights[67]), .rectangle3_x(rectangle3_xs[67]), .rectangle3_y(rectangle3_ys[67]), .rectangle3_width(rectangle3_widths[67]), .rectangle3_height(rectangle3_heights[67]), .rectangle3_weight(rectangle3_weights[67]), .feature_threshold(feature_thresholds[67]), .feature_above(feature_aboves[67]), .feature_below(feature_belows[67]), .scan_win_std_dev(scan_win_std_dev[67]), .feature_accum(feature_accums[67]));
  accum_calculator ac68(.scan_win(scan_win68), .rectangle1_x(rectangle1_xs[68]), .rectangle1_y(rectangle1_ys[68]), .rectangle1_width(rectangle1_widths[68]), .rectangle1_height(rectangle1_heights[68]), .rectangle1_weight(rectangle1_weights[68]), .rectangle2_x(rectangle2_xs[68]), .rectangle2_y(rectangle2_ys[68]), .rectangle2_width(rectangle2_widths[68]), .rectangle2_height(rectangle2_heights[68]), .rectangle2_weight(rectangle2_weights[68]), .rectangle3_x(rectangle3_xs[68]), .rectangle3_y(rectangle3_ys[68]), .rectangle3_width(rectangle3_widths[68]), .rectangle3_height(rectangle3_heights[68]), .rectangle3_weight(rectangle3_weights[68]), .feature_threshold(feature_thresholds[68]), .feature_above(feature_aboves[68]), .feature_below(feature_belows[68]), .scan_win_std_dev(scan_win_std_dev[68]), .feature_accum(feature_accums[68]));
  accum_calculator ac69(.scan_win(scan_win69), .rectangle1_x(rectangle1_xs[69]), .rectangle1_y(rectangle1_ys[69]), .rectangle1_width(rectangle1_widths[69]), .rectangle1_height(rectangle1_heights[69]), .rectangle1_weight(rectangle1_weights[69]), .rectangle2_x(rectangle2_xs[69]), .rectangle2_y(rectangle2_ys[69]), .rectangle2_width(rectangle2_widths[69]), .rectangle2_height(rectangle2_heights[69]), .rectangle2_weight(rectangle2_weights[69]), .rectangle3_x(rectangle3_xs[69]), .rectangle3_y(rectangle3_ys[69]), .rectangle3_width(rectangle3_widths[69]), .rectangle3_height(rectangle3_heights[69]), .rectangle3_weight(rectangle3_weights[69]), .feature_threshold(feature_thresholds[69]), .feature_above(feature_aboves[69]), .feature_below(feature_belows[69]), .scan_win_std_dev(scan_win_std_dev[69]), .feature_accum(feature_accums[69]));
  accum_calculator ac70(.scan_win(scan_win70), .rectangle1_x(rectangle1_xs[70]), .rectangle1_y(rectangle1_ys[70]), .rectangle1_width(rectangle1_widths[70]), .rectangle1_height(rectangle1_heights[70]), .rectangle1_weight(rectangle1_weights[70]), .rectangle2_x(rectangle2_xs[70]), .rectangle2_y(rectangle2_ys[70]), .rectangle2_width(rectangle2_widths[70]), .rectangle2_height(rectangle2_heights[70]), .rectangle2_weight(rectangle2_weights[70]), .rectangle3_x(rectangle3_xs[70]), .rectangle3_y(rectangle3_ys[70]), .rectangle3_width(rectangle3_widths[70]), .rectangle3_height(rectangle3_heights[70]), .rectangle3_weight(rectangle3_weights[70]), .feature_threshold(feature_thresholds[70]), .feature_above(feature_aboves[70]), .feature_below(feature_belows[70]), .scan_win_std_dev(scan_win_std_dev[70]), .feature_accum(feature_accums[70]));
  accum_calculator ac71(.scan_win(scan_win71), .rectangle1_x(rectangle1_xs[71]), .rectangle1_y(rectangle1_ys[71]), .rectangle1_width(rectangle1_widths[71]), .rectangle1_height(rectangle1_heights[71]), .rectangle1_weight(rectangle1_weights[71]), .rectangle2_x(rectangle2_xs[71]), .rectangle2_y(rectangle2_ys[71]), .rectangle2_width(rectangle2_widths[71]), .rectangle2_height(rectangle2_heights[71]), .rectangle2_weight(rectangle2_weights[71]), .rectangle3_x(rectangle3_xs[71]), .rectangle3_y(rectangle3_ys[71]), .rectangle3_width(rectangle3_widths[71]), .rectangle3_height(rectangle3_heights[71]), .rectangle3_weight(rectangle3_weights[71]), .feature_threshold(feature_thresholds[71]), .feature_above(feature_aboves[71]), .feature_below(feature_belows[71]), .scan_win_std_dev(scan_win_std_dev[71]), .feature_accum(feature_accums[71]));
  accum_calculator ac72(.scan_win(scan_win72), .rectangle1_x(rectangle1_xs[72]), .rectangle1_y(rectangle1_ys[72]), .rectangle1_width(rectangle1_widths[72]), .rectangle1_height(rectangle1_heights[72]), .rectangle1_weight(rectangle1_weights[72]), .rectangle2_x(rectangle2_xs[72]), .rectangle2_y(rectangle2_ys[72]), .rectangle2_width(rectangle2_widths[72]), .rectangle2_height(rectangle2_heights[72]), .rectangle2_weight(rectangle2_weights[72]), .rectangle3_x(rectangle3_xs[72]), .rectangle3_y(rectangle3_ys[72]), .rectangle3_width(rectangle3_widths[72]), .rectangle3_height(rectangle3_heights[72]), .rectangle3_weight(rectangle3_weights[72]), .feature_threshold(feature_thresholds[72]), .feature_above(feature_aboves[72]), .feature_below(feature_belows[72]), .scan_win_std_dev(scan_win_std_dev[72]), .feature_accum(feature_accums[72]));
  accum_calculator ac73(.scan_win(scan_win73), .rectangle1_x(rectangle1_xs[73]), .rectangle1_y(rectangle1_ys[73]), .rectangle1_width(rectangle1_widths[73]), .rectangle1_height(rectangle1_heights[73]), .rectangle1_weight(rectangle1_weights[73]), .rectangle2_x(rectangle2_xs[73]), .rectangle2_y(rectangle2_ys[73]), .rectangle2_width(rectangle2_widths[73]), .rectangle2_height(rectangle2_heights[73]), .rectangle2_weight(rectangle2_weights[73]), .rectangle3_x(rectangle3_xs[73]), .rectangle3_y(rectangle3_ys[73]), .rectangle3_width(rectangle3_widths[73]), .rectangle3_height(rectangle3_heights[73]), .rectangle3_weight(rectangle3_weights[73]), .feature_threshold(feature_thresholds[73]), .feature_above(feature_aboves[73]), .feature_below(feature_belows[73]), .scan_win_std_dev(scan_win_std_dev[73]), .feature_accum(feature_accums[73]));
  accum_calculator ac74(.scan_win(scan_win74), .rectangle1_x(rectangle1_xs[74]), .rectangle1_y(rectangle1_ys[74]), .rectangle1_width(rectangle1_widths[74]), .rectangle1_height(rectangle1_heights[74]), .rectangle1_weight(rectangle1_weights[74]), .rectangle2_x(rectangle2_xs[74]), .rectangle2_y(rectangle2_ys[74]), .rectangle2_width(rectangle2_widths[74]), .rectangle2_height(rectangle2_heights[74]), .rectangle2_weight(rectangle2_weights[74]), .rectangle3_x(rectangle3_xs[74]), .rectangle3_y(rectangle3_ys[74]), .rectangle3_width(rectangle3_widths[74]), .rectangle3_height(rectangle3_heights[74]), .rectangle3_weight(rectangle3_weights[74]), .feature_threshold(feature_thresholds[74]), .feature_above(feature_aboves[74]), .feature_below(feature_belows[74]), .scan_win_std_dev(scan_win_std_dev[74]), .feature_accum(feature_accums[74]));
  accum_calculator ac75(.scan_win(scan_win75), .rectangle1_x(rectangle1_xs[75]), .rectangle1_y(rectangle1_ys[75]), .rectangle1_width(rectangle1_widths[75]), .rectangle1_height(rectangle1_heights[75]), .rectangle1_weight(rectangle1_weights[75]), .rectangle2_x(rectangle2_xs[75]), .rectangle2_y(rectangle2_ys[75]), .rectangle2_width(rectangle2_widths[75]), .rectangle2_height(rectangle2_heights[75]), .rectangle2_weight(rectangle2_weights[75]), .rectangle3_x(rectangle3_xs[75]), .rectangle3_y(rectangle3_ys[75]), .rectangle3_width(rectangle3_widths[75]), .rectangle3_height(rectangle3_heights[75]), .rectangle3_weight(rectangle3_weights[75]), .feature_threshold(feature_thresholds[75]), .feature_above(feature_aboves[75]), .feature_below(feature_belows[75]), .scan_win_std_dev(scan_win_std_dev[75]), .feature_accum(feature_accums[75]));
  accum_calculator ac76(.scan_win(scan_win76), .rectangle1_x(rectangle1_xs[76]), .rectangle1_y(rectangle1_ys[76]), .rectangle1_width(rectangle1_widths[76]), .rectangle1_height(rectangle1_heights[76]), .rectangle1_weight(rectangle1_weights[76]), .rectangle2_x(rectangle2_xs[76]), .rectangle2_y(rectangle2_ys[76]), .rectangle2_width(rectangle2_widths[76]), .rectangle2_height(rectangle2_heights[76]), .rectangle2_weight(rectangle2_weights[76]), .rectangle3_x(rectangle3_xs[76]), .rectangle3_y(rectangle3_ys[76]), .rectangle3_width(rectangle3_widths[76]), .rectangle3_height(rectangle3_heights[76]), .rectangle3_weight(rectangle3_weights[76]), .feature_threshold(feature_thresholds[76]), .feature_above(feature_aboves[76]), .feature_below(feature_belows[76]), .scan_win_std_dev(scan_win_std_dev[76]), .feature_accum(feature_accums[76]));
  accum_calculator ac77(.scan_win(scan_win77), .rectangle1_x(rectangle1_xs[77]), .rectangle1_y(rectangle1_ys[77]), .rectangle1_width(rectangle1_widths[77]), .rectangle1_height(rectangle1_heights[77]), .rectangle1_weight(rectangle1_weights[77]), .rectangle2_x(rectangle2_xs[77]), .rectangle2_y(rectangle2_ys[77]), .rectangle2_width(rectangle2_widths[77]), .rectangle2_height(rectangle2_heights[77]), .rectangle2_weight(rectangle2_weights[77]), .rectangle3_x(rectangle3_xs[77]), .rectangle3_y(rectangle3_ys[77]), .rectangle3_width(rectangle3_widths[77]), .rectangle3_height(rectangle3_heights[77]), .rectangle3_weight(rectangle3_weights[77]), .feature_threshold(feature_thresholds[77]), .feature_above(feature_aboves[77]), .feature_below(feature_belows[77]), .scan_win_std_dev(scan_win_std_dev[77]), .feature_accum(feature_accums[77]));
  accum_calculator ac78(.scan_win(scan_win78), .rectangle1_x(rectangle1_xs[78]), .rectangle1_y(rectangle1_ys[78]), .rectangle1_width(rectangle1_widths[78]), .rectangle1_height(rectangle1_heights[78]), .rectangle1_weight(rectangle1_weights[78]), .rectangle2_x(rectangle2_xs[78]), .rectangle2_y(rectangle2_ys[78]), .rectangle2_width(rectangle2_widths[78]), .rectangle2_height(rectangle2_heights[78]), .rectangle2_weight(rectangle2_weights[78]), .rectangle3_x(rectangle3_xs[78]), .rectangle3_y(rectangle3_ys[78]), .rectangle3_width(rectangle3_widths[78]), .rectangle3_height(rectangle3_heights[78]), .rectangle3_weight(rectangle3_weights[78]), .feature_threshold(feature_thresholds[78]), .feature_above(feature_aboves[78]), .feature_below(feature_belows[78]), .scan_win_std_dev(scan_win_std_dev[78]), .feature_accum(feature_accums[78]));
  accum_calculator ac79(.scan_win(scan_win79), .rectangle1_x(rectangle1_xs[79]), .rectangle1_y(rectangle1_ys[79]), .rectangle1_width(rectangle1_widths[79]), .rectangle1_height(rectangle1_heights[79]), .rectangle1_weight(rectangle1_weights[79]), .rectangle2_x(rectangle2_xs[79]), .rectangle2_y(rectangle2_ys[79]), .rectangle2_width(rectangle2_widths[79]), .rectangle2_height(rectangle2_heights[79]), .rectangle2_weight(rectangle2_weights[79]), .rectangle3_x(rectangle3_xs[79]), .rectangle3_y(rectangle3_ys[79]), .rectangle3_width(rectangle3_widths[79]), .rectangle3_height(rectangle3_heights[79]), .rectangle3_weight(rectangle3_weights[79]), .feature_threshold(feature_thresholds[79]), .feature_above(feature_aboves[79]), .feature_below(feature_belows[79]), .scan_win_std_dev(scan_win_std_dev[79]), .feature_accum(feature_accums[79]));
  accum_calculator ac80(.scan_win(scan_win80), .rectangle1_x(rectangle1_xs[80]), .rectangle1_y(rectangle1_ys[80]), .rectangle1_width(rectangle1_widths[80]), .rectangle1_height(rectangle1_heights[80]), .rectangle1_weight(rectangle1_weights[80]), .rectangle2_x(rectangle2_xs[80]), .rectangle2_y(rectangle2_ys[80]), .rectangle2_width(rectangle2_widths[80]), .rectangle2_height(rectangle2_heights[80]), .rectangle2_weight(rectangle2_weights[80]), .rectangle3_x(rectangle3_xs[80]), .rectangle3_y(rectangle3_ys[80]), .rectangle3_width(rectangle3_widths[80]), .rectangle3_height(rectangle3_heights[80]), .rectangle3_weight(rectangle3_weights[80]), .feature_threshold(feature_thresholds[80]), .feature_above(feature_aboves[80]), .feature_below(feature_belows[80]), .scan_win_std_dev(scan_win_std_dev[80]), .feature_accum(feature_accums[80]));
  accum_calculator ac81(.scan_win(scan_win81), .rectangle1_x(rectangle1_xs[81]), .rectangle1_y(rectangle1_ys[81]), .rectangle1_width(rectangle1_widths[81]), .rectangle1_height(rectangle1_heights[81]), .rectangle1_weight(rectangle1_weights[81]), .rectangle2_x(rectangle2_xs[81]), .rectangle2_y(rectangle2_ys[81]), .rectangle2_width(rectangle2_widths[81]), .rectangle2_height(rectangle2_heights[81]), .rectangle2_weight(rectangle2_weights[81]), .rectangle3_x(rectangle3_xs[81]), .rectangle3_y(rectangle3_ys[81]), .rectangle3_width(rectangle3_widths[81]), .rectangle3_height(rectangle3_heights[81]), .rectangle3_weight(rectangle3_weights[81]), .feature_threshold(feature_thresholds[81]), .feature_above(feature_aboves[81]), .feature_below(feature_belows[81]), .scan_win_std_dev(scan_win_std_dev[81]), .feature_accum(feature_accums[81]));
  accum_calculator ac82(.scan_win(scan_win82), .rectangle1_x(rectangle1_xs[82]), .rectangle1_y(rectangle1_ys[82]), .rectangle1_width(rectangle1_widths[82]), .rectangle1_height(rectangle1_heights[82]), .rectangle1_weight(rectangle1_weights[82]), .rectangle2_x(rectangle2_xs[82]), .rectangle2_y(rectangle2_ys[82]), .rectangle2_width(rectangle2_widths[82]), .rectangle2_height(rectangle2_heights[82]), .rectangle2_weight(rectangle2_weights[82]), .rectangle3_x(rectangle3_xs[82]), .rectangle3_y(rectangle3_ys[82]), .rectangle3_width(rectangle3_widths[82]), .rectangle3_height(rectangle3_heights[82]), .rectangle3_weight(rectangle3_weights[82]), .feature_threshold(feature_thresholds[82]), .feature_above(feature_aboves[82]), .feature_below(feature_belows[82]), .scan_win_std_dev(scan_win_std_dev[82]), .feature_accum(feature_accums[82]));
  accum_calculator ac83(.scan_win(scan_win83), .rectangle1_x(rectangle1_xs[83]), .rectangle1_y(rectangle1_ys[83]), .rectangle1_width(rectangle1_widths[83]), .rectangle1_height(rectangle1_heights[83]), .rectangle1_weight(rectangle1_weights[83]), .rectangle2_x(rectangle2_xs[83]), .rectangle2_y(rectangle2_ys[83]), .rectangle2_width(rectangle2_widths[83]), .rectangle2_height(rectangle2_heights[83]), .rectangle2_weight(rectangle2_weights[83]), .rectangle3_x(rectangle3_xs[83]), .rectangle3_y(rectangle3_ys[83]), .rectangle3_width(rectangle3_widths[83]), .rectangle3_height(rectangle3_heights[83]), .rectangle3_weight(rectangle3_weights[83]), .feature_threshold(feature_thresholds[83]), .feature_above(feature_aboves[83]), .feature_below(feature_belows[83]), .scan_win_std_dev(scan_win_std_dev[83]), .feature_accum(feature_accums[83]));
  accum_calculator ac84(.scan_win(scan_win84), .rectangle1_x(rectangle1_xs[84]), .rectangle1_y(rectangle1_ys[84]), .rectangle1_width(rectangle1_widths[84]), .rectangle1_height(rectangle1_heights[84]), .rectangle1_weight(rectangle1_weights[84]), .rectangle2_x(rectangle2_xs[84]), .rectangle2_y(rectangle2_ys[84]), .rectangle2_width(rectangle2_widths[84]), .rectangle2_height(rectangle2_heights[84]), .rectangle2_weight(rectangle2_weights[84]), .rectangle3_x(rectangle3_xs[84]), .rectangle3_y(rectangle3_ys[84]), .rectangle3_width(rectangle3_widths[84]), .rectangle3_height(rectangle3_heights[84]), .rectangle3_weight(rectangle3_weights[84]), .feature_threshold(feature_thresholds[84]), .feature_above(feature_aboves[84]), .feature_below(feature_belows[84]), .scan_win_std_dev(scan_win_std_dev[84]), .feature_accum(feature_accums[84]));
  accum_calculator ac85(.scan_win(scan_win85), .rectangle1_x(rectangle1_xs[85]), .rectangle1_y(rectangle1_ys[85]), .rectangle1_width(rectangle1_widths[85]), .rectangle1_height(rectangle1_heights[85]), .rectangle1_weight(rectangle1_weights[85]), .rectangle2_x(rectangle2_xs[85]), .rectangle2_y(rectangle2_ys[85]), .rectangle2_width(rectangle2_widths[85]), .rectangle2_height(rectangle2_heights[85]), .rectangle2_weight(rectangle2_weights[85]), .rectangle3_x(rectangle3_xs[85]), .rectangle3_y(rectangle3_ys[85]), .rectangle3_width(rectangle3_widths[85]), .rectangle3_height(rectangle3_heights[85]), .rectangle3_weight(rectangle3_weights[85]), .feature_threshold(feature_thresholds[85]), .feature_above(feature_aboves[85]), .feature_below(feature_belows[85]), .scan_win_std_dev(scan_win_std_dev[85]), .feature_accum(feature_accums[85]));
  accum_calculator ac86(.scan_win(scan_win86), .rectangle1_x(rectangle1_xs[86]), .rectangle1_y(rectangle1_ys[86]), .rectangle1_width(rectangle1_widths[86]), .rectangle1_height(rectangle1_heights[86]), .rectangle1_weight(rectangle1_weights[86]), .rectangle2_x(rectangle2_xs[86]), .rectangle2_y(rectangle2_ys[86]), .rectangle2_width(rectangle2_widths[86]), .rectangle2_height(rectangle2_heights[86]), .rectangle2_weight(rectangle2_weights[86]), .rectangle3_x(rectangle3_xs[86]), .rectangle3_y(rectangle3_ys[86]), .rectangle3_width(rectangle3_widths[86]), .rectangle3_height(rectangle3_heights[86]), .rectangle3_weight(rectangle3_weights[86]), .feature_threshold(feature_thresholds[86]), .feature_above(feature_aboves[86]), .feature_below(feature_belows[86]), .scan_win_std_dev(scan_win_std_dev[86]), .feature_accum(feature_accums[86]));
  accum_calculator ac87(.scan_win(scan_win87), .rectangle1_x(rectangle1_xs[87]), .rectangle1_y(rectangle1_ys[87]), .rectangle1_width(rectangle1_widths[87]), .rectangle1_height(rectangle1_heights[87]), .rectangle1_weight(rectangle1_weights[87]), .rectangle2_x(rectangle2_xs[87]), .rectangle2_y(rectangle2_ys[87]), .rectangle2_width(rectangle2_widths[87]), .rectangle2_height(rectangle2_heights[87]), .rectangle2_weight(rectangle2_weights[87]), .rectangle3_x(rectangle3_xs[87]), .rectangle3_y(rectangle3_ys[87]), .rectangle3_width(rectangle3_widths[87]), .rectangle3_height(rectangle3_heights[87]), .rectangle3_weight(rectangle3_weights[87]), .feature_threshold(feature_thresholds[87]), .feature_above(feature_aboves[87]), .feature_below(feature_belows[87]), .scan_win_std_dev(scan_win_std_dev[87]), .feature_accum(feature_accums[87]));
  accum_calculator ac88(.scan_win(scan_win88), .rectangle1_x(rectangle1_xs[88]), .rectangle1_y(rectangle1_ys[88]), .rectangle1_width(rectangle1_widths[88]), .rectangle1_height(rectangle1_heights[88]), .rectangle1_weight(rectangle1_weights[88]), .rectangle2_x(rectangle2_xs[88]), .rectangle2_y(rectangle2_ys[88]), .rectangle2_width(rectangle2_widths[88]), .rectangle2_height(rectangle2_heights[88]), .rectangle2_weight(rectangle2_weights[88]), .rectangle3_x(rectangle3_xs[88]), .rectangle3_y(rectangle3_ys[88]), .rectangle3_width(rectangle3_widths[88]), .rectangle3_height(rectangle3_heights[88]), .rectangle3_weight(rectangle3_weights[88]), .feature_threshold(feature_thresholds[88]), .feature_above(feature_aboves[88]), .feature_below(feature_belows[88]), .scan_win_std_dev(scan_win_std_dev[88]), .feature_accum(feature_accums[88]));
  accum_calculator ac89(.scan_win(scan_win89), .rectangle1_x(rectangle1_xs[89]), .rectangle1_y(rectangle1_ys[89]), .rectangle1_width(rectangle1_widths[89]), .rectangle1_height(rectangle1_heights[89]), .rectangle1_weight(rectangle1_weights[89]), .rectangle2_x(rectangle2_xs[89]), .rectangle2_y(rectangle2_ys[89]), .rectangle2_width(rectangle2_widths[89]), .rectangle2_height(rectangle2_heights[89]), .rectangle2_weight(rectangle2_weights[89]), .rectangle3_x(rectangle3_xs[89]), .rectangle3_y(rectangle3_ys[89]), .rectangle3_width(rectangle3_widths[89]), .rectangle3_height(rectangle3_heights[89]), .rectangle3_weight(rectangle3_weights[89]), .feature_threshold(feature_thresholds[89]), .feature_above(feature_aboves[89]), .feature_below(feature_belows[89]), .scan_win_std_dev(scan_win_std_dev[89]), .feature_accum(feature_accums[89]));
  accum_calculator ac90(.scan_win(scan_win90), .rectangle1_x(rectangle1_xs[90]), .rectangle1_y(rectangle1_ys[90]), .rectangle1_width(rectangle1_widths[90]), .rectangle1_height(rectangle1_heights[90]), .rectangle1_weight(rectangle1_weights[90]), .rectangle2_x(rectangle2_xs[90]), .rectangle2_y(rectangle2_ys[90]), .rectangle2_width(rectangle2_widths[90]), .rectangle2_height(rectangle2_heights[90]), .rectangle2_weight(rectangle2_weights[90]), .rectangle3_x(rectangle3_xs[90]), .rectangle3_y(rectangle3_ys[90]), .rectangle3_width(rectangle3_widths[90]), .rectangle3_height(rectangle3_heights[90]), .rectangle3_weight(rectangle3_weights[90]), .feature_threshold(feature_thresholds[90]), .feature_above(feature_aboves[90]), .feature_below(feature_belows[90]), .scan_win_std_dev(scan_win_std_dev[90]), .feature_accum(feature_accums[90]));
  accum_calculator ac91(.scan_win(scan_win91), .rectangle1_x(rectangle1_xs[91]), .rectangle1_y(rectangle1_ys[91]), .rectangle1_width(rectangle1_widths[91]), .rectangle1_height(rectangle1_heights[91]), .rectangle1_weight(rectangle1_weights[91]), .rectangle2_x(rectangle2_xs[91]), .rectangle2_y(rectangle2_ys[91]), .rectangle2_width(rectangle2_widths[91]), .rectangle2_height(rectangle2_heights[91]), .rectangle2_weight(rectangle2_weights[91]), .rectangle3_x(rectangle3_xs[91]), .rectangle3_y(rectangle3_ys[91]), .rectangle3_width(rectangle3_widths[91]), .rectangle3_height(rectangle3_heights[91]), .rectangle3_weight(rectangle3_weights[91]), .feature_threshold(feature_thresholds[91]), .feature_above(feature_aboves[91]), .feature_below(feature_belows[91]), .scan_win_std_dev(scan_win_std_dev[91]), .feature_accum(feature_accums[91]));
  accum_calculator ac92(.scan_win(scan_win92), .rectangle1_x(rectangle1_xs[92]), .rectangle1_y(rectangle1_ys[92]), .rectangle1_width(rectangle1_widths[92]), .rectangle1_height(rectangle1_heights[92]), .rectangle1_weight(rectangle1_weights[92]), .rectangle2_x(rectangle2_xs[92]), .rectangle2_y(rectangle2_ys[92]), .rectangle2_width(rectangle2_widths[92]), .rectangle2_height(rectangle2_heights[92]), .rectangle2_weight(rectangle2_weights[92]), .rectangle3_x(rectangle3_xs[92]), .rectangle3_y(rectangle3_ys[92]), .rectangle3_width(rectangle3_widths[92]), .rectangle3_height(rectangle3_heights[92]), .rectangle3_weight(rectangle3_weights[92]), .feature_threshold(feature_thresholds[92]), .feature_above(feature_aboves[92]), .feature_below(feature_belows[92]), .scan_win_std_dev(scan_win_std_dev[92]), .feature_accum(feature_accums[92]));
  accum_calculator ac93(.scan_win(scan_win93), .rectangle1_x(rectangle1_xs[93]), .rectangle1_y(rectangle1_ys[93]), .rectangle1_width(rectangle1_widths[93]), .rectangle1_height(rectangle1_heights[93]), .rectangle1_weight(rectangle1_weights[93]), .rectangle2_x(rectangle2_xs[93]), .rectangle2_y(rectangle2_ys[93]), .rectangle2_width(rectangle2_widths[93]), .rectangle2_height(rectangle2_heights[93]), .rectangle2_weight(rectangle2_weights[93]), .rectangle3_x(rectangle3_xs[93]), .rectangle3_y(rectangle3_ys[93]), .rectangle3_width(rectangle3_widths[93]), .rectangle3_height(rectangle3_heights[93]), .rectangle3_weight(rectangle3_weights[93]), .feature_threshold(feature_thresholds[93]), .feature_above(feature_aboves[93]), .feature_below(feature_belows[93]), .scan_win_std_dev(scan_win_std_dev[93]), .feature_accum(feature_accums[93]));
  accum_calculator ac94(.scan_win(scan_win94), .rectangle1_x(rectangle1_xs[94]), .rectangle1_y(rectangle1_ys[94]), .rectangle1_width(rectangle1_widths[94]), .rectangle1_height(rectangle1_heights[94]), .rectangle1_weight(rectangle1_weights[94]), .rectangle2_x(rectangle2_xs[94]), .rectangle2_y(rectangle2_ys[94]), .rectangle2_width(rectangle2_widths[94]), .rectangle2_height(rectangle2_heights[94]), .rectangle2_weight(rectangle2_weights[94]), .rectangle3_x(rectangle3_xs[94]), .rectangle3_y(rectangle3_ys[94]), .rectangle3_width(rectangle3_widths[94]), .rectangle3_height(rectangle3_heights[94]), .rectangle3_weight(rectangle3_weights[94]), .feature_threshold(feature_thresholds[94]), .feature_above(feature_aboves[94]), .feature_below(feature_belows[94]), .scan_win_std_dev(scan_win_std_dev[94]), .feature_accum(feature_accums[94]));
  accum_calculator ac95(.scan_win(scan_win95), .rectangle1_x(rectangle1_xs[95]), .rectangle1_y(rectangle1_ys[95]), .rectangle1_width(rectangle1_widths[95]), .rectangle1_height(rectangle1_heights[95]), .rectangle1_weight(rectangle1_weights[95]), .rectangle2_x(rectangle2_xs[95]), .rectangle2_y(rectangle2_ys[95]), .rectangle2_width(rectangle2_widths[95]), .rectangle2_height(rectangle2_heights[95]), .rectangle2_weight(rectangle2_weights[95]), .rectangle3_x(rectangle3_xs[95]), .rectangle3_y(rectangle3_ys[95]), .rectangle3_width(rectangle3_widths[95]), .rectangle3_height(rectangle3_heights[95]), .rectangle3_weight(rectangle3_weights[95]), .feature_threshold(feature_thresholds[95]), .feature_above(feature_aboves[95]), .feature_below(feature_belows[95]), .scan_win_std_dev(scan_win_std_dev[95]), .feature_accum(feature_accums[95]));
  accum_calculator ac96(.scan_win(scan_win96), .rectangle1_x(rectangle1_xs[96]), .rectangle1_y(rectangle1_ys[96]), .rectangle1_width(rectangle1_widths[96]), .rectangle1_height(rectangle1_heights[96]), .rectangle1_weight(rectangle1_weights[96]), .rectangle2_x(rectangle2_xs[96]), .rectangle2_y(rectangle2_ys[96]), .rectangle2_width(rectangle2_widths[96]), .rectangle2_height(rectangle2_heights[96]), .rectangle2_weight(rectangle2_weights[96]), .rectangle3_x(rectangle3_xs[96]), .rectangle3_y(rectangle3_ys[96]), .rectangle3_width(rectangle3_widths[96]), .rectangle3_height(rectangle3_heights[96]), .rectangle3_weight(rectangle3_weights[96]), .feature_threshold(feature_thresholds[96]), .feature_above(feature_aboves[96]), .feature_below(feature_belows[96]), .scan_win_std_dev(scan_win_std_dev[96]), .feature_accum(feature_accums[96]));
  accum_calculator ac97(.scan_win(scan_win97), .rectangle1_x(rectangle1_xs[97]), .rectangle1_y(rectangle1_ys[97]), .rectangle1_width(rectangle1_widths[97]), .rectangle1_height(rectangle1_heights[97]), .rectangle1_weight(rectangle1_weights[97]), .rectangle2_x(rectangle2_xs[97]), .rectangle2_y(rectangle2_ys[97]), .rectangle2_width(rectangle2_widths[97]), .rectangle2_height(rectangle2_heights[97]), .rectangle2_weight(rectangle2_weights[97]), .rectangle3_x(rectangle3_xs[97]), .rectangle3_y(rectangle3_ys[97]), .rectangle3_width(rectangle3_widths[97]), .rectangle3_height(rectangle3_heights[97]), .rectangle3_weight(rectangle3_weights[97]), .feature_threshold(feature_thresholds[97]), .feature_above(feature_aboves[97]), .feature_below(feature_belows[97]), .scan_win_std_dev(scan_win_std_dev[97]), .feature_accum(feature_accums[97]));
  accum_calculator ac98(.scan_win(scan_win98), .rectangle1_x(rectangle1_xs[98]), .rectangle1_y(rectangle1_ys[98]), .rectangle1_width(rectangle1_widths[98]), .rectangle1_height(rectangle1_heights[98]), .rectangle1_weight(rectangle1_weights[98]), .rectangle2_x(rectangle2_xs[98]), .rectangle2_y(rectangle2_ys[98]), .rectangle2_width(rectangle2_widths[98]), .rectangle2_height(rectangle2_heights[98]), .rectangle2_weight(rectangle2_weights[98]), .rectangle3_x(rectangle3_xs[98]), .rectangle3_y(rectangle3_ys[98]), .rectangle3_width(rectangle3_widths[98]), .rectangle3_height(rectangle3_heights[98]), .rectangle3_weight(rectangle3_weights[98]), .feature_threshold(feature_thresholds[98]), .feature_above(feature_aboves[98]), .feature_below(feature_belows[98]), .scan_win_std_dev(scan_win_std_dev[98]), .feature_accum(feature_accums[98]));
  accum_calculator ac99(.scan_win(scan_win99), .rectangle1_x(rectangle1_xs[99]), .rectangle1_y(rectangle1_ys[99]), .rectangle1_width(rectangle1_widths[99]), .rectangle1_height(rectangle1_heights[99]), .rectangle1_weight(rectangle1_weights[99]), .rectangle2_x(rectangle2_xs[99]), .rectangle2_y(rectangle2_ys[99]), .rectangle2_width(rectangle2_widths[99]), .rectangle2_height(rectangle2_heights[99]), .rectangle2_weight(rectangle2_weights[99]), .rectangle3_x(rectangle3_xs[99]), .rectangle3_y(rectangle3_ys[99]), .rectangle3_width(rectangle3_widths[99]), .rectangle3_height(rectangle3_heights[99]), .rectangle3_weight(rectangle3_weights[99]), .feature_threshold(feature_thresholds[99]), .feature_above(feature_aboves[99]), .feature_below(feature_belows[99]), .scan_win_std_dev(scan_win_std_dev[99]), .feature_accum(feature_accums[99]));
  accum_calculator ac100(.scan_win(scan_win100), .rectangle1_x(rectangle1_xs[100]), .rectangle1_y(rectangle1_ys[100]), .rectangle1_width(rectangle1_widths[100]), .rectangle1_height(rectangle1_heights[100]), .rectangle1_weight(rectangle1_weights[100]), .rectangle2_x(rectangle2_xs[100]), .rectangle2_y(rectangle2_ys[100]), .rectangle2_width(rectangle2_widths[100]), .rectangle2_height(rectangle2_heights[100]), .rectangle2_weight(rectangle2_weights[100]), .rectangle3_x(rectangle3_xs[100]), .rectangle3_y(rectangle3_ys[100]), .rectangle3_width(rectangle3_widths[100]), .rectangle3_height(rectangle3_heights[100]), .rectangle3_weight(rectangle3_weights[100]), .feature_threshold(feature_thresholds[100]), .feature_above(feature_aboves[100]), .feature_below(feature_belows[100]), .scan_win_std_dev(scan_win_std_dev[100]), .feature_accum(feature_accums[100]));
  accum_calculator ac101(.scan_win(scan_win101), .rectangle1_x(rectangle1_xs[101]), .rectangle1_y(rectangle1_ys[101]), .rectangle1_width(rectangle1_widths[101]), .rectangle1_height(rectangle1_heights[101]), .rectangle1_weight(rectangle1_weights[101]), .rectangle2_x(rectangle2_xs[101]), .rectangle2_y(rectangle2_ys[101]), .rectangle2_width(rectangle2_widths[101]), .rectangle2_height(rectangle2_heights[101]), .rectangle2_weight(rectangle2_weights[101]), .rectangle3_x(rectangle3_xs[101]), .rectangle3_y(rectangle3_ys[101]), .rectangle3_width(rectangle3_widths[101]), .rectangle3_height(rectangle3_heights[101]), .rectangle3_weight(rectangle3_weights[101]), .feature_threshold(feature_thresholds[101]), .feature_above(feature_aboves[101]), .feature_below(feature_belows[101]), .scan_win_std_dev(scan_win_std_dev[101]), .feature_accum(feature_accums[101]));
  accum_calculator ac102(.scan_win(scan_win102), .rectangle1_x(rectangle1_xs[102]), .rectangle1_y(rectangle1_ys[102]), .rectangle1_width(rectangle1_widths[102]), .rectangle1_height(rectangle1_heights[102]), .rectangle1_weight(rectangle1_weights[102]), .rectangle2_x(rectangle2_xs[102]), .rectangle2_y(rectangle2_ys[102]), .rectangle2_width(rectangle2_widths[102]), .rectangle2_height(rectangle2_heights[102]), .rectangle2_weight(rectangle2_weights[102]), .rectangle3_x(rectangle3_xs[102]), .rectangle3_y(rectangle3_ys[102]), .rectangle3_width(rectangle3_widths[102]), .rectangle3_height(rectangle3_heights[102]), .rectangle3_weight(rectangle3_weights[102]), .feature_threshold(feature_thresholds[102]), .feature_above(feature_aboves[102]), .feature_below(feature_belows[102]), .scan_win_std_dev(scan_win_std_dev[102]), .feature_accum(feature_accums[102]));
  accum_calculator ac103(.scan_win(scan_win103), .rectangle1_x(rectangle1_xs[103]), .rectangle1_y(rectangle1_ys[103]), .rectangle1_width(rectangle1_widths[103]), .rectangle1_height(rectangle1_heights[103]), .rectangle1_weight(rectangle1_weights[103]), .rectangle2_x(rectangle2_xs[103]), .rectangle2_y(rectangle2_ys[103]), .rectangle2_width(rectangle2_widths[103]), .rectangle2_height(rectangle2_heights[103]), .rectangle2_weight(rectangle2_weights[103]), .rectangle3_x(rectangle3_xs[103]), .rectangle3_y(rectangle3_ys[103]), .rectangle3_width(rectangle3_widths[103]), .rectangle3_height(rectangle3_heights[103]), .rectangle3_weight(rectangle3_weights[103]), .feature_threshold(feature_thresholds[103]), .feature_above(feature_aboves[103]), .feature_below(feature_belows[103]), .scan_win_std_dev(scan_win_std_dev[103]), .feature_accum(feature_accums[103]));
  accum_calculator ac104(.scan_win(scan_win104), .rectangle1_x(rectangle1_xs[104]), .rectangle1_y(rectangle1_ys[104]), .rectangle1_width(rectangle1_widths[104]), .rectangle1_height(rectangle1_heights[104]), .rectangle1_weight(rectangle1_weights[104]), .rectangle2_x(rectangle2_xs[104]), .rectangle2_y(rectangle2_ys[104]), .rectangle2_width(rectangle2_widths[104]), .rectangle2_height(rectangle2_heights[104]), .rectangle2_weight(rectangle2_weights[104]), .rectangle3_x(rectangle3_xs[104]), .rectangle3_y(rectangle3_ys[104]), .rectangle3_width(rectangle3_widths[104]), .rectangle3_height(rectangle3_heights[104]), .rectangle3_weight(rectangle3_weights[104]), .feature_threshold(feature_thresholds[104]), .feature_above(feature_aboves[104]), .feature_below(feature_belows[104]), .scan_win_std_dev(scan_win_std_dev[104]), .feature_accum(feature_accums[104]));
  accum_calculator ac105(.scan_win(scan_win105), .rectangle1_x(rectangle1_xs[105]), .rectangle1_y(rectangle1_ys[105]), .rectangle1_width(rectangle1_widths[105]), .rectangle1_height(rectangle1_heights[105]), .rectangle1_weight(rectangle1_weights[105]), .rectangle2_x(rectangle2_xs[105]), .rectangle2_y(rectangle2_ys[105]), .rectangle2_width(rectangle2_widths[105]), .rectangle2_height(rectangle2_heights[105]), .rectangle2_weight(rectangle2_weights[105]), .rectangle3_x(rectangle3_xs[105]), .rectangle3_y(rectangle3_ys[105]), .rectangle3_width(rectangle3_widths[105]), .rectangle3_height(rectangle3_heights[105]), .rectangle3_weight(rectangle3_weights[105]), .feature_threshold(feature_thresholds[105]), .feature_above(feature_aboves[105]), .feature_below(feature_belows[105]), .scan_win_std_dev(scan_win_std_dev[105]), .feature_accum(feature_accums[105]));
  accum_calculator ac106(.scan_win(scan_win106), .rectangle1_x(rectangle1_xs[106]), .rectangle1_y(rectangle1_ys[106]), .rectangle1_width(rectangle1_widths[106]), .rectangle1_height(rectangle1_heights[106]), .rectangle1_weight(rectangle1_weights[106]), .rectangle2_x(rectangle2_xs[106]), .rectangle2_y(rectangle2_ys[106]), .rectangle2_width(rectangle2_widths[106]), .rectangle2_height(rectangle2_heights[106]), .rectangle2_weight(rectangle2_weights[106]), .rectangle3_x(rectangle3_xs[106]), .rectangle3_y(rectangle3_ys[106]), .rectangle3_width(rectangle3_widths[106]), .rectangle3_height(rectangle3_heights[106]), .rectangle3_weight(rectangle3_weights[106]), .feature_threshold(feature_thresholds[106]), .feature_above(feature_aboves[106]), .feature_below(feature_belows[106]), .scan_win_std_dev(scan_win_std_dev[106]), .feature_accum(feature_accums[106]));
  accum_calculator ac107(.scan_win(scan_win107), .rectangle1_x(rectangle1_xs[107]), .rectangle1_y(rectangle1_ys[107]), .rectangle1_width(rectangle1_widths[107]), .rectangle1_height(rectangle1_heights[107]), .rectangle1_weight(rectangle1_weights[107]), .rectangle2_x(rectangle2_xs[107]), .rectangle2_y(rectangle2_ys[107]), .rectangle2_width(rectangle2_widths[107]), .rectangle2_height(rectangle2_heights[107]), .rectangle2_weight(rectangle2_weights[107]), .rectangle3_x(rectangle3_xs[107]), .rectangle3_y(rectangle3_ys[107]), .rectangle3_width(rectangle3_widths[107]), .rectangle3_height(rectangle3_heights[107]), .rectangle3_weight(rectangle3_weights[107]), .feature_threshold(feature_thresholds[107]), .feature_above(feature_aboves[107]), .feature_below(feature_belows[107]), .scan_win_std_dev(scan_win_std_dev[107]), .feature_accum(feature_accums[107]));
  accum_calculator ac108(.scan_win(scan_win108), .rectangle1_x(rectangle1_xs[108]), .rectangle1_y(rectangle1_ys[108]), .rectangle1_width(rectangle1_widths[108]), .rectangle1_height(rectangle1_heights[108]), .rectangle1_weight(rectangle1_weights[108]), .rectangle2_x(rectangle2_xs[108]), .rectangle2_y(rectangle2_ys[108]), .rectangle2_width(rectangle2_widths[108]), .rectangle2_height(rectangle2_heights[108]), .rectangle2_weight(rectangle2_weights[108]), .rectangle3_x(rectangle3_xs[108]), .rectangle3_y(rectangle3_ys[108]), .rectangle3_width(rectangle3_widths[108]), .rectangle3_height(rectangle3_heights[108]), .rectangle3_weight(rectangle3_weights[108]), .feature_threshold(feature_thresholds[108]), .feature_above(feature_aboves[108]), .feature_below(feature_belows[108]), .scan_win_std_dev(scan_win_std_dev[108]), .feature_accum(feature_accums[108]));
  accum_calculator ac109(.scan_win(scan_win109), .rectangle1_x(rectangle1_xs[109]), .rectangle1_y(rectangle1_ys[109]), .rectangle1_width(rectangle1_widths[109]), .rectangle1_height(rectangle1_heights[109]), .rectangle1_weight(rectangle1_weights[109]), .rectangle2_x(rectangle2_xs[109]), .rectangle2_y(rectangle2_ys[109]), .rectangle2_width(rectangle2_widths[109]), .rectangle2_height(rectangle2_heights[109]), .rectangle2_weight(rectangle2_weights[109]), .rectangle3_x(rectangle3_xs[109]), .rectangle3_y(rectangle3_ys[109]), .rectangle3_width(rectangle3_widths[109]), .rectangle3_height(rectangle3_heights[109]), .rectangle3_weight(rectangle3_weights[109]), .feature_threshold(feature_thresholds[109]), .feature_above(feature_aboves[109]), .feature_below(feature_belows[109]), .scan_win_std_dev(scan_win_std_dev[109]), .feature_accum(feature_accums[109]));
  accum_calculator ac110(.scan_win(scan_win110), .rectangle1_x(rectangle1_xs[110]), .rectangle1_y(rectangle1_ys[110]), .rectangle1_width(rectangle1_widths[110]), .rectangle1_height(rectangle1_heights[110]), .rectangle1_weight(rectangle1_weights[110]), .rectangle2_x(rectangle2_xs[110]), .rectangle2_y(rectangle2_ys[110]), .rectangle2_width(rectangle2_widths[110]), .rectangle2_height(rectangle2_heights[110]), .rectangle2_weight(rectangle2_weights[110]), .rectangle3_x(rectangle3_xs[110]), .rectangle3_y(rectangle3_ys[110]), .rectangle3_width(rectangle3_widths[110]), .rectangle3_height(rectangle3_heights[110]), .rectangle3_weight(rectangle3_weights[110]), .feature_threshold(feature_thresholds[110]), .feature_above(feature_aboves[110]), .feature_below(feature_belows[110]), .scan_win_std_dev(scan_win_std_dev[110]), .feature_accum(feature_accums[110]));
  accum_calculator ac111(.scan_win(scan_win111), .rectangle1_x(rectangle1_xs[111]), .rectangle1_y(rectangle1_ys[111]), .rectangle1_width(rectangle1_widths[111]), .rectangle1_height(rectangle1_heights[111]), .rectangle1_weight(rectangle1_weights[111]), .rectangle2_x(rectangle2_xs[111]), .rectangle2_y(rectangle2_ys[111]), .rectangle2_width(rectangle2_widths[111]), .rectangle2_height(rectangle2_heights[111]), .rectangle2_weight(rectangle2_weights[111]), .rectangle3_x(rectangle3_xs[111]), .rectangle3_y(rectangle3_ys[111]), .rectangle3_width(rectangle3_widths[111]), .rectangle3_height(rectangle3_heights[111]), .rectangle3_weight(rectangle3_weights[111]), .feature_threshold(feature_thresholds[111]), .feature_above(feature_aboves[111]), .feature_below(feature_belows[111]), .scan_win_std_dev(scan_win_std_dev[111]), .feature_accum(feature_accums[111]));
  accum_calculator ac112(.scan_win(scan_win112), .rectangle1_x(rectangle1_xs[112]), .rectangle1_y(rectangle1_ys[112]), .rectangle1_width(rectangle1_widths[112]), .rectangle1_height(rectangle1_heights[112]), .rectangle1_weight(rectangle1_weights[112]), .rectangle2_x(rectangle2_xs[112]), .rectangle2_y(rectangle2_ys[112]), .rectangle2_width(rectangle2_widths[112]), .rectangle2_height(rectangle2_heights[112]), .rectangle2_weight(rectangle2_weights[112]), .rectangle3_x(rectangle3_xs[112]), .rectangle3_y(rectangle3_ys[112]), .rectangle3_width(rectangle3_widths[112]), .rectangle3_height(rectangle3_heights[112]), .rectangle3_weight(rectangle3_weights[112]), .feature_threshold(feature_thresholds[112]), .feature_above(feature_aboves[112]), .feature_below(feature_belows[112]), .scan_win_std_dev(scan_win_std_dev[112]), .feature_accum(feature_accums[112]));
  accum_calculator ac113(.scan_win(scan_win113), .rectangle1_x(rectangle1_xs[113]), .rectangle1_y(rectangle1_ys[113]), .rectangle1_width(rectangle1_widths[113]), .rectangle1_height(rectangle1_heights[113]), .rectangle1_weight(rectangle1_weights[113]), .rectangle2_x(rectangle2_xs[113]), .rectangle2_y(rectangle2_ys[113]), .rectangle2_width(rectangle2_widths[113]), .rectangle2_height(rectangle2_heights[113]), .rectangle2_weight(rectangle2_weights[113]), .rectangle3_x(rectangle3_xs[113]), .rectangle3_y(rectangle3_ys[113]), .rectangle3_width(rectangle3_widths[113]), .rectangle3_height(rectangle3_heights[113]), .rectangle3_weight(rectangle3_weights[113]), .feature_threshold(feature_thresholds[113]), .feature_above(feature_aboves[113]), .feature_below(feature_belows[113]), .scan_win_std_dev(scan_win_std_dev[113]), .feature_accum(feature_accums[113]));
  accum_calculator ac114(.scan_win(scan_win114), .rectangle1_x(rectangle1_xs[114]), .rectangle1_y(rectangle1_ys[114]), .rectangle1_width(rectangle1_widths[114]), .rectangle1_height(rectangle1_heights[114]), .rectangle1_weight(rectangle1_weights[114]), .rectangle2_x(rectangle2_xs[114]), .rectangle2_y(rectangle2_ys[114]), .rectangle2_width(rectangle2_widths[114]), .rectangle2_height(rectangle2_heights[114]), .rectangle2_weight(rectangle2_weights[114]), .rectangle3_x(rectangle3_xs[114]), .rectangle3_y(rectangle3_ys[114]), .rectangle3_width(rectangle3_widths[114]), .rectangle3_height(rectangle3_heights[114]), .rectangle3_weight(rectangle3_weights[114]), .feature_threshold(feature_thresholds[114]), .feature_above(feature_aboves[114]), .feature_below(feature_belows[114]), .scan_win_std_dev(scan_win_std_dev[114]), .feature_accum(feature_accums[114]));
  accum_calculator ac115(.scan_win(scan_win115), .rectangle1_x(rectangle1_xs[115]), .rectangle1_y(rectangle1_ys[115]), .rectangle1_width(rectangle1_widths[115]), .rectangle1_height(rectangle1_heights[115]), .rectangle1_weight(rectangle1_weights[115]), .rectangle2_x(rectangle2_xs[115]), .rectangle2_y(rectangle2_ys[115]), .rectangle2_width(rectangle2_widths[115]), .rectangle2_height(rectangle2_heights[115]), .rectangle2_weight(rectangle2_weights[115]), .rectangle3_x(rectangle3_xs[115]), .rectangle3_y(rectangle3_ys[115]), .rectangle3_width(rectangle3_widths[115]), .rectangle3_height(rectangle3_heights[115]), .rectangle3_weight(rectangle3_weights[115]), .feature_threshold(feature_thresholds[115]), .feature_above(feature_aboves[115]), .feature_below(feature_belows[115]), .scan_win_std_dev(scan_win_std_dev[115]), .feature_accum(feature_accums[115]));
  accum_calculator ac116(.scan_win(scan_win116), .rectangle1_x(rectangle1_xs[116]), .rectangle1_y(rectangle1_ys[116]), .rectangle1_width(rectangle1_widths[116]), .rectangle1_height(rectangle1_heights[116]), .rectangle1_weight(rectangle1_weights[116]), .rectangle2_x(rectangle2_xs[116]), .rectangle2_y(rectangle2_ys[116]), .rectangle2_width(rectangle2_widths[116]), .rectangle2_height(rectangle2_heights[116]), .rectangle2_weight(rectangle2_weights[116]), .rectangle3_x(rectangle3_xs[116]), .rectangle3_y(rectangle3_ys[116]), .rectangle3_width(rectangle3_widths[116]), .rectangle3_height(rectangle3_heights[116]), .rectangle3_weight(rectangle3_weights[116]), .feature_threshold(feature_thresholds[116]), .feature_above(feature_aboves[116]), .feature_below(feature_belows[116]), .scan_win_std_dev(scan_win_std_dev[116]), .feature_accum(feature_accums[116]));
  accum_calculator ac117(.scan_win(scan_win117), .rectangle1_x(rectangle1_xs[117]), .rectangle1_y(rectangle1_ys[117]), .rectangle1_width(rectangle1_widths[117]), .rectangle1_height(rectangle1_heights[117]), .rectangle1_weight(rectangle1_weights[117]), .rectangle2_x(rectangle2_xs[117]), .rectangle2_y(rectangle2_ys[117]), .rectangle2_width(rectangle2_widths[117]), .rectangle2_height(rectangle2_heights[117]), .rectangle2_weight(rectangle2_weights[117]), .rectangle3_x(rectangle3_xs[117]), .rectangle3_y(rectangle3_ys[117]), .rectangle3_width(rectangle3_widths[117]), .rectangle3_height(rectangle3_heights[117]), .rectangle3_weight(rectangle3_weights[117]), .feature_threshold(feature_thresholds[117]), .feature_above(feature_aboves[117]), .feature_below(feature_belows[117]), .scan_win_std_dev(scan_win_std_dev[117]), .feature_accum(feature_accums[117]));
  accum_calculator ac118(.scan_win(scan_win118), .rectangle1_x(rectangle1_xs[118]), .rectangle1_y(rectangle1_ys[118]), .rectangle1_width(rectangle1_widths[118]), .rectangle1_height(rectangle1_heights[118]), .rectangle1_weight(rectangle1_weights[118]), .rectangle2_x(rectangle2_xs[118]), .rectangle2_y(rectangle2_ys[118]), .rectangle2_width(rectangle2_widths[118]), .rectangle2_height(rectangle2_heights[118]), .rectangle2_weight(rectangle2_weights[118]), .rectangle3_x(rectangle3_xs[118]), .rectangle3_y(rectangle3_ys[118]), .rectangle3_width(rectangle3_widths[118]), .rectangle3_height(rectangle3_heights[118]), .rectangle3_weight(rectangle3_weights[118]), .feature_threshold(feature_thresholds[118]), .feature_above(feature_aboves[118]), .feature_below(feature_belows[118]), .scan_win_std_dev(scan_win_std_dev[118]), .feature_accum(feature_accums[118]));
  accum_calculator ac119(.scan_win(scan_win119), .rectangle1_x(rectangle1_xs[119]), .rectangle1_y(rectangle1_ys[119]), .rectangle1_width(rectangle1_widths[119]), .rectangle1_height(rectangle1_heights[119]), .rectangle1_weight(rectangle1_weights[119]), .rectangle2_x(rectangle2_xs[119]), .rectangle2_y(rectangle2_ys[119]), .rectangle2_width(rectangle2_widths[119]), .rectangle2_height(rectangle2_heights[119]), .rectangle2_weight(rectangle2_weights[119]), .rectangle3_x(rectangle3_xs[119]), .rectangle3_y(rectangle3_ys[119]), .rectangle3_width(rectangle3_widths[119]), .rectangle3_height(rectangle3_heights[119]), .rectangle3_weight(rectangle3_weights[119]), .feature_threshold(feature_thresholds[119]), .feature_above(feature_aboves[119]), .feature_below(feature_belows[119]), .scan_win_std_dev(scan_win_std_dev[119]), .feature_accum(feature_accums[119]));
  accum_calculator ac120(.scan_win(scan_win120), .rectangle1_x(rectangle1_xs[120]), .rectangle1_y(rectangle1_ys[120]), .rectangle1_width(rectangle1_widths[120]), .rectangle1_height(rectangle1_heights[120]), .rectangle1_weight(rectangle1_weights[120]), .rectangle2_x(rectangle2_xs[120]), .rectangle2_y(rectangle2_ys[120]), .rectangle2_width(rectangle2_widths[120]), .rectangle2_height(rectangle2_heights[120]), .rectangle2_weight(rectangle2_weights[120]), .rectangle3_x(rectangle3_xs[120]), .rectangle3_y(rectangle3_ys[120]), .rectangle3_width(rectangle3_widths[120]), .rectangle3_height(rectangle3_heights[120]), .rectangle3_weight(rectangle3_weights[120]), .feature_threshold(feature_thresholds[120]), .feature_above(feature_aboves[120]), .feature_below(feature_belows[120]), .scan_win_std_dev(scan_win_std_dev[120]), .feature_accum(feature_accums[120]));
  accum_calculator ac121(.scan_win(scan_win121), .rectangle1_x(rectangle1_xs[121]), .rectangle1_y(rectangle1_ys[121]), .rectangle1_width(rectangle1_widths[121]), .rectangle1_height(rectangle1_heights[121]), .rectangle1_weight(rectangle1_weights[121]), .rectangle2_x(rectangle2_xs[121]), .rectangle2_y(rectangle2_ys[121]), .rectangle2_width(rectangle2_widths[121]), .rectangle2_height(rectangle2_heights[121]), .rectangle2_weight(rectangle2_weights[121]), .rectangle3_x(rectangle3_xs[121]), .rectangle3_y(rectangle3_ys[121]), .rectangle3_width(rectangle3_widths[121]), .rectangle3_height(rectangle3_heights[121]), .rectangle3_weight(rectangle3_weights[121]), .feature_threshold(feature_thresholds[121]), .feature_above(feature_aboves[121]), .feature_below(feature_belows[121]), .scan_win_std_dev(scan_win_std_dev[121]), .feature_accum(feature_accums[121]));
  accum_calculator ac122(.scan_win(scan_win122), .rectangle1_x(rectangle1_xs[122]), .rectangle1_y(rectangle1_ys[122]), .rectangle1_width(rectangle1_widths[122]), .rectangle1_height(rectangle1_heights[122]), .rectangle1_weight(rectangle1_weights[122]), .rectangle2_x(rectangle2_xs[122]), .rectangle2_y(rectangle2_ys[122]), .rectangle2_width(rectangle2_widths[122]), .rectangle2_height(rectangle2_heights[122]), .rectangle2_weight(rectangle2_weights[122]), .rectangle3_x(rectangle3_xs[122]), .rectangle3_y(rectangle3_ys[122]), .rectangle3_width(rectangle3_widths[122]), .rectangle3_height(rectangle3_heights[122]), .rectangle3_weight(rectangle3_weights[122]), .feature_threshold(feature_thresholds[122]), .feature_above(feature_aboves[122]), .feature_below(feature_belows[122]), .scan_win_std_dev(scan_win_std_dev[122]), .feature_accum(feature_accums[122]));
  accum_calculator ac123(.scan_win(scan_win123), .rectangle1_x(rectangle1_xs[123]), .rectangle1_y(rectangle1_ys[123]), .rectangle1_width(rectangle1_widths[123]), .rectangle1_height(rectangle1_heights[123]), .rectangle1_weight(rectangle1_weights[123]), .rectangle2_x(rectangle2_xs[123]), .rectangle2_y(rectangle2_ys[123]), .rectangle2_width(rectangle2_widths[123]), .rectangle2_height(rectangle2_heights[123]), .rectangle2_weight(rectangle2_weights[123]), .rectangle3_x(rectangle3_xs[123]), .rectangle3_y(rectangle3_ys[123]), .rectangle3_width(rectangle3_widths[123]), .rectangle3_height(rectangle3_heights[123]), .rectangle3_weight(rectangle3_weights[123]), .feature_threshold(feature_thresholds[123]), .feature_above(feature_aboves[123]), .feature_below(feature_belows[123]), .scan_win_std_dev(scan_win_std_dev[123]), .feature_accum(feature_accums[123]));
  accum_calculator ac124(.scan_win(scan_win124), .rectangle1_x(rectangle1_xs[124]), .rectangle1_y(rectangle1_ys[124]), .rectangle1_width(rectangle1_widths[124]), .rectangle1_height(rectangle1_heights[124]), .rectangle1_weight(rectangle1_weights[124]), .rectangle2_x(rectangle2_xs[124]), .rectangle2_y(rectangle2_ys[124]), .rectangle2_width(rectangle2_widths[124]), .rectangle2_height(rectangle2_heights[124]), .rectangle2_weight(rectangle2_weights[124]), .rectangle3_x(rectangle3_xs[124]), .rectangle3_y(rectangle3_ys[124]), .rectangle3_width(rectangle3_widths[124]), .rectangle3_height(rectangle3_heights[124]), .rectangle3_weight(rectangle3_weights[124]), .feature_threshold(feature_thresholds[124]), .feature_above(feature_aboves[124]), .feature_below(feature_belows[124]), .scan_win_std_dev(scan_win_std_dev[124]), .feature_accum(feature_accums[124]));
  accum_calculator ac125(.scan_win(scan_win125), .rectangle1_x(rectangle1_xs[125]), .rectangle1_y(rectangle1_ys[125]), .rectangle1_width(rectangle1_widths[125]), .rectangle1_height(rectangle1_heights[125]), .rectangle1_weight(rectangle1_weights[125]), .rectangle2_x(rectangle2_xs[125]), .rectangle2_y(rectangle2_ys[125]), .rectangle2_width(rectangle2_widths[125]), .rectangle2_height(rectangle2_heights[125]), .rectangle2_weight(rectangle2_weights[125]), .rectangle3_x(rectangle3_xs[125]), .rectangle3_y(rectangle3_ys[125]), .rectangle3_width(rectangle3_widths[125]), .rectangle3_height(rectangle3_heights[125]), .rectangle3_weight(rectangle3_weights[125]), .feature_threshold(feature_thresholds[125]), .feature_above(feature_aboves[125]), .feature_below(feature_belows[125]), .scan_win_std_dev(scan_win_std_dev[125]), .feature_accum(feature_accums[125]));
  accum_calculator ac126(.scan_win(scan_win126), .rectangle1_x(rectangle1_xs[126]), .rectangle1_y(rectangle1_ys[126]), .rectangle1_width(rectangle1_widths[126]), .rectangle1_height(rectangle1_heights[126]), .rectangle1_weight(rectangle1_weights[126]), .rectangle2_x(rectangle2_xs[126]), .rectangle2_y(rectangle2_ys[126]), .rectangle2_width(rectangle2_widths[126]), .rectangle2_height(rectangle2_heights[126]), .rectangle2_weight(rectangle2_weights[126]), .rectangle3_x(rectangle3_xs[126]), .rectangle3_y(rectangle3_ys[126]), .rectangle3_width(rectangle3_widths[126]), .rectangle3_height(rectangle3_heights[126]), .rectangle3_weight(rectangle3_weights[126]), .feature_threshold(feature_thresholds[126]), .feature_above(feature_aboves[126]), .feature_below(feature_belows[126]), .scan_win_std_dev(scan_win_std_dev[126]), .feature_accum(feature_accums[126]));
  accum_calculator ac127(.scan_win(scan_win127), .rectangle1_x(rectangle1_xs[127]), .rectangle1_y(rectangle1_ys[127]), .rectangle1_width(rectangle1_widths[127]), .rectangle1_height(rectangle1_heights[127]), .rectangle1_weight(rectangle1_weights[127]), .rectangle2_x(rectangle2_xs[127]), .rectangle2_y(rectangle2_ys[127]), .rectangle2_width(rectangle2_widths[127]), .rectangle2_height(rectangle2_heights[127]), .rectangle2_weight(rectangle2_weights[127]), .rectangle3_x(rectangle3_xs[127]), .rectangle3_y(rectangle3_ys[127]), .rectangle3_width(rectangle3_widths[127]), .rectangle3_height(rectangle3_heights[127]), .rectangle3_weight(rectangle3_weights[127]), .feature_threshold(feature_thresholds[127]), .feature_above(feature_aboves[127]), .feature_below(feature_belows[127]), .scan_win_std_dev(scan_win_std_dev[127]), .feature_accum(feature_accums[127]));
  accum_calculator ac128(.scan_win(scan_win128), .rectangle1_x(rectangle1_xs[128]), .rectangle1_y(rectangle1_ys[128]), .rectangle1_width(rectangle1_widths[128]), .rectangle1_height(rectangle1_heights[128]), .rectangle1_weight(rectangle1_weights[128]), .rectangle2_x(rectangle2_xs[128]), .rectangle2_y(rectangle2_ys[128]), .rectangle2_width(rectangle2_widths[128]), .rectangle2_height(rectangle2_heights[128]), .rectangle2_weight(rectangle2_weights[128]), .rectangle3_x(rectangle3_xs[128]), .rectangle3_y(rectangle3_ys[128]), .rectangle3_width(rectangle3_widths[128]), .rectangle3_height(rectangle3_heights[128]), .rectangle3_weight(rectangle3_weights[128]), .feature_threshold(feature_thresholds[128]), .feature_above(feature_aboves[128]), .feature_below(feature_belows[128]), .scan_win_std_dev(scan_win_std_dev[128]), .feature_accum(feature_accums[128]));
  accum_calculator ac129(.scan_win(scan_win129), .rectangle1_x(rectangle1_xs[129]), .rectangle1_y(rectangle1_ys[129]), .rectangle1_width(rectangle1_widths[129]), .rectangle1_height(rectangle1_heights[129]), .rectangle1_weight(rectangle1_weights[129]), .rectangle2_x(rectangle2_xs[129]), .rectangle2_y(rectangle2_ys[129]), .rectangle2_width(rectangle2_widths[129]), .rectangle2_height(rectangle2_heights[129]), .rectangle2_weight(rectangle2_weights[129]), .rectangle3_x(rectangle3_xs[129]), .rectangle3_y(rectangle3_ys[129]), .rectangle3_width(rectangle3_widths[129]), .rectangle3_height(rectangle3_heights[129]), .rectangle3_weight(rectangle3_weights[129]), .feature_threshold(feature_thresholds[129]), .feature_above(feature_aboves[129]), .feature_below(feature_belows[129]), .scan_win_std_dev(scan_win_std_dev[129]), .feature_accum(feature_accums[129]));
  accum_calculator ac130(.scan_win(scan_win130), .rectangle1_x(rectangle1_xs[130]), .rectangle1_y(rectangle1_ys[130]), .rectangle1_width(rectangle1_widths[130]), .rectangle1_height(rectangle1_heights[130]), .rectangle1_weight(rectangle1_weights[130]), .rectangle2_x(rectangle2_xs[130]), .rectangle2_y(rectangle2_ys[130]), .rectangle2_width(rectangle2_widths[130]), .rectangle2_height(rectangle2_heights[130]), .rectangle2_weight(rectangle2_weights[130]), .rectangle3_x(rectangle3_xs[130]), .rectangle3_y(rectangle3_ys[130]), .rectangle3_width(rectangle3_widths[130]), .rectangle3_height(rectangle3_heights[130]), .rectangle3_weight(rectangle3_weights[130]), .feature_threshold(feature_thresholds[130]), .feature_above(feature_aboves[130]), .feature_below(feature_belows[130]), .scan_win_std_dev(scan_win_std_dev[130]), .feature_accum(feature_accums[130]));
  accum_calculator ac131(.scan_win(scan_win131), .rectangle1_x(rectangle1_xs[131]), .rectangle1_y(rectangle1_ys[131]), .rectangle1_width(rectangle1_widths[131]), .rectangle1_height(rectangle1_heights[131]), .rectangle1_weight(rectangle1_weights[131]), .rectangle2_x(rectangle2_xs[131]), .rectangle2_y(rectangle2_ys[131]), .rectangle2_width(rectangle2_widths[131]), .rectangle2_height(rectangle2_heights[131]), .rectangle2_weight(rectangle2_weights[131]), .rectangle3_x(rectangle3_xs[131]), .rectangle3_y(rectangle3_ys[131]), .rectangle3_width(rectangle3_widths[131]), .rectangle3_height(rectangle3_heights[131]), .rectangle3_weight(rectangle3_weights[131]), .feature_threshold(feature_thresholds[131]), .feature_above(feature_aboves[131]), .feature_below(feature_belows[131]), .scan_win_std_dev(scan_win_std_dev[131]), .feature_accum(feature_accums[131]));
  accum_calculator ac132(.scan_win(scan_win132), .rectangle1_x(rectangle1_xs[132]), .rectangle1_y(rectangle1_ys[132]), .rectangle1_width(rectangle1_widths[132]), .rectangle1_height(rectangle1_heights[132]), .rectangle1_weight(rectangle1_weights[132]), .rectangle2_x(rectangle2_xs[132]), .rectangle2_y(rectangle2_ys[132]), .rectangle2_width(rectangle2_widths[132]), .rectangle2_height(rectangle2_heights[132]), .rectangle2_weight(rectangle2_weights[132]), .rectangle3_x(rectangle3_xs[132]), .rectangle3_y(rectangle3_ys[132]), .rectangle3_width(rectangle3_widths[132]), .rectangle3_height(rectangle3_heights[132]), .rectangle3_weight(rectangle3_weights[132]), .feature_threshold(feature_thresholds[132]), .feature_above(feature_aboves[132]), .feature_below(feature_belows[132]), .scan_win_std_dev(scan_win_std_dev[132]), .feature_accum(feature_accums[132]));
  accum_calculator ac133(.scan_win(scan_win133), .rectangle1_x(rectangle1_xs[133]), .rectangle1_y(rectangle1_ys[133]), .rectangle1_width(rectangle1_widths[133]), .rectangle1_height(rectangle1_heights[133]), .rectangle1_weight(rectangle1_weights[133]), .rectangle2_x(rectangle2_xs[133]), .rectangle2_y(rectangle2_ys[133]), .rectangle2_width(rectangle2_widths[133]), .rectangle2_height(rectangle2_heights[133]), .rectangle2_weight(rectangle2_weights[133]), .rectangle3_x(rectangle3_xs[133]), .rectangle3_y(rectangle3_ys[133]), .rectangle3_width(rectangle3_widths[133]), .rectangle3_height(rectangle3_heights[133]), .rectangle3_weight(rectangle3_weights[133]), .feature_threshold(feature_thresholds[133]), .feature_above(feature_aboves[133]), .feature_below(feature_belows[133]), .scan_win_std_dev(scan_win_std_dev[133]), .feature_accum(feature_accums[133]));
  accum_calculator ac134(.scan_win(scan_win134), .rectangle1_x(rectangle1_xs[134]), .rectangle1_y(rectangle1_ys[134]), .rectangle1_width(rectangle1_widths[134]), .rectangle1_height(rectangle1_heights[134]), .rectangle1_weight(rectangle1_weights[134]), .rectangle2_x(rectangle2_xs[134]), .rectangle2_y(rectangle2_ys[134]), .rectangle2_width(rectangle2_widths[134]), .rectangle2_height(rectangle2_heights[134]), .rectangle2_weight(rectangle2_weights[134]), .rectangle3_x(rectangle3_xs[134]), .rectangle3_y(rectangle3_ys[134]), .rectangle3_width(rectangle3_widths[134]), .rectangle3_height(rectangle3_heights[134]), .rectangle3_weight(rectangle3_weights[134]), .feature_threshold(feature_thresholds[134]), .feature_above(feature_aboves[134]), .feature_below(feature_belows[134]), .scan_win_std_dev(scan_win_std_dev[134]), .feature_accum(feature_accums[134]));
  accum_calculator ac135(.scan_win(scan_win135), .rectangle1_x(rectangle1_xs[135]), .rectangle1_y(rectangle1_ys[135]), .rectangle1_width(rectangle1_widths[135]), .rectangle1_height(rectangle1_heights[135]), .rectangle1_weight(rectangle1_weights[135]), .rectangle2_x(rectangle2_xs[135]), .rectangle2_y(rectangle2_ys[135]), .rectangle2_width(rectangle2_widths[135]), .rectangle2_height(rectangle2_heights[135]), .rectangle2_weight(rectangle2_weights[135]), .rectangle3_x(rectangle3_xs[135]), .rectangle3_y(rectangle3_ys[135]), .rectangle3_width(rectangle3_widths[135]), .rectangle3_height(rectangle3_heights[135]), .rectangle3_weight(rectangle3_weights[135]), .feature_threshold(feature_thresholds[135]), .feature_above(feature_aboves[135]), .feature_below(feature_belows[135]), .scan_win_std_dev(scan_win_std_dev[135]), .feature_accum(feature_accums[135]));
  accum_calculator ac136(.scan_win(scan_win136), .rectangle1_x(rectangle1_xs[136]), .rectangle1_y(rectangle1_ys[136]), .rectangle1_width(rectangle1_widths[136]), .rectangle1_height(rectangle1_heights[136]), .rectangle1_weight(rectangle1_weights[136]), .rectangle2_x(rectangle2_xs[136]), .rectangle2_y(rectangle2_ys[136]), .rectangle2_width(rectangle2_widths[136]), .rectangle2_height(rectangle2_heights[136]), .rectangle2_weight(rectangle2_weights[136]), .rectangle3_x(rectangle3_xs[136]), .rectangle3_y(rectangle3_ys[136]), .rectangle3_width(rectangle3_widths[136]), .rectangle3_height(rectangle3_heights[136]), .rectangle3_weight(rectangle3_weights[136]), .feature_threshold(feature_thresholds[136]), .feature_above(feature_aboves[136]), .feature_below(feature_belows[136]), .scan_win_std_dev(scan_win_std_dev[136]), .feature_accum(feature_accums[136]));
  accum_calculator ac137(.scan_win(scan_win137), .rectangle1_x(rectangle1_xs[137]), .rectangle1_y(rectangle1_ys[137]), .rectangle1_width(rectangle1_widths[137]), .rectangle1_height(rectangle1_heights[137]), .rectangle1_weight(rectangle1_weights[137]), .rectangle2_x(rectangle2_xs[137]), .rectangle2_y(rectangle2_ys[137]), .rectangle2_width(rectangle2_widths[137]), .rectangle2_height(rectangle2_heights[137]), .rectangle2_weight(rectangle2_weights[137]), .rectangle3_x(rectangle3_xs[137]), .rectangle3_y(rectangle3_ys[137]), .rectangle3_width(rectangle3_widths[137]), .rectangle3_height(rectangle3_heights[137]), .rectangle3_weight(rectangle3_weights[137]), .feature_threshold(feature_thresholds[137]), .feature_above(feature_aboves[137]), .feature_below(feature_belows[137]), .scan_win_std_dev(scan_win_std_dev[137]), .feature_accum(feature_accums[137]));
  accum_calculator ac138(.scan_win(scan_win138), .rectangle1_x(rectangle1_xs[138]), .rectangle1_y(rectangle1_ys[138]), .rectangle1_width(rectangle1_widths[138]), .rectangle1_height(rectangle1_heights[138]), .rectangle1_weight(rectangle1_weights[138]), .rectangle2_x(rectangle2_xs[138]), .rectangle2_y(rectangle2_ys[138]), .rectangle2_width(rectangle2_widths[138]), .rectangle2_height(rectangle2_heights[138]), .rectangle2_weight(rectangle2_weights[138]), .rectangle3_x(rectangle3_xs[138]), .rectangle3_y(rectangle3_ys[138]), .rectangle3_width(rectangle3_widths[138]), .rectangle3_height(rectangle3_heights[138]), .rectangle3_weight(rectangle3_weights[138]), .feature_threshold(feature_thresholds[138]), .feature_above(feature_aboves[138]), .feature_below(feature_belows[138]), .scan_win_std_dev(scan_win_std_dev[138]), .feature_accum(feature_accums[138]));
  accum_calculator ac139(.scan_win(scan_win139), .rectangle1_x(rectangle1_xs[139]), .rectangle1_y(rectangle1_ys[139]), .rectangle1_width(rectangle1_widths[139]), .rectangle1_height(rectangle1_heights[139]), .rectangle1_weight(rectangle1_weights[139]), .rectangle2_x(rectangle2_xs[139]), .rectangle2_y(rectangle2_ys[139]), .rectangle2_width(rectangle2_widths[139]), .rectangle2_height(rectangle2_heights[139]), .rectangle2_weight(rectangle2_weights[139]), .rectangle3_x(rectangle3_xs[139]), .rectangle3_y(rectangle3_ys[139]), .rectangle3_width(rectangle3_widths[139]), .rectangle3_height(rectangle3_heights[139]), .rectangle3_weight(rectangle3_weights[139]), .feature_threshold(feature_thresholds[139]), .feature_above(feature_aboves[139]), .feature_below(feature_belows[139]), .scan_win_std_dev(scan_win_std_dev[139]), .feature_accum(feature_accums[139]));
  accum_calculator ac140(.scan_win(scan_win140), .rectangle1_x(rectangle1_xs[140]), .rectangle1_y(rectangle1_ys[140]), .rectangle1_width(rectangle1_widths[140]), .rectangle1_height(rectangle1_heights[140]), .rectangle1_weight(rectangle1_weights[140]), .rectangle2_x(rectangle2_xs[140]), .rectangle2_y(rectangle2_ys[140]), .rectangle2_width(rectangle2_widths[140]), .rectangle2_height(rectangle2_heights[140]), .rectangle2_weight(rectangle2_weights[140]), .rectangle3_x(rectangle3_xs[140]), .rectangle3_y(rectangle3_ys[140]), .rectangle3_width(rectangle3_widths[140]), .rectangle3_height(rectangle3_heights[140]), .rectangle3_weight(rectangle3_weights[140]), .feature_threshold(feature_thresholds[140]), .feature_above(feature_aboves[140]), .feature_below(feature_belows[140]), .scan_win_std_dev(scan_win_std_dev[140]), .feature_accum(feature_accums[140]));
  accum_calculator ac141(.scan_win(scan_win141), .rectangle1_x(rectangle1_xs[141]), .rectangle1_y(rectangle1_ys[141]), .rectangle1_width(rectangle1_widths[141]), .rectangle1_height(rectangle1_heights[141]), .rectangle1_weight(rectangle1_weights[141]), .rectangle2_x(rectangle2_xs[141]), .rectangle2_y(rectangle2_ys[141]), .rectangle2_width(rectangle2_widths[141]), .rectangle2_height(rectangle2_heights[141]), .rectangle2_weight(rectangle2_weights[141]), .rectangle3_x(rectangle3_xs[141]), .rectangle3_y(rectangle3_ys[141]), .rectangle3_width(rectangle3_widths[141]), .rectangle3_height(rectangle3_heights[141]), .rectangle3_weight(rectangle3_weights[141]), .feature_threshold(feature_thresholds[141]), .feature_above(feature_aboves[141]), .feature_below(feature_belows[141]), .scan_win_std_dev(scan_win_std_dev[141]), .feature_accum(feature_accums[141]));
  accum_calculator ac142(.scan_win(scan_win142), .rectangle1_x(rectangle1_xs[142]), .rectangle1_y(rectangle1_ys[142]), .rectangle1_width(rectangle1_widths[142]), .rectangle1_height(rectangle1_heights[142]), .rectangle1_weight(rectangle1_weights[142]), .rectangle2_x(rectangle2_xs[142]), .rectangle2_y(rectangle2_ys[142]), .rectangle2_width(rectangle2_widths[142]), .rectangle2_height(rectangle2_heights[142]), .rectangle2_weight(rectangle2_weights[142]), .rectangle3_x(rectangle3_xs[142]), .rectangle3_y(rectangle3_ys[142]), .rectangle3_width(rectangle3_widths[142]), .rectangle3_height(rectangle3_heights[142]), .rectangle3_weight(rectangle3_weights[142]), .feature_threshold(feature_thresholds[142]), .feature_above(feature_aboves[142]), .feature_below(feature_belows[142]), .scan_win_std_dev(scan_win_std_dev[142]), .feature_accum(feature_accums[142]));
  accum_calculator ac143(.scan_win(scan_win143), .rectangle1_x(rectangle1_xs[143]), .rectangle1_y(rectangle1_ys[143]), .rectangle1_width(rectangle1_widths[143]), .rectangle1_height(rectangle1_heights[143]), .rectangle1_weight(rectangle1_weights[143]), .rectangle2_x(rectangle2_xs[143]), .rectangle2_y(rectangle2_ys[143]), .rectangle2_width(rectangle2_widths[143]), .rectangle2_height(rectangle2_heights[143]), .rectangle2_weight(rectangle2_weights[143]), .rectangle3_x(rectangle3_xs[143]), .rectangle3_y(rectangle3_ys[143]), .rectangle3_width(rectangle3_widths[143]), .rectangle3_height(rectangle3_heights[143]), .rectangle3_weight(rectangle3_weights[143]), .feature_threshold(feature_thresholds[143]), .feature_above(feature_aboves[143]), .feature_below(feature_belows[143]), .scan_win_std_dev(scan_win_std_dev[143]), .feature_accum(feature_accums[143]));
  accum_calculator ac144(.scan_win(scan_win144), .rectangle1_x(rectangle1_xs[144]), .rectangle1_y(rectangle1_ys[144]), .rectangle1_width(rectangle1_widths[144]), .rectangle1_height(rectangle1_heights[144]), .rectangle1_weight(rectangle1_weights[144]), .rectangle2_x(rectangle2_xs[144]), .rectangle2_y(rectangle2_ys[144]), .rectangle2_width(rectangle2_widths[144]), .rectangle2_height(rectangle2_heights[144]), .rectangle2_weight(rectangle2_weights[144]), .rectangle3_x(rectangle3_xs[144]), .rectangle3_y(rectangle3_ys[144]), .rectangle3_width(rectangle3_widths[144]), .rectangle3_height(rectangle3_heights[144]), .rectangle3_weight(rectangle3_weights[144]), .feature_threshold(feature_thresholds[144]), .feature_above(feature_aboves[144]), .feature_below(feature_belows[144]), .scan_win_std_dev(scan_win_std_dev[144]), .feature_accum(feature_accums[144]));
  accum_calculator ac145(.scan_win(scan_win145), .rectangle1_x(rectangle1_xs[145]), .rectangle1_y(rectangle1_ys[145]), .rectangle1_width(rectangle1_widths[145]), .rectangle1_height(rectangle1_heights[145]), .rectangle1_weight(rectangle1_weights[145]), .rectangle2_x(rectangle2_xs[145]), .rectangle2_y(rectangle2_ys[145]), .rectangle2_width(rectangle2_widths[145]), .rectangle2_height(rectangle2_heights[145]), .rectangle2_weight(rectangle2_weights[145]), .rectangle3_x(rectangle3_xs[145]), .rectangle3_y(rectangle3_ys[145]), .rectangle3_width(rectangle3_widths[145]), .rectangle3_height(rectangle3_heights[145]), .rectangle3_weight(rectangle3_weights[145]), .feature_threshold(feature_thresholds[145]), .feature_above(feature_aboves[145]), .feature_below(feature_belows[145]), .scan_win_std_dev(scan_win_std_dev[145]), .feature_accum(feature_accums[145]));
  accum_calculator ac146(.scan_win(scan_win146), .rectangle1_x(rectangle1_xs[146]), .rectangle1_y(rectangle1_ys[146]), .rectangle1_width(rectangle1_widths[146]), .rectangle1_height(rectangle1_heights[146]), .rectangle1_weight(rectangle1_weights[146]), .rectangle2_x(rectangle2_xs[146]), .rectangle2_y(rectangle2_ys[146]), .rectangle2_width(rectangle2_widths[146]), .rectangle2_height(rectangle2_heights[146]), .rectangle2_weight(rectangle2_weights[146]), .rectangle3_x(rectangle3_xs[146]), .rectangle3_y(rectangle3_ys[146]), .rectangle3_width(rectangle3_widths[146]), .rectangle3_height(rectangle3_heights[146]), .rectangle3_weight(rectangle3_weights[146]), .feature_threshold(feature_thresholds[146]), .feature_above(feature_aboves[146]), .feature_below(feature_belows[146]), .scan_win_std_dev(scan_win_std_dev[146]), .feature_accum(feature_accums[146]));
  accum_calculator ac147(.scan_win(scan_win147), .rectangle1_x(rectangle1_xs[147]), .rectangle1_y(rectangle1_ys[147]), .rectangle1_width(rectangle1_widths[147]), .rectangle1_height(rectangle1_heights[147]), .rectangle1_weight(rectangle1_weights[147]), .rectangle2_x(rectangle2_xs[147]), .rectangle2_y(rectangle2_ys[147]), .rectangle2_width(rectangle2_widths[147]), .rectangle2_height(rectangle2_heights[147]), .rectangle2_weight(rectangle2_weights[147]), .rectangle3_x(rectangle3_xs[147]), .rectangle3_y(rectangle3_ys[147]), .rectangle3_width(rectangle3_widths[147]), .rectangle3_height(rectangle3_heights[147]), .rectangle3_weight(rectangle3_weights[147]), .feature_threshold(feature_thresholds[147]), .feature_above(feature_aboves[147]), .feature_below(feature_belows[147]), .scan_win_std_dev(scan_win_std_dev[147]), .feature_accum(feature_accums[147]));
  accum_calculator ac148(.scan_win(scan_win148), .rectangle1_x(rectangle1_xs[148]), .rectangle1_y(rectangle1_ys[148]), .rectangle1_width(rectangle1_widths[148]), .rectangle1_height(rectangle1_heights[148]), .rectangle1_weight(rectangle1_weights[148]), .rectangle2_x(rectangle2_xs[148]), .rectangle2_y(rectangle2_ys[148]), .rectangle2_width(rectangle2_widths[148]), .rectangle2_height(rectangle2_heights[148]), .rectangle2_weight(rectangle2_weights[148]), .rectangle3_x(rectangle3_xs[148]), .rectangle3_y(rectangle3_ys[148]), .rectangle3_width(rectangle3_widths[148]), .rectangle3_height(rectangle3_heights[148]), .rectangle3_weight(rectangle3_weights[148]), .feature_threshold(feature_thresholds[148]), .feature_above(feature_aboves[148]), .feature_below(feature_belows[148]), .scan_win_std_dev(scan_win_std_dev[148]), .feature_accum(feature_accums[148]));
  accum_calculator ac149(.scan_win(scan_win149), .rectangle1_x(rectangle1_xs[149]), .rectangle1_y(rectangle1_ys[149]), .rectangle1_width(rectangle1_widths[149]), .rectangle1_height(rectangle1_heights[149]), .rectangle1_weight(rectangle1_weights[149]), .rectangle2_x(rectangle2_xs[149]), .rectangle2_y(rectangle2_ys[149]), .rectangle2_width(rectangle2_widths[149]), .rectangle2_height(rectangle2_heights[149]), .rectangle2_weight(rectangle2_weights[149]), .rectangle3_x(rectangle3_xs[149]), .rectangle3_y(rectangle3_ys[149]), .rectangle3_width(rectangle3_widths[149]), .rectangle3_height(rectangle3_heights[149]), .rectangle3_weight(rectangle3_weights[149]), .feature_threshold(feature_thresholds[149]), .feature_above(feature_aboves[149]), .feature_below(feature_belows[149]), .scan_win_std_dev(scan_win_std_dev[149]), .feature_accum(feature_accums[149]));
  accum_calculator ac150(.scan_win(scan_win150), .rectangle1_x(rectangle1_xs[150]), .rectangle1_y(rectangle1_ys[150]), .rectangle1_width(rectangle1_widths[150]), .rectangle1_height(rectangle1_heights[150]), .rectangle1_weight(rectangle1_weights[150]), .rectangle2_x(rectangle2_xs[150]), .rectangle2_y(rectangle2_ys[150]), .rectangle2_width(rectangle2_widths[150]), .rectangle2_height(rectangle2_heights[150]), .rectangle2_weight(rectangle2_weights[150]), .rectangle3_x(rectangle3_xs[150]), .rectangle3_y(rectangle3_ys[150]), .rectangle3_width(rectangle3_widths[150]), .rectangle3_height(rectangle3_heights[150]), .rectangle3_weight(rectangle3_weights[150]), .feature_threshold(feature_thresholds[150]), .feature_above(feature_aboves[150]), .feature_below(feature_belows[150]), .scan_win_std_dev(scan_win_std_dev[150]), .feature_accum(feature_accums[150]));
  accum_calculator ac151(.scan_win(scan_win151), .rectangle1_x(rectangle1_xs[151]), .rectangle1_y(rectangle1_ys[151]), .rectangle1_width(rectangle1_widths[151]), .rectangle1_height(rectangle1_heights[151]), .rectangle1_weight(rectangle1_weights[151]), .rectangle2_x(rectangle2_xs[151]), .rectangle2_y(rectangle2_ys[151]), .rectangle2_width(rectangle2_widths[151]), .rectangle2_height(rectangle2_heights[151]), .rectangle2_weight(rectangle2_weights[151]), .rectangle3_x(rectangle3_xs[151]), .rectangle3_y(rectangle3_ys[151]), .rectangle3_width(rectangle3_widths[151]), .rectangle3_height(rectangle3_heights[151]), .rectangle3_weight(rectangle3_weights[151]), .feature_threshold(feature_thresholds[151]), .feature_above(feature_aboves[151]), .feature_below(feature_belows[151]), .scan_win_std_dev(scan_win_std_dev[151]), .feature_accum(feature_accums[151]));
  accum_calculator ac152(.scan_win(scan_win152), .rectangle1_x(rectangle1_xs[152]), .rectangle1_y(rectangle1_ys[152]), .rectangle1_width(rectangle1_widths[152]), .rectangle1_height(rectangle1_heights[152]), .rectangle1_weight(rectangle1_weights[152]), .rectangle2_x(rectangle2_xs[152]), .rectangle2_y(rectangle2_ys[152]), .rectangle2_width(rectangle2_widths[152]), .rectangle2_height(rectangle2_heights[152]), .rectangle2_weight(rectangle2_weights[152]), .rectangle3_x(rectangle3_xs[152]), .rectangle3_y(rectangle3_ys[152]), .rectangle3_width(rectangle3_widths[152]), .rectangle3_height(rectangle3_heights[152]), .rectangle3_weight(rectangle3_weights[152]), .feature_threshold(feature_thresholds[152]), .feature_above(feature_aboves[152]), .feature_below(feature_belows[152]), .scan_win_std_dev(scan_win_std_dev[152]), .feature_accum(feature_accums[152]));
  accum_calculator ac153(.scan_win(scan_win153), .rectangle1_x(rectangle1_xs[153]), .rectangle1_y(rectangle1_ys[153]), .rectangle1_width(rectangle1_widths[153]), .rectangle1_height(rectangle1_heights[153]), .rectangle1_weight(rectangle1_weights[153]), .rectangle2_x(rectangle2_xs[153]), .rectangle2_y(rectangle2_ys[153]), .rectangle2_width(rectangle2_widths[153]), .rectangle2_height(rectangle2_heights[153]), .rectangle2_weight(rectangle2_weights[153]), .rectangle3_x(rectangle3_xs[153]), .rectangle3_y(rectangle3_ys[153]), .rectangle3_width(rectangle3_widths[153]), .rectangle3_height(rectangle3_heights[153]), .rectangle3_weight(rectangle3_weights[153]), .feature_threshold(feature_thresholds[153]), .feature_above(feature_aboves[153]), .feature_below(feature_belows[153]), .scan_win_std_dev(scan_win_std_dev[153]), .feature_accum(feature_accums[153]));
  accum_calculator ac154(.scan_win(scan_win154), .rectangle1_x(rectangle1_xs[154]), .rectangle1_y(rectangle1_ys[154]), .rectangle1_width(rectangle1_widths[154]), .rectangle1_height(rectangle1_heights[154]), .rectangle1_weight(rectangle1_weights[154]), .rectangle2_x(rectangle2_xs[154]), .rectangle2_y(rectangle2_ys[154]), .rectangle2_width(rectangle2_widths[154]), .rectangle2_height(rectangle2_heights[154]), .rectangle2_weight(rectangle2_weights[154]), .rectangle3_x(rectangle3_xs[154]), .rectangle3_y(rectangle3_ys[154]), .rectangle3_width(rectangle3_widths[154]), .rectangle3_height(rectangle3_heights[154]), .rectangle3_weight(rectangle3_weights[154]), .feature_threshold(feature_thresholds[154]), .feature_above(feature_aboves[154]), .feature_below(feature_belows[154]), .scan_win_std_dev(scan_win_std_dev[154]), .feature_accum(feature_accums[154]));
  accum_calculator ac155(.scan_win(scan_win155), .rectangle1_x(rectangle1_xs[155]), .rectangle1_y(rectangle1_ys[155]), .rectangle1_width(rectangle1_widths[155]), .rectangle1_height(rectangle1_heights[155]), .rectangle1_weight(rectangle1_weights[155]), .rectangle2_x(rectangle2_xs[155]), .rectangle2_y(rectangle2_ys[155]), .rectangle2_width(rectangle2_widths[155]), .rectangle2_height(rectangle2_heights[155]), .rectangle2_weight(rectangle2_weights[155]), .rectangle3_x(rectangle3_xs[155]), .rectangle3_y(rectangle3_ys[155]), .rectangle3_width(rectangle3_widths[155]), .rectangle3_height(rectangle3_heights[155]), .rectangle3_weight(rectangle3_weights[155]), .feature_threshold(feature_thresholds[155]), .feature_above(feature_aboves[155]), .feature_below(feature_belows[155]), .scan_win_std_dev(scan_win_std_dev[155]), .feature_accum(feature_accums[155]));
  accum_calculator ac156(.scan_win(scan_win156), .rectangle1_x(rectangle1_xs[156]), .rectangle1_y(rectangle1_ys[156]), .rectangle1_width(rectangle1_widths[156]), .rectangle1_height(rectangle1_heights[156]), .rectangle1_weight(rectangle1_weights[156]), .rectangle2_x(rectangle2_xs[156]), .rectangle2_y(rectangle2_ys[156]), .rectangle2_width(rectangle2_widths[156]), .rectangle2_height(rectangle2_heights[156]), .rectangle2_weight(rectangle2_weights[156]), .rectangle3_x(rectangle3_xs[156]), .rectangle3_y(rectangle3_ys[156]), .rectangle3_width(rectangle3_widths[156]), .rectangle3_height(rectangle3_heights[156]), .rectangle3_weight(rectangle3_weights[156]), .feature_threshold(feature_thresholds[156]), .feature_above(feature_aboves[156]), .feature_below(feature_belows[156]), .scan_win_std_dev(scan_win_std_dev[156]), .feature_accum(feature_accums[156]));
  accum_calculator ac157(.scan_win(scan_win157), .rectangle1_x(rectangle1_xs[157]), .rectangle1_y(rectangle1_ys[157]), .rectangle1_width(rectangle1_widths[157]), .rectangle1_height(rectangle1_heights[157]), .rectangle1_weight(rectangle1_weights[157]), .rectangle2_x(rectangle2_xs[157]), .rectangle2_y(rectangle2_ys[157]), .rectangle2_width(rectangle2_widths[157]), .rectangle2_height(rectangle2_heights[157]), .rectangle2_weight(rectangle2_weights[157]), .rectangle3_x(rectangle3_xs[157]), .rectangle3_y(rectangle3_ys[157]), .rectangle3_width(rectangle3_widths[157]), .rectangle3_height(rectangle3_heights[157]), .rectangle3_weight(rectangle3_weights[157]), .feature_threshold(feature_thresholds[157]), .feature_above(feature_aboves[157]), .feature_below(feature_belows[157]), .scan_win_std_dev(scan_win_std_dev[157]), .feature_accum(feature_accums[157]));
  accum_calculator ac158(.scan_win(scan_win158), .rectangle1_x(rectangle1_xs[158]), .rectangle1_y(rectangle1_ys[158]), .rectangle1_width(rectangle1_widths[158]), .rectangle1_height(rectangle1_heights[158]), .rectangle1_weight(rectangle1_weights[158]), .rectangle2_x(rectangle2_xs[158]), .rectangle2_y(rectangle2_ys[158]), .rectangle2_width(rectangle2_widths[158]), .rectangle2_height(rectangle2_heights[158]), .rectangle2_weight(rectangle2_weights[158]), .rectangle3_x(rectangle3_xs[158]), .rectangle3_y(rectangle3_ys[158]), .rectangle3_width(rectangle3_widths[158]), .rectangle3_height(rectangle3_heights[158]), .rectangle3_weight(rectangle3_weights[158]), .feature_threshold(feature_thresholds[158]), .feature_above(feature_aboves[158]), .feature_below(feature_belows[158]), .scan_win_std_dev(scan_win_std_dev[158]), .feature_accum(feature_accums[158]));
  accum_calculator ac159(.scan_win(scan_win159), .rectangle1_x(rectangle1_xs[159]), .rectangle1_y(rectangle1_ys[159]), .rectangle1_width(rectangle1_widths[159]), .rectangle1_height(rectangle1_heights[159]), .rectangle1_weight(rectangle1_weights[159]), .rectangle2_x(rectangle2_xs[159]), .rectangle2_y(rectangle2_ys[159]), .rectangle2_width(rectangle2_widths[159]), .rectangle2_height(rectangle2_heights[159]), .rectangle2_weight(rectangle2_weights[159]), .rectangle3_x(rectangle3_xs[159]), .rectangle3_y(rectangle3_ys[159]), .rectangle3_width(rectangle3_widths[159]), .rectangle3_height(rectangle3_heights[159]), .rectangle3_weight(rectangle3_weights[159]), .feature_threshold(feature_thresholds[159]), .feature_above(feature_aboves[159]), .feature_below(feature_belows[159]), .scan_win_std_dev(scan_win_std_dev[159]), .feature_accum(feature_accums[159]));
  accum_calculator ac160(.scan_win(scan_win160), .rectangle1_x(rectangle1_xs[160]), .rectangle1_y(rectangle1_ys[160]), .rectangle1_width(rectangle1_widths[160]), .rectangle1_height(rectangle1_heights[160]), .rectangle1_weight(rectangle1_weights[160]), .rectangle2_x(rectangle2_xs[160]), .rectangle2_y(rectangle2_ys[160]), .rectangle2_width(rectangle2_widths[160]), .rectangle2_height(rectangle2_heights[160]), .rectangle2_weight(rectangle2_weights[160]), .rectangle3_x(rectangle3_xs[160]), .rectangle3_y(rectangle3_ys[160]), .rectangle3_width(rectangle3_widths[160]), .rectangle3_height(rectangle3_heights[160]), .rectangle3_weight(rectangle3_weights[160]), .feature_threshold(feature_thresholds[160]), .feature_above(feature_aboves[160]), .feature_below(feature_belows[160]), .scan_win_std_dev(scan_win_std_dev[160]), .feature_accum(feature_accums[160]));
  accum_calculator ac161(.scan_win(scan_win161), .rectangle1_x(rectangle1_xs[161]), .rectangle1_y(rectangle1_ys[161]), .rectangle1_width(rectangle1_widths[161]), .rectangle1_height(rectangle1_heights[161]), .rectangle1_weight(rectangle1_weights[161]), .rectangle2_x(rectangle2_xs[161]), .rectangle2_y(rectangle2_ys[161]), .rectangle2_width(rectangle2_widths[161]), .rectangle2_height(rectangle2_heights[161]), .rectangle2_weight(rectangle2_weights[161]), .rectangle3_x(rectangle3_xs[161]), .rectangle3_y(rectangle3_ys[161]), .rectangle3_width(rectangle3_widths[161]), .rectangle3_height(rectangle3_heights[161]), .rectangle3_weight(rectangle3_weights[161]), .feature_threshold(feature_thresholds[161]), .feature_above(feature_aboves[161]), .feature_below(feature_belows[161]), .scan_win_std_dev(scan_win_std_dev[161]), .feature_accum(feature_accums[161]));
  accum_calculator ac162(.scan_win(scan_win162), .rectangle1_x(rectangle1_xs[162]), .rectangle1_y(rectangle1_ys[162]), .rectangle1_width(rectangle1_widths[162]), .rectangle1_height(rectangle1_heights[162]), .rectangle1_weight(rectangle1_weights[162]), .rectangle2_x(rectangle2_xs[162]), .rectangle2_y(rectangle2_ys[162]), .rectangle2_width(rectangle2_widths[162]), .rectangle2_height(rectangle2_heights[162]), .rectangle2_weight(rectangle2_weights[162]), .rectangle3_x(rectangle3_xs[162]), .rectangle3_y(rectangle3_ys[162]), .rectangle3_width(rectangle3_widths[162]), .rectangle3_height(rectangle3_heights[162]), .rectangle3_weight(rectangle3_weights[162]), .feature_threshold(feature_thresholds[162]), .feature_above(feature_aboves[162]), .feature_below(feature_belows[162]), .scan_win_std_dev(scan_win_std_dev[162]), .feature_accum(feature_accums[162]));
  accum_calculator ac163(.scan_win(scan_win163), .rectangle1_x(rectangle1_xs[163]), .rectangle1_y(rectangle1_ys[163]), .rectangle1_width(rectangle1_widths[163]), .rectangle1_height(rectangle1_heights[163]), .rectangle1_weight(rectangle1_weights[163]), .rectangle2_x(rectangle2_xs[163]), .rectangle2_y(rectangle2_ys[163]), .rectangle2_width(rectangle2_widths[163]), .rectangle2_height(rectangle2_heights[163]), .rectangle2_weight(rectangle2_weights[163]), .rectangle3_x(rectangle3_xs[163]), .rectangle3_y(rectangle3_ys[163]), .rectangle3_width(rectangle3_widths[163]), .rectangle3_height(rectangle3_heights[163]), .rectangle3_weight(rectangle3_weights[163]), .feature_threshold(feature_thresholds[163]), .feature_above(feature_aboves[163]), .feature_below(feature_belows[163]), .scan_win_std_dev(scan_win_std_dev[163]), .feature_accum(feature_accums[163]));
  accum_calculator ac164(.scan_win(scan_win164), .rectangle1_x(rectangle1_xs[164]), .rectangle1_y(rectangle1_ys[164]), .rectangle1_width(rectangle1_widths[164]), .rectangle1_height(rectangle1_heights[164]), .rectangle1_weight(rectangle1_weights[164]), .rectangle2_x(rectangle2_xs[164]), .rectangle2_y(rectangle2_ys[164]), .rectangle2_width(rectangle2_widths[164]), .rectangle2_height(rectangle2_heights[164]), .rectangle2_weight(rectangle2_weights[164]), .rectangle3_x(rectangle3_xs[164]), .rectangle3_y(rectangle3_ys[164]), .rectangle3_width(rectangle3_widths[164]), .rectangle3_height(rectangle3_heights[164]), .rectangle3_weight(rectangle3_weights[164]), .feature_threshold(feature_thresholds[164]), .feature_above(feature_aboves[164]), .feature_below(feature_belows[164]), .scan_win_std_dev(scan_win_std_dev[164]), .feature_accum(feature_accums[164]));
  accum_calculator ac165(.scan_win(scan_win165), .rectangle1_x(rectangle1_xs[165]), .rectangle1_y(rectangle1_ys[165]), .rectangle1_width(rectangle1_widths[165]), .rectangle1_height(rectangle1_heights[165]), .rectangle1_weight(rectangle1_weights[165]), .rectangle2_x(rectangle2_xs[165]), .rectangle2_y(rectangle2_ys[165]), .rectangle2_width(rectangle2_widths[165]), .rectangle2_height(rectangle2_heights[165]), .rectangle2_weight(rectangle2_weights[165]), .rectangle3_x(rectangle3_xs[165]), .rectangle3_y(rectangle3_ys[165]), .rectangle3_width(rectangle3_widths[165]), .rectangle3_height(rectangle3_heights[165]), .rectangle3_weight(rectangle3_weights[165]), .feature_threshold(feature_thresholds[165]), .feature_above(feature_aboves[165]), .feature_below(feature_belows[165]), .scan_win_std_dev(scan_win_std_dev[165]), .feature_accum(feature_accums[165]));
  accum_calculator ac166(.scan_win(scan_win166), .rectangle1_x(rectangle1_xs[166]), .rectangle1_y(rectangle1_ys[166]), .rectangle1_width(rectangle1_widths[166]), .rectangle1_height(rectangle1_heights[166]), .rectangle1_weight(rectangle1_weights[166]), .rectangle2_x(rectangle2_xs[166]), .rectangle2_y(rectangle2_ys[166]), .rectangle2_width(rectangle2_widths[166]), .rectangle2_height(rectangle2_heights[166]), .rectangle2_weight(rectangle2_weights[166]), .rectangle3_x(rectangle3_xs[166]), .rectangle3_y(rectangle3_ys[166]), .rectangle3_width(rectangle3_widths[166]), .rectangle3_height(rectangle3_heights[166]), .rectangle3_weight(rectangle3_weights[166]), .feature_threshold(feature_thresholds[166]), .feature_above(feature_aboves[166]), .feature_below(feature_belows[166]), .scan_win_std_dev(scan_win_std_dev[166]), .feature_accum(feature_accums[166]));
  accum_calculator ac167(.scan_win(scan_win167), .rectangle1_x(rectangle1_xs[167]), .rectangle1_y(rectangle1_ys[167]), .rectangle1_width(rectangle1_widths[167]), .rectangle1_height(rectangle1_heights[167]), .rectangle1_weight(rectangle1_weights[167]), .rectangle2_x(rectangle2_xs[167]), .rectangle2_y(rectangle2_ys[167]), .rectangle2_width(rectangle2_widths[167]), .rectangle2_height(rectangle2_heights[167]), .rectangle2_weight(rectangle2_weights[167]), .rectangle3_x(rectangle3_xs[167]), .rectangle3_y(rectangle3_ys[167]), .rectangle3_width(rectangle3_widths[167]), .rectangle3_height(rectangle3_heights[167]), .rectangle3_weight(rectangle3_weights[167]), .feature_threshold(feature_thresholds[167]), .feature_above(feature_aboves[167]), .feature_below(feature_belows[167]), .scan_win_std_dev(scan_win_std_dev[167]), .feature_accum(feature_accums[167]));
  accum_calculator ac168(.scan_win(scan_win168), .rectangle1_x(rectangle1_xs[168]), .rectangle1_y(rectangle1_ys[168]), .rectangle1_width(rectangle1_widths[168]), .rectangle1_height(rectangle1_heights[168]), .rectangle1_weight(rectangle1_weights[168]), .rectangle2_x(rectangle2_xs[168]), .rectangle2_y(rectangle2_ys[168]), .rectangle2_width(rectangle2_widths[168]), .rectangle2_height(rectangle2_heights[168]), .rectangle2_weight(rectangle2_weights[168]), .rectangle3_x(rectangle3_xs[168]), .rectangle3_y(rectangle3_ys[168]), .rectangle3_width(rectangle3_widths[168]), .rectangle3_height(rectangle3_heights[168]), .rectangle3_weight(rectangle3_weights[168]), .feature_threshold(feature_thresholds[168]), .feature_above(feature_aboves[168]), .feature_below(feature_belows[168]), .scan_win_std_dev(scan_win_std_dev[168]), .feature_accum(feature_accums[168]));
  accum_calculator ac169(.scan_win(scan_win169), .rectangle1_x(rectangle1_xs[169]), .rectangle1_y(rectangle1_ys[169]), .rectangle1_width(rectangle1_widths[169]), .rectangle1_height(rectangle1_heights[169]), .rectangle1_weight(rectangle1_weights[169]), .rectangle2_x(rectangle2_xs[169]), .rectangle2_y(rectangle2_ys[169]), .rectangle2_width(rectangle2_widths[169]), .rectangle2_height(rectangle2_heights[169]), .rectangle2_weight(rectangle2_weights[169]), .rectangle3_x(rectangle3_xs[169]), .rectangle3_y(rectangle3_ys[169]), .rectangle3_width(rectangle3_widths[169]), .rectangle3_height(rectangle3_heights[169]), .rectangle3_weight(rectangle3_weights[169]), .feature_threshold(feature_thresholds[169]), .feature_above(feature_aboves[169]), .feature_below(feature_belows[169]), .scan_win_std_dev(scan_win_std_dev[169]), .feature_accum(feature_accums[169]));
  accum_calculator ac170(.scan_win(scan_win170), .rectangle1_x(rectangle1_xs[170]), .rectangle1_y(rectangle1_ys[170]), .rectangle1_width(rectangle1_widths[170]), .rectangle1_height(rectangle1_heights[170]), .rectangle1_weight(rectangle1_weights[170]), .rectangle2_x(rectangle2_xs[170]), .rectangle2_y(rectangle2_ys[170]), .rectangle2_width(rectangle2_widths[170]), .rectangle2_height(rectangle2_heights[170]), .rectangle2_weight(rectangle2_weights[170]), .rectangle3_x(rectangle3_xs[170]), .rectangle3_y(rectangle3_ys[170]), .rectangle3_width(rectangle3_widths[170]), .rectangle3_height(rectangle3_heights[170]), .rectangle3_weight(rectangle3_weights[170]), .feature_threshold(feature_thresholds[170]), .feature_above(feature_aboves[170]), .feature_below(feature_belows[170]), .scan_win_std_dev(scan_win_std_dev[170]), .feature_accum(feature_accums[170]));
  accum_calculator ac171(.scan_win(scan_win171), .rectangle1_x(rectangle1_xs[171]), .rectangle1_y(rectangle1_ys[171]), .rectangle1_width(rectangle1_widths[171]), .rectangle1_height(rectangle1_heights[171]), .rectangle1_weight(rectangle1_weights[171]), .rectangle2_x(rectangle2_xs[171]), .rectangle2_y(rectangle2_ys[171]), .rectangle2_width(rectangle2_widths[171]), .rectangle2_height(rectangle2_heights[171]), .rectangle2_weight(rectangle2_weights[171]), .rectangle3_x(rectangle3_xs[171]), .rectangle3_y(rectangle3_ys[171]), .rectangle3_width(rectangle3_widths[171]), .rectangle3_height(rectangle3_heights[171]), .rectangle3_weight(rectangle3_weights[171]), .feature_threshold(feature_thresholds[171]), .feature_above(feature_aboves[171]), .feature_below(feature_belows[171]), .scan_win_std_dev(scan_win_std_dev[171]), .feature_accum(feature_accums[171]));
  accum_calculator ac172(.scan_win(scan_win172), .rectangle1_x(rectangle1_xs[172]), .rectangle1_y(rectangle1_ys[172]), .rectangle1_width(rectangle1_widths[172]), .rectangle1_height(rectangle1_heights[172]), .rectangle1_weight(rectangle1_weights[172]), .rectangle2_x(rectangle2_xs[172]), .rectangle2_y(rectangle2_ys[172]), .rectangle2_width(rectangle2_widths[172]), .rectangle2_height(rectangle2_heights[172]), .rectangle2_weight(rectangle2_weights[172]), .rectangle3_x(rectangle3_xs[172]), .rectangle3_y(rectangle3_ys[172]), .rectangle3_width(rectangle3_widths[172]), .rectangle3_height(rectangle3_heights[172]), .rectangle3_weight(rectangle3_weights[172]), .feature_threshold(feature_thresholds[172]), .feature_above(feature_aboves[172]), .feature_below(feature_belows[172]), .scan_win_std_dev(scan_win_std_dev[172]), .feature_accum(feature_accums[172]));
  accum_calculator ac173(.scan_win(scan_win173), .rectangle1_x(rectangle1_xs[173]), .rectangle1_y(rectangle1_ys[173]), .rectangle1_width(rectangle1_widths[173]), .rectangle1_height(rectangle1_heights[173]), .rectangle1_weight(rectangle1_weights[173]), .rectangle2_x(rectangle2_xs[173]), .rectangle2_y(rectangle2_ys[173]), .rectangle2_width(rectangle2_widths[173]), .rectangle2_height(rectangle2_heights[173]), .rectangle2_weight(rectangle2_weights[173]), .rectangle3_x(rectangle3_xs[173]), .rectangle3_y(rectangle3_ys[173]), .rectangle3_width(rectangle3_widths[173]), .rectangle3_height(rectangle3_heights[173]), .rectangle3_weight(rectangle3_weights[173]), .feature_threshold(feature_thresholds[173]), .feature_above(feature_aboves[173]), .feature_below(feature_belows[173]), .scan_win_std_dev(scan_win_std_dev[173]), .feature_accum(feature_accums[173]));
  accum_calculator ac174(.scan_win(scan_win174), .rectangle1_x(rectangle1_xs[174]), .rectangle1_y(rectangle1_ys[174]), .rectangle1_width(rectangle1_widths[174]), .rectangle1_height(rectangle1_heights[174]), .rectangle1_weight(rectangle1_weights[174]), .rectangle2_x(rectangle2_xs[174]), .rectangle2_y(rectangle2_ys[174]), .rectangle2_width(rectangle2_widths[174]), .rectangle2_height(rectangle2_heights[174]), .rectangle2_weight(rectangle2_weights[174]), .rectangle3_x(rectangle3_xs[174]), .rectangle3_y(rectangle3_ys[174]), .rectangle3_width(rectangle3_widths[174]), .rectangle3_height(rectangle3_heights[174]), .rectangle3_weight(rectangle3_weights[174]), .feature_threshold(feature_thresholds[174]), .feature_above(feature_aboves[174]), .feature_below(feature_belows[174]), .scan_win_std_dev(scan_win_std_dev[174]), .feature_accum(feature_accums[174]));
  accum_calculator ac175(.scan_win(scan_win175), .rectangle1_x(rectangle1_xs[175]), .rectangle1_y(rectangle1_ys[175]), .rectangle1_width(rectangle1_widths[175]), .rectangle1_height(rectangle1_heights[175]), .rectangle1_weight(rectangle1_weights[175]), .rectangle2_x(rectangle2_xs[175]), .rectangle2_y(rectangle2_ys[175]), .rectangle2_width(rectangle2_widths[175]), .rectangle2_height(rectangle2_heights[175]), .rectangle2_weight(rectangle2_weights[175]), .rectangle3_x(rectangle3_xs[175]), .rectangle3_y(rectangle3_ys[175]), .rectangle3_width(rectangle3_widths[175]), .rectangle3_height(rectangle3_heights[175]), .rectangle3_weight(rectangle3_weights[175]), .feature_threshold(feature_thresholds[175]), .feature_above(feature_aboves[175]), .feature_below(feature_belows[175]), .scan_win_std_dev(scan_win_std_dev[175]), .feature_accum(feature_accums[175]));
  accum_calculator ac176(.scan_win(scan_win176), .rectangle1_x(rectangle1_xs[176]), .rectangle1_y(rectangle1_ys[176]), .rectangle1_width(rectangle1_widths[176]), .rectangle1_height(rectangle1_heights[176]), .rectangle1_weight(rectangle1_weights[176]), .rectangle2_x(rectangle2_xs[176]), .rectangle2_y(rectangle2_ys[176]), .rectangle2_width(rectangle2_widths[176]), .rectangle2_height(rectangle2_heights[176]), .rectangle2_weight(rectangle2_weights[176]), .rectangle3_x(rectangle3_xs[176]), .rectangle3_y(rectangle3_ys[176]), .rectangle3_width(rectangle3_widths[176]), .rectangle3_height(rectangle3_heights[176]), .rectangle3_weight(rectangle3_weights[176]), .feature_threshold(feature_thresholds[176]), .feature_above(feature_aboves[176]), .feature_below(feature_belows[176]), .scan_win_std_dev(scan_win_std_dev[176]), .feature_accum(feature_accums[176]));
  accum_calculator ac177(.scan_win(scan_win177), .rectangle1_x(rectangle1_xs[177]), .rectangle1_y(rectangle1_ys[177]), .rectangle1_width(rectangle1_widths[177]), .rectangle1_height(rectangle1_heights[177]), .rectangle1_weight(rectangle1_weights[177]), .rectangle2_x(rectangle2_xs[177]), .rectangle2_y(rectangle2_ys[177]), .rectangle2_width(rectangle2_widths[177]), .rectangle2_height(rectangle2_heights[177]), .rectangle2_weight(rectangle2_weights[177]), .rectangle3_x(rectangle3_xs[177]), .rectangle3_y(rectangle3_ys[177]), .rectangle3_width(rectangle3_widths[177]), .rectangle3_height(rectangle3_heights[177]), .rectangle3_weight(rectangle3_weights[177]), .feature_threshold(feature_thresholds[177]), .feature_above(feature_aboves[177]), .feature_below(feature_belows[177]), .scan_win_std_dev(scan_win_std_dev[177]), .feature_accum(feature_accums[177]));
  accum_calculator ac178(.scan_win(scan_win178), .rectangle1_x(rectangle1_xs[178]), .rectangle1_y(rectangle1_ys[178]), .rectangle1_width(rectangle1_widths[178]), .rectangle1_height(rectangle1_heights[178]), .rectangle1_weight(rectangle1_weights[178]), .rectangle2_x(rectangle2_xs[178]), .rectangle2_y(rectangle2_ys[178]), .rectangle2_width(rectangle2_widths[178]), .rectangle2_height(rectangle2_heights[178]), .rectangle2_weight(rectangle2_weights[178]), .rectangle3_x(rectangle3_xs[178]), .rectangle3_y(rectangle3_ys[178]), .rectangle3_width(rectangle3_widths[178]), .rectangle3_height(rectangle3_heights[178]), .rectangle3_weight(rectangle3_weights[178]), .feature_threshold(feature_thresholds[178]), .feature_above(feature_aboves[178]), .feature_below(feature_belows[178]), .scan_win_std_dev(scan_win_std_dev[178]), .feature_accum(feature_accums[178]));
  accum_calculator ac179(.scan_win(scan_win179), .rectangle1_x(rectangle1_xs[179]), .rectangle1_y(rectangle1_ys[179]), .rectangle1_width(rectangle1_widths[179]), .rectangle1_height(rectangle1_heights[179]), .rectangle1_weight(rectangle1_weights[179]), .rectangle2_x(rectangle2_xs[179]), .rectangle2_y(rectangle2_ys[179]), .rectangle2_width(rectangle2_widths[179]), .rectangle2_height(rectangle2_heights[179]), .rectangle2_weight(rectangle2_weights[179]), .rectangle3_x(rectangle3_xs[179]), .rectangle3_y(rectangle3_ys[179]), .rectangle3_width(rectangle3_widths[179]), .rectangle3_height(rectangle3_heights[179]), .rectangle3_weight(rectangle3_weights[179]), .feature_threshold(feature_thresholds[179]), .feature_above(feature_aboves[179]), .feature_below(feature_belows[179]), .scan_win_std_dev(scan_win_std_dev[179]), .feature_accum(feature_accums[179]));
  accum_calculator ac180(.scan_win(scan_win180), .rectangle1_x(rectangle1_xs[180]), .rectangle1_y(rectangle1_ys[180]), .rectangle1_width(rectangle1_widths[180]), .rectangle1_height(rectangle1_heights[180]), .rectangle1_weight(rectangle1_weights[180]), .rectangle2_x(rectangle2_xs[180]), .rectangle2_y(rectangle2_ys[180]), .rectangle2_width(rectangle2_widths[180]), .rectangle2_height(rectangle2_heights[180]), .rectangle2_weight(rectangle2_weights[180]), .rectangle3_x(rectangle3_xs[180]), .rectangle3_y(rectangle3_ys[180]), .rectangle3_width(rectangle3_widths[180]), .rectangle3_height(rectangle3_heights[180]), .rectangle3_weight(rectangle3_weights[180]), .feature_threshold(feature_thresholds[180]), .feature_above(feature_aboves[180]), .feature_below(feature_belows[180]), .scan_win_std_dev(scan_win_std_dev[180]), .feature_accum(feature_accums[180]));
  accum_calculator ac181(.scan_win(scan_win181), .rectangle1_x(rectangle1_xs[181]), .rectangle1_y(rectangle1_ys[181]), .rectangle1_width(rectangle1_widths[181]), .rectangle1_height(rectangle1_heights[181]), .rectangle1_weight(rectangle1_weights[181]), .rectangle2_x(rectangle2_xs[181]), .rectangle2_y(rectangle2_ys[181]), .rectangle2_width(rectangle2_widths[181]), .rectangle2_height(rectangle2_heights[181]), .rectangle2_weight(rectangle2_weights[181]), .rectangle3_x(rectangle3_xs[181]), .rectangle3_y(rectangle3_ys[181]), .rectangle3_width(rectangle3_widths[181]), .rectangle3_height(rectangle3_heights[181]), .rectangle3_weight(rectangle3_weights[181]), .feature_threshold(feature_thresholds[181]), .feature_above(feature_aboves[181]), .feature_below(feature_belows[181]), .scan_win_std_dev(scan_win_std_dev[181]), .feature_accum(feature_accums[181]));
  accum_calculator ac182(.scan_win(scan_win182), .rectangle1_x(rectangle1_xs[182]), .rectangle1_y(rectangle1_ys[182]), .rectangle1_width(rectangle1_widths[182]), .rectangle1_height(rectangle1_heights[182]), .rectangle1_weight(rectangle1_weights[182]), .rectangle2_x(rectangle2_xs[182]), .rectangle2_y(rectangle2_ys[182]), .rectangle2_width(rectangle2_widths[182]), .rectangle2_height(rectangle2_heights[182]), .rectangle2_weight(rectangle2_weights[182]), .rectangle3_x(rectangle3_xs[182]), .rectangle3_y(rectangle3_ys[182]), .rectangle3_width(rectangle3_widths[182]), .rectangle3_height(rectangle3_heights[182]), .rectangle3_weight(rectangle3_weights[182]), .feature_threshold(feature_thresholds[182]), .feature_above(feature_aboves[182]), .feature_below(feature_belows[182]), .scan_win_std_dev(scan_win_std_dev[182]), .feature_accum(feature_accums[182]));
  accum_calculator ac183(.scan_win(scan_win183), .rectangle1_x(rectangle1_xs[183]), .rectangle1_y(rectangle1_ys[183]), .rectangle1_width(rectangle1_widths[183]), .rectangle1_height(rectangle1_heights[183]), .rectangle1_weight(rectangle1_weights[183]), .rectangle2_x(rectangle2_xs[183]), .rectangle2_y(rectangle2_ys[183]), .rectangle2_width(rectangle2_widths[183]), .rectangle2_height(rectangle2_heights[183]), .rectangle2_weight(rectangle2_weights[183]), .rectangle3_x(rectangle3_xs[183]), .rectangle3_y(rectangle3_ys[183]), .rectangle3_width(rectangle3_widths[183]), .rectangle3_height(rectangle3_heights[183]), .rectangle3_weight(rectangle3_weights[183]), .feature_threshold(feature_thresholds[183]), .feature_above(feature_aboves[183]), .feature_below(feature_belows[183]), .scan_win_std_dev(scan_win_std_dev[183]), .feature_accum(feature_accums[183]));
  accum_calculator ac184(.scan_win(scan_win184), .rectangle1_x(rectangle1_xs[184]), .rectangle1_y(rectangle1_ys[184]), .rectangle1_width(rectangle1_widths[184]), .rectangle1_height(rectangle1_heights[184]), .rectangle1_weight(rectangle1_weights[184]), .rectangle2_x(rectangle2_xs[184]), .rectangle2_y(rectangle2_ys[184]), .rectangle2_width(rectangle2_widths[184]), .rectangle2_height(rectangle2_heights[184]), .rectangle2_weight(rectangle2_weights[184]), .rectangle3_x(rectangle3_xs[184]), .rectangle3_y(rectangle3_ys[184]), .rectangle3_width(rectangle3_widths[184]), .rectangle3_height(rectangle3_heights[184]), .rectangle3_weight(rectangle3_weights[184]), .feature_threshold(feature_thresholds[184]), .feature_above(feature_aboves[184]), .feature_below(feature_belows[184]), .scan_win_std_dev(scan_win_std_dev[184]), .feature_accum(feature_accums[184]));
  accum_calculator ac185(.scan_win(scan_win185), .rectangle1_x(rectangle1_xs[185]), .rectangle1_y(rectangle1_ys[185]), .rectangle1_width(rectangle1_widths[185]), .rectangle1_height(rectangle1_heights[185]), .rectangle1_weight(rectangle1_weights[185]), .rectangle2_x(rectangle2_xs[185]), .rectangle2_y(rectangle2_ys[185]), .rectangle2_width(rectangle2_widths[185]), .rectangle2_height(rectangle2_heights[185]), .rectangle2_weight(rectangle2_weights[185]), .rectangle3_x(rectangle3_xs[185]), .rectangle3_y(rectangle3_ys[185]), .rectangle3_width(rectangle3_widths[185]), .rectangle3_height(rectangle3_heights[185]), .rectangle3_weight(rectangle3_weights[185]), .feature_threshold(feature_thresholds[185]), .feature_above(feature_aboves[185]), .feature_below(feature_belows[185]), .scan_win_std_dev(scan_win_std_dev[185]), .feature_accum(feature_accums[185]));
  accum_calculator ac186(.scan_win(scan_win186), .rectangle1_x(rectangle1_xs[186]), .rectangle1_y(rectangle1_ys[186]), .rectangle1_width(rectangle1_widths[186]), .rectangle1_height(rectangle1_heights[186]), .rectangle1_weight(rectangle1_weights[186]), .rectangle2_x(rectangle2_xs[186]), .rectangle2_y(rectangle2_ys[186]), .rectangle2_width(rectangle2_widths[186]), .rectangle2_height(rectangle2_heights[186]), .rectangle2_weight(rectangle2_weights[186]), .rectangle3_x(rectangle3_xs[186]), .rectangle3_y(rectangle3_ys[186]), .rectangle3_width(rectangle3_widths[186]), .rectangle3_height(rectangle3_heights[186]), .rectangle3_weight(rectangle3_weights[186]), .feature_threshold(feature_thresholds[186]), .feature_above(feature_aboves[186]), .feature_below(feature_belows[186]), .scan_win_std_dev(scan_win_std_dev[186]), .feature_accum(feature_accums[186]));
  accum_calculator ac187(.scan_win(scan_win187), .rectangle1_x(rectangle1_xs[187]), .rectangle1_y(rectangle1_ys[187]), .rectangle1_width(rectangle1_widths[187]), .rectangle1_height(rectangle1_heights[187]), .rectangle1_weight(rectangle1_weights[187]), .rectangle2_x(rectangle2_xs[187]), .rectangle2_y(rectangle2_ys[187]), .rectangle2_width(rectangle2_widths[187]), .rectangle2_height(rectangle2_heights[187]), .rectangle2_weight(rectangle2_weights[187]), .rectangle3_x(rectangle3_xs[187]), .rectangle3_y(rectangle3_ys[187]), .rectangle3_width(rectangle3_widths[187]), .rectangle3_height(rectangle3_heights[187]), .rectangle3_weight(rectangle3_weights[187]), .feature_threshold(feature_thresholds[187]), .feature_above(feature_aboves[187]), .feature_below(feature_belows[187]), .scan_win_std_dev(scan_win_std_dev[187]), .feature_accum(feature_accums[187]));
  accum_calculator ac188(.scan_win(scan_win188), .rectangle1_x(rectangle1_xs[188]), .rectangle1_y(rectangle1_ys[188]), .rectangle1_width(rectangle1_widths[188]), .rectangle1_height(rectangle1_heights[188]), .rectangle1_weight(rectangle1_weights[188]), .rectangle2_x(rectangle2_xs[188]), .rectangle2_y(rectangle2_ys[188]), .rectangle2_width(rectangle2_widths[188]), .rectangle2_height(rectangle2_heights[188]), .rectangle2_weight(rectangle2_weights[188]), .rectangle3_x(rectangle3_xs[188]), .rectangle3_y(rectangle3_ys[188]), .rectangle3_width(rectangle3_widths[188]), .rectangle3_height(rectangle3_heights[188]), .rectangle3_weight(rectangle3_weights[188]), .feature_threshold(feature_thresholds[188]), .feature_above(feature_aboves[188]), .feature_below(feature_belows[188]), .scan_win_std_dev(scan_win_std_dev[188]), .feature_accum(feature_accums[188]));
  accum_calculator ac189(.scan_win(scan_win189), .rectangle1_x(rectangle1_xs[189]), .rectangle1_y(rectangle1_ys[189]), .rectangle1_width(rectangle1_widths[189]), .rectangle1_height(rectangle1_heights[189]), .rectangle1_weight(rectangle1_weights[189]), .rectangle2_x(rectangle2_xs[189]), .rectangle2_y(rectangle2_ys[189]), .rectangle2_width(rectangle2_widths[189]), .rectangle2_height(rectangle2_heights[189]), .rectangle2_weight(rectangle2_weights[189]), .rectangle3_x(rectangle3_xs[189]), .rectangle3_y(rectangle3_ys[189]), .rectangle3_width(rectangle3_widths[189]), .rectangle3_height(rectangle3_heights[189]), .rectangle3_weight(rectangle3_weights[189]), .feature_threshold(feature_thresholds[189]), .feature_above(feature_aboves[189]), .feature_below(feature_belows[189]), .scan_win_std_dev(scan_win_std_dev[189]), .feature_accum(feature_accums[189]));
  accum_calculator ac190(.scan_win(scan_win190), .rectangle1_x(rectangle1_xs[190]), .rectangle1_y(rectangle1_ys[190]), .rectangle1_width(rectangle1_widths[190]), .rectangle1_height(rectangle1_heights[190]), .rectangle1_weight(rectangle1_weights[190]), .rectangle2_x(rectangle2_xs[190]), .rectangle2_y(rectangle2_ys[190]), .rectangle2_width(rectangle2_widths[190]), .rectangle2_height(rectangle2_heights[190]), .rectangle2_weight(rectangle2_weights[190]), .rectangle3_x(rectangle3_xs[190]), .rectangle3_y(rectangle3_ys[190]), .rectangle3_width(rectangle3_widths[190]), .rectangle3_height(rectangle3_heights[190]), .rectangle3_weight(rectangle3_weights[190]), .feature_threshold(feature_thresholds[190]), .feature_above(feature_aboves[190]), .feature_below(feature_belows[190]), .scan_win_std_dev(scan_win_std_dev[190]), .feature_accum(feature_accums[190]));
  accum_calculator ac191(.scan_win(scan_win191), .rectangle1_x(rectangle1_xs[191]), .rectangle1_y(rectangle1_ys[191]), .rectangle1_width(rectangle1_widths[191]), .rectangle1_height(rectangle1_heights[191]), .rectangle1_weight(rectangle1_weights[191]), .rectangle2_x(rectangle2_xs[191]), .rectangle2_y(rectangle2_ys[191]), .rectangle2_width(rectangle2_widths[191]), .rectangle2_height(rectangle2_heights[191]), .rectangle2_weight(rectangle2_weights[191]), .rectangle3_x(rectangle3_xs[191]), .rectangle3_y(rectangle3_ys[191]), .rectangle3_width(rectangle3_widths[191]), .rectangle3_height(rectangle3_heights[191]), .rectangle3_weight(rectangle3_weights[191]), .feature_threshold(feature_thresholds[191]), .feature_above(feature_aboves[191]), .feature_below(feature_belows[191]), .scan_win_std_dev(scan_win_std_dev[191]), .feature_accum(feature_accums[191]));
  accum_calculator ac192(.scan_win(scan_win192), .rectangle1_x(rectangle1_xs[192]), .rectangle1_y(rectangle1_ys[192]), .rectangle1_width(rectangle1_widths[192]), .rectangle1_height(rectangle1_heights[192]), .rectangle1_weight(rectangle1_weights[192]), .rectangle2_x(rectangle2_xs[192]), .rectangle2_y(rectangle2_ys[192]), .rectangle2_width(rectangle2_widths[192]), .rectangle2_height(rectangle2_heights[192]), .rectangle2_weight(rectangle2_weights[192]), .rectangle3_x(rectangle3_xs[192]), .rectangle3_y(rectangle3_ys[192]), .rectangle3_width(rectangle3_widths[192]), .rectangle3_height(rectangle3_heights[192]), .rectangle3_weight(rectangle3_weights[192]), .feature_threshold(feature_thresholds[192]), .feature_above(feature_aboves[192]), .feature_below(feature_belows[192]), .scan_win_std_dev(scan_win_std_dev[192]), .feature_accum(feature_accums[192]));
  accum_calculator ac193(.scan_win(scan_win193), .rectangle1_x(rectangle1_xs[193]), .rectangle1_y(rectangle1_ys[193]), .rectangle1_width(rectangle1_widths[193]), .rectangle1_height(rectangle1_heights[193]), .rectangle1_weight(rectangle1_weights[193]), .rectangle2_x(rectangle2_xs[193]), .rectangle2_y(rectangle2_ys[193]), .rectangle2_width(rectangle2_widths[193]), .rectangle2_height(rectangle2_heights[193]), .rectangle2_weight(rectangle2_weights[193]), .rectangle3_x(rectangle3_xs[193]), .rectangle3_y(rectangle3_ys[193]), .rectangle3_width(rectangle3_widths[193]), .rectangle3_height(rectangle3_heights[193]), .rectangle3_weight(rectangle3_weights[193]), .feature_threshold(feature_thresholds[193]), .feature_above(feature_aboves[193]), .feature_below(feature_belows[193]), .scan_win_std_dev(scan_win_std_dev[193]), .feature_accum(feature_accums[193]));
  accum_calculator ac194(.scan_win(scan_win194), .rectangle1_x(rectangle1_xs[194]), .rectangle1_y(rectangle1_ys[194]), .rectangle1_width(rectangle1_widths[194]), .rectangle1_height(rectangle1_heights[194]), .rectangle1_weight(rectangle1_weights[194]), .rectangle2_x(rectangle2_xs[194]), .rectangle2_y(rectangle2_ys[194]), .rectangle2_width(rectangle2_widths[194]), .rectangle2_height(rectangle2_heights[194]), .rectangle2_weight(rectangle2_weights[194]), .rectangle3_x(rectangle3_xs[194]), .rectangle3_y(rectangle3_ys[194]), .rectangle3_width(rectangle3_widths[194]), .rectangle3_height(rectangle3_heights[194]), .rectangle3_weight(rectangle3_weights[194]), .feature_threshold(feature_thresholds[194]), .feature_above(feature_aboves[194]), .feature_below(feature_belows[194]), .scan_win_std_dev(scan_win_std_dev[194]), .feature_accum(feature_accums[194]));
  accum_calculator ac195(.scan_win(scan_win195), .rectangle1_x(rectangle1_xs[195]), .rectangle1_y(rectangle1_ys[195]), .rectangle1_width(rectangle1_widths[195]), .rectangle1_height(rectangle1_heights[195]), .rectangle1_weight(rectangle1_weights[195]), .rectangle2_x(rectangle2_xs[195]), .rectangle2_y(rectangle2_ys[195]), .rectangle2_width(rectangle2_widths[195]), .rectangle2_height(rectangle2_heights[195]), .rectangle2_weight(rectangle2_weights[195]), .rectangle3_x(rectangle3_xs[195]), .rectangle3_y(rectangle3_ys[195]), .rectangle3_width(rectangle3_widths[195]), .rectangle3_height(rectangle3_heights[195]), .rectangle3_weight(rectangle3_weights[195]), .feature_threshold(feature_thresholds[195]), .feature_above(feature_aboves[195]), .feature_below(feature_belows[195]), .scan_win_std_dev(scan_win_std_dev[195]), .feature_accum(feature_accums[195]));
  accum_calculator ac196(.scan_win(scan_win196), .rectangle1_x(rectangle1_xs[196]), .rectangle1_y(rectangle1_ys[196]), .rectangle1_width(rectangle1_widths[196]), .rectangle1_height(rectangle1_heights[196]), .rectangle1_weight(rectangle1_weights[196]), .rectangle2_x(rectangle2_xs[196]), .rectangle2_y(rectangle2_ys[196]), .rectangle2_width(rectangle2_widths[196]), .rectangle2_height(rectangle2_heights[196]), .rectangle2_weight(rectangle2_weights[196]), .rectangle3_x(rectangle3_xs[196]), .rectangle3_y(rectangle3_ys[196]), .rectangle3_width(rectangle3_widths[196]), .rectangle3_height(rectangle3_heights[196]), .rectangle3_weight(rectangle3_weights[196]), .feature_threshold(feature_thresholds[196]), .feature_above(feature_aboves[196]), .feature_below(feature_belows[196]), .scan_win_std_dev(scan_win_std_dev[196]), .feature_accum(feature_accums[196]));
  accum_calculator ac197(.scan_win(scan_win197), .rectangle1_x(rectangle1_xs[197]), .rectangle1_y(rectangle1_ys[197]), .rectangle1_width(rectangle1_widths[197]), .rectangle1_height(rectangle1_heights[197]), .rectangle1_weight(rectangle1_weights[197]), .rectangle2_x(rectangle2_xs[197]), .rectangle2_y(rectangle2_ys[197]), .rectangle2_width(rectangle2_widths[197]), .rectangle2_height(rectangle2_heights[197]), .rectangle2_weight(rectangle2_weights[197]), .rectangle3_x(rectangle3_xs[197]), .rectangle3_y(rectangle3_ys[197]), .rectangle3_width(rectangle3_widths[197]), .rectangle3_height(rectangle3_heights[197]), .rectangle3_weight(rectangle3_weights[197]), .feature_threshold(feature_thresholds[197]), .feature_above(feature_aboves[197]), .feature_below(feature_belows[197]), .scan_win_std_dev(scan_win_std_dev[197]), .feature_accum(feature_accums[197]));
  accum_calculator ac198(.scan_win(scan_win198), .rectangle1_x(rectangle1_xs[198]), .rectangle1_y(rectangle1_ys[198]), .rectangle1_width(rectangle1_widths[198]), .rectangle1_height(rectangle1_heights[198]), .rectangle1_weight(rectangle1_weights[198]), .rectangle2_x(rectangle2_xs[198]), .rectangle2_y(rectangle2_ys[198]), .rectangle2_width(rectangle2_widths[198]), .rectangle2_height(rectangle2_heights[198]), .rectangle2_weight(rectangle2_weights[198]), .rectangle3_x(rectangle3_xs[198]), .rectangle3_y(rectangle3_ys[198]), .rectangle3_width(rectangle3_widths[198]), .rectangle3_height(rectangle3_heights[198]), .rectangle3_weight(rectangle3_weights[198]), .feature_threshold(feature_thresholds[198]), .feature_above(feature_aboves[198]), .feature_below(feature_belows[198]), .scan_win_std_dev(scan_win_std_dev[198]), .feature_accum(feature_accums[198]));
  accum_calculator ac199(.scan_win(scan_win199), .rectangle1_x(rectangle1_xs[199]), .rectangle1_y(rectangle1_ys[199]), .rectangle1_width(rectangle1_widths[199]), .rectangle1_height(rectangle1_heights[199]), .rectangle1_weight(rectangle1_weights[199]), .rectangle2_x(rectangle2_xs[199]), .rectangle2_y(rectangle2_ys[199]), .rectangle2_width(rectangle2_widths[199]), .rectangle2_height(rectangle2_heights[199]), .rectangle2_weight(rectangle2_weights[199]), .rectangle3_x(rectangle3_xs[199]), .rectangle3_y(rectangle3_ys[199]), .rectangle3_width(rectangle3_widths[199]), .rectangle3_height(rectangle3_heights[199]), .rectangle3_weight(rectangle3_weights[199]), .feature_threshold(feature_thresholds[199]), .feature_above(feature_aboves[199]), .feature_below(feature_belows[199]), .scan_win_std_dev(scan_win_std_dev[199]), .feature_accum(feature_accums[199]));
  accum_calculator ac200(.scan_win(scan_win200), .rectangle1_x(rectangle1_xs[200]), .rectangle1_y(rectangle1_ys[200]), .rectangle1_width(rectangle1_widths[200]), .rectangle1_height(rectangle1_heights[200]), .rectangle1_weight(rectangle1_weights[200]), .rectangle2_x(rectangle2_xs[200]), .rectangle2_y(rectangle2_ys[200]), .rectangle2_width(rectangle2_widths[200]), .rectangle2_height(rectangle2_heights[200]), .rectangle2_weight(rectangle2_weights[200]), .rectangle3_x(rectangle3_xs[200]), .rectangle3_y(rectangle3_ys[200]), .rectangle3_width(rectangle3_widths[200]), .rectangle3_height(rectangle3_heights[200]), .rectangle3_weight(rectangle3_weights[200]), .feature_threshold(feature_thresholds[200]), .feature_above(feature_aboves[200]), .feature_below(feature_belows[200]), .scan_win_std_dev(scan_win_std_dev[200]), .feature_accum(feature_accums[200]));
  accum_calculator ac201(.scan_win(scan_win201), .rectangle1_x(rectangle1_xs[201]), .rectangle1_y(rectangle1_ys[201]), .rectangle1_width(rectangle1_widths[201]), .rectangle1_height(rectangle1_heights[201]), .rectangle1_weight(rectangle1_weights[201]), .rectangle2_x(rectangle2_xs[201]), .rectangle2_y(rectangle2_ys[201]), .rectangle2_width(rectangle2_widths[201]), .rectangle2_height(rectangle2_heights[201]), .rectangle2_weight(rectangle2_weights[201]), .rectangle3_x(rectangle3_xs[201]), .rectangle3_y(rectangle3_ys[201]), .rectangle3_width(rectangle3_widths[201]), .rectangle3_height(rectangle3_heights[201]), .rectangle3_weight(rectangle3_weights[201]), .feature_threshold(feature_thresholds[201]), .feature_above(feature_aboves[201]), .feature_below(feature_belows[201]), .scan_win_std_dev(scan_win_std_dev[201]), .feature_accum(feature_accums[201]));
  accum_calculator ac202(.scan_win(scan_win202), .rectangle1_x(rectangle1_xs[202]), .rectangle1_y(rectangle1_ys[202]), .rectangle1_width(rectangle1_widths[202]), .rectangle1_height(rectangle1_heights[202]), .rectangle1_weight(rectangle1_weights[202]), .rectangle2_x(rectangle2_xs[202]), .rectangle2_y(rectangle2_ys[202]), .rectangle2_width(rectangle2_widths[202]), .rectangle2_height(rectangle2_heights[202]), .rectangle2_weight(rectangle2_weights[202]), .rectangle3_x(rectangle3_xs[202]), .rectangle3_y(rectangle3_ys[202]), .rectangle3_width(rectangle3_widths[202]), .rectangle3_height(rectangle3_heights[202]), .rectangle3_weight(rectangle3_weights[202]), .feature_threshold(feature_thresholds[202]), .feature_above(feature_aboves[202]), .feature_below(feature_belows[202]), .scan_win_std_dev(scan_win_std_dev[202]), .feature_accum(feature_accums[202]));
  accum_calculator ac203(.scan_win(scan_win203), .rectangle1_x(rectangle1_xs[203]), .rectangle1_y(rectangle1_ys[203]), .rectangle1_width(rectangle1_widths[203]), .rectangle1_height(rectangle1_heights[203]), .rectangle1_weight(rectangle1_weights[203]), .rectangle2_x(rectangle2_xs[203]), .rectangle2_y(rectangle2_ys[203]), .rectangle2_width(rectangle2_widths[203]), .rectangle2_height(rectangle2_heights[203]), .rectangle2_weight(rectangle2_weights[203]), .rectangle3_x(rectangle3_xs[203]), .rectangle3_y(rectangle3_ys[203]), .rectangle3_width(rectangle3_widths[203]), .rectangle3_height(rectangle3_heights[203]), .rectangle3_weight(rectangle3_weights[203]), .feature_threshold(feature_thresholds[203]), .feature_above(feature_aboves[203]), .feature_below(feature_belows[203]), .scan_win_std_dev(scan_win_std_dev[203]), .feature_accum(feature_accums[203]));
  accum_calculator ac204(.scan_win(scan_win204), .rectangle1_x(rectangle1_xs[204]), .rectangle1_y(rectangle1_ys[204]), .rectangle1_width(rectangle1_widths[204]), .rectangle1_height(rectangle1_heights[204]), .rectangle1_weight(rectangle1_weights[204]), .rectangle2_x(rectangle2_xs[204]), .rectangle2_y(rectangle2_ys[204]), .rectangle2_width(rectangle2_widths[204]), .rectangle2_height(rectangle2_heights[204]), .rectangle2_weight(rectangle2_weights[204]), .rectangle3_x(rectangle3_xs[204]), .rectangle3_y(rectangle3_ys[204]), .rectangle3_width(rectangle3_widths[204]), .rectangle3_height(rectangle3_heights[204]), .rectangle3_weight(rectangle3_weights[204]), .feature_threshold(feature_thresholds[204]), .feature_above(feature_aboves[204]), .feature_below(feature_belows[204]), .scan_win_std_dev(scan_win_std_dev[204]), .feature_accum(feature_accums[204]));
  accum_calculator ac205(.scan_win(scan_win205), .rectangle1_x(rectangle1_xs[205]), .rectangle1_y(rectangle1_ys[205]), .rectangle1_width(rectangle1_widths[205]), .rectangle1_height(rectangle1_heights[205]), .rectangle1_weight(rectangle1_weights[205]), .rectangle2_x(rectangle2_xs[205]), .rectangle2_y(rectangle2_ys[205]), .rectangle2_width(rectangle2_widths[205]), .rectangle2_height(rectangle2_heights[205]), .rectangle2_weight(rectangle2_weights[205]), .rectangle3_x(rectangle3_xs[205]), .rectangle3_y(rectangle3_ys[205]), .rectangle3_width(rectangle3_widths[205]), .rectangle3_height(rectangle3_heights[205]), .rectangle3_weight(rectangle3_weights[205]), .feature_threshold(feature_thresholds[205]), .feature_above(feature_aboves[205]), .feature_below(feature_belows[205]), .scan_win_std_dev(scan_win_std_dev[205]), .feature_accum(feature_accums[205]));
  accum_calculator ac206(.scan_win(scan_win206), .rectangle1_x(rectangle1_xs[206]), .rectangle1_y(rectangle1_ys[206]), .rectangle1_width(rectangle1_widths[206]), .rectangle1_height(rectangle1_heights[206]), .rectangle1_weight(rectangle1_weights[206]), .rectangle2_x(rectangle2_xs[206]), .rectangle2_y(rectangle2_ys[206]), .rectangle2_width(rectangle2_widths[206]), .rectangle2_height(rectangle2_heights[206]), .rectangle2_weight(rectangle2_weights[206]), .rectangle3_x(rectangle3_xs[206]), .rectangle3_y(rectangle3_ys[206]), .rectangle3_width(rectangle3_widths[206]), .rectangle3_height(rectangle3_heights[206]), .rectangle3_weight(rectangle3_weights[206]), .feature_threshold(feature_thresholds[206]), .feature_above(feature_aboves[206]), .feature_below(feature_belows[206]), .scan_win_std_dev(scan_win_std_dev[206]), .feature_accum(feature_accums[206]));
  accum_calculator ac207(.scan_win(scan_win207), .rectangle1_x(rectangle1_xs[207]), .rectangle1_y(rectangle1_ys[207]), .rectangle1_width(rectangle1_widths[207]), .rectangle1_height(rectangle1_heights[207]), .rectangle1_weight(rectangle1_weights[207]), .rectangle2_x(rectangle2_xs[207]), .rectangle2_y(rectangle2_ys[207]), .rectangle2_width(rectangle2_widths[207]), .rectangle2_height(rectangle2_heights[207]), .rectangle2_weight(rectangle2_weights[207]), .rectangle3_x(rectangle3_xs[207]), .rectangle3_y(rectangle3_ys[207]), .rectangle3_width(rectangle3_widths[207]), .rectangle3_height(rectangle3_heights[207]), .rectangle3_weight(rectangle3_weights[207]), .feature_threshold(feature_thresholds[207]), .feature_above(feature_aboves[207]), .feature_below(feature_belows[207]), .scan_win_std_dev(scan_win_std_dev[207]), .feature_accum(feature_accums[207]));
  accum_calculator ac208(.scan_win(scan_win208), .rectangle1_x(rectangle1_xs[208]), .rectangle1_y(rectangle1_ys[208]), .rectangle1_width(rectangle1_widths[208]), .rectangle1_height(rectangle1_heights[208]), .rectangle1_weight(rectangle1_weights[208]), .rectangle2_x(rectangle2_xs[208]), .rectangle2_y(rectangle2_ys[208]), .rectangle2_width(rectangle2_widths[208]), .rectangle2_height(rectangle2_heights[208]), .rectangle2_weight(rectangle2_weights[208]), .rectangle3_x(rectangle3_xs[208]), .rectangle3_y(rectangle3_ys[208]), .rectangle3_width(rectangle3_widths[208]), .rectangle3_height(rectangle3_heights[208]), .rectangle3_weight(rectangle3_weights[208]), .feature_threshold(feature_thresholds[208]), .feature_above(feature_aboves[208]), .feature_below(feature_belows[208]), .scan_win_std_dev(scan_win_std_dev[208]), .feature_accum(feature_accums[208]));
  accum_calculator ac209(.scan_win(scan_win209), .rectangle1_x(rectangle1_xs[209]), .rectangle1_y(rectangle1_ys[209]), .rectangle1_width(rectangle1_widths[209]), .rectangle1_height(rectangle1_heights[209]), .rectangle1_weight(rectangle1_weights[209]), .rectangle2_x(rectangle2_xs[209]), .rectangle2_y(rectangle2_ys[209]), .rectangle2_width(rectangle2_widths[209]), .rectangle2_height(rectangle2_heights[209]), .rectangle2_weight(rectangle2_weights[209]), .rectangle3_x(rectangle3_xs[209]), .rectangle3_y(rectangle3_ys[209]), .rectangle3_width(rectangle3_widths[209]), .rectangle3_height(rectangle3_heights[209]), .rectangle3_weight(rectangle3_weights[209]), .feature_threshold(feature_thresholds[209]), .feature_above(feature_aboves[209]), .feature_below(feature_belows[209]), .scan_win_std_dev(scan_win_std_dev[209]), .feature_accum(feature_accums[209]));
  accum_calculator ac210(.scan_win(scan_win210), .rectangle1_x(rectangle1_xs[210]), .rectangle1_y(rectangle1_ys[210]), .rectangle1_width(rectangle1_widths[210]), .rectangle1_height(rectangle1_heights[210]), .rectangle1_weight(rectangle1_weights[210]), .rectangle2_x(rectangle2_xs[210]), .rectangle2_y(rectangle2_ys[210]), .rectangle2_width(rectangle2_widths[210]), .rectangle2_height(rectangle2_heights[210]), .rectangle2_weight(rectangle2_weights[210]), .rectangle3_x(rectangle3_xs[210]), .rectangle3_y(rectangle3_ys[210]), .rectangle3_width(rectangle3_widths[210]), .rectangle3_height(rectangle3_heights[210]), .rectangle3_weight(rectangle3_weights[210]), .feature_threshold(feature_thresholds[210]), .feature_above(feature_aboves[210]), .feature_below(feature_belows[210]), .scan_win_std_dev(scan_win_std_dev[210]), .feature_accum(feature_accums[210]));
  accum_calculator ac211(.scan_win(scan_win211), .rectangle1_x(rectangle1_xs[211]), .rectangle1_y(rectangle1_ys[211]), .rectangle1_width(rectangle1_widths[211]), .rectangle1_height(rectangle1_heights[211]), .rectangle1_weight(rectangle1_weights[211]), .rectangle2_x(rectangle2_xs[211]), .rectangle2_y(rectangle2_ys[211]), .rectangle2_width(rectangle2_widths[211]), .rectangle2_height(rectangle2_heights[211]), .rectangle2_weight(rectangle2_weights[211]), .rectangle3_x(rectangle3_xs[211]), .rectangle3_y(rectangle3_ys[211]), .rectangle3_width(rectangle3_widths[211]), .rectangle3_height(rectangle3_heights[211]), .rectangle3_weight(rectangle3_weights[211]), .feature_threshold(feature_thresholds[211]), .feature_above(feature_aboves[211]), .feature_below(feature_belows[211]), .scan_win_std_dev(scan_win_std_dev[211]), .feature_accum(feature_accums[211]));
  accum_calculator ac212(.scan_win(scan_win212), .rectangle1_x(rectangle1_xs[212]), .rectangle1_y(rectangle1_ys[212]), .rectangle1_width(rectangle1_widths[212]), .rectangle1_height(rectangle1_heights[212]), .rectangle1_weight(rectangle1_weights[212]), .rectangle2_x(rectangle2_xs[212]), .rectangle2_y(rectangle2_ys[212]), .rectangle2_width(rectangle2_widths[212]), .rectangle2_height(rectangle2_heights[212]), .rectangle2_weight(rectangle2_weights[212]), .rectangle3_x(rectangle3_xs[212]), .rectangle3_y(rectangle3_ys[212]), .rectangle3_width(rectangle3_widths[212]), .rectangle3_height(rectangle3_heights[212]), .rectangle3_weight(rectangle3_weights[212]), .feature_threshold(feature_thresholds[212]), .feature_above(feature_aboves[212]), .feature_below(feature_belows[212]), .scan_win_std_dev(scan_win_std_dev[212]), .feature_accum(feature_accums[212]));
  accum_calculator ac213(.scan_win(scan_win213), .rectangle1_x(rectangle1_xs[213]), .rectangle1_y(rectangle1_ys[213]), .rectangle1_width(rectangle1_widths[213]), .rectangle1_height(rectangle1_heights[213]), .rectangle1_weight(rectangle1_weights[213]), .rectangle2_x(rectangle2_xs[213]), .rectangle2_y(rectangle2_ys[213]), .rectangle2_width(rectangle2_widths[213]), .rectangle2_height(rectangle2_heights[213]), .rectangle2_weight(rectangle2_weights[213]), .rectangle3_x(rectangle3_xs[213]), .rectangle3_y(rectangle3_ys[213]), .rectangle3_width(rectangle3_widths[213]), .rectangle3_height(rectangle3_heights[213]), .rectangle3_weight(rectangle3_weights[213]), .feature_threshold(feature_thresholds[213]), .feature_above(feature_aboves[213]), .feature_below(feature_belows[213]), .scan_win_std_dev(scan_win_std_dev[213]), .feature_accum(feature_accums[213]));
  accum_calculator ac214(.scan_win(scan_win214), .rectangle1_x(rectangle1_xs[214]), .rectangle1_y(rectangle1_ys[214]), .rectangle1_width(rectangle1_widths[214]), .rectangle1_height(rectangle1_heights[214]), .rectangle1_weight(rectangle1_weights[214]), .rectangle2_x(rectangle2_xs[214]), .rectangle2_y(rectangle2_ys[214]), .rectangle2_width(rectangle2_widths[214]), .rectangle2_height(rectangle2_heights[214]), .rectangle2_weight(rectangle2_weights[214]), .rectangle3_x(rectangle3_xs[214]), .rectangle3_y(rectangle3_ys[214]), .rectangle3_width(rectangle3_widths[214]), .rectangle3_height(rectangle3_heights[214]), .rectangle3_weight(rectangle3_weights[214]), .feature_threshold(feature_thresholds[214]), .feature_above(feature_aboves[214]), .feature_below(feature_belows[214]), .scan_win_std_dev(scan_win_std_dev[214]), .feature_accum(feature_accums[214]));
  accum_calculator ac215(.scan_win(scan_win215), .rectangle1_x(rectangle1_xs[215]), .rectangle1_y(rectangle1_ys[215]), .rectangle1_width(rectangle1_widths[215]), .rectangle1_height(rectangle1_heights[215]), .rectangle1_weight(rectangle1_weights[215]), .rectangle2_x(rectangle2_xs[215]), .rectangle2_y(rectangle2_ys[215]), .rectangle2_width(rectangle2_widths[215]), .rectangle2_height(rectangle2_heights[215]), .rectangle2_weight(rectangle2_weights[215]), .rectangle3_x(rectangle3_xs[215]), .rectangle3_y(rectangle3_ys[215]), .rectangle3_width(rectangle3_widths[215]), .rectangle3_height(rectangle3_heights[215]), .rectangle3_weight(rectangle3_weights[215]), .feature_threshold(feature_thresholds[215]), .feature_above(feature_aboves[215]), .feature_below(feature_belows[215]), .scan_win_std_dev(scan_win_std_dev[215]), .feature_accum(feature_accums[215]));
  accum_calculator ac216(.scan_win(scan_win216), .rectangle1_x(rectangle1_xs[216]), .rectangle1_y(rectangle1_ys[216]), .rectangle1_width(rectangle1_widths[216]), .rectangle1_height(rectangle1_heights[216]), .rectangle1_weight(rectangle1_weights[216]), .rectangle2_x(rectangle2_xs[216]), .rectangle2_y(rectangle2_ys[216]), .rectangle2_width(rectangle2_widths[216]), .rectangle2_height(rectangle2_heights[216]), .rectangle2_weight(rectangle2_weights[216]), .rectangle3_x(rectangle3_xs[216]), .rectangle3_y(rectangle3_ys[216]), .rectangle3_width(rectangle3_widths[216]), .rectangle3_height(rectangle3_heights[216]), .rectangle3_weight(rectangle3_weights[216]), .feature_threshold(feature_thresholds[216]), .feature_above(feature_aboves[216]), .feature_below(feature_belows[216]), .scan_win_std_dev(scan_win_std_dev[216]), .feature_accum(feature_accums[216]));
  accum_calculator ac217(.scan_win(scan_win217), .rectangle1_x(rectangle1_xs[217]), .rectangle1_y(rectangle1_ys[217]), .rectangle1_width(rectangle1_widths[217]), .rectangle1_height(rectangle1_heights[217]), .rectangle1_weight(rectangle1_weights[217]), .rectangle2_x(rectangle2_xs[217]), .rectangle2_y(rectangle2_ys[217]), .rectangle2_width(rectangle2_widths[217]), .rectangle2_height(rectangle2_heights[217]), .rectangle2_weight(rectangle2_weights[217]), .rectangle3_x(rectangle3_xs[217]), .rectangle3_y(rectangle3_ys[217]), .rectangle3_width(rectangle3_widths[217]), .rectangle3_height(rectangle3_heights[217]), .rectangle3_weight(rectangle3_weights[217]), .feature_threshold(feature_thresholds[217]), .feature_above(feature_aboves[217]), .feature_below(feature_belows[217]), .scan_win_std_dev(scan_win_std_dev[217]), .feature_accum(feature_accums[217]));
  accum_calculator ac218(.scan_win(scan_win218), .rectangle1_x(rectangle1_xs[218]), .rectangle1_y(rectangle1_ys[218]), .rectangle1_width(rectangle1_widths[218]), .rectangle1_height(rectangle1_heights[218]), .rectangle1_weight(rectangle1_weights[218]), .rectangle2_x(rectangle2_xs[218]), .rectangle2_y(rectangle2_ys[218]), .rectangle2_width(rectangle2_widths[218]), .rectangle2_height(rectangle2_heights[218]), .rectangle2_weight(rectangle2_weights[218]), .rectangle3_x(rectangle3_xs[218]), .rectangle3_y(rectangle3_ys[218]), .rectangle3_width(rectangle3_widths[218]), .rectangle3_height(rectangle3_heights[218]), .rectangle3_weight(rectangle3_weights[218]), .feature_threshold(feature_thresholds[218]), .feature_above(feature_aboves[218]), .feature_below(feature_belows[218]), .scan_win_std_dev(scan_win_std_dev[218]), .feature_accum(feature_accums[218]));
  accum_calculator ac219(.scan_win(scan_win219), .rectangle1_x(rectangle1_xs[219]), .rectangle1_y(rectangle1_ys[219]), .rectangle1_width(rectangle1_widths[219]), .rectangle1_height(rectangle1_heights[219]), .rectangle1_weight(rectangle1_weights[219]), .rectangle2_x(rectangle2_xs[219]), .rectangle2_y(rectangle2_ys[219]), .rectangle2_width(rectangle2_widths[219]), .rectangle2_height(rectangle2_heights[219]), .rectangle2_weight(rectangle2_weights[219]), .rectangle3_x(rectangle3_xs[219]), .rectangle3_y(rectangle3_ys[219]), .rectangle3_width(rectangle3_widths[219]), .rectangle3_height(rectangle3_heights[219]), .rectangle3_weight(rectangle3_weights[219]), .feature_threshold(feature_thresholds[219]), .feature_above(feature_aboves[219]), .feature_below(feature_belows[219]), .scan_win_std_dev(scan_win_std_dev[219]), .feature_accum(feature_accums[219]));
  accum_calculator ac220(.scan_win(scan_win220), .rectangle1_x(rectangle1_xs[220]), .rectangle1_y(rectangle1_ys[220]), .rectangle1_width(rectangle1_widths[220]), .rectangle1_height(rectangle1_heights[220]), .rectangle1_weight(rectangle1_weights[220]), .rectangle2_x(rectangle2_xs[220]), .rectangle2_y(rectangle2_ys[220]), .rectangle2_width(rectangle2_widths[220]), .rectangle2_height(rectangle2_heights[220]), .rectangle2_weight(rectangle2_weights[220]), .rectangle3_x(rectangle3_xs[220]), .rectangle3_y(rectangle3_ys[220]), .rectangle3_width(rectangle3_widths[220]), .rectangle3_height(rectangle3_heights[220]), .rectangle3_weight(rectangle3_weights[220]), .feature_threshold(feature_thresholds[220]), .feature_above(feature_aboves[220]), .feature_below(feature_belows[220]), .scan_win_std_dev(scan_win_std_dev[220]), .feature_accum(feature_accums[220]));
  accum_calculator ac221(.scan_win(scan_win221), .rectangle1_x(rectangle1_xs[221]), .rectangle1_y(rectangle1_ys[221]), .rectangle1_width(rectangle1_widths[221]), .rectangle1_height(rectangle1_heights[221]), .rectangle1_weight(rectangle1_weights[221]), .rectangle2_x(rectangle2_xs[221]), .rectangle2_y(rectangle2_ys[221]), .rectangle2_width(rectangle2_widths[221]), .rectangle2_height(rectangle2_heights[221]), .rectangle2_weight(rectangle2_weights[221]), .rectangle3_x(rectangle3_xs[221]), .rectangle3_y(rectangle3_ys[221]), .rectangle3_width(rectangle3_widths[221]), .rectangle3_height(rectangle3_heights[221]), .rectangle3_weight(rectangle3_weights[221]), .feature_threshold(feature_thresholds[221]), .feature_above(feature_aboves[221]), .feature_below(feature_belows[221]), .scan_win_std_dev(scan_win_std_dev[221]), .feature_accum(feature_accums[221]));
  accum_calculator ac222(.scan_win(scan_win222), .rectangle1_x(rectangle1_xs[222]), .rectangle1_y(rectangle1_ys[222]), .rectangle1_width(rectangle1_widths[222]), .rectangle1_height(rectangle1_heights[222]), .rectangle1_weight(rectangle1_weights[222]), .rectangle2_x(rectangle2_xs[222]), .rectangle2_y(rectangle2_ys[222]), .rectangle2_width(rectangle2_widths[222]), .rectangle2_height(rectangle2_heights[222]), .rectangle2_weight(rectangle2_weights[222]), .rectangle3_x(rectangle3_xs[222]), .rectangle3_y(rectangle3_ys[222]), .rectangle3_width(rectangle3_widths[222]), .rectangle3_height(rectangle3_heights[222]), .rectangle3_weight(rectangle3_weights[222]), .feature_threshold(feature_thresholds[222]), .feature_above(feature_aboves[222]), .feature_below(feature_belows[222]), .scan_win_std_dev(scan_win_std_dev[222]), .feature_accum(feature_accums[222]));
  accum_calculator ac223(.scan_win(scan_win223), .rectangle1_x(rectangle1_xs[223]), .rectangle1_y(rectangle1_ys[223]), .rectangle1_width(rectangle1_widths[223]), .rectangle1_height(rectangle1_heights[223]), .rectangle1_weight(rectangle1_weights[223]), .rectangle2_x(rectangle2_xs[223]), .rectangle2_y(rectangle2_ys[223]), .rectangle2_width(rectangle2_widths[223]), .rectangle2_height(rectangle2_heights[223]), .rectangle2_weight(rectangle2_weights[223]), .rectangle3_x(rectangle3_xs[223]), .rectangle3_y(rectangle3_ys[223]), .rectangle3_width(rectangle3_widths[223]), .rectangle3_height(rectangle3_heights[223]), .rectangle3_weight(rectangle3_weights[223]), .feature_threshold(feature_thresholds[223]), .feature_above(feature_aboves[223]), .feature_below(feature_belows[223]), .scan_win_std_dev(scan_win_std_dev[223]), .feature_accum(feature_accums[223]));
  accum_calculator ac224(.scan_win(scan_win224), .rectangle1_x(rectangle1_xs[224]), .rectangle1_y(rectangle1_ys[224]), .rectangle1_width(rectangle1_widths[224]), .rectangle1_height(rectangle1_heights[224]), .rectangle1_weight(rectangle1_weights[224]), .rectangle2_x(rectangle2_xs[224]), .rectangle2_y(rectangle2_ys[224]), .rectangle2_width(rectangle2_widths[224]), .rectangle2_height(rectangle2_heights[224]), .rectangle2_weight(rectangle2_weights[224]), .rectangle3_x(rectangle3_xs[224]), .rectangle3_y(rectangle3_ys[224]), .rectangle3_width(rectangle3_widths[224]), .rectangle3_height(rectangle3_heights[224]), .rectangle3_weight(rectangle3_weights[224]), .feature_threshold(feature_thresholds[224]), .feature_above(feature_aboves[224]), .feature_below(feature_belows[224]), .scan_win_std_dev(scan_win_std_dev[224]), .feature_accum(feature_accums[224]));
  accum_calculator ac225(.scan_win(scan_win225), .rectangle1_x(rectangle1_xs[225]), .rectangle1_y(rectangle1_ys[225]), .rectangle1_width(rectangle1_widths[225]), .rectangle1_height(rectangle1_heights[225]), .rectangle1_weight(rectangle1_weights[225]), .rectangle2_x(rectangle2_xs[225]), .rectangle2_y(rectangle2_ys[225]), .rectangle2_width(rectangle2_widths[225]), .rectangle2_height(rectangle2_heights[225]), .rectangle2_weight(rectangle2_weights[225]), .rectangle3_x(rectangle3_xs[225]), .rectangle3_y(rectangle3_ys[225]), .rectangle3_width(rectangle3_widths[225]), .rectangle3_height(rectangle3_heights[225]), .rectangle3_weight(rectangle3_weights[225]), .feature_threshold(feature_thresholds[225]), .feature_above(feature_aboves[225]), .feature_below(feature_belows[225]), .scan_win_std_dev(scan_win_std_dev[225]), .feature_accum(feature_accums[225]));
  accum_calculator ac226(.scan_win(scan_win226), .rectangle1_x(rectangle1_xs[226]), .rectangle1_y(rectangle1_ys[226]), .rectangle1_width(rectangle1_widths[226]), .rectangle1_height(rectangle1_heights[226]), .rectangle1_weight(rectangle1_weights[226]), .rectangle2_x(rectangle2_xs[226]), .rectangle2_y(rectangle2_ys[226]), .rectangle2_width(rectangle2_widths[226]), .rectangle2_height(rectangle2_heights[226]), .rectangle2_weight(rectangle2_weights[226]), .rectangle3_x(rectangle3_xs[226]), .rectangle3_y(rectangle3_ys[226]), .rectangle3_width(rectangle3_widths[226]), .rectangle3_height(rectangle3_heights[226]), .rectangle3_weight(rectangle3_weights[226]), .feature_threshold(feature_thresholds[226]), .feature_above(feature_aboves[226]), .feature_below(feature_belows[226]), .scan_win_std_dev(scan_win_std_dev[226]), .feature_accum(feature_accums[226]));
  accum_calculator ac227(.scan_win(scan_win227), .rectangle1_x(rectangle1_xs[227]), .rectangle1_y(rectangle1_ys[227]), .rectangle1_width(rectangle1_widths[227]), .rectangle1_height(rectangle1_heights[227]), .rectangle1_weight(rectangle1_weights[227]), .rectangle2_x(rectangle2_xs[227]), .rectangle2_y(rectangle2_ys[227]), .rectangle2_width(rectangle2_widths[227]), .rectangle2_height(rectangle2_heights[227]), .rectangle2_weight(rectangle2_weights[227]), .rectangle3_x(rectangle3_xs[227]), .rectangle3_y(rectangle3_ys[227]), .rectangle3_width(rectangle3_widths[227]), .rectangle3_height(rectangle3_heights[227]), .rectangle3_weight(rectangle3_weights[227]), .feature_threshold(feature_thresholds[227]), .feature_above(feature_aboves[227]), .feature_below(feature_belows[227]), .scan_win_std_dev(scan_win_std_dev[227]), .feature_accum(feature_accums[227]));
  accum_calculator ac228(.scan_win(scan_win228), .rectangle1_x(rectangle1_xs[228]), .rectangle1_y(rectangle1_ys[228]), .rectangle1_width(rectangle1_widths[228]), .rectangle1_height(rectangle1_heights[228]), .rectangle1_weight(rectangle1_weights[228]), .rectangle2_x(rectangle2_xs[228]), .rectangle2_y(rectangle2_ys[228]), .rectangle2_width(rectangle2_widths[228]), .rectangle2_height(rectangle2_heights[228]), .rectangle2_weight(rectangle2_weights[228]), .rectangle3_x(rectangle3_xs[228]), .rectangle3_y(rectangle3_ys[228]), .rectangle3_width(rectangle3_widths[228]), .rectangle3_height(rectangle3_heights[228]), .rectangle3_weight(rectangle3_weights[228]), .feature_threshold(feature_thresholds[228]), .feature_above(feature_aboves[228]), .feature_below(feature_belows[228]), .scan_win_std_dev(scan_win_std_dev[228]), .feature_accum(feature_accums[228]));
  accum_calculator ac229(.scan_win(scan_win229), .rectangle1_x(rectangle1_xs[229]), .rectangle1_y(rectangle1_ys[229]), .rectangle1_width(rectangle1_widths[229]), .rectangle1_height(rectangle1_heights[229]), .rectangle1_weight(rectangle1_weights[229]), .rectangle2_x(rectangle2_xs[229]), .rectangle2_y(rectangle2_ys[229]), .rectangle2_width(rectangle2_widths[229]), .rectangle2_height(rectangle2_heights[229]), .rectangle2_weight(rectangle2_weights[229]), .rectangle3_x(rectangle3_xs[229]), .rectangle3_y(rectangle3_ys[229]), .rectangle3_width(rectangle3_widths[229]), .rectangle3_height(rectangle3_heights[229]), .rectangle3_weight(rectangle3_weights[229]), .feature_threshold(feature_thresholds[229]), .feature_above(feature_aboves[229]), .feature_below(feature_belows[229]), .scan_win_std_dev(scan_win_std_dev[229]), .feature_accum(feature_accums[229]));
  accum_calculator ac230(.scan_win(scan_win230), .rectangle1_x(rectangle1_xs[230]), .rectangle1_y(rectangle1_ys[230]), .rectangle1_width(rectangle1_widths[230]), .rectangle1_height(rectangle1_heights[230]), .rectangle1_weight(rectangle1_weights[230]), .rectangle2_x(rectangle2_xs[230]), .rectangle2_y(rectangle2_ys[230]), .rectangle2_width(rectangle2_widths[230]), .rectangle2_height(rectangle2_heights[230]), .rectangle2_weight(rectangle2_weights[230]), .rectangle3_x(rectangle3_xs[230]), .rectangle3_y(rectangle3_ys[230]), .rectangle3_width(rectangle3_widths[230]), .rectangle3_height(rectangle3_heights[230]), .rectangle3_weight(rectangle3_weights[230]), .feature_threshold(feature_thresholds[230]), .feature_above(feature_aboves[230]), .feature_below(feature_belows[230]), .scan_win_std_dev(scan_win_std_dev[230]), .feature_accum(feature_accums[230]));
  accum_calculator ac231(.scan_win(scan_win231), .rectangle1_x(rectangle1_xs[231]), .rectangle1_y(rectangle1_ys[231]), .rectangle1_width(rectangle1_widths[231]), .rectangle1_height(rectangle1_heights[231]), .rectangle1_weight(rectangle1_weights[231]), .rectangle2_x(rectangle2_xs[231]), .rectangle2_y(rectangle2_ys[231]), .rectangle2_width(rectangle2_widths[231]), .rectangle2_height(rectangle2_heights[231]), .rectangle2_weight(rectangle2_weights[231]), .rectangle3_x(rectangle3_xs[231]), .rectangle3_y(rectangle3_ys[231]), .rectangle3_width(rectangle3_widths[231]), .rectangle3_height(rectangle3_heights[231]), .rectangle3_weight(rectangle3_weights[231]), .feature_threshold(feature_thresholds[231]), .feature_above(feature_aboves[231]), .feature_below(feature_belows[231]), .scan_win_std_dev(scan_win_std_dev[231]), .feature_accum(feature_accums[231]));
  accum_calculator ac232(.scan_win(scan_win232), .rectangle1_x(rectangle1_xs[232]), .rectangle1_y(rectangle1_ys[232]), .rectangle1_width(rectangle1_widths[232]), .rectangle1_height(rectangle1_heights[232]), .rectangle1_weight(rectangle1_weights[232]), .rectangle2_x(rectangle2_xs[232]), .rectangle2_y(rectangle2_ys[232]), .rectangle2_width(rectangle2_widths[232]), .rectangle2_height(rectangle2_heights[232]), .rectangle2_weight(rectangle2_weights[232]), .rectangle3_x(rectangle3_xs[232]), .rectangle3_y(rectangle3_ys[232]), .rectangle3_width(rectangle3_widths[232]), .rectangle3_height(rectangle3_heights[232]), .rectangle3_weight(rectangle3_weights[232]), .feature_threshold(feature_thresholds[232]), .feature_above(feature_aboves[232]), .feature_below(feature_belows[232]), .scan_win_std_dev(scan_win_std_dev[232]), .feature_accum(feature_accums[232]));
  accum_calculator ac233(.scan_win(scan_win233), .rectangle1_x(rectangle1_xs[233]), .rectangle1_y(rectangle1_ys[233]), .rectangle1_width(rectangle1_widths[233]), .rectangle1_height(rectangle1_heights[233]), .rectangle1_weight(rectangle1_weights[233]), .rectangle2_x(rectangle2_xs[233]), .rectangle2_y(rectangle2_ys[233]), .rectangle2_width(rectangle2_widths[233]), .rectangle2_height(rectangle2_heights[233]), .rectangle2_weight(rectangle2_weights[233]), .rectangle3_x(rectangle3_xs[233]), .rectangle3_y(rectangle3_ys[233]), .rectangle3_width(rectangle3_widths[233]), .rectangle3_height(rectangle3_heights[233]), .rectangle3_weight(rectangle3_weights[233]), .feature_threshold(feature_thresholds[233]), .feature_above(feature_aboves[233]), .feature_below(feature_belows[233]), .scan_win_std_dev(scan_win_std_dev[233]), .feature_accum(feature_accums[233]));
  accum_calculator ac234(.scan_win(scan_win234), .rectangle1_x(rectangle1_xs[234]), .rectangle1_y(rectangle1_ys[234]), .rectangle1_width(rectangle1_widths[234]), .rectangle1_height(rectangle1_heights[234]), .rectangle1_weight(rectangle1_weights[234]), .rectangle2_x(rectangle2_xs[234]), .rectangle2_y(rectangle2_ys[234]), .rectangle2_width(rectangle2_widths[234]), .rectangle2_height(rectangle2_heights[234]), .rectangle2_weight(rectangle2_weights[234]), .rectangle3_x(rectangle3_xs[234]), .rectangle3_y(rectangle3_ys[234]), .rectangle3_width(rectangle3_widths[234]), .rectangle3_height(rectangle3_heights[234]), .rectangle3_weight(rectangle3_weights[234]), .feature_threshold(feature_thresholds[234]), .feature_above(feature_aboves[234]), .feature_below(feature_belows[234]), .scan_win_std_dev(scan_win_std_dev[234]), .feature_accum(feature_accums[234]));
  accum_calculator ac235(.scan_win(scan_win235), .rectangle1_x(rectangle1_xs[235]), .rectangle1_y(rectangle1_ys[235]), .rectangle1_width(rectangle1_widths[235]), .rectangle1_height(rectangle1_heights[235]), .rectangle1_weight(rectangle1_weights[235]), .rectangle2_x(rectangle2_xs[235]), .rectangle2_y(rectangle2_ys[235]), .rectangle2_width(rectangle2_widths[235]), .rectangle2_height(rectangle2_heights[235]), .rectangle2_weight(rectangle2_weights[235]), .rectangle3_x(rectangle3_xs[235]), .rectangle3_y(rectangle3_ys[235]), .rectangle3_width(rectangle3_widths[235]), .rectangle3_height(rectangle3_heights[235]), .rectangle3_weight(rectangle3_weights[235]), .feature_threshold(feature_thresholds[235]), .feature_above(feature_aboves[235]), .feature_below(feature_belows[235]), .scan_win_std_dev(scan_win_std_dev[235]), .feature_accum(feature_accums[235]));
  accum_calculator ac236(.scan_win(scan_win236), .rectangle1_x(rectangle1_xs[236]), .rectangle1_y(rectangle1_ys[236]), .rectangle1_width(rectangle1_widths[236]), .rectangle1_height(rectangle1_heights[236]), .rectangle1_weight(rectangle1_weights[236]), .rectangle2_x(rectangle2_xs[236]), .rectangle2_y(rectangle2_ys[236]), .rectangle2_width(rectangle2_widths[236]), .rectangle2_height(rectangle2_heights[236]), .rectangle2_weight(rectangle2_weights[236]), .rectangle3_x(rectangle3_xs[236]), .rectangle3_y(rectangle3_ys[236]), .rectangle3_width(rectangle3_widths[236]), .rectangle3_height(rectangle3_heights[236]), .rectangle3_weight(rectangle3_weights[236]), .feature_threshold(feature_thresholds[236]), .feature_above(feature_aboves[236]), .feature_below(feature_belows[236]), .scan_win_std_dev(scan_win_std_dev[236]), .feature_accum(feature_accums[236]));
  accum_calculator ac237(.scan_win(scan_win237), .rectangle1_x(rectangle1_xs[237]), .rectangle1_y(rectangle1_ys[237]), .rectangle1_width(rectangle1_widths[237]), .rectangle1_height(rectangle1_heights[237]), .rectangle1_weight(rectangle1_weights[237]), .rectangle2_x(rectangle2_xs[237]), .rectangle2_y(rectangle2_ys[237]), .rectangle2_width(rectangle2_widths[237]), .rectangle2_height(rectangle2_heights[237]), .rectangle2_weight(rectangle2_weights[237]), .rectangle3_x(rectangle3_xs[237]), .rectangle3_y(rectangle3_ys[237]), .rectangle3_width(rectangle3_widths[237]), .rectangle3_height(rectangle3_heights[237]), .rectangle3_weight(rectangle3_weights[237]), .feature_threshold(feature_thresholds[237]), .feature_above(feature_aboves[237]), .feature_below(feature_belows[237]), .scan_win_std_dev(scan_win_std_dev[237]), .feature_accum(feature_accums[237]));
  accum_calculator ac238(.scan_win(scan_win238), .rectangle1_x(rectangle1_xs[238]), .rectangle1_y(rectangle1_ys[238]), .rectangle1_width(rectangle1_widths[238]), .rectangle1_height(rectangle1_heights[238]), .rectangle1_weight(rectangle1_weights[238]), .rectangle2_x(rectangle2_xs[238]), .rectangle2_y(rectangle2_ys[238]), .rectangle2_width(rectangle2_widths[238]), .rectangle2_height(rectangle2_heights[238]), .rectangle2_weight(rectangle2_weights[238]), .rectangle3_x(rectangle3_xs[238]), .rectangle3_y(rectangle3_ys[238]), .rectangle3_width(rectangle3_widths[238]), .rectangle3_height(rectangle3_heights[238]), .rectangle3_weight(rectangle3_weights[238]), .feature_threshold(feature_thresholds[238]), .feature_above(feature_aboves[238]), .feature_below(feature_belows[238]), .scan_win_std_dev(scan_win_std_dev[238]), .feature_accum(feature_accums[238]));
  accum_calculator ac239(.scan_win(scan_win239), .rectangle1_x(rectangle1_xs[239]), .rectangle1_y(rectangle1_ys[239]), .rectangle1_width(rectangle1_widths[239]), .rectangle1_height(rectangle1_heights[239]), .rectangle1_weight(rectangle1_weights[239]), .rectangle2_x(rectangle2_xs[239]), .rectangle2_y(rectangle2_ys[239]), .rectangle2_width(rectangle2_widths[239]), .rectangle2_height(rectangle2_heights[239]), .rectangle2_weight(rectangle2_weights[239]), .rectangle3_x(rectangle3_xs[239]), .rectangle3_y(rectangle3_ys[239]), .rectangle3_width(rectangle3_widths[239]), .rectangle3_height(rectangle3_heights[239]), .rectangle3_weight(rectangle3_weights[239]), .feature_threshold(feature_thresholds[239]), .feature_above(feature_aboves[239]), .feature_below(feature_belows[239]), .scan_win_std_dev(scan_win_std_dev[239]), .feature_accum(feature_accums[239]));
  accum_calculator ac240(.scan_win(scan_win240), .rectangle1_x(rectangle1_xs[240]), .rectangle1_y(rectangle1_ys[240]), .rectangle1_width(rectangle1_widths[240]), .rectangle1_height(rectangle1_heights[240]), .rectangle1_weight(rectangle1_weights[240]), .rectangle2_x(rectangle2_xs[240]), .rectangle2_y(rectangle2_ys[240]), .rectangle2_width(rectangle2_widths[240]), .rectangle2_height(rectangle2_heights[240]), .rectangle2_weight(rectangle2_weights[240]), .rectangle3_x(rectangle3_xs[240]), .rectangle3_y(rectangle3_ys[240]), .rectangle3_width(rectangle3_widths[240]), .rectangle3_height(rectangle3_heights[240]), .rectangle3_weight(rectangle3_weights[240]), .feature_threshold(feature_thresholds[240]), .feature_above(feature_aboves[240]), .feature_below(feature_belows[240]), .scan_win_std_dev(scan_win_std_dev[240]), .feature_accum(feature_accums[240]));
  accum_calculator ac241(.scan_win(scan_win241), .rectangle1_x(rectangle1_xs[241]), .rectangle1_y(rectangle1_ys[241]), .rectangle1_width(rectangle1_widths[241]), .rectangle1_height(rectangle1_heights[241]), .rectangle1_weight(rectangle1_weights[241]), .rectangle2_x(rectangle2_xs[241]), .rectangle2_y(rectangle2_ys[241]), .rectangle2_width(rectangle2_widths[241]), .rectangle2_height(rectangle2_heights[241]), .rectangle2_weight(rectangle2_weights[241]), .rectangle3_x(rectangle3_xs[241]), .rectangle3_y(rectangle3_ys[241]), .rectangle3_width(rectangle3_widths[241]), .rectangle3_height(rectangle3_heights[241]), .rectangle3_weight(rectangle3_weights[241]), .feature_threshold(feature_thresholds[241]), .feature_above(feature_aboves[241]), .feature_below(feature_belows[241]), .scan_win_std_dev(scan_win_std_dev[241]), .feature_accum(feature_accums[241]));
  accum_calculator ac242(.scan_win(scan_win242), .rectangle1_x(rectangle1_xs[242]), .rectangle1_y(rectangle1_ys[242]), .rectangle1_width(rectangle1_widths[242]), .rectangle1_height(rectangle1_heights[242]), .rectangle1_weight(rectangle1_weights[242]), .rectangle2_x(rectangle2_xs[242]), .rectangle2_y(rectangle2_ys[242]), .rectangle2_width(rectangle2_widths[242]), .rectangle2_height(rectangle2_heights[242]), .rectangle2_weight(rectangle2_weights[242]), .rectangle3_x(rectangle3_xs[242]), .rectangle3_y(rectangle3_ys[242]), .rectangle3_width(rectangle3_widths[242]), .rectangle3_height(rectangle3_heights[242]), .rectangle3_weight(rectangle3_weights[242]), .feature_threshold(feature_thresholds[242]), .feature_above(feature_aboves[242]), .feature_below(feature_belows[242]), .scan_win_std_dev(scan_win_std_dev[242]), .feature_accum(feature_accums[242]));
  accum_calculator ac243(.scan_win(scan_win243), .rectangle1_x(rectangle1_xs[243]), .rectangle1_y(rectangle1_ys[243]), .rectangle1_width(rectangle1_widths[243]), .rectangle1_height(rectangle1_heights[243]), .rectangle1_weight(rectangle1_weights[243]), .rectangle2_x(rectangle2_xs[243]), .rectangle2_y(rectangle2_ys[243]), .rectangle2_width(rectangle2_widths[243]), .rectangle2_height(rectangle2_heights[243]), .rectangle2_weight(rectangle2_weights[243]), .rectangle3_x(rectangle3_xs[243]), .rectangle3_y(rectangle3_ys[243]), .rectangle3_width(rectangle3_widths[243]), .rectangle3_height(rectangle3_heights[243]), .rectangle3_weight(rectangle3_weights[243]), .feature_threshold(feature_thresholds[243]), .feature_above(feature_aboves[243]), .feature_below(feature_belows[243]), .scan_win_std_dev(scan_win_std_dev[243]), .feature_accum(feature_accums[243]));
  accum_calculator ac244(.scan_win(scan_win244), .rectangle1_x(rectangle1_xs[244]), .rectangle1_y(rectangle1_ys[244]), .rectangle1_width(rectangle1_widths[244]), .rectangle1_height(rectangle1_heights[244]), .rectangle1_weight(rectangle1_weights[244]), .rectangle2_x(rectangle2_xs[244]), .rectangle2_y(rectangle2_ys[244]), .rectangle2_width(rectangle2_widths[244]), .rectangle2_height(rectangle2_heights[244]), .rectangle2_weight(rectangle2_weights[244]), .rectangle3_x(rectangle3_xs[244]), .rectangle3_y(rectangle3_ys[244]), .rectangle3_width(rectangle3_widths[244]), .rectangle3_height(rectangle3_heights[244]), .rectangle3_weight(rectangle3_weights[244]), .feature_threshold(feature_thresholds[244]), .feature_above(feature_aboves[244]), .feature_below(feature_belows[244]), .scan_win_std_dev(scan_win_std_dev[244]), .feature_accum(feature_accums[244]));
  accum_calculator ac245(.scan_win(scan_win245), .rectangle1_x(rectangle1_xs[245]), .rectangle1_y(rectangle1_ys[245]), .rectangle1_width(rectangle1_widths[245]), .rectangle1_height(rectangle1_heights[245]), .rectangle1_weight(rectangle1_weights[245]), .rectangle2_x(rectangle2_xs[245]), .rectangle2_y(rectangle2_ys[245]), .rectangle2_width(rectangle2_widths[245]), .rectangle2_height(rectangle2_heights[245]), .rectangle2_weight(rectangle2_weights[245]), .rectangle3_x(rectangle3_xs[245]), .rectangle3_y(rectangle3_ys[245]), .rectangle3_width(rectangle3_widths[245]), .rectangle3_height(rectangle3_heights[245]), .rectangle3_weight(rectangle3_weights[245]), .feature_threshold(feature_thresholds[245]), .feature_above(feature_aboves[245]), .feature_below(feature_belows[245]), .scan_win_std_dev(scan_win_std_dev[245]), .feature_accum(feature_accums[245]));
  accum_calculator ac246(.scan_win(scan_win246), .rectangle1_x(rectangle1_xs[246]), .rectangle1_y(rectangle1_ys[246]), .rectangle1_width(rectangle1_widths[246]), .rectangle1_height(rectangle1_heights[246]), .rectangle1_weight(rectangle1_weights[246]), .rectangle2_x(rectangle2_xs[246]), .rectangle2_y(rectangle2_ys[246]), .rectangle2_width(rectangle2_widths[246]), .rectangle2_height(rectangle2_heights[246]), .rectangle2_weight(rectangle2_weights[246]), .rectangle3_x(rectangle3_xs[246]), .rectangle3_y(rectangle3_ys[246]), .rectangle3_width(rectangle3_widths[246]), .rectangle3_height(rectangle3_heights[246]), .rectangle3_weight(rectangle3_weights[246]), .feature_threshold(feature_thresholds[246]), .feature_above(feature_aboves[246]), .feature_below(feature_belows[246]), .scan_win_std_dev(scan_win_std_dev[246]), .feature_accum(feature_accums[246]));
  accum_calculator ac247(.scan_win(scan_win247), .rectangle1_x(rectangle1_xs[247]), .rectangle1_y(rectangle1_ys[247]), .rectangle1_width(rectangle1_widths[247]), .rectangle1_height(rectangle1_heights[247]), .rectangle1_weight(rectangle1_weights[247]), .rectangle2_x(rectangle2_xs[247]), .rectangle2_y(rectangle2_ys[247]), .rectangle2_width(rectangle2_widths[247]), .rectangle2_height(rectangle2_heights[247]), .rectangle2_weight(rectangle2_weights[247]), .rectangle3_x(rectangle3_xs[247]), .rectangle3_y(rectangle3_ys[247]), .rectangle3_width(rectangle3_widths[247]), .rectangle3_height(rectangle3_heights[247]), .rectangle3_weight(rectangle3_weights[247]), .feature_threshold(feature_thresholds[247]), .feature_above(feature_aboves[247]), .feature_below(feature_belows[247]), .scan_win_std_dev(scan_win_std_dev[247]), .feature_accum(feature_accums[247]));
  accum_calculator ac248(.scan_win(scan_win248), .rectangle1_x(rectangle1_xs[248]), .rectangle1_y(rectangle1_ys[248]), .rectangle1_width(rectangle1_widths[248]), .rectangle1_height(rectangle1_heights[248]), .rectangle1_weight(rectangle1_weights[248]), .rectangle2_x(rectangle2_xs[248]), .rectangle2_y(rectangle2_ys[248]), .rectangle2_width(rectangle2_widths[248]), .rectangle2_height(rectangle2_heights[248]), .rectangle2_weight(rectangle2_weights[248]), .rectangle3_x(rectangle3_xs[248]), .rectangle3_y(rectangle3_ys[248]), .rectangle3_width(rectangle3_widths[248]), .rectangle3_height(rectangle3_heights[248]), .rectangle3_weight(rectangle3_weights[248]), .feature_threshold(feature_thresholds[248]), .feature_above(feature_aboves[248]), .feature_below(feature_belows[248]), .scan_win_std_dev(scan_win_std_dev[248]), .feature_accum(feature_accums[248]));
  accum_calculator ac249(.scan_win(scan_win249), .rectangle1_x(rectangle1_xs[249]), .rectangle1_y(rectangle1_ys[249]), .rectangle1_width(rectangle1_widths[249]), .rectangle1_height(rectangle1_heights[249]), .rectangle1_weight(rectangle1_weights[249]), .rectangle2_x(rectangle2_xs[249]), .rectangle2_y(rectangle2_ys[249]), .rectangle2_width(rectangle2_widths[249]), .rectangle2_height(rectangle2_heights[249]), .rectangle2_weight(rectangle2_weights[249]), .rectangle3_x(rectangle3_xs[249]), .rectangle3_y(rectangle3_ys[249]), .rectangle3_width(rectangle3_widths[249]), .rectangle3_height(rectangle3_heights[249]), .rectangle3_weight(rectangle3_weights[249]), .feature_threshold(feature_thresholds[249]), .feature_above(feature_aboves[249]), .feature_below(feature_belows[249]), .scan_win_std_dev(scan_win_std_dev[249]), .feature_accum(feature_accums[249]));
  accum_calculator ac250(.scan_win(scan_win250), .rectangle1_x(rectangle1_xs[250]), .rectangle1_y(rectangle1_ys[250]), .rectangle1_width(rectangle1_widths[250]), .rectangle1_height(rectangle1_heights[250]), .rectangle1_weight(rectangle1_weights[250]), .rectangle2_x(rectangle2_xs[250]), .rectangle2_y(rectangle2_ys[250]), .rectangle2_width(rectangle2_widths[250]), .rectangle2_height(rectangle2_heights[250]), .rectangle2_weight(rectangle2_weights[250]), .rectangle3_x(rectangle3_xs[250]), .rectangle3_y(rectangle3_ys[250]), .rectangle3_width(rectangle3_widths[250]), .rectangle3_height(rectangle3_heights[250]), .rectangle3_weight(rectangle3_weights[250]), .feature_threshold(feature_thresholds[250]), .feature_above(feature_aboves[250]), .feature_below(feature_belows[250]), .scan_win_std_dev(scan_win_std_dev[250]), .feature_accum(feature_accums[250]));
  accum_calculator ac251(.scan_win(scan_win251), .rectangle1_x(rectangle1_xs[251]), .rectangle1_y(rectangle1_ys[251]), .rectangle1_width(rectangle1_widths[251]), .rectangle1_height(rectangle1_heights[251]), .rectangle1_weight(rectangle1_weights[251]), .rectangle2_x(rectangle2_xs[251]), .rectangle2_y(rectangle2_ys[251]), .rectangle2_width(rectangle2_widths[251]), .rectangle2_height(rectangle2_heights[251]), .rectangle2_weight(rectangle2_weights[251]), .rectangle3_x(rectangle3_xs[251]), .rectangle3_y(rectangle3_ys[251]), .rectangle3_width(rectangle3_widths[251]), .rectangle3_height(rectangle3_heights[251]), .rectangle3_weight(rectangle3_weights[251]), .feature_threshold(feature_thresholds[251]), .feature_above(feature_aboves[251]), .feature_below(feature_belows[251]), .scan_win_std_dev(scan_win_std_dev[251]), .feature_accum(feature_accums[251]));
  accum_calculator ac252(.scan_win(scan_win252), .rectangle1_x(rectangle1_xs[252]), .rectangle1_y(rectangle1_ys[252]), .rectangle1_width(rectangle1_widths[252]), .rectangle1_height(rectangle1_heights[252]), .rectangle1_weight(rectangle1_weights[252]), .rectangle2_x(rectangle2_xs[252]), .rectangle2_y(rectangle2_ys[252]), .rectangle2_width(rectangle2_widths[252]), .rectangle2_height(rectangle2_heights[252]), .rectangle2_weight(rectangle2_weights[252]), .rectangle3_x(rectangle3_xs[252]), .rectangle3_y(rectangle3_ys[252]), .rectangle3_width(rectangle3_widths[252]), .rectangle3_height(rectangle3_heights[252]), .rectangle3_weight(rectangle3_weights[252]), .feature_threshold(feature_thresholds[252]), .feature_above(feature_aboves[252]), .feature_below(feature_belows[252]), .scan_win_std_dev(scan_win_std_dev[252]), .feature_accum(feature_accums[252]));
  accum_calculator ac253(.scan_win(scan_win253), .rectangle1_x(rectangle1_xs[253]), .rectangle1_y(rectangle1_ys[253]), .rectangle1_width(rectangle1_widths[253]), .rectangle1_height(rectangle1_heights[253]), .rectangle1_weight(rectangle1_weights[253]), .rectangle2_x(rectangle2_xs[253]), .rectangle2_y(rectangle2_ys[253]), .rectangle2_width(rectangle2_widths[253]), .rectangle2_height(rectangle2_heights[253]), .rectangle2_weight(rectangle2_weights[253]), .rectangle3_x(rectangle3_xs[253]), .rectangle3_y(rectangle3_ys[253]), .rectangle3_width(rectangle3_widths[253]), .rectangle3_height(rectangle3_heights[253]), .rectangle3_weight(rectangle3_weights[253]), .feature_threshold(feature_thresholds[253]), .feature_above(feature_aboves[253]), .feature_below(feature_belows[253]), .scan_win_std_dev(scan_win_std_dev[253]), .feature_accum(feature_accums[253]));
  accum_calculator ac254(.scan_win(scan_win254), .rectangle1_x(rectangle1_xs[254]), .rectangle1_y(rectangle1_ys[254]), .rectangle1_width(rectangle1_widths[254]), .rectangle1_height(rectangle1_heights[254]), .rectangle1_weight(rectangle1_weights[254]), .rectangle2_x(rectangle2_xs[254]), .rectangle2_y(rectangle2_ys[254]), .rectangle2_width(rectangle2_widths[254]), .rectangle2_height(rectangle2_heights[254]), .rectangle2_weight(rectangle2_weights[254]), .rectangle3_x(rectangle3_xs[254]), .rectangle3_y(rectangle3_ys[254]), .rectangle3_width(rectangle3_widths[254]), .rectangle3_height(rectangle3_heights[254]), .rectangle3_weight(rectangle3_weights[254]), .feature_threshold(feature_thresholds[254]), .feature_above(feature_aboves[254]), .feature_below(feature_belows[254]), .scan_win_std_dev(scan_win_std_dev[254]), .feature_accum(feature_accums[254]));
  accum_calculator ac255(.scan_win(scan_win255), .rectangle1_x(rectangle1_xs[255]), .rectangle1_y(rectangle1_ys[255]), .rectangle1_width(rectangle1_widths[255]), .rectangle1_height(rectangle1_heights[255]), .rectangle1_weight(rectangle1_weights[255]), .rectangle2_x(rectangle2_xs[255]), .rectangle2_y(rectangle2_ys[255]), .rectangle2_width(rectangle2_widths[255]), .rectangle2_height(rectangle2_heights[255]), .rectangle2_weight(rectangle2_weights[255]), .rectangle3_x(rectangle3_xs[255]), .rectangle3_y(rectangle3_ys[255]), .rectangle3_width(rectangle3_widths[255]), .rectangle3_height(rectangle3_heights[255]), .rectangle3_weight(rectangle3_weights[255]), .feature_threshold(feature_thresholds[255]), .feature_above(feature_aboves[255]), .feature_below(feature_belows[255]), .scan_win_std_dev(scan_win_std_dev[255]), .feature_accum(feature_accums[255]));
  accum_calculator ac256(.scan_win(scan_win256), .rectangle1_x(rectangle1_xs[256]), .rectangle1_y(rectangle1_ys[256]), .rectangle1_width(rectangle1_widths[256]), .rectangle1_height(rectangle1_heights[256]), .rectangle1_weight(rectangle1_weights[256]), .rectangle2_x(rectangle2_xs[256]), .rectangle2_y(rectangle2_ys[256]), .rectangle2_width(rectangle2_widths[256]), .rectangle2_height(rectangle2_heights[256]), .rectangle2_weight(rectangle2_weights[256]), .rectangle3_x(rectangle3_xs[256]), .rectangle3_y(rectangle3_ys[256]), .rectangle3_width(rectangle3_widths[256]), .rectangle3_height(rectangle3_heights[256]), .rectangle3_weight(rectangle3_weights[256]), .feature_threshold(feature_thresholds[256]), .feature_above(feature_aboves[256]), .feature_below(feature_belows[256]), .scan_win_std_dev(scan_win_std_dev[256]), .feature_accum(feature_accums[256]));
  accum_calculator ac257(.scan_win(scan_win257), .rectangle1_x(rectangle1_xs[257]), .rectangle1_y(rectangle1_ys[257]), .rectangle1_width(rectangle1_widths[257]), .rectangle1_height(rectangle1_heights[257]), .rectangle1_weight(rectangle1_weights[257]), .rectangle2_x(rectangle2_xs[257]), .rectangle2_y(rectangle2_ys[257]), .rectangle2_width(rectangle2_widths[257]), .rectangle2_height(rectangle2_heights[257]), .rectangle2_weight(rectangle2_weights[257]), .rectangle3_x(rectangle3_xs[257]), .rectangle3_y(rectangle3_ys[257]), .rectangle3_width(rectangle3_widths[257]), .rectangle3_height(rectangle3_heights[257]), .rectangle3_weight(rectangle3_weights[257]), .feature_threshold(feature_thresholds[257]), .feature_above(feature_aboves[257]), .feature_below(feature_belows[257]), .scan_win_std_dev(scan_win_std_dev[257]), .feature_accum(feature_accums[257]));
  accum_calculator ac258(.scan_win(scan_win258), .rectangle1_x(rectangle1_xs[258]), .rectangle1_y(rectangle1_ys[258]), .rectangle1_width(rectangle1_widths[258]), .rectangle1_height(rectangle1_heights[258]), .rectangle1_weight(rectangle1_weights[258]), .rectangle2_x(rectangle2_xs[258]), .rectangle2_y(rectangle2_ys[258]), .rectangle2_width(rectangle2_widths[258]), .rectangle2_height(rectangle2_heights[258]), .rectangle2_weight(rectangle2_weights[258]), .rectangle3_x(rectangle3_xs[258]), .rectangle3_y(rectangle3_ys[258]), .rectangle3_width(rectangle3_widths[258]), .rectangle3_height(rectangle3_heights[258]), .rectangle3_weight(rectangle3_weights[258]), .feature_threshold(feature_thresholds[258]), .feature_above(feature_aboves[258]), .feature_below(feature_belows[258]), .scan_win_std_dev(scan_win_std_dev[258]), .feature_accum(feature_accums[258]));
  accum_calculator ac259(.scan_win(scan_win259), .rectangle1_x(rectangle1_xs[259]), .rectangle1_y(rectangle1_ys[259]), .rectangle1_width(rectangle1_widths[259]), .rectangle1_height(rectangle1_heights[259]), .rectangle1_weight(rectangle1_weights[259]), .rectangle2_x(rectangle2_xs[259]), .rectangle2_y(rectangle2_ys[259]), .rectangle2_width(rectangle2_widths[259]), .rectangle2_height(rectangle2_heights[259]), .rectangle2_weight(rectangle2_weights[259]), .rectangle3_x(rectangle3_xs[259]), .rectangle3_y(rectangle3_ys[259]), .rectangle3_width(rectangle3_widths[259]), .rectangle3_height(rectangle3_heights[259]), .rectangle3_weight(rectangle3_weights[259]), .feature_threshold(feature_thresholds[259]), .feature_above(feature_aboves[259]), .feature_below(feature_belows[259]), .scan_win_std_dev(scan_win_std_dev[259]), .feature_accum(feature_accums[259]));
  accum_calculator ac260(.scan_win(scan_win260), .rectangle1_x(rectangle1_xs[260]), .rectangle1_y(rectangle1_ys[260]), .rectangle1_width(rectangle1_widths[260]), .rectangle1_height(rectangle1_heights[260]), .rectangle1_weight(rectangle1_weights[260]), .rectangle2_x(rectangle2_xs[260]), .rectangle2_y(rectangle2_ys[260]), .rectangle2_width(rectangle2_widths[260]), .rectangle2_height(rectangle2_heights[260]), .rectangle2_weight(rectangle2_weights[260]), .rectangle3_x(rectangle3_xs[260]), .rectangle3_y(rectangle3_ys[260]), .rectangle3_width(rectangle3_widths[260]), .rectangle3_height(rectangle3_heights[260]), .rectangle3_weight(rectangle3_weights[260]), .feature_threshold(feature_thresholds[260]), .feature_above(feature_aboves[260]), .feature_below(feature_belows[260]), .scan_win_std_dev(scan_win_std_dev[260]), .feature_accum(feature_accums[260]));
  accum_calculator ac261(.scan_win(scan_win261), .rectangle1_x(rectangle1_xs[261]), .rectangle1_y(rectangle1_ys[261]), .rectangle1_width(rectangle1_widths[261]), .rectangle1_height(rectangle1_heights[261]), .rectangle1_weight(rectangle1_weights[261]), .rectangle2_x(rectangle2_xs[261]), .rectangle2_y(rectangle2_ys[261]), .rectangle2_width(rectangle2_widths[261]), .rectangle2_height(rectangle2_heights[261]), .rectangle2_weight(rectangle2_weights[261]), .rectangle3_x(rectangle3_xs[261]), .rectangle3_y(rectangle3_ys[261]), .rectangle3_width(rectangle3_widths[261]), .rectangle3_height(rectangle3_heights[261]), .rectangle3_weight(rectangle3_weights[261]), .feature_threshold(feature_thresholds[261]), .feature_above(feature_aboves[261]), .feature_below(feature_belows[261]), .scan_win_std_dev(scan_win_std_dev[261]), .feature_accum(feature_accums[261]));
  accum_calculator ac262(.scan_win(scan_win262), .rectangle1_x(rectangle1_xs[262]), .rectangle1_y(rectangle1_ys[262]), .rectangle1_width(rectangle1_widths[262]), .rectangle1_height(rectangle1_heights[262]), .rectangle1_weight(rectangle1_weights[262]), .rectangle2_x(rectangle2_xs[262]), .rectangle2_y(rectangle2_ys[262]), .rectangle2_width(rectangle2_widths[262]), .rectangle2_height(rectangle2_heights[262]), .rectangle2_weight(rectangle2_weights[262]), .rectangle3_x(rectangle3_xs[262]), .rectangle3_y(rectangle3_ys[262]), .rectangle3_width(rectangle3_widths[262]), .rectangle3_height(rectangle3_heights[262]), .rectangle3_weight(rectangle3_weights[262]), .feature_threshold(feature_thresholds[262]), .feature_above(feature_aboves[262]), .feature_below(feature_belows[262]), .scan_win_std_dev(scan_win_std_dev[262]), .feature_accum(feature_accums[262]));
  accum_calculator ac263(.scan_win(scan_win263), .rectangle1_x(rectangle1_xs[263]), .rectangle1_y(rectangle1_ys[263]), .rectangle1_width(rectangle1_widths[263]), .rectangle1_height(rectangle1_heights[263]), .rectangle1_weight(rectangle1_weights[263]), .rectangle2_x(rectangle2_xs[263]), .rectangle2_y(rectangle2_ys[263]), .rectangle2_width(rectangle2_widths[263]), .rectangle2_height(rectangle2_heights[263]), .rectangle2_weight(rectangle2_weights[263]), .rectangle3_x(rectangle3_xs[263]), .rectangle3_y(rectangle3_ys[263]), .rectangle3_width(rectangle3_widths[263]), .rectangle3_height(rectangle3_heights[263]), .rectangle3_weight(rectangle3_weights[263]), .feature_threshold(feature_thresholds[263]), .feature_above(feature_aboves[263]), .feature_below(feature_belows[263]), .scan_win_std_dev(scan_win_std_dev[263]), .feature_accum(feature_accums[263]));
  accum_calculator ac264(.scan_win(scan_win264), .rectangle1_x(rectangle1_xs[264]), .rectangle1_y(rectangle1_ys[264]), .rectangle1_width(rectangle1_widths[264]), .rectangle1_height(rectangle1_heights[264]), .rectangle1_weight(rectangle1_weights[264]), .rectangle2_x(rectangle2_xs[264]), .rectangle2_y(rectangle2_ys[264]), .rectangle2_width(rectangle2_widths[264]), .rectangle2_height(rectangle2_heights[264]), .rectangle2_weight(rectangle2_weights[264]), .rectangle3_x(rectangle3_xs[264]), .rectangle3_y(rectangle3_ys[264]), .rectangle3_width(rectangle3_widths[264]), .rectangle3_height(rectangle3_heights[264]), .rectangle3_weight(rectangle3_weights[264]), .feature_threshold(feature_thresholds[264]), .feature_above(feature_aboves[264]), .feature_below(feature_belows[264]), .scan_win_std_dev(scan_win_std_dev[264]), .feature_accum(feature_accums[264]));
  accum_calculator ac265(.scan_win(scan_win265), .rectangle1_x(rectangle1_xs[265]), .rectangle1_y(rectangle1_ys[265]), .rectangle1_width(rectangle1_widths[265]), .rectangle1_height(rectangle1_heights[265]), .rectangle1_weight(rectangle1_weights[265]), .rectangle2_x(rectangle2_xs[265]), .rectangle2_y(rectangle2_ys[265]), .rectangle2_width(rectangle2_widths[265]), .rectangle2_height(rectangle2_heights[265]), .rectangle2_weight(rectangle2_weights[265]), .rectangle3_x(rectangle3_xs[265]), .rectangle3_y(rectangle3_ys[265]), .rectangle3_width(rectangle3_widths[265]), .rectangle3_height(rectangle3_heights[265]), .rectangle3_weight(rectangle3_weights[265]), .feature_threshold(feature_thresholds[265]), .feature_above(feature_aboves[265]), .feature_below(feature_belows[265]), .scan_win_std_dev(scan_win_std_dev[265]), .feature_accum(feature_accums[265]));
  accum_calculator ac266(.scan_win(scan_win266), .rectangle1_x(rectangle1_xs[266]), .rectangle1_y(rectangle1_ys[266]), .rectangle1_width(rectangle1_widths[266]), .rectangle1_height(rectangle1_heights[266]), .rectangle1_weight(rectangle1_weights[266]), .rectangle2_x(rectangle2_xs[266]), .rectangle2_y(rectangle2_ys[266]), .rectangle2_width(rectangle2_widths[266]), .rectangle2_height(rectangle2_heights[266]), .rectangle2_weight(rectangle2_weights[266]), .rectangle3_x(rectangle3_xs[266]), .rectangle3_y(rectangle3_ys[266]), .rectangle3_width(rectangle3_widths[266]), .rectangle3_height(rectangle3_heights[266]), .rectangle3_weight(rectangle3_weights[266]), .feature_threshold(feature_thresholds[266]), .feature_above(feature_aboves[266]), .feature_below(feature_belows[266]), .scan_win_std_dev(scan_win_std_dev[266]), .feature_accum(feature_accums[266]));
  accum_calculator ac267(.scan_win(scan_win267), .rectangle1_x(rectangle1_xs[267]), .rectangle1_y(rectangle1_ys[267]), .rectangle1_width(rectangle1_widths[267]), .rectangle1_height(rectangle1_heights[267]), .rectangle1_weight(rectangle1_weights[267]), .rectangle2_x(rectangle2_xs[267]), .rectangle2_y(rectangle2_ys[267]), .rectangle2_width(rectangle2_widths[267]), .rectangle2_height(rectangle2_heights[267]), .rectangle2_weight(rectangle2_weights[267]), .rectangle3_x(rectangle3_xs[267]), .rectangle3_y(rectangle3_ys[267]), .rectangle3_width(rectangle3_widths[267]), .rectangle3_height(rectangle3_heights[267]), .rectangle3_weight(rectangle3_weights[267]), .feature_threshold(feature_thresholds[267]), .feature_above(feature_aboves[267]), .feature_below(feature_belows[267]), .scan_win_std_dev(scan_win_std_dev[267]), .feature_accum(feature_accums[267]));
  accum_calculator ac268(.scan_win(scan_win268), .rectangle1_x(rectangle1_xs[268]), .rectangle1_y(rectangle1_ys[268]), .rectangle1_width(rectangle1_widths[268]), .rectangle1_height(rectangle1_heights[268]), .rectangle1_weight(rectangle1_weights[268]), .rectangle2_x(rectangle2_xs[268]), .rectangle2_y(rectangle2_ys[268]), .rectangle2_width(rectangle2_widths[268]), .rectangle2_height(rectangle2_heights[268]), .rectangle2_weight(rectangle2_weights[268]), .rectangle3_x(rectangle3_xs[268]), .rectangle3_y(rectangle3_ys[268]), .rectangle3_width(rectangle3_widths[268]), .rectangle3_height(rectangle3_heights[268]), .rectangle3_weight(rectangle3_weights[268]), .feature_threshold(feature_thresholds[268]), .feature_above(feature_aboves[268]), .feature_below(feature_belows[268]), .scan_win_std_dev(scan_win_std_dev[268]), .feature_accum(feature_accums[268]));
  accum_calculator ac269(.scan_win(scan_win269), .rectangle1_x(rectangle1_xs[269]), .rectangle1_y(rectangle1_ys[269]), .rectangle1_width(rectangle1_widths[269]), .rectangle1_height(rectangle1_heights[269]), .rectangle1_weight(rectangle1_weights[269]), .rectangle2_x(rectangle2_xs[269]), .rectangle2_y(rectangle2_ys[269]), .rectangle2_width(rectangle2_widths[269]), .rectangle2_height(rectangle2_heights[269]), .rectangle2_weight(rectangle2_weights[269]), .rectangle3_x(rectangle3_xs[269]), .rectangle3_y(rectangle3_ys[269]), .rectangle3_width(rectangle3_widths[269]), .rectangle3_height(rectangle3_heights[269]), .rectangle3_weight(rectangle3_weights[269]), .feature_threshold(feature_thresholds[269]), .feature_above(feature_aboves[269]), .feature_below(feature_belows[269]), .scan_win_std_dev(scan_win_std_dev[269]), .feature_accum(feature_accums[269]));
  accum_calculator ac270(.scan_win(scan_win270), .rectangle1_x(rectangle1_xs[270]), .rectangle1_y(rectangle1_ys[270]), .rectangle1_width(rectangle1_widths[270]), .rectangle1_height(rectangle1_heights[270]), .rectangle1_weight(rectangle1_weights[270]), .rectangle2_x(rectangle2_xs[270]), .rectangle2_y(rectangle2_ys[270]), .rectangle2_width(rectangle2_widths[270]), .rectangle2_height(rectangle2_heights[270]), .rectangle2_weight(rectangle2_weights[270]), .rectangle3_x(rectangle3_xs[270]), .rectangle3_y(rectangle3_ys[270]), .rectangle3_width(rectangle3_widths[270]), .rectangle3_height(rectangle3_heights[270]), .rectangle3_weight(rectangle3_weights[270]), .feature_threshold(feature_thresholds[270]), .feature_above(feature_aboves[270]), .feature_below(feature_belows[270]), .scan_win_std_dev(scan_win_std_dev[270]), .feature_accum(feature_accums[270]));
  accum_calculator ac271(.scan_win(scan_win271), .rectangle1_x(rectangle1_xs[271]), .rectangle1_y(rectangle1_ys[271]), .rectangle1_width(rectangle1_widths[271]), .rectangle1_height(rectangle1_heights[271]), .rectangle1_weight(rectangle1_weights[271]), .rectangle2_x(rectangle2_xs[271]), .rectangle2_y(rectangle2_ys[271]), .rectangle2_width(rectangle2_widths[271]), .rectangle2_height(rectangle2_heights[271]), .rectangle2_weight(rectangle2_weights[271]), .rectangle3_x(rectangle3_xs[271]), .rectangle3_y(rectangle3_ys[271]), .rectangle3_width(rectangle3_widths[271]), .rectangle3_height(rectangle3_heights[271]), .rectangle3_weight(rectangle3_weights[271]), .feature_threshold(feature_thresholds[271]), .feature_above(feature_aboves[271]), .feature_below(feature_belows[271]), .scan_win_std_dev(scan_win_std_dev[271]), .feature_accum(feature_accums[271]));
  accum_calculator ac272(.scan_win(scan_win272), .rectangle1_x(rectangle1_xs[272]), .rectangle1_y(rectangle1_ys[272]), .rectangle1_width(rectangle1_widths[272]), .rectangle1_height(rectangle1_heights[272]), .rectangle1_weight(rectangle1_weights[272]), .rectangle2_x(rectangle2_xs[272]), .rectangle2_y(rectangle2_ys[272]), .rectangle2_width(rectangle2_widths[272]), .rectangle2_height(rectangle2_heights[272]), .rectangle2_weight(rectangle2_weights[272]), .rectangle3_x(rectangle3_xs[272]), .rectangle3_y(rectangle3_ys[272]), .rectangle3_width(rectangle3_widths[272]), .rectangle3_height(rectangle3_heights[272]), .rectangle3_weight(rectangle3_weights[272]), .feature_threshold(feature_thresholds[272]), .feature_above(feature_aboves[272]), .feature_below(feature_belows[272]), .scan_win_std_dev(scan_win_std_dev[272]), .feature_accum(feature_accums[272]));
  accum_calculator ac273(.scan_win(scan_win273), .rectangle1_x(rectangle1_xs[273]), .rectangle1_y(rectangle1_ys[273]), .rectangle1_width(rectangle1_widths[273]), .rectangle1_height(rectangle1_heights[273]), .rectangle1_weight(rectangle1_weights[273]), .rectangle2_x(rectangle2_xs[273]), .rectangle2_y(rectangle2_ys[273]), .rectangle2_width(rectangle2_widths[273]), .rectangle2_height(rectangle2_heights[273]), .rectangle2_weight(rectangle2_weights[273]), .rectangle3_x(rectangle3_xs[273]), .rectangle3_y(rectangle3_ys[273]), .rectangle3_width(rectangle3_widths[273]), .rectangle3_height(rectangle3_heights[273]), .rectangle3_weight(rectangle3_weights[273]), .feature_threshold(feature_thresholds[273]), .feature_above(feature_aboves[273]), .feature_below(feature_belows[273]), .scan_win_std_dev(scan_win_std_dev[273]), .feature_accum(feature_accums[273]));
  accum_calculator ac274(.scan_win(scan_win274), .rectangle1_x(rectangle1_xs[274]), .rectangle1_y(rectangle1_ys[274]), .rectangle1_width(rectangle1_widths[274]), .rectangle1_height(rectangle1_heights[274]), .rectangle1_weight(rectangle1_weights[274]), .rectangle2_x(rectangle2_xs[274]), .rectangle2_y(rectangle2_ys[274]), .rectangle2_width(rectangle2_widths[274]), .rectangle2_height(rectangle2_heights[274]), .rectangle2_weight(rectangle2_weights[274]), .rectangle3_x(rectangle3_xs[274]), .rectangle3_y(rectangle3_ys[274]), .rectangle3_width(rectangle3_widths[274]), .rectangle3_height(rectangle3_heights[274]), .rectangle3_weight(rectangle3_weights[274]), .feature_threshold(feature_thresholds[274]), .feature_above(feature_aboves[274]), .feature_below(feature_belows[274]), .scan_win_std_dev(scan_win_std_dev[274]), .feature_accum(feature_accums[274]));
  accum_calculator ac275(.scan_win(scan_win275), .rectangle1_x(rectangle1_xs[275]), .rectangle1_y(rectangle1_ys[275]), .rectangle1_width(rectangle1_widths[275]), .rectangle1_height(rectangle1_heights[275]), .rectangle1_weight(rectangle1_weights[275]), .rectangle2_x(rectangle2_xs[275]), .rectangle2_y(rectangle2_ys[275]), .rectangle2_width(rectangle2_widths[275]), .rectangle2_height(rectangle2_heights[275]), .rectangle2_weight(rectangle2_weights[275]), .rectangle3_x(rectangle3_xs[275]), .rectangle3_y(rectangle3_ys[275]), .rectangle3_width(rectangle3_widths[275]), .rectangle3_height(rectangle3_heights[275]), .rectangle3_weight(rectangle3_weights[275]), .feature_threshold(feature_thresholds[275]), .feature_above(feature_aboves[275]), .feature_below(feature_belows[275]), .scan_win_std_dev(scan_win_std_dev[275]), .feature_accum(feature_accums[275]));
  accum_calculator ac276(.scan_win(scan_win276), .rectangle1_x(rectangle1_xs[276]), .rectangle1_y(rectangle1_ys[276]), .rectangle1_width(rectangle1_widths[276]), .rectangle1_height(rectangle1_heights[276]), .rectangle1_weight(rectangle1_weights[276]), .rectangle2_x(rectangle2_xs[276]), .rectangle2_y(rectangle2_ys[276]), .rectangle2_width(rectangle2_widths[276]), .rectangle2_height(rectangle2_heights[276]), .rectangle2_weight(rectangle2_weights[276]), .rectangle3_x(rectangle3_xs[276]), .rectangle3_y(rectangle3_ys[276]), .rectangle3_width(rectangle3_widths[276]), .rectangle3_height(rectangle3_heights[276]), .rectangle3_weight(rectangle3_weights[276]), .feature_threshold(feature_thresholds[276]), .feature_above(feature_aboves[276]), .feature_below(feature_belows[276]), .scan_win_std_dev(scan_win_std_dev[276]), .feature_accum(feature_accums[276]));
  accum_calculator ac277(.scan_win(scan_win277), .rectangle1_x(rectangle1_xs[277]), .rectangle1_y(rectangle1_ys[277]), .rectangle1_width(rectangle1_widths[277]), .rectangle1_height(rectangle1_heights[277]), .rectangle1_weight(rectangle1_weights[277]), .rectangle2_x(rectangle2_xs[277]), .rectangle2_y(rectangle2_ys[277]), .rectangle2_width(rectangle2_widths[277]), .rectangle2_height(rectangle2_heights[277]), .rectangle2_weight(rectangle2_weights[277]), .rectangle3_x(rectangle3_xs[277]), .rectangle3_y(rectangle3_ys[277]), .rectangle3_width(rectangle3_widths[277]), .rectangle3_height(rectangle3_heights[277]), .rectangle3_weight(rectangle3_weights[277]), .feature_threshold(feature_thresholds[277]), .feature_above(feature_aboves[277]), .feature_below(feature_belows[277]), .scan_win_std_dev(scan_win_std_dev[277]), .feature_accum(feature_accums[277]));
  accum_calculator ac278(.scan_win(scan_win278), .rectangle1_x(rectangle1_xs[278]), .rectangle1_y(rectangle1_ys[278]), .rectangle1_width(rectangle1_widths[278]), .rectangle1_height(rectangle1_heights[278]), .rectangle1_weight(rectangle1_weights[278]), .rectangle2_x(rectangle2_xs[278]), .rectangle2_y(rectangle2_ys[278]), .rectangle2_width(rectangle2_widths[278]), .rectangle2_height(rectangle2_heights[278]), .rectangle2_weight(rectangle2_weights[278]), .rectangle3_x(rectangle3_xs[278]), .rectangle3_y(rectangle3_ys[278]), .rectangle3_width(rectangle3_widths[278]), .rectangle3_height(rectangle3_heights[278]), .rectangle3_weight(rectangle3_weights[278]), .feature_threshold(feature_thresholds[278]), .feature_above(feature_aboves[278]), .feature_below(feature_belows[278]), .scan_win_std_dev(scan_win_std_dev[278]), .feature_accum(feature_accums[278]));
  accum_calculator ac279(.scan_win(scan_win279), .rectangle1_x(rectangle1_xs[279]), .rectangle1_y(rectangle1_ys[279]), .rectangle1_width(rectangle1_widths[279]), .rectangle1_height(rectangle1_heights[279]), .rectangle1_weight(rectangle1_weights[279]), .rectangle2_x(rectangle2_xs[279]), .rectangle2_y(rectangle2_ys[279]), .rectangle2_width(rectangle2_widths[279]), .rectangle2_height(rectangle2_heights[279]), .rectangle2_weight(rectangle2_weights[279]), .rectangle3_x(rectangle3_xs[279]), .rectangle3_y(rectangle3_ys[279]), .rectangle3_width(rectangle3_widths[279]), .rectangle3_height(rectangle3_heights[279]), .rectangle3_weight(rectangle3_weights[279]), .feature_threshold(feature_thresholds[279]), .feature_above(feature_aboves[279]), .feature_below(feature_belows[279]), .scan_win_std_dev(scan_win_std_dev[279]), .feature_accum(feature_accums[279]));
  accum_calculator ac280(.scan_win(scan_win280), .rectangle1_x(rectangle1_xs[280]), .rectangle1_y(rectangle1_ys[280]), .rectangle1_width(rectangle1_widths[280]), .rectangle1_height(rectangle1_heights[280]), .rectangle1_weight(rectangle1_weights[280]), .rectangle2_x(rectangle2_xs[280]), .rectangle2_y(rectangle2_ys[280]), .rectangle2_width(rectangle2_widths[280]), .rectangle2_height(rectangle2_heights[280]), .rectangle2_weight(rectangle2_weights[280]), .rectangle3_x(rectangle3_xs[280]), .rectangle3_y(rectangle3_ys[280]), .rectangle3_width(rectangle3_widths[280]), .rectangle3_height(rectangle3_heights[280]), .rectangle3_weight(rectangle3_weights[280]), .feature_threshold(feature_thresholds[280]), .feature_above(feature_aboves[280]), .feature_below(feature_belows[280]), .scan_win_std_dev(scan_win_std_dev[280]), .feature_accum(feature_accums[280]));
  accum_calculator ac281(.scan_win(scan_win281), .rectangle1_x(rectangle1_xs[281]), .rectangle1_y(rectangle1_ys[281]), .rectangle1_width(rectangle1_widths[281]), .rectangle1_height(rectangle1_heights[281]), .rectangle1_weight(rectangle1_weights[281]), .rectangle2_x(rectangle2_xs[281]), .rectangle2_y(rectangle2_ys[281]), .rectangle2_width(rectangle2_widths[281]), .rectangle2_height(rectangle2_heights[281]), .rectangle2_weight(rectangle2_weights[281]), .rectangle3_x(rectangle3_xs[281]), .rectangle3_y(rectangle3_ys[281]), .rectangle3_width(rectangle3_widths[281]), .rectangle3_height(rectangle3_heights[281]), .rectangle3_weight(rectangle3_weights[281]), .feature_threshold(feature_thresholds[281]), .feature_above(feature_aboves[281]), .feature_below(feature_belows[281]), .scan_win_std_dev(scan_win_std_dev[281]), .feature_accum(feature_accums[281]));
  accum_calculator ac282(.scan_win(scan_win282), .rectangle1_x(rectangle1_xs[282]), .rectangle1_y(rectangle1_ys[282]), .rectangle1_width(rectangle1_widths[282]), .rectangle1_height(rectangle1_heights[282]), .rectangle1_weight(rectangle1_weights[282]), .rectangle2_x(rectangle2_xs[282]), .rectangle2_y(rectangle2_ys[282]), .rectangle2_width(rectangle2_widths[282]), .rectangle2_height(rectangle2_heights[282]), .rectangle2_weight(rectangle2_weights[282]), .rectangle3_x(rectangle3_xs[282]), .rectangle3_y(rectangle3_ys[282]), .rectangle3_width(rectangle3_widths[282]), .rectangle3_height(rectangle3_heights[282]), .rectangle3_weight(rectangle3_weights[282]), .feature_threshold(feature_thresholds[282]), .feature_above(feature_aboves[282]), .feature_below(feature_belows[282]), .scan_win_std_dev(scan_win_std_dev[282]), .feature_accum(feature_accums[282]));
  accum_calculator ac283(.scan_win(scan_win283), .rectangle1_x(rectangle1_xs[283]), .rectangle1_y(rectangle1_ys[283]), .rectangle1_width(rectangle1_widths[283]), .rectangle1_height(rectangle1_heights[283]), .rectangle1_weight(rectangle1_weights[283]), .rectangle2_x(rectangle2_xs[283]), .rectangle2_y(rectangle2_ys[283]), .rectangle2_width(rectangle2_widths[283]), .rectangle2_height(rectangle2_heights[283]), .rectangle2_weight(rectangle2_weights[283]), .rectangle3_x(rectangle3_xs[283]), .rectangle3_y(rectangle3_ys[283]), .rectangle3_width(rectangle3_widths[283]), .rectangle3_height(rectangle3_heights[283]), .rectangle3_weight(rectangle3_weights[283]), .feature_threshold(feature_thresholds[283]), .feature_above(feature_aboves[283]), .feature_below(feature_belows[283]), .scan_win_std_dev(scan_win_std_dev[283]), .feature_accum(feature_accums[283]));
  accum_calculator ac284(.scan_win(scan_win284), .rectangle1_x(rectangle1_xs[284]), .rectangle1_y(rectangle1_ys[284]), .rectangle1_width(rectangle1_widths[284]), .rectangle1_height(rectangle1_heights[284]), .rectangle1_weight(rectangle1_weights[284]), .rectangle2_x(rectangle2_xs[284]), .rectangle2_y(rectangle2_ys[284]), .rectangle2_width(rectangle2_widths[284]), .rectangle2_height(rectangle2_heights[284]), .rectangle2_weight(rectangle2_weights[284]), .rectangle3_x(rectangle3_xs[284]), .rectangle3_y(rectangle3_ys[284]), .rectangle3_width(rectangle3_widths[284]), .rectangle3_height(rectangle3_heights[284]), .rectangle3_weight(rectangle3_weights[284]), .feature_threshold(feature_thresholds[284]), .feature_above(feature_aboves[284]), .feature_below(feature_belows[284]), .scan_win_std_dev(scan_win_std_dev[284]), .feature_accum(feature_accums[284]));
  accum_calculator ac285(.scan_win(scan_win285), .rectangle1_x(rectangle1_xs[285]), .rectangle1_y(rectangle1_ys[285]), .rectangle1_width(rectangle1_widths[285]), .rectangle1_height(rectangle1_heights[285]), .rectangle1_weight(rectangle1_weights[285]), .rectangle2_x(rectangle2_xs[285]), .rectangle2_y(rectangle2_ys[285]), .rectangle2_width(rectangle2_widths[285]), .rectangle2_height(rectangle2_heights[285]), .rectangle2_weight(rectangle2_weights[285]), .rectangle3_x(rectangle3_xs[285]), .rectangle3_y(rectangle3_ys[285]), .rectangle3_width(rectangle3_widths[285]), .rectangle3_height(rectangle3_heights[285]), .rectangle3_weight(rectangle3_weights[285]), .feature_threshold(feature_thresholds[285]), .feature_above(feature_aboves[285]), .feature_below(feature_belows[285]), .scan_win_std_dev(scan_win_std_dev[285]), .feature_accum(feature_accums[285]));
  accum_calculator ac286(.scan_win(scan_win286), .rectangle1_x(rectangle1_xs[286]), .rectangle1_y(rectangle1_ys[286]), .rectangle1_width(rectangle1_widths[286]), .rectangle1_height(rectangle1_heights[286]), .rectangle1_weight(rectangle1_weights[286]), .rectangle2_x(rectangle2_xs[286]), .rectangle2_y(rectangle2_ys[286]), .rectangle2_width(rectangle2_widths[286]), .rectangle2_height(rectangle2_heights[286]), .rectangle2_weight(rectangle2_weights[286]), .rectangle3_x(rectangle3_xs[286]), .rectangle3_y(rectangle3_ys[286]), .rectangle3_width(rectangle3_widths[286]), .rectangle3_height(rectangle3_heights[286]), .rectangle3_weight(rectangle3_weights[286]), .feature_threshold(feature_thresholds[286]), .feature_above(feature_aboves[286]), .feature_below(feature_belows[286]), .scan_win_std_dev(scan_win_std_dev[286]), .feature_accum(feature_accums[286]));
  accum_calculator ac287(.scan_win(scan_win287), .rectangle1_x(rectangle1_xs[287]), .rectangle1_y(rectangle1_ys[287]), .rectangle1_width(rectangle1_widths[287]), .rectangle1_height(rectangle1_heights[287]), .rectangle1_weight(rectangle1_weights[287]), .rectangle2_x(rectangle2_xs[287]), .rectangle2_y(rectangle2_ys[287]), .rectangle2_width(rectangle2_widths[287]), .rectangle2_height(rectangle2_heights[287]), .rectangle2_weight(rectangle2_weights[287]), .rectangle3_x(rectangle3_xs[287]), .rectangle3_y(rectangle3_ys[287]), .rectangle3_width(rectangle3_widths[287]), .rectangle3_height(rectangle3_heights[287]), .rectangle3_weight(rectangle3_weights[287]), .feature_threshold(feature_thresholds[287]), .feature_above(feature_aboves[287]), .feature_below(feature_belows[287]), .scan_win_std_dev(scan_win_std_dev[287]), .feature_accum(feature_accums[287]));
  accum_calculator ac288(.scan_win(scan_win288), .rectangle1_x(rectangle1_xs[288]), .rectangle1_y(rectangle1_ys[288]), .rectangle1_width(rectangle1_widths[288]), .rectangle1_height(rectangle1_heights[288]), .rectangle1_weight(rectangle1_weights[288]), .rectangle2_x(rectangle2_xs[288]), .rectangle2_y(rectangle2_ys[288]), .rectangle2_width(rectangle2_widths[288]), .rectangle2_height(rectangle2_heights[288]), .rectangle2_weight(rectangle2_weights[288]), .rectangle3_x(rectangle3_xs[288]), .rectangle3_y(rectangle3_ys[288]), .rectangle3_width(rectangle3_widths[288]), .rectangle3_height(rectangle3_heights[288]), .rectangle3_weight(rectangle3_weights[288]), .feature_threshold(feature_thresholds[288]), .feature_above(feature_aboves[288]), .feature_below(feature_belows[288]), .scan_win_std_dev(scan_win_std_dev[288]), .feature_accum(feature_accums[288]));
  accum_calculator ac289(.scan_win(scan_win289), .rectangle1_x(rectangle1_xs[289]), .rectangle1_y(rectangle1_ys[289]), .rectangle1_width(rectangle1_widths[289]), .rectangle1_height(rectangle1_heights[289]), .rectangle1_weight(rectangle1_weights[289]), .rectangle2_x(rectangle2_xs[289]), .rectangle2_y(rectangle2_ys[289]), .rectangle2_width(rectangle2_widths[289]), .rectangle2_height(rectangle2_heights[289]), .rectangle2_weight(rectangle2_weights[289]), .rectangle3_x(rectangle3_xs[289]), .rectangle3_y(rectangle3_ys[289]), .rectangle3_width(rectangle3_widths[289]), .rectangle3_height(rectangle3_heights[289]), .rectangle3_weight(rectangle3_weights[289]), .feature_threshold(feature_thresholds[289]), .feature_above(feature_aboves[289]), .feature_below(feature_belows[289]), .scan_win_std_dev(scan_win_std_dev[289]), .feature_accum(feature_accums[289]));
  accum_calculator ac290(.scan_win(scan_win290), .rectangle1_x(rectangle1_xs[290]), .rectangle1_y(rectangle1_ys[290]), .rectangle1_width(rectangle1_widths[290]), .rectangle1_height(rectangle1_heights[290]), .rectangle1_weight(rectangle1_weights[290]), .rectangle2_x(rectangle2_xs[290]), .rectangle2_y(rectangle2_ys[290]), .rectangle2_width(rectangle2_widths[290]), .rectangle2_height(rectangle2_heights[290]), .rectangle2_weight(rectangle2_weights[290]), .rectangle3_x(rectangle3_xs[290]), .rectangle3_y(rectangle3_ys[290]), .rectangle3_width(rectangle3_widths[290]), .rectangle3_height(rectangle3_heights[290]), .rectangle3_weight(rectangle3_weights[290]), .feature_threshold(feature_thresholds[290]), .feature_above(feature_aboves[290]), .feature_below(feature_belows[290]), .scan_win_std_dev(scan_win_std_dev[290]), .feature_accum(feature_accums[290]));
  accum_calculator ac291(.scan_win(scan_win291), .rectangle1_x(rectangle1_xs[291]), .rectangle1_y(rectangle1_ys[291]), .rectangle1_width(rectangle1_widths[291]), .rectangle1_height(rectangle1_heights[291]), .rectangle1_weight(rectangle1_weights[291]), .rectangle2_x(rectangle2_xs[291]), .rectangle2_y(rectangle2_ys[291]), .rectangle2_width(rectangle2_widths[291]), .rectangle2_height(rectangle2_heights[291]), .rectangle2_weight(rectangle2_weights[291]), .rectangle3_x(rectangle3_xs[291]), .rectangle3_y(rectangle3_ys[291]), .rectangle3_width(rectangle3_widths[291]), .rectangle3_height(rectangle3_heights[291]), .rectangle3_weight(rectangle3_weights[291]), .feature_threshold(feature_thresholds[291]), .feature_above(feature_aboves[291]), .feature_below(feature_belows[291]), .scan_win_std_dev(scan_win_std_dev[291]), .feature_accum(feature_accums[291]));
  accum_calculator ac292(.scan_win(scan_win292), .rectangle1_x(rectangle1_xs[292]), .rectangle1_y(rectangle1_ys[292]), .rectangle1_width(rectangle1_widths[292]), .rectangle1_height(rectangle1_heights[292]), .rectangle1_weight(rectangle1_weights[292]), .rectangle2_x(rectangle2_xs[292]), .rectangle2_y(rectangle2_ys[292]), .rectangle2_width(rectangle2_widths[292]), .rectangle2_height(rectangle2_heights[292]), .rectangle2_weight(rectangle2_weights[292]), .rectangle3_x(rectangle3_xs[292]), .rectangle3_y(rectangle3_ys[292]), .rectangle3_width(rectangle3_widths[292]), .rectangle3_height(rectangle3_heights[292]), .rectangle3_weight(rectangle3_weights[292]), .feature_threshold(feature_thresholds[292]), .feature_above(feature_aboves[292]), .feature_below(feature_belows[292]), .scan_win_std_dev(scan_win_std_dev[292]), .feature_accum(feature_accums[292]));
  accum_calculator ac293(.scan_win(scan_win293), .rectangle1_x(rectangle1_xs[293]), .rectangle1_y(rectangle1_ys[293]), .rectangle1_width(rectangle1_widths[293]), .rectangle1_height(rectangle1_heights[293]), .rectangle1_weight(rectangle1_weights[293]), .rectangle2_x(rectangle2_xs[293]), .rectangle2_y(rectangle2_ys[293]), .rectangle2_width(rectangle2_widths[293]), .rectangle2_height(rectangle2_heights[293]), .rectangle2_weight(rectangle2_weights[293]), .rectangle3_x(rectangle3_xs[293]), .rectangle3_y(rectangle3_ys[293]), .rectangle3_width(rectangle3_widths[293]), .rectangle3_height(rectangle3_heights[293]), .rectangle3_weight(rectangle3_weights[293]), .feature_threshold(feature_thresholds[293]), .feature_above(feature_aboves[293]), .feature_below(feature_belows[293]), .scan_win_std_dev(scan_win_std_dev[293]), .feature_accum(feature_accums[293]));
  accum_calculator ac294(.scan_win(scan_win294), .rectangle1_x(rectangle1_xs[294]), .rectangle1_y(rectangle1_ys[294]), .rectangle1_width(rectangle1_widths[294]), .rectangle1_height(rectangle1_heights[294]), .rectangle1_weight(rectangle1_weights[294]), .rectangle2_x(rectangle2_xs[294]), .rectangle2_y(rectangle2_ys[294]), .rectangle2_width(rectangle2_widths[294]), .rectangle2_height(rectangle2_heights[294]), .rectangle2_weight(rectangle2_weights[294]), .rectangle3_x(rectangle3_xs[294]), .rectangle3_y(rectangle3_ys[294]), .rectangle3_width(rectangle3_widths[294]), .rectangle3_height(rectangle3_heights[294]), .rectangle3_weight(rectangle3_weights[294]), .feature_threshold(feature_thresholds[294]), .feature_above(feature_aboves[294]), .feature_below(feature_belows[294]), .scan_win_std_dev(scan_win_std_dev[294]), .feature_accum(feature_accums[294]));
  accum_calculator ac295(.scan_win(scan_win295), .rectangle1_x(rectangle1_xs[295]), .rectangle1_y(rectangle1_ys[295]), .rectangle1_width(rectangle1_widths[295]), .rectangle1_height(rectangle1_heights[295]), .rectangle1_weight(rectangle1_weights[295]), .rectangle2_x(rectangle2_xs[295]), .rectangle2_y(rectangle2_ys[295]), .rectangle2_width(rectangle2_widths[295]), .rectangle2_height(rectangle2_heights[295]), .rectangle2_weight(rectangle2_weights[295]), .rectangle3_x(rectangle3_xs[295]), .rectangle3_y(rectangle3_ys[295]), .rectangle3_width(rectangle3_widths[295]), .rectangle3_height(rectangle3_heights[295]), .rectangle3_weight(rectangle3_weights[295]), .feature_threshold(feature_thresholds[295]), .feature_above(feature_aboves[295]), .feature_below(feature_belows[295]), .scan_win_std_dev(scan_win_std_dev[295]), .feature_accum(feature_accums[295]));
  accum_calculator ac296(.scan_win(scan_win296), .rectangle1_x(rectangle1_xs[296]), .rectangle1_y(rectangle1_ys[296]), .rectangle1_width(rectangle1_widths[296]), .rectangle1_height(rectangle1_heights[296]), .rectangle1_weight(rectangle1_weights[296]), .rectangle2_x(rectangle2_xs[296]), .rectangle2_y(rectangle2_ys[296]), .rectangle2_width(rectangle2_widths[296]), .rectangle2_height(rectangle2_heights[296]), .rectangle2_weight(rectangle2_weights[296]), .rectangle3_x(rectangle3_xs[296]), .rectangle3_y(rectangle3_ys[296]), .rectangle3_width(rectangle3_widths[296]), .rectangle3_height(rectangle3_heights[296]), .rectangle3_weight(rectangle3_weights[296]), .feature_threshold(feature_thresholds[296]), .feature_above(feature_aboves[296]), .feature_below(feature_belows[296]), .scan_win_std_dev(scan_win_std_dev[296]), .feature_accum(feature_accums[296]));
  accum_calculator ac297(.scan_win(scan_win297), .rectangle1_x(rectangle1_xs[297]), .rectangle1_y(rectangle1_ys[297]), .rectangle1_width(rectangle1_widths[297]), .rectangle1_height(rectangle1_heights[297]), .rectangle1_weight(rectangle1_weights[297]), .rectangle2_x(rectangle2_xs[297]), .rectangle2_y(rectangle2_ys[297]), .rectangle2_width(rectangle2_widths[297]), .rectangle2_height(rectangle2_heights[297]), .rectangle2_weight(rectangle2_weights[297]), .rectangle3_x(rectangle3_xs[297]), .rectangle3_y(rectangle3_ys[297]), .rectangle3_width(rectangle3_widths[297]), .rectangle3_height(rectangle3_heights[297]), .rectangle3_weight(rectangle3_weights[297]), .feature_threshold(feature_thresholds[297]), .feature_above(feature_aboves[297]), .feature_below(feature_belows[297]), .scan_win_std_dev(scan_win_std_dev[297]), .feature_accum(feature_accums[297]));
  accum_calculator ac298(.scan_win(scan_win298), .rectangle1_x(rectangle1_xs[298]), .rectangle1_y(rectangle1_ys[298]), .rectangle1_width(rectangle1_widths[298]), .rectangle1_height(rectangle1_heights[298]), .rectangle1_weight(rectangle1_weights[298]), .rectangle2_x(rectangle2_xs[298]), .rectangle2_y(rectangle2_ys[298]), .rectangle2_width(rectangle2_widths[298]), .rectangle2_height(rectangle2_heights[298]), .rectangle2_weight(rectangle2_weights[298]), .rectangle3_x(rectangle3_xs[298]), .rectangle3_y(rectangle3_ys[298]), .rectangle3_width(rectangle3_widths[298]), .rectangle3_height(rectangle3_heights[298]), .rectangle3_weight(rectangle3_weights[298]), .feature_threshold(feature_thresholds[298]), .feature_above(feature_aboves[298]), .feature_below(feature_belows[298]), .scan_win_std_dev(scan_win_std_dev[298]), .feature_accum(feature_accums[298]));
  accum_calculator ac299(.scan_win(scan_win299), .rectangle1_x(rectangle1_xs[299]), .rectangle1_y(rectangle1_ys[299]), .rectangle1_width(rectangle1_widths[299]), .rectangle1_height(rectangle1_heights[299]), .rectangle1_weight(rectangle1_weights[299]), .rectangle2_x(rectangle2_xs[299]), .rectangle2_y(rectangle2_ys[299]), .rectangle2_width(rectangle2_widths[299]), .rectangle2_height(rectangle2_heights[299]), .rectangle2_weight(rectangle2_weights[299]), .rectangle3_x(rectangle3_xs[299]), .rectangle3_y(rectangle3_ys[299]), .rectangle3_width(rectangle3_widths[299]), .rectangle3_height(rectangle3_heights[299]), .rectangle3_weight(rectangle3_weights[299]), .feature_threshold(feature_thresholds[299]), .feature_above(feature_aboves[299]), .feature_below(feature_belows[299]), .scan_win_std_dev(scan_win_std_dev[299]), .feature_accum(feature_accums[299]));
  accum_calculator ac300(.scan_win(scan_win300), .rectangle1_x(rectangle1_xs[300]), .rectangle1_y(rectangle1_ys[300]), .rectangle1_width(rectangle1_widths[300]), .rectangle1_height(rectangle1_heights[300]), .rectangle1_weight(rectangle1_weights[300]), .rectangle2_x(rectangle2_xs[300]), .rectangle2_y(rectangle2_ys[300]), .rectangle2_width(rectangle2_widths[300]), .rectangle2_height(rectangle2_heights[300]), .rectangle2_weight(rectangle2_weights[300]), .rectangle3_x(rectangle3_xs[300]), .rectangle3_y(rectangle3_ys[300]), .rectangle3_width(rectangle3_widths[300]), .rectangle3_height(rectangle3_heights[300]), .rectangle3_weight(rectangle3_weights[300]), .feature_threshold(feature_thresholds[300]), .feature_above(feature_aboves[300]), .feature_below(feature_belows[300]), .scan_win_std_dev(scan_win_std_dev[300]), .feature_accum(feature_accums[300]));
  accum_calculator ac301(.scan_win(scan_win301), .rectangle1_x(rectangle1_xs[301]), .rectangle1_y(rectangle1_ys[301]), .rectangle1_width(rectangle1_widths[301]), .rectangle1_height(rectangle1_heights[301]), .rectangle1_weight(rectangle1_weights[301]), .rectangle2_x(rectangle2_xs[301]), .rectangle2_y(rectangle2_ys[301]), .rectangle2_width(rectangle2_widths[301]), .rectangle2_height(rectangle2_heights[301]), .rectangle2_weight(rectangle2_weights[301]), .rectangle3_x(rectangle3_xs[301]), .rectangle3_y(rectangle3_ys[301]), .rectangle3_width(rectangle3_widths[301]), .rectangle3_height(rectangle3_heights[301]), .rectangle3_weight(rectangle3_weights[301]), .feature_threshold(feature_thresholds[301]), .feature_above(feature_aboves[301]), .feature_below(feature_belows[301]), .scan_win_std_dev(scan_win_std_dev[301]), .feature_accum(feature_accums[301]));
  accum_calculator ac302(.scan_win(scan_win302), .rectangle1_x(rectangle1_xs[302]), .rectangle1_y(rectangle1_ys[302]), .rectangle1_width(rectangle1_widths[302]), .rectangle1_height(rectangle1_heights[302]), .rectangle1_weight(rectangle1_weights[302]), .rectangle2_x(rectangle2_xs[302]), .rectangle2_y(rectangle2_ys[302]), .rectangle2_width(rectangle2_widths[302]), .rectangle2_height(rectangle2_heights[302]), .rectangle2_weight(rectangle2_weights[302]), .rectangle3_x(rectangle3_xs[302]), .rectangle3_y(rectangle3_ys[302]), .rectangle3_width(rectangle3_widths[302]), .rectangle3_height(rectangle3_heights[302]), .rectangle3_weight(rectangle3_weights[302]), .feature_threshold(feature_thresholds[302]), .feature_above(feature_aboves[302]), .feature_below(feature_belows[302]), .scan_win_std_dev(scan_win_std_dev[302]), .feature_accum(feature_accums[302]));
  accum_calculator ac303(.scan_win(scan_win303), .rectangle1_x(rectangle1_xs[303]), .rectangle1_y(rectangle1_ys[303]), .rectangle1_width(rectangle1_widths[303]), .rectangle1_height(rectangle1_heights[303]), .rectangle1_weight(rectangle1_weights[303]), .rectangle2_x(rectangle2_xs[303]), .rectangle2_y(rectangle2_ys[303]), .rectangle2_width(rectangle2_widths[303]), .rectangle2_height(rectangle2_heights[303]), .rectangle2_weight(rectangle2_weights[303]), .rectangle3_x(rectangle3_xs[303]), .rectangle3_y(rectangle3_ys[303]), .rectangle3_width(rectangle3_widths[303]), .rectangle3_height(rectangle3_heights[303]), .rectangle3_weight(rectangle3_weights[303]), .feature_threshold(feature_thresholds[303]), .feature_above(feature_aboves[303]), .feature_below(feature_belows[303]), .scan_win_std_dev(scan_win_std_dev[303]), .feature_accum(feature_accums[303]));
  accum_calculator ac304(.scan_win(scan_win304), .rectangle1_x(rectangle1_xs[304]), .rectangle1_y(rectangle1_ys[304]), .rectangle1_width(rectangle1_widths[304]), .rectangle1_height(rectangle1_heights[304]), .rectangle1_weight(rectangle1_weights[304]), .rectangle2_x(rectangle2_xs[304]), .rectangle2_y(rectangle2_ys[304]), .rectangle2_width(rectangle2_widths[304]), .rectangle2_height(rectangle2_heights[304]), .rectangle2_weight(rectangle2_weights[304]), .rectangle3_x(rectangle3_xs[304]), .rectangle3_y(rectangle3_ys[304]), .rectangle3_width(rectangle3_widths[304]), .rectangle3_height(rectangle3_heights[304]), .rectangle3_weight(rectangle3_weights[304]), .feature_threshold(feature_thresholds[304]), .feature_above(feature_aboves[304]), .feature_below(feature_belows[304]), .scan_win_std_dev(scan_win_std_dev[304]), .feature_accum(feature_accums[304]));
  accum_calculator ac305(.scan_win(scan_win305), .rectangle1_x(rectangle1_xs[305]), .rectangle1_y(rectangle1_ys[305]), .rectangle1_width(rectangle1_widths[305]), .rectangle1_height(rectangle1_heights[305]), .rectangle1_weight(rectangle1_weights[305]), .rectangle2_x(rectangle2_xs[305]), .rectangle2_y(rectangle2_ys[305]), .rectangle2_width(rectangle2_widths[305]), .rectangle2_height(rectangle2_heights[305]), .rectangle2_weight(rectangle2_weights[305]), .rectangle3_x(rectangle3_xs[305]), .rectangle3_y(rectangle3_ys[305]), .rectangle3_width(rectangle3_widths[305]), .rectangle3_height(rectangle3_heights[305]), .rectangle3_weight(rectangle3_weights[305]), .feature_threshold(feature_thresholds[305]), .feature_above(feature_aboves[305]), .feature_below(feature_belows[305]), .scan_win_std_dev(scan_win_std_dev[305]), .feature_accum(feature_accums[305]));
  accum_calculator ac306(.scan_win(scan_win306), .rectangle1_x(rectangle1_xs[306]), .rectangle1_y(rectangle1_ys[306]), .rectangle1_width(rectangle1_widths[306]), .rectangle1_height(rectangle1_heights[306]), .rectangle1_weight(rectangle1_weights[306]), .rectangle2_x(rectangle2_xs[306]), .rectangle2_y(rectangle2_ys[306]), .rectangle2_width(rectangle2_widths[306]), .rectangle2_height(rectangle2_heights[306]), .rectangle2_weight(rectangle2_weights[306]), .rectangle3_x(rectangle3_xs[306]), .rectangle3_y(rectangle3_ys[306]), .rectangle3_width(rectangle3_widths[306]), .rectangle3_height(rectangle3_heights[306]), .rectangle3_weight(rectangle3_weights[306]), .feature_threshold(feature_thresholds[306]), .feature_above(feature_aboves[306]), .feature_below(feature_belows[306]), .scan_win_std_dev(scan_win_std_dev[306]), .feature_accum(feature_accums[306]));
  accum_calculator ac307(.scan_win(scan_win307), .rectangle1_x(rectangle1_xs[307]), .rectangle1_y(rectangle1_ys[307]), .rectangle1_width(rectangle1_widths[307]), .rectangle1_height(rectangle1_heights[307]), .rectangle1_weight(rectangle1_weights[307]), .rectangle2_x(rectangle2_xs[307]), .rectangle2_y(rectangle2_ys[307]), .rectangle2_width(rectangle2_widths[307]), .rectangle2_height(rectangle2_heights[307]), .rectangle2_weight(rectangle2_weights[307]), .rectangle3_x(rectangle3_xs[307]), .rectangle3_y(rectangle3_ys[307]), .rectangle3_width(rectangle3_widths[307]), .rectangle3_height(rectangle3_heights[307]), .rectangle3_weight(rectangle3_weights[307]), .feature_threshold(feature_thresholds[307]), .feature_above(feature_aboves[307]), .feature_below(feature_belows[307]), .scan_win_std_dev(scan_win_std_dev[307]), .feature_accum(feature_accums[307]));
  accum_calculator ac308(.scan_win(scan_win308), .rectangle1_x(rectangle1_xs[308]), .rectangle1_y(rectangle1_ys[308]), .rectangle1_width(rectangle1_widths[308]), .rectangle1_height(rectangle1_heights[308]), .rectangle1_weight(rectangle1_weights[308]), .rectangle2_x(rectangle2_xs[308]), .rectangle2_y(rectangle2_ys[308]), .rectangle2_width(rectangle2_widths[308]), .rectangle2_height(rectangle2_heights[308]), .rectangle2_weight(rectangle2_weights[308]), .rectangle3_x(rectangle3_xs[308]), .rectangle3_y(rectangle3_ys[308]), .rectangle3_width(rectangle3_widths[308]), .rectangle3_height(rectangle3_heights[308]), .rectangle3_weight(rectangle3_weights[308]), .feature_threshold(feature_thresholds[308]), .feature_above(feature_aboves[308]), .feature_below(feature_belows[308]), .scan_win_std_dev(scan_win_std_dev[308]), .feature_accum(feature_accums[308]));
  accum_calculator ac309(.scan_win(scan_win309), .rectangle1_x(rectangle1_xs[309]), .rectangle1_y(rectangle1_ys[309]), .rectangle1_width(rectangle1_widths[309]), .rectangle1_height(rectangle1_heights[309]), .rectangle1_weight(rectangle1_weights[309]), .rectangle2_x(rectangle2_xs[309]), .rectangle2_y(rectangle2_ys[309]), .rectangle2_width(rectangle2_widths[309]), .rectangle2_height(rectangle2_heights[309]), .rectangle2_weight(rectangle2_weights[309]), .rectangle3_x(rectangle3_xs[309]), .rectangle3_y(rectangle3_ys[309]), .rectangle3_width(rectangle3_widths[309]), .rectangle3_height(rectangle3_heights[309]), .rectangle3_weight(rectangle3_weights[309]), .feature_threshold(feature_thresholds[309]), .feature_above(feature_aboves[309]), .feature_below(feature_belows[309]), .scan_win_std_dev(scan_win_std_dev[309]), .feature_accum(feature_accums[309]));
  accum_calculator ac310(.scan_win(scan_win310), .rectangle1_x(rectangle1_xs[310]), .rectangle1_y(rectangle1_ys[310]), .rectangle1_width(rectangle1_widths[310]), .rectangle1_height(rectangle1_heights[310]), .rectangle1_weight(rectangle1_weights[310]), .rectangle2_x(rectangle2_xs[310]), .rectangle2_y(rectangle2_ys[310]), .rectangle2_width(rectangle2_widths[310]), .rectangle2_height(rectangle2_heights[310]), .rectangle2_weight(rectangle2_weights[310]), .rectangle3_x(rectangle3_xs[310]), .rectangle3_y(rectangle3_ys[310]), .rectangle3_width(rectangle3_widths[310]), .rectangle3_height(rectangle3_heights[310]), .rectangle3_weight(rectangle3_weights[310]), .feature_threshold(feature_thresholds[310]), .feature_above(feature_aboves[310]), .feature_below(feature_belows[310]), .scan_win_std_dev(scan_win_std_dev[310]), .feature_accum(feature_accums[310]));
  accum_calculator ac311(.scan_win(scan_win311), .rectangle1_x(rectangle1_xs[311]), .rectangle1_y(rectangle1_ys[311]), .rectangle1_width(rectangle1_widths[311]), .rectangle1_height(rectangle1_heights[311]), .rectangle1_weight(rectangle1_weights[311]), .rectangle2_x(rectangle2_xs[311]), .rectangle2_y(rectangle2_ys[311]), .rectangle2_width(rectangle2_widths[311]), .rectangle2_height(rectangle2_heights[311]), .rectangle2_weight(rectangle2_weights[311]), .rectangle3_x(rectangle3_xs[311]), .rectangle3_y(rectangle3_ys[311]), .rectangle3_width(rectangle3_widths[311]), .rectangle3_height(rectangle3_heights[311]), .rectangle3_weight(rectangle3_weights[311]), .feature_threshold(feature_thresholds[311]), .feature_above(feature_aboves[311]), .feature_below(feature_belows[311]), .scan_win_std_dev(scan_win_std_dev[311]), .feature_accum(feature_accums[311]));
  accum_calculator ac312(.scan_win(scan_win312), .rectangle1_x(rectangle1_xs[312]), .rectangle1_y(rectangle1_ys[312]), .rectangle1_width(rectangle1_widths[312]), .rectangle1_height(rectangle1_heights[312]), .rectangle1_weight(rectangle1_weights[312]), .rectangle2_x(rectangle2_xs[312]), .rectangle2_y(rectangle2_ys[312]), .rectangle2_width(rectangle2_widths[312]), .rectangle2_height(rectangle2_heights[312]), .rectangle2_weight(rectangle2_weights[312]), .rectangle3_x(rectangle3_xs[312]), .rectangle3_y(rectangle3_ys[312]), .rectangle3_width(rectangle3_widths[312]), .rectangle3_height(rectangle3_heights[312]), .rectangle3_weight(rectangle3_weights[312]), .feature_threshold(feature_thresholds[312]), .feature_above(feature_aboves[312]), .feature_below(feature_belows[312]), .scan_win_std_dev(scan_win_std_dev[312]), .feature_accum(feature_accums[312]));
  accum_calculator ac313(.scan_win(scan_win313), .rectangle1_x(rectangle1_xs[313]), .rectangle1_y(rectangle1_ys[313]), .rectangle1_width(rectangle1_widths[313]), .rectangle1_height(rectangle1_heights[313]), .rectangle1_weight(rectangle1_weights[313]), .rectangle2_x(rectangle2_xs[313]), .rectangle2_y(rectangle2_ys[313]), .rectangle2_width(rectangle2_widths[313]), .rectangle2_height(rectangle2_heights[313]), .rectangle2_weight(rectangle2_weights[313]), .rectangle3_x(rectangle3_xs[313]), .rectangle3_y(rectangle3_ys[313]), .rectangle3_width(rectangle3_widths[313]), .rectangle3_height(rectangle3_heights[313]), .rectangle3_weight(rectangle3_weights[313]), .feature_threshold(feature_thresholds[313]), .feature_above(feature_aboves[313]), .feature_below(feature_belows[313]), .scan_win_std_dev(scan_win_std_dev[313]), .feature_accum(feature_accums[313]));
  accum_calculator ac314(.scan_win(scan_win314), .rectangle1_x(rectangle1_xs[314]), .rectangle1_y(rectangle1_ys[314]), .rectangle1_width(rectangle1_widths[314]), .rectangle1_height(rectangle1_heights[314]), .rectangle1_weight(rectangle1_weights[314]), .rectangle2_x(rectangle2_xs[314]), .rectangle2_y(rectangle2_ys[314]), .rectangle2_width(rectangle2_widths[314]), .rectangle2_height(rectangle2_heights[314]), .rectangle2_weight(rectangle2_weights[314]), .rectangle3_x(rectangle3_xs[314]), .rectangle3_y(rectangle3_ys[314]), .rectangle3_width(rectangle3_widths[314]), .rectangle3_height(rectangle3_heights[314]), .rectangle3_weight(rectangle3_weights[314]), .feature_threshold(feature_thresholds[314]), .feature_above(feature_aboves[314]), .feature_below(feature_belows[314]), .scan_win_std_dev(scan_win_std_dev[314]), .feature_accum(feature_accums[314]));
  accum_calculator ac315(.scan_win(scan_win315), .rectangle1_x(rectangle1_xs[315]), .rectangle1_y(rectangle1_ys[315]), .rectangle1_width(rectangle1_widths[315]), .rectangle1_height(rectangle1_heights[315]), .rectangle1_weight(rectangle1_weights[315]), .rectangle2_x(rectangle2_xs[315]), .rectangle2_y(rectangle2_ys[315]), .rectangle2_width(rectangle2_widths[315]), .rectangle2_height(rectangle2_heights[315]), .rectangle2_weight(rectangle2_weights[315]), .rectangle3_x(rectangle3_xs[315]), .rectangle3_y(rectangle3_ys[315]), .rectangle3_width(rectangle3_widths[315]), .rectangle3_height(rectangle3_heights[315]), .rectangle3_weight(rectangle3_weights[315]), .feature_threshold(feature_thresholds[315]), .feature_above(feature_aboves[315]), .feature_below(feature_belows[315]), .scan_win_std_dev(scan_win_std_dev[315]), .feature_accum(feature_accums[315]));
  accum_calculator ac316(.scan_win(scan_win316), .rectangle1_x(rectangle1_xs[316]), .rectangle1_y(rectangle1_ys[316]), .rectangle1_width(rectangle1_widths[316]), .rectangle1_height(rectangle1_heights[316]), .rectangle1_weight(rectangle1_weights[316]), .rectangle2_x(rectangle2_xs[316]), .rectangle2_y(rectangle2_ys[316]), .rectangle2_width(rectangle2_widths[316]), .rectangle2_height(rectangle2_heights[316]), .rectangle2_weight(rectangle2_weights[316]), .rectangle3_x(rectangle3_xs[316]), .rectangle3_y(rectangle3_ys[316]), .rectangle3_width(rectangle3_widths[316]), .rectangle3_height(rectangle3_heights[316]), .rectangle3_weight(rectangle3_weights[316]), .feature_threshold(feature_thresholds[316]), .feature_above(feature_aboves[316]), .feature_below(feature_belows[316]), .scan_win_std_dev(scan_win_std_dev[316]), .feature_accum(feature_accums[316]));
  accum_calculator ac317(.scan_win(scan_win317), .rectangle1_x(rectangle1_xs[317]), .rectangle1_y(rectangle1_ys[317]), .rectangle1_width(rectangle1_widths[317]), .rectangle1_height(rectangle1_heights[317]), .rectangle1_weight(rectangle1_weights[317]), .rectangle2_x(rectangle2_xs[317]), .rectangle2_y(rectangle2_ys[317]), .rectangle2_width(rectangle2_widths[317]), .rectangle2_height(rectangle2_heights[317]), .rectangle2_weight(rectangle2_weights[317]), .rectangle3_x(rectangle3_xs[317]), .rectangle3_y(rectangle3_ys[317]), .rectangle3_width(rectangle3_widths[317]), .rectangle3_height(rectangle3_heights[317]), .rectangle3_weight(rectangle3_weights[317]), .feature_threshold(feature_thresholds[317]), .feature_above(feature_aboves[317]), .feature_below(feature_belows[317]), .scan_win_std_dev(scan_win_std_dev[317]), .feature_accum(feature_accums[317]));
  accum_calculator ac318(.scan_win(scan_win318), .rectangle1_x(rectangle1_xs[318]), .rectangle1_y(rectangle1_ys[318]), .rectangle1_width(rectangle1_widths[318]), .rectangle1_height(rectangle1_heights[318]), .rectangle1_weight(rectangle1_weights[318]), .rectangle2_x(rectangle2_xs[318]), .rectangle2_y(rectangle2_ys[318]), .rectangle2_width(rectangle2_widths[318]), .rectangle2_height(rectangle2_heights[318]), .rectangle2_weight(rectangle2_weights[318]), .rectangle3_x(rectangle3_xs[318]), .rectangle3_y(rectangle3_ys[318]), .rectangle3_width(rectangle3_widths[318]), .rectangle3_height(rectangle3_heights[318]), .rectangle3_weight(rectangle3_weights[318]), .feature_threshold(feature_thresholds[318]), .feature_above(feature_aboves[318]), .feature_below(feature_belows[318]), .scan_win_std_dev(scan_win_std_dev[318]), .feature_accum(feature_accums[318]));
  accum_calculator ac319(.scan_win(scan_win319), .rectangle1_x(rectangle1_xs[319]), .rectangle1_y(rectangle1_ys[319]), .rectangle1_width(rectangle1_widths[319]), .rectangle1_height(rectangle1_heights[319]), .rectangle1_weight(rectangle1_weights[319]), .rectangle2_x(rectangle2_xs[319]), .rectangle2_y(rectangle2_ys[319]), .rectangle2_width(rectangle2_widths[319]), .rectangle2_height(rectangle2_heights[319]), .rectangle2_weight(rectangle2_weights[319]), .rectangle3_x(rectangle3_xs[319]), .rectangle3_y(rectangle3_ys[319]), .rectangle3_width(rectangle3_widths[319]), .rectangle3_height(rectangle3_heights[319]), .rectangle3_weight(rectangle3_weights[319]), .feature_threshold(feature_thresholds[319]), .feature_above(feature_aboves[319]), .feature_below(feature_belows[319]), .scan_win_std_dev(scan_win_std_dev[319]), .feature_accum(feature_accums[319]));
  accum_calculator ac320(.scan_win(scan_win320), .rectangle1_x(rectangle1_xs[320]), .rectangle1_y(rectangle1_ys[320]), .rectangle1_width(rectangle1_widths[320]), .rectangle1_height(rectangle1_heights[320]), .rectangle1_weight(rectangle1_weights[320]), .rectangle2_x(rectangle2_xs[320]), .rectangle2_y(rectangle2_ys[320]), .rectangle2_width(rectangle2_widths[320]), .rectangle2_height(rectangle2_heights[320]), .rectangle2_weight(rectangle2_weights[320]), .rectangle3_x(rectangle3_xs[320]), .rectangle3_y(rectangle3_ys[320]), .rectangle3_width(rectangle3_widths[320]), .rectangle3_height(rectangle3_heights[320]), .rectangle3_weight(rectangle3_weights[320]), .feature_threshold(feature_thresholds[320]), .feature_above(feature_aboves[320]), .feature_below(feature_belows[320]), .scan_win_std_dev(scan_win_std_dev[320]), .feature_accum(feature_accums[320]));
  accum_calculator ac321(.scan_win(scan_win321), .rectangle1_x(rectangle1_xs[321]), .rectangle1_y(rectangle1_ys[321]), .rectangle1_width(rectangle1_widths[321]), .rectangle1_height(rectangle1_heights[321]), .rectangle1_weight(rectangle1_weights[321]), .rectangle2_x(rectangle2_xs[321]), .rectangle2_y(rectangle2_ys[321]), .rectangle2_width(rectangle2_widths[321]), .rectangle2_height(rectangle2_heights[321]), .rectangle2_weight(rectangle2_weights[321]), .rectangle3_x(rectangle3_xs[321]), .rectangle3_y(rectangle3_ys[321]), .rectangle3_width(rectangle3_widths[321]), .rectangle3_height(rectangle3_heights[321]), .rectangle3_weight(rectangle3_weights[321]), .feature_threshold(feature_thresholds[321]), .feature_above(feature_aboves[321]), .feature_below(feature_belows[321]), .scan_win_std_dev(scan_win_std_dev[321]), .feature_accum(feature_accums[321]));
  accum_calculator ac322(.scan_win(scan_win322), .rectangle1_x(rectangle1_xs[322]), .rectangle1_y(rectangle1_ys[322]), .rectangle1_width(rectangle1_widths[322]), .rectangle1_height(rectangle1_heights[322]), .rectangle1_weight(rectangle1_weights[322]), .rectangle2_x(rectangle2_xs[322]), .rectangle2_y(rectangle2_ys[322]), .rectangle2_width(rectangle2_widths[322]), .rectangle2_height(rectangle2_heights[322]), .rectangle2_weight(rectangle2_weights[322]), .rectangle3_x(rectangle3_xs[322]), .rectangle3_y(rectangle3_ys[322]), .rectangle3_width(rectangle3_widths[322]), .rectangle3_height(rectangle3_heights[322]), .rectangle3_weight(rectangle3_weights[322]), .feature_threshold(feature_thresholds[322]), .feature_above(feature_aboves[322]), .feature_below(feature_belows[322]), .scan_win_std_dev(scan_win_std_dev[322]), .feature_accum(feature_accums[322]));
  accum_calculator ac323(.scan_win(scan_win323), .rectangle1_x(rectangle1_xs[323]), .rectangle1_y(rectangle1_ys[323]), .rectangle1_width(rectangle1_widths[323]), .rectangle1_height(rectangle1_heights[323]), .rectangle1_weight(rectangle1_weights[323]), .rectangle2_x(rectangle2_xs[323]), .rectangle2_y(rectangle2_ys[323]), .rectangle2_width(rectangle2_widths[323]), .rectangle2_height(rectangle2_heights[323]), .rectangle2_weight(rectangle2_weights[323]), .rectangle3_x(rectangle3_xs[323]), .rectangle3_y(rectangle3_ys[323]), .rectangle3_width(rectangle3_widths[323]), .rectangle3_height(rectangle3_heights[323]), .rectangle3_weight(rectangle3_weights[323]), .feature_threshold(feature_thresholds[323]), .feature_above(feature_aboves[323]), .feature_below(feature_belows[323]), .scan_win_std_dev(scan_win_std_dev[323]), .feature_accum(feature_accums[323]));
  accum_calculator ac324(.scan_win(scan_win324), .rectangle1_x(rectangle1_xs[324]), .rectangle1_y(rectangle1_ys[324]), .rectangle1_width(rectangle1_widths[324]), .rectangle1_height(rectangle1_heights[324]), .rectangle1_weight(rectangle1_weights[324]), .rectangle2_x(rectangle2_xs[324]), .rectangle2_y(rectangle2_ys[324]), .rectangle2_width(rectangle2_widths[324]), .rectangle2_height(rectangle2_heights[324]), .rectangle2_weight(rectangle2_weights[324]), .rectangle3_x(rectangle3_xs[324]), .rectangle3_y(rectangle3_ys[324]), .rectangle3_width(rectangle3_widths[324]), .rectangle3_height(rectangle3_heights[324]), .rectangle3_weight(rectangle3_weights[324]), .feature_threshold(feature_thresholds[324]), .feature_above(feature_aboves[324]), .feature_below(feature_belows[324]), .scan_win_std_dev(scan_win_std_dev[324]), .feature_accum(feature_accums[324]));
  accum_calculator ac325(.scan_win(scan_win325), .rectangle1_x(rectangle1_xs[325]), .rectangle1_y(rectangle1_ys[325]), .rectangle1_width(rectangle1_widths[325]), .rectangle1_height(rectangle1_heights[325]), .rectangle1_weight(rectangle1_weights[325]), .rectangle2_x(rectangle2_xs[325]), .rectangle2_y(rectangle2_ys[325]), .rectangle2_width(rectangle2_widths[325]), .rectangle2_height(rectangle2_heights[325]), .rectangle2_weight(rectangle2_weights[325]), .rectangle3_x(rectangle3_xs[325]), .rectangle3_y(rectangle3_ys[325]), .rectangle3_width(rectangle3_widths[325]), .rectangle3_height(rectangle3_heights[325]), .rectangle3_weight(rectangle3_weights[325]), .feature_threshold(feature_thresholds[325]), .feature_above(feature_aboves[325]), .feature_below(feature_belows[325]), .scan_win_std_dev(scan_win_std_dev[325]), .feature_accum(feature_accums[325]));
  accum_calculator ac326(.scan_win(scan_win326), .rectangle1_x(rectangle1_xs[326]), .rectangle1_y(rectangle1_ys[326]), .rectangle1_width(rectangle1_widths[326]), .rectangle1_height(rectangle1_heights[326]), .rectangle1_weight(rectangle1_weights[326]), .rectangle2_x(rectangle2_xs[326]), .rectangle2_y(rectangle2_ys[326]), .rectangle2_width(rectangle2_widths[326]), .rectangle2_height(rectangle2_heights[326]), .rectangle2_weight(rectangle2_weights[326]), .rectangle3_x(rectangle3_xs[326]), .rectangle3_y(rectangle3_ys[326]), .rectangle3_width(rectangle3_widths[326]), .rectangle3_height(rectangle3_heights[326]), .rectangle3_weight(rectangle3_weights[326]), .feature_threshold(feature_thresholds[326]), .feature_above(feature_aboves[326]), .feature_below(feature_belows[326]), .scan_win_std_dev(scan_win_std_dev[326]), .feature_accum(feature_accums[326]));
  accum_calculator ac327(.scan_win(scan_win327), .rectangle1_x(rectangle1_xs[327]), .rectangle1_y(rectangle1_ys[327]), .rectangle1_width(rectangle1_widths[327]), .rectangle1_height(rectangle1_heights[327]), .rectangle1_weight(rectangle1_weights[327]), .rectangle2_x(rectangle2_xs[327]), .rectangle2_y(rectangle2_ys[327]), .rectangle2_width(rectangle2_widths[327]), .rectangle2_height(rectangle2_heights[327]), .rectangle2_weight(rectangle2_weights[327]), .rectangle3_x(rectangle3_xs[327]), .rectangle3_y(rectangle3_ys[327]), .rectangle3_width(rectangle3_widths[327]), .rectangle3_height(rectangle3_heights[327]), .rectangle3_weight(rectangle3_weights[327]), .feature_threshold(feature_thresholds[327]), .feature_above(feature_aboves[327]), .feature_below(feature_belows[327]), .scan_win_std_dev(scan_win_std_dev[327]), .feature_accum(feature_accums[327]));
  accum_calculator ac328(.scan_win(scan_win328), .rectangle1_x(rectangle1_xs[328]), .rectangle1_y(rectangle1_ys[328]), .rectangle1_width(rectangle1_widths[328]), .rectangle1_height(rectangle1_heights[328]), .rectangle1_weight(rectangle1_weights[328]), .rectangle2_x(rectangle2_xs[328]), .rectangle2_y(rectangle2_ys[328]), .rectangle2_width(rectangle2_widths[328]), .rectangle2_height(rectangle2_heights[328]), .rectangle2_weight(rectangle2_weights[328]), .rectangle3_x(rectangle3_xs[328]), .rectangle3_y(rectangle3_ys[328]), .rectangle3_width(rectangle3_widths[328]), .rectangle3_height(rectangle3_heights[328]), .rectangle3_weight(rectangle3_weights[328]), .feature_threshold(feature_thresholds[328]), .feature_above(feature_aboves[328]), .feature_below(feature_belows[328]), .scan_win_std_dev(scan_win_std_dev[328]), .feature_accum(feature_accums[328]));
  accum_calculator ac329(.scan_win(scan_win329), .rectangle1_x(rectangle1_xs[329]), .rectangle1_y(rectangle1_ys[329]), .rectangle1_width(rectangle1_widths[329]), .rectangle1_height(rectangle1_heights[329]), .rectangle1_weight(rectangle1_weights[329]), .rectangle2_x(rectangle2_xs[329]), .rectangle2_y(rectangle2_ys[329]), .rectangle2_width(rectangle2_widths[329]), .rectangle2_height(rectangle2_heights[329]), .rectangle2_weight(rectangle2_weights[329]), .rectangle3_x(rectangle3_xs[329]), .rectangle3_y(rectangle3_ys[329]), .rectangle3_width(rectangle3_widths[329]), .rectangle3_height(rectangle3_heights[329]), .rectangle3_weight(rectangle3_weights[329]), .feature_threshold(feature_thresholds[329]), .feature_above(feature_aboves[329]), .feature_below(feature_belows[329]), .scan_win_std_dev(scan_win_std_dev[329]), .feature_accum(feature_accums[329]));
  accum_calculator ac330(.scan_win(scan_win330), .rectangle1_x(rectangle1_xs[330]), .rectangle1_y(rectangle1_ys[330]), .rectangle1_width(rectangle1_widths[330]), .rectangle1_height(rectangle1_heights[330]), .rectangle1_weight(rectangle1_weights[330]), .rectangle2_x(rectangle2_xs[330]), .rectangle2_y(rectangle2_ys[330]), .rectangle2_width(rectangle2_widths[330]), .rectangle2_height(rectangle2_heights[330]), .rectangle2_weight(rectangle2_weights[330]), .rectangle3_x(rectangle3_xs[330]), .rectangle3_y(rectangle3_ys[330]), .rectangle3_width(rectangle3_widths[330]), .rectangle3_height(rectangle3_heights[330]), .rectangle3_weight(rectangle3_weights[330]), .feature_threshold(feature_thresholds[330]), .feature_above(feature_aboves[330]), .feature_below(feature_belows[330]), .scan_win_std_dev(scan_win_std_dev[330]), .feature_accum(feature_accums[330]));
  accum_calculator ac331(.scan_win(scan_win331), .rectangle1_x(rectangle1_xs[331]), .rectangle1_y(rectangle1_ys[331]), .rectangle1_width(rectangle1_widths[331]), .rectangle1_height(rectangle1_heights[331]), .rectangle1_weight(rectangle1_weights[331]), .rectangle2_x(rectangle2_xs[331]), .rectangle2_y(rectangle2_ys[331]), .rectangle2_width(rectangle2_widths[331]), .rectangle2_height(rectangle2_heights[331]), .rectangle2_weight(rectangle2_weights[331]), .rectangle3_x(rectangle3_xs[331]), .rectangle3_y(rectangle3_ys[331]), .rectangle3_width(rectangle3_widths[331]), .rectangle3_height(rectangle3_heights[331]), .rectangle3_weight(rectangle3_weights[331]), .feature_threshold(feature_thresholds[331]), .feature_above(feature_aboves[331]), .feature_below(feature_belows[331]), .scan_win_std_dev(scan_win_std_dev[331]), .feature_accum(feature_accums[331]));
  accum_calculator ac332(.scan_win(scan_win332), .rectangle1_x(rectangle1_xs[332]), .rectangle1_y(rectangle1_ys[332]), .rectangle1_width(rectangle1_widths[332]), .rectangle1_height(rectangle1_heights[332]), .rectangle1_weight(rectangle1_weights[332]), .rectangle2_x(rectangle2_xs[332]), .rectangle2_y(rectangle2_ys[332]), .rectangle2_width(rectangle2_widths[332]), .rectangle2_height(rectangle2_heights[332]), .rectangle2_weight(rectangle2_weights[332]), .rectangle3_x(rectangle3_xs[332]), .rectangle3_y(rectangle3_ys[332]), .rectangle3_width(rectangle3_widths[332]), .rectangle3_height(rectangle3_heights[332]), .rectangle3_weight(rectangle3_weights[332]), .feature_threshold(feature_thresholds[332]), .feature_above(feature_aboves[332]), .feature_below(feature_belows[332]), .scan_win_std_dev(scan_win_std_dev[332]), .feature_accum(feature_accums[332]));
  accum_calculator ac333(.scan_win(scan_win333), .rectangle1_x(rectangle1_xs[333]), .rectangle1_y(rectangle1_ys[333]), .rectangle1_width(rectangle1_widths[333]), .rectangle1_height(rectangle1_heights[333]), .rectangle1_weight(rectangle1_weights[333]), .rectangle2_x(rectangle2_xs[333]), .rectangle2_y(rectangle2_ys[333]), .rectangle2_width(rectangle2_widths[333]), .rectangle2_height(rectangle2_heights[333]), .rectangle2_weight(rectangle2_weights[333]), .rectangle3_x(rectangle3_xs[333]), .rectangle3_y(rectangle3_ys[333]), .rectangle3_width(rectangle3_widths[333]), .rectangle3_height(rectangle3_heights[333]), .rectangle3_weight(rectangle3_weights[333]), .feature_threshold(feature_thresholds[333]), .feature_above(feature_aboves[333]), .feature_below(feature_belows[333]), .scan_win_std_dev(scan_win_std_dev[333]), .feature_accum(feature_accums[333]));
  accum_calculator ac334(.scan_win(scan_win334), .rectangle1_x(rectangle1_xs[334]), .rectangle1_y(rectangle1_ys[334]), .rectangle1_width(rectangle1_widths[334]), .rectangle1_height(rectangle1_heights[334]), .rectangle1_weight(rectangle1_weights[334]), .rectangle2_x(rectangle2_xs[334]), .rectangle2_y(rectangle2_ys[334]), .rectangle2_width(rectangle2_widths[334]), .rectangle2_height(rectangle2_heights[334]), .rectangle2_weight(rectangle2_weights[334]), .rectangle3_x(rectangle3_xs[334]), .rectangle3_y(rectangle3_ys[334]), .rectangle3_width(rectangle3_widths[334]), .rectangle3_height(rectangle3_heights[334]), .rectangle3_weight(rectangle3_weights[334]), .feature_threshold(feature_thresholds[334]), .feature_above(feature_aboves[334]), .feature_below(feature_belows[334]), .scan_win_std_dev(scan_win_std_dev[334]), .feature_accum(feature_accums[334]));
  accum_calculator ac335(.scan_win(scan_win335), .rectangle1_x(rectangle1_xs[335]), .rectangle1_y(rectangle1_ys[335]), .rectangle1_width(rectangle1_widths[335]), .rectangle1_height(rectangle1_heights[335]), .rectangle1_weight(rectangle1_weights[335]), .rectangle2_x(rectangle2_xs[335]), .rectangle2_y(rectangle2_ys[335]), .rectangle2_width(rectangle2_widths[335]), .rectangle2_height(rectangle2_heights[335]), .rectangle2_weight(rectangle2_weights[335]), .rectangle3_x(rectangle3_xs[335]), .rectangle3_y(rectangle3_ys[335]), .rectangle3_width(rectangle3_widths[335]), .rectangle3_height(rectangle3_heights[335]), .rectangle3_weight(rectangle3_weights[335]), .feature_threshold(feature_thresholds[335]), .feature_above(feature_aboves[335]), .feature_below(feature_belows[335]), .scan_win_std_dev(scan_win_std_dev[335]), .feature_accum(feature_accums[335]));
  accum_calculator ac336(.scan_win(scan_win336), .rectangle1_x(rectangle1_xs[336]), .rectangle1_y(rectangle1_ys[336]), .rectangle1_width(rectangle1_widths[336]), .rectangle1_height(rectangle1_heights[336]), .rectangle1_weight(rectangle1_weights[336]), .rectangle2_x(rectangle2_xs[336]), .rectangle2_y(rectangle2_ys[336]), .rectangle2_width(rectangle2_widths[336]), .rectangle2_height(rectangle2_heights[336]), .rectangle2_weight(rectangle2_weights[336]), .rectangle3_x(rectangle3_xs[336]), .rectangle3_y(rectangle3_ys[336]), .rectangle3_width(rectangle3_widths[336]), .rectangle3_height(rectangle3_heights[336]), .rectangle3_weight(rectangle3_weights[336]), .feature_threshold(feature_thresholds[336]), .feature_above(feature_aboves[336]), .feature_below(feature_belows[336]), .scan_win_std_dev(scan_win_std_dev[336]), .feature_accum(feature_accums[336]));
  accum_calculator ac337(.scan_win(scan_win337), .rectangle1_x(rectangle1_xs[337]), .rectangle1_y(rectangle1_ys[337]), .rectangle1_width(rectangle1_widths[337]), .rectangle1_height(rectangle1_heights[337]), .rectangle1_weight(rectangle1_weights[337]), .rectangle2_x(rectangle2_xs[337]), .rectangle2_y(rectangle2_ys[337]), .rectangle2_width(rectangle2_widths[337]), .rectangle2_height(rectangle2_heights[337]), .rectangle2_weight(rectangle2_weights[337]), .rectangle3_x(rectangle3_xs[337]), .rectangle3_y(rectangle3_ys[337]), .rectangle3_width(rectangle3_widths[337]), .rectangle3_height(rectangle3_heights[337]), .rectangle3_weight(rectangle3_weights[337]), .feature_threshold(feature_thresholds[337]), .feature_above(feature_aboves[337]), .feature_below(feature_belows[337]), .scan_win_std_dev(scan_win_std_dev[337]), .feature_accum(feature_accums[337]));
  accum_calculator ac338(.scan_win(scan_win338), .rectangle1_x(rectangle1_xs[338]), .rectangle1_y(rectangle1_ys[338]), .rectangle1_width(rectangle1_widths[338]), .rectangle1_height(rectangle1_heights[338]), .rectangle1_weight(rectangle1_weights[338]), .rectangle2_x(rectangle2_xs[338]), .rectangle2_y(rectangle2_ys[338]), .rectangle2_width(rectangle2_widths[338]), .rectangle2_height(rectangle2_heights[338]), .rectangle2_weight(rectangle2_weights[338]), .rectangle3_x(rectangle3_xs[338]), .rectangle3_y(rectangle3_ys[338]), .rectangle3_width(rectangle3_widths[338]), .rectangle3_height(rectangle3_heights[338]), .rectangle3_weight(rectangle3_weights[338]), .feature_threshold(feature_thresholds[338]), .feature_above(feature_aboves[338]), .feature_below(feature_belows[338]), .scan_win_std_dev(scan_win_std_dev[338]), .feature_accum(feature_accums[338]));
  accum_calculator ac339(.scan_win(scan_win339), .rectangle1_x(rectangle1_xs[339]), .rectangle1_y(rectangle1_ys[339]), .rectangle1_width(rectangle1_widths[339]), .rectangle1_height(rectangle1_heights[339]), .rectangle1_weight(rectangle1_weights[339]), .rectangle2_x(rectangle2_xs[339]), .rectangle2_y(rectangle2_ys[339]), .rectangle2_width(rectangle2_widths[339]), .rectangle2_height(rectangle2_heights[339]), .rectangle2_weight(rectangle2_weights[339]), .rectangle3_x(rectangle3_xs[339]), .rectangle3_y(rectangle3_ys[339]), .rectangle3_width(rectangle3_widths[339]), .rectangle3_height(rectangle3_heights[339]), .rectangle3_weight(rectangle3_weights[339]), .feature_threshold(feature_thresholds[339]), .feature_above(feature_aboves[339]), .feature_below(feature_belows[339]), .scan_win_std_dev(scan_win_std_dev[339]), .feature_accum(feature_accums[339]));
  accum_calculator ac340(.scan_win(scan_win340), .rectangle1_x(rectangle1_xs[340]), .rectangle1_y(rectangle1_ys[340]), .rectangle1_width(rectangle1_widths[340]), .rectangle1_height(rectangle1_heights[340]), .rectangle1_weight(rectangle1_weights[340]), .rectangle2_x(rectangle2_xs[340]), .rectangle2_y(rectangle2_ys[340]), .rectangle2_width(rectangle2_widths[340]), .rectangle2_height(rectangle2_heights[340]), .rectangle2_weight(rectangle2_weights[340]), .rectangle3_x(rectangle3_xs[340]), .rectangle3_y(rectangle3_ys[340]), .rectangle3_width(rectangle3_widths[340]), .rectangle3_height(rectangle3_heights[340]), .rectangle3_weight(rectangle3_weights[340]), .feature_threshold(feature_thresholds[340]), .feature_above(feature_aboves[340]), .feature_below(feature_belows[340]), .scan_win_std_dev(scan_win_std_dev[340]), .feature_accum(feature_accums[340]));
  accum_calculator ac341(.scan_win(scan_win341), .rectangle1_x(rectangle1_xs[341]), .rectangle1_y(rectangle1_ys[341]), .rectangle1_width(rectangle1_widths[341]), .rectangle1_height(rectangle1_heights[341]), .rectangle1_weight(rectangle1_weights[341]), .rectangle2_x(rectangle2_xs[341]), .rectangle2_y(rectangle2_ys[341]), .rectangle2_width(rectangle2_widths[341]), .rectangle2_height(rectangle2_heights[341]), .rectangle2_weight(rectangle2_weights[341]), .rectangle3_x(rectangle3_xs[341]), .rectangle3_y(rectangle3_ys[341]), .rectangle3_width(rectangle3_widths[341]), .rectangle3_height(rectangle3_heights[341]), .rectangle3_weight(rectangle3_weights[341]), .feature_threshold(feature_thresholds[341]), .feature_above(feature_aboves[341]), .feature_below(feature_belows[341]), .scan_win_std_dev(scan_win_std_dev[341]), .feature_accum(feature_accums[341]));
  accum_calculator ac342(.scan_win(scan_win342), .rectangle1_x(rectangle1_xs[342]), .rectangle1_y(rectangle1_ys[342]), .rectangle1_width(rectangle1_widths[342]), .rectangle1_height(rectangle1_heights[342]), .rectangle1_weight(rectangle1_weights[342]), .rectangle2_x(rectangle2_xs[342]), .rectangle2_y(rectangle2_ys[342]), .rectangle2_width(rectangle2_widths[342]), .rectangle2_height(rectangle2_heights[342]), .rectangle2_weight(rectangle2_weights[342]), .rectangle3_x(rectangle3_xs[342]), .rectangle3_y(rectangle3_ys[342]), .rectangle3_width(rectangle3_widths[342]), .rectangle3_height(rectangle3_heights[342]), .rectangle3_weight(rectangle3_weights[342]), .feature_threshold(feature_thresholds[342]), .feature_above(feature_aboves[342]), .feature_below(feature_belows[342]), .scan_win_std_dev(scan_win_std_dev[342]), .feature_accum(feature_accums[342]));
  accum_calculator ac343(.scan_win(scan_win343), .rectangle1_x(rectangle1_xs[343]), .rectangle1_y(rectangle1_ys[343]), .rectangle1_width(rectangle1_widths[343]), .rectangle1_height(rectangle1_heights[343]), .rectangle1_weight(rectangle1_weights[343]), .rectangle2_x(rectangle2_xs[343]), .rectangle2_y(rectangle2_ys[343]), .rectangle2_width(rectangle2_widths[343]), .rectangle2_height(rectangle2_heights[343]), .rectangle2_weight(rectangle2_weights[343]), .rectangle3_x(rectangle3_xs[343]), .rectangle3_y(rectangle3_ys[343]), .rectangle3_width(rectangle3_widths[343]), .rectangle3_height(rectangle3_heights[343]), .rectangle3_weight(rectangle3_weights[343]), .feature_threshold(feature_thresholds[343]), .feature_above(feature_aboves[343]), .feature_below(feature_belows[343]), .scan_win_std_dev(scan_win_std_dev[343]), .feature_accum(feature_accums[343]));
  accum_calculator ac344(.scan_win(scan_win344), .rectangle1_x(rectangle1_xs[344]), .rectangle1_y(rectangle1_ys[344]), .rectangle1_width(rectangle1_widths[344]), .rectangle1_height(rectangle1_heights[344]), .rectangle1_weight(rectangle1_weights[344]), .rectangle2_x(rectangle2_xs[344]), .rectangle2_y(rectangle2_ys[344]), .rectangle2_width(rectangle2_widths[344]), .rectangle2_height(rectangle2_heights[344]), .rectangle2_weight(rectangle2_weights[344]), .rectangle3_x(rectangle3_xs[344]), .rectangle3_y(rectangle3_ys[344]), .rectangle3_width(rectangle3_widths[344]), .rectangle3_height(rectangle3_heights[344]), .rectangle3_weight(rectangle3_weights[344]), .feature_threshold(feature_thresholds[344]), .feature_above(feature_aboves[344]), .feature_below(feature_belows[344]), .scan_win_std_dev(scan_win_std_dev[344]), .feature_accum(feature_accums[344]));
  accum_calculator ac345(.scan_win(scan_win345), .rectangle1_x(rectangle1_xs[345]), .rectangle1_y(rectangle1_ys[345]), .rectangle1_width(rectangle1_widths[345]), .rectangle1_height(rectangle1_heights[345]), .rectangle1_weight(rectangle1_weights[345]), .rectangle2_x(rectangle2_xs[345]), .rectangle2_y(rectangle2_ys[345]), .rectangle2_width(rectangle2_widths[345]), .rectangle2_height(rectangle2_heights[345]), .rectangle2_weight(rectangle2_weights[345]), .rectangle3_x(rectangle3_xs[345]), .rectangle3_y(rectangle3_ys[345]), .rectangle3_width(rectangle3_widths[345]), .rectangle3_height(rectangle3_heights[345]), .rectangle3_weight(rectangle3_weights[345]), .feature_threshold(feature_thresholds[345]), .feature_above(feature_aboves[345]), .feature_below(feature_belows[345]), .scan_win_std_dev(scan_win_std_dev[345]), .feature_accum(feature_accums[345]));
  accum_calculator ac346(.scan_win(scan_win346), .rectangle1_x(rectangle1_xs[346]), .rectangle1_y(rectangle1_ys[346]), .rectangle1_width(rectangle1_widths[346]), .rectangle1_height(rectangle1_heights[346]), .rectangle1_weight(rectangle1_weights[346]), .rectangle2_x(rectangle2_xs[346]), .rectangle2_y(rectangle2_ys[346]), .rectangle2_width(rectangle2_widths[346]), .rectangle2_height(rectangle2_heights[346]), .rectangle2_weight(rectangle2_weights[346]), .rectangle3_x(rectangle3_xs[346]), .rectangle3_y(rectangle3_ys[346]), .rectangle3_width(rectangle3_widths[346]), .rectangle3_height(rectangle3_heights[346]), .rectangle3_weight(rectangle3_weights[346]), .feature_threshold(feature_thresholds[346]), .feature_above(feature_aboves[346]), .feature_below(feature_belows[346]), .scan_win_std_dev(scan_win_std_dev[346]), .feature_accum(feature_accums[346]));
  accum_calculator ac347(.scan_win(scan_win347), .rectangle1_x(rectangle1_xs[347]), .rectangle1_y(rectangle1_ys[347]), .rectangle1_width(rectangle1_widths[347]), .rectangle1_height(rectangle1_heights[347]), .rectangle1_weight(rectangle1_weights[347]), .rectangle2_x(rectangle2_xs[347]), .rectangle2_y(rectangle2_ys[347]), .rectangle2_width(rectangle2_widths[347]), .rectangle2_height(rectangle2_heights[347]), .rectangle2_weight(rectangle2_weights[347]), .rectangle3_x(rectangle3_xs[347]), .rectangle3_y(rectangle3_ys[347]), .rectangle3_width(rectangle3_widths[347]), .rectangle3_height(rectangle3_heights[347]), .rectangle3_weight(rectangle3_weights[347]), .feature_threshold(feature_thresholds[347]), .feature_above(feature_aboves[347]), .feature_below(feature_belows[347]), .scan_win_std_dev(scan_win_std_dev[347]), .feature_accum(feature_accums[347]));
  accum_calculator ac348(.scan_win(scan_win348), .rectangle1_x(rectangle1_xs[348]), .rectangle1_y(rectangle1_ys[348]), .rectangle1_width(rectangle1_widths[348]), .rectangle1_height(rectangle1_heights[348]), .rectangle1_weight(rectangle1_weights[348]), .rectangle2_x(rectangle2_xs[348]), .rectangle2_y(rectangle2_ys[348]), .rectangle2_width(rectangle2_widths[348]), .rectangle2_height(rectangle2_heights[348]), .rectangle2_weight(rectangle2_weights[348]), .rectangle3_x(rectangle3_xs[348]), .rectangle3_y(rectangle3_ys[348]), .rectangle3_width(rectangle3_widths[348]), .rectangle3_height(rectangle3_heights[348]), .rectangle3_weight(rectangle3_weights[348]), .feature_threshold(feature_thresholds[348]), .feature_above(feature_aboves[348]), .feature_below(feature_belows[348]), .scan_win_std_dev(scan_win_std_dev[348]), .feature_accum(feature_accums[348]));
  accum_calculator ac349(.scan_win(scan_win349), .rectangle1_x(rectangle1_xs[349]), .rectangle1_y(rectangle1_ys[349]), .rectangle1_width(rectangle1_widths[349]), .rectangle1_height(rectangle1_heights[349]), .rectangle1_weight(rectangle1_weights[349]), .rectangle2_x(rectangle2_xs[349]), .rectangle2_y(rectangle2_ys[349]), .rectangle2_width(rectangle2_widths[349]), .rectangle2_height(rectangle2_heights[349]), .rectangle2_weight(rectangle2_weights[349]), .rectangle3_x(rectangle3_xs[349]), .rectangle3_y(rectangle3_ys[349]), .rectangle3_width(rectangle3_widths[349]), .rectangle3_height(rectangle3_heights[349]), .rectangle3_weight(rectangle3_weights[349]), .feature_threshold(feature_thresholds[349]), .feature_above(feature_aboves[349]), .feature_below(feature_belows[349]), .scan_win_std_dev(scan_win_std_dev[349]), .feature_accum(feature_accums[349]));
  accum_calculator ac350(.scan_win(scan_win350), .rectangle1_x(rectangle1_xs[350]), .rectangle1_y(rectangle1_ys[350]), .rectangle1_width(rectangle1_widths[350]), .rectangle1_height(rectangle1_heights[350]), .rectangle1_weight(rectangle1_weights[350]), .rectangle2_x(rectangle2_xs[350]), .rectangle2_y(rectangle2_ys[350]), .rectangle2_width(rectangle2_widths[350]), .rectangle2_height(rectangle2_heights[350]), .rectangle2_weight(rectangle2_weights[350]), .rectangle3_x(rectangle3_xs[350]), .rectangle3_y(rectangle3_ys[350]), .rectangle3_width(rectangle3_widths[350]), .rectangle3_height(rectangle3_heights[350]), .rectangle3_weight(rectangle3_weights[350]), .feature_threshold(feature_thresholds[350]), .feature_above(feature_aboves[350]), .feature_below(feature_belows[350]), .scan_win_std_dev(scan_win_std_dev[350]), .feature_accum(feature_accums[350]));
  accum_calculator ac351(.scan_win(scan_win351), .rectangle1_x(rectangle1_xs[351]), .rectangle1_y(rectangle1_ys[351]), .rectangle1_width(rectangle1_widths[351]), .rectangle1_height(rectangle1_heights[351]), .rectangle1_weight(rectangle1_weights[351]), .rectangle2_x(rectangle2_xs[351]), .rectangle2_y(rectangle2_ys[351]), .rectangle2_width(rectangle2_widths[351]), .rectangle2_height(rectangle2_heights[351]), .rectangle2_weight(rectangle2_weights[351]), .rectangle3_x(rectangle3_xs[351]), .rectangle3_y(rectangle3_ys[351]), .rectangle3_width(rectangle3_widths[351]), .rectangle3_height(rectangle3_heights[351]), .rectangle3_weight(rectangle3_weights[351]), .feature_threshold(feature_thresholds[351]), .feature_above(feature_aboves[351]), .feature_below(feature_belows[351]), .scan_win_std_dev(scan_win_std_dev[351]), .feature_accum(feature_accums[351]));
  accum_calculator ac352(.scan_win(scan_win352), .rectangle1_x(rectangle1_xs[352]), .rectangle1_y(rectangle1_ys[352]), .rectangle1_width(rectangle1_widths[352]), .rectangle1_height(rectangle1_heights[352]), .rectangle1_weight(rectangle1_weights[352]), .rectangle2_x(rectangle2_xs[352]), .rectangle2_y(rectangle2_ys[352]), .rectangle2_width(rectangle2_widths[352]), .rectangle2_height(rectangle2_heights[352]), .rectangle2_weight(rectangle2_weights[352]), .rectangle3_x(rectangle3_xs[352]), .rectangle3_y(rectangle3_ys[352]), .rectangle3_width(rectangle3_widths[352]), .rectangle3_height(rectangle3_heights[352]), .rectangle3_weight(rectangle3_weights[352]), .feature_threshold(feature_thresholds[352]), .feature_above(feature_aboves[352]), .feature_below(feature_belows[352]), .scan_win_std_dev(scan_win_std_dev[352]), .feature_accum(feature_accums[352]));
  accum_calculator ac353(.scan_win(scan_win353), .rectangle1_x(rectangle1_xs[353]), .rectangle1_y(rectangle1_ys[353]), .rectangle1_width(rectangle1_widths[353]), .rectangle1_height(rectangle1_heights[353]), .rectangle1_weight(rectangle1_weights[353]), .rectangle2_x(rectangle2_xs[353]), .rectangle2_y(rectangle2_ys[353]), .rectangle2_width(rectangle2_widths[353]), .rectangle2_height(rectangle2_heights[353]), .rectangle2_weight(rectangle2_weights[353]), .rectangle3_x(rectangle3_xs[353]), .rectangle3_y(rectangle3_ys[353]), .rectangle3_width(rectangle3_widths[353]), .rectangle3_height(rectangle3_heights[353]), .rectangle3_weight(rectangle3_weights[353]), .feature_threshold(feature_thresholds[353]), .feature_above(feature_aboves[353]), .feature_below(feature_belows[353]), .scan_win_std_dev(scan_win_std_dev[353]), .feature_accum(feature_accums[353]));
  accum_calculator ac354(.scan_win(scan_win354), .rectangle1_x(rectangle1_xs[354]), .rectangle1_y(rectangle1_ys[354]), .rectangle1_width(rectangle1_widths[354]), .rectangle1_height(rectangle1_heights[354]), .rectangle1_weight(rectangle1_weights[354]), .rectangle2_x(rectangle2_xs[354]), .rectangle2_y(rectangle2_ys[354]), .rectangle2_width(rectangle2_widths[354]), .rectangle2_height(rectangle2_heights[354]), .rectangle2_weight(rectangle2_weights[354]), .rectangle3_x(rectangle3_xs[354]), .rectangle3_y(rectangle3_ys[354]), .rectangle3_width(rectangle3_widths[354]), .rectangle3_height(rectangle3_heights[354]), .rectangle3_weight(rectangle3_weights[354]), .feature_threshold(feature_thresholds[354]), .feature_above(feature_aboves[354]), .feature_below(feature_belows[354]), .scan_win_std_dev(scan_win_std_dev[354]), .feature_accum(feature_accums[354]));
  accum_calculator ac355(.scan_win(scan_win355), .rectangle1_x(rectangle1_xs[355]), .rectangle1_y(rectangle1_ys[355]), .rectangle1_width(rectangle1_widths[355]), .rectangle1_height(rectangle1_heights[355]), .rectangle1_weight(rectangle1_weights[355]), .rectangle2_x(rectangle2_xs[355]), .rectangle2_y(rectangle2_ys[355]), .rectangle2_width(rectangle2_widths[355]), .rectangle2_height(rectangle2_heights[355]), .rectangle2_weight(rectangle2_weights[355]), .rectangle3_x(rectangle3_xs[355]), .rectangle3_y(rectangle3_ys[355]), .rectangle3_width(rectangle3_widths[355]), .rectangle3_height(rectangle3_heights[355]), .rectangle3_weight(rectangle3_weights[355]), .feature_threshold(feature_thresholds[355]), .feature_above(feature_aboves[355]), .feature_below(feature_belows[355]), .scan_win_std_dev(scan_win_std_dev[355]), .feature_accum(feature_accums[355]));
  accum_calculator ac356(.scan_win(scan_win356), .rectangle1_x(rectangle1_xs[356]), .rectangle1_y(rectangle1_ys[356]), .rectangle1_width(rectangle1_widths[356]), .rectangle1_height(rectangle1_heights[356]), .rectangle1_weight(rectangle1_weights[356]), .rectangle2_x(rectangle2_xs[356]), .rectangle2_y(rectangle2_ys[356]), .rectangle2_width(rectangle2_widths[356]), .rectangle2_height(rectangle2_heights[356]), .rectangle2_weight(rectangle2_weights[356]), .rectangle3_x(rectangle3_xs[356]), .rectangle3_y(rectangle3_ys[356]), .rectangle3_width(rectangle3_widths[356]), .rectangle3_height(rectangle3_heights[356]), .rectangle3_weight(rectangle3_weights[356]), .feature_threshold(feature_thresholds[356]), .feature_above(feature_aboves[356]), .feature_below(feature_belows[356]), .scan_win_std_dev(scan_win_std_dev[356]), .feature_accum(feature_accums[356]));
  accum_calculator ac357(.scan_win(scan_win357), .rectangle1_x(rectangle1_xs[357]), .rectangle1_y(rectangle1_ys[357]), .rectangle1_width(rectangle1_widths[357]), .rectangle1_height(rectangle1_heights[357]), .rectangle1_weight(rectangle1_weights[357]), .rectangle2_x(rectangle2_xs[357]), .rectangle2_y(rectangle2_ys[357]), .rectangle2_width(rectangle2_widths[357]), .rectangle2_height(rectangle2_heights[357]), .rectangle2_weight(rectangle2_weights[357]), .rectangle3_x(rectangle3_xs[357]), .rectangle3_y(rectangle3_ys[357]), .rectangle3_width(rectangle3_widths[357]), .rectangle3_height(rectangle3_heights[357]), .rectangle3_weight(rectangle3_weights[357]), .feature_threshold(feature_thresholds[357]), .feature_above(feature_aboves[357]), .feature_below(feature_belows[357]), .scan_win_std_dev(scan_win_std_dev[357]), .feature_accum(feature_accums[357]));
  accum_calculator ac358(.scan_win(scan_win358), .rectangle1_x(rectangle1_xs[358]), .rectangle1_y(rectangle1_ys[358]), .rectangle1_width(rectangle1_widths[358]), .rectangle1_height(rectangle1_heights[358]), .rectangle1_weight(rectangle1_weights[358]), .rectangle2_x(rectangle2_xs[358]), .rectangle2_y(rectangle2_ys[358]), .rectangle2_width(rectangle2_widths[358]), .rectangle2_height(rectangle2_heights[358]), .rectangle2_weight(rectangle2_weights[358]), .rectangle3_x(rectangle3_xs[358]), .rectangle3_y(rectangle3_ys[358]), .rectangle3_width(rectangle3_widths[358]), .rectangle3_height(rectangle3_heights[358]), .rectangle3_weight(rectangle3_weights[358]), .feature_threshold(feature_thresholds[358]), .feature_above(feature_aboves[358]), .feature_below(feature_belows[358]), .scan_win_std_dev(scan_win_std_dev[358]), .feature_accum(feature_accums[358]));
  accum_calculator ac359(.scan_win(scan_win359), .rectangle1_x(rectangle1_xs[359]), .rectangle1_y(rectangle1_ys[359]), .rectangle1_width(rectangle1_widths[359]), .rectangle1_height(rectangle1_heights[359]), .rectangle1_weight(rectangle1_weights[359]), .rectangle2_x(rectangle2_xs[359]), .rectangle2_y(rectangle2_ys[359]), .rectangle2_width(rectangle2_widths[359]), .rectangle2_height(rectangle2_heights[359]), .rectangle2_weight(rectangle2_weights[359]), .rectangle3_x(rectangle3_xs[359]), .rectangle3_y(rectangle3_ys[359]), .rectangle3_width(rectangle3_widths[359]), .rectangle3_height(rectangle3_heights[359]), .rectangle3_weight(rectangle3_weights[359]), .feature_threshold(feature_thresholds[359]), .feature_above(feature_aboves[359]), .feature_below(feature_belows[359]), .scan_win_std_dev(scan_win_std_dev[359]), .feature_accum(feature_accums[359]));
  accum_calculator ac360(.scan_win(scan_win360), .rectangle1_x(rectangle1_xs[360]), .rectangle1_y(rectangle1_ys[360]), .rectangle1_width(rectangle1_widths[360]), .rectangle1_height(rectangle1_heights[360]), .rectangle1_weight(rectangle1_weights[360]), .rectangle2_x(rectangle2_xs[360]), .rectangle2_y(rectangle2_ys[360]), .rectangle2_width(rectangle2_widths[360]), .rectangle2_height(rectangle2_heights[360]), .rectangle2_weight(rectangle2_weights[360]), .rectangle3_x(rectangle3_xs[360]), .rectangle3_y(rectangle3_ys[360]), .rectangle3_width(rectangle3_widths[360]), .rectangle3_height(rectangle3_heights[360]), .rectangle3_weight(rectangle3_weights[360]), .feature_threshold(feature_thresholds[360]), .feature_above(feature_aboves[360]), .feature_below(feature_belows[360]), .scan_win_std_dev(scan_win_std_dev[360]), .feature_accum(feature_accums[360]));
  accum_calculator ac361(.scan_win(scan_win361), .rectangle1_x(rectangle1_xs[361]), .rectangle1_y(rectangle1_ys[361]), .rectangle1_width(rectangle1_widths[361]), .rectangle1_height(rectangle1_heights[361]), .rectangle1_weight(rectangle1_weights[361]), .rectangle2_x(rectangle2_xs[361]), .rectangle2_y(rectangle2_ys[361]), .rectangle2_width(rectangle2_widths[361]), .rectangle2_height(rectangle2_heights[361]), .rectangle2_weight(rectangle2_weights[361]), .rectangle3_x(rectangle3_xs[361]), .rectangle3_y(rectangle3_ys[361]), .rectangle3_width(rectangle3_widths[361]), .rectangle3_height(rectangle3_heights[361]), .rectangle3_weight(rectangle3_weights[361]), .feature_threshold(feature_thresholds[361]), .feature_above(feature_aboves[361]), .feature_below(feature_belows[361]), .scan_win_std_dev(scan_win_std_dev[361]), .feature_accum(feature_accums[361]));
  accum_calculator ac362(.scan_win(scan_win362), .rectangle1_x(rectangle1_xs[362]), .rectangle1_y(rectangle1_ys[362]), .rectangle1_width(rectangle1_widths[362]), .rectangle1_height(rectangle1_heights[362]), .rectangle1_weight(rectangle1_weights[362]), .rectangle2_x(rectangle2_xs[362]), .rectangle2_y(rectangle2_ys[362]), .rectangle2_width(rectangle2_widths[362]), .rectangle2_height(rectangle2_heights[362]), .rectangle2_weight(rectangle2_weights[362]), .rectangle3_x(rectangle3_xs[362]), .rectangle3_y(rectangle3_ys[362]), .rectangle3_width(rectangle3_widths[362]), .rectangle3_height(rectangle3_heights[362]), .rectangle3_weight(rectangle3_weights[362]), .feature_threshold(feature_thresholds[362]), .feature_above(feature_aboves[362]), .feature_below(feature_belows[362]), .scan_win_std_dev(scan_win_std_dev[362]), .feature_accum(feature_accums[362]));
  accum_calculator ac363(.scan_win(scan_win363), .rectangle1_x(rectangle1_xs[363]), .rectangle1_y(rectangle1_ys[363]), .rectangle1_width(rectangle1_widths[363]), .rectangle1_height(rectangle1_heights[363]), .rectangle1_weight(rectangle1_weights[363]), .rectangle2_x(rectangle2_xs[363]), .rectangle2_y(rectangle2_ys[363]), .rectangle2_width(rectangle2_widths[363]), .rectangle2_height(rectangle2_heights[363]), .rectangle2_weight(rectangle2_weights[363]), .rectangle3_x(rectangle3_xs[363]), .rectangle3_y(rectangle3_ys[363]), .rectangle3_width(rectangle3_widths[363]), .rectangle3_height(rectangle3_heights[363]), .rectangle3_weight(rectangle3_weights[363]), .feature_threshold(feature_thresholds[363]), .feature_above(feature_aboves[363]), .feature_below(feature_belows[363]), .scan_win_std_dev(scan_win_std_dev[363]), .feature_accum(feature_accums[363]));
  accum_calculator ac364(.scan_win(scan_win364), .rectangle1_x(rectangle1_xs[364]), .rectangle1_y(rectangle1_ys[364]), .rectangle1_width(rectangle1_widths[364]), .rectangle1_height(rectangle1_heights[364]), .rectangle1_weight(rectangle1_weights[364]), .rectangle2_x(rectangle2_xs[364]), .rectangle2_y(rectangle2_ys[364]), .rectangle2_width(rectangle2_widths[364]), .rectangle2_height(rectangle2_heights[364]), .rectangle2_weight(rectangle2_weights[364]), .rectangle3_x(rectangle3_xs[364]), .rectangle3_y(rectangle3_ys[364]), .rectangle3_width(rectangle3_widths[364]), .rectangle3_height(rectangle3_heights[364]), .rectangle3_weight(rectangle3_weights[364]), .feature_threshold(feature_thresholds[364]), .feature_above(feature_aboves[364]), .feature_below(feature_belows[364]), .scan_win_std_dev(scan_win_std_dev[364]), .feature_accum(feature_accums[364]));
  accum_calculator ac365(.scan_win(scan_win365), .rectangle1_x(rectangle1_xs[365]), .rectangle1_y(rectangle1_ys[365]), .rectangle1_width(rectangle1_widths[365]), .rectangle1_height(rectangle1_heights[365]), .rectangle1_weight(rectangle1_weights[365]), .rectangle2_x(rectangle2_xs[365]), .rectangle2_y(rectangle2_ys[365]), .rectangle2_width(rectangle2_widths[365]), .rectangle2_height(rectangle2_heights[365]), .rectangle2_weight(rectangle2_weights[365]), .rectangle3_x(rectangle3_xs[365]), .rectangle3_y(rectangle3_ys[365]), .rectangle3_width(rectangle3_widths[365]), .rectangle3_height(rectangle3_heights[365]), .rectangle3_weight(rectangle3_weights[365]), .feature_threshold(feature_thresholds[365]), .feature_above(feature_aboves[365]), .feature_below(feature_belows[365]), .scan_win_std_dev(scan_win_std_dev[365]), .feature_accum(feature_accums[365]));
  accum_calculator ac366(.scan_win(scan_win366), .rectangle1_x(rectangle1_xs[366]), .rectangle1_y(rectangle1_ys[366]), .rectangle1_width(rectangle1_widths[366]), .rectangle1_height(rectangle1_heights[366]), .rectangle1_weight(rectangle1_weights[366]), .rectangle2_x(rectangle2_xs[366]), .rectangle2_y(rectangle2_ys[366]), .rectangle2_width(rectangle2_widths[366]), .rectangle2_height(rectangle2_heights[366]), .rectangle2_weight(rectangle2_weights[366]), .rectangle3_x(rectangle3_xs[366]), .rectangle3_y(rectangle3_ys[366]), .rectangle3_width(rectangle3_widths[366]), .rectangle3_height(rectangle3_heights[366]), .rectangle3_weight(rectangle3_weights[366]), .feature_threshold(feature_thresholds[366]), .feature_above(feature_aboves[366]), .feature_below(feature_belows[366]), .scan_win_std_dev(scan_win_std_dev[366]), .feature_accum(feature_accums[366]));
  accum_calculator ac367(.scan_win(scan_win367), .rectangle1_x(rectangle1_xs[367]), .rectangle1_y(rectangle1_ys[367]), .rectangle1_width(rectangle1_widths[367]), .rectangle1_height(rectangle1_heights[367]), .rectangle1_weight(rectangle1_weights[367]), .rectangle2_x(rectangle2_xs[367]), .rectangle2_y(rectangle2_ys[367]), .rectangle2_width(rectangle2_widths[367]), .rectangle2_height(rectangle2_heights[367]), .rectangle2_weight(rectangle2_weights[367]), .rectangle3_x(rectangle3_xs[367]), .rectangle3_y(rectangle3_ys[367]), .rectangle3_width(rectangle3_widths[367]), .rectangle3_height(rectangle3_heights[367]), .rectangle3_weight(rectangle3_weights[367]), .feature_threshold(feature_thresholds[367]), .feature_above(feature_aboves[367]), .feature_below(feature_belows[367]), .scan_win_std_dev(scan_win_std_dev[367]), .feature_accum(feature_accums[367]));
  accum_calculator ac368(.scan_win(scan_win368), .rectangle1_x(rectangle1_xs[368]), .rectangle1_y(rectangle1_ys[368]), .rectangle1_width(rectangle1_widths[368]), .rectangle1_height(rectangle1_heights[368]), .rectangle1_weight(rectangle1_weights[368]), .rectangle2_x(rectangle2_xs[368]), .rectangle2_y(rectangle2_ys[368]), .rectangle2_width(rectangle2_widths[368]), .rectangle2_height(rectangle2_heights[368]), .rectangle2_weight(rectangle2_weights[368]), .rectangle3_x(rectangle3_xs[368]), .rectangle3_y(rectangle3_ys[368]), .rectangle3_width(rectangle3_widths[368]), .rectangle3_height(rectangle3_heights[368]), .rectangle3_weight(rectangle3_weights[368]), .feature_threshold(feature_thresholds[368]), .feature_above(feature_aboves[368]), .feature_below(feature_belows[368]), .scan_win_std_dev(scan_win_std_dev[368]), .feature_accum(feature_accums[368]));
  accum_calculator ac369(.scan_win(scan_win369), .rectangle1_x(rectangle1_xs[369]), .rectangle1_y(rectangle1_ys[369]), .rectangle1_width(rectangle1_widths[369]), .rectangle1_height(rectangle1_heights[369]), .rectangle1_weight(rectangle1_weights[369]), .rectangle2_x(rectangle2_xs[369]), .rectangle2_y(rectangle2_ys[369]), .rectangle2_width(rectangle2_widths[369]), .rectangle2_height(rectangle2_heights[369]), .rectangle2_weight(rectangle2_weights[369]), .rectangle3_x(rectangle3_xs[369]), .rectangle3_y(rectangle3_ys[369]), .rectangle3_width(rectangle3_widths[369]), .rectangle3_height(rectangle3_heights[369]), .rectangle3_weight(rectangle3_weights[369]), .feature_threshold(feature_thresholds[369]), .feature_above(feature_aboves[369]), .feature_below(feature_belows[369]), .scan_win_std_dev(scan_win_std_dev[369]), .feature_accum(feature_accums[369]));
  accum_calculator ac370(.scan_win(scan_win370), .rectangle1_x(rectangle1_xs[370]), .rectangle1_y(rectangle1_ys[370]), .rectangle1_width(rectangle1_widths[370]), .rectangle1_height(rectangle1_heights[370]), .rectangle1_weight(rectangle1_weights[370]), .rectangle2_x(rectangle2_xs[370]), .rectangle2_y(rectangle2_ys[370]), .rectangle2_width(rectangle2_widths[370]), .rectangle2_height(rectangle2_heights[370]), .rectangle2_weight(rectangle2_weights[370]), .rectangle3_x(rectangle3_xs[370]), .rectangle3_y(rectangle3_ys[370]), .rectangle3_width(rectangle3_widths[370]), .rectangle3_height(rectangle3_heights[370]), .rectangle3_weight(rectangle3_weights[370]), .feature_threshold(feature_thresholds[370]), .feature_above(feature_aboves[370]), .feature_below(feature_belows[370]), .scan_win_std_dev(scan_win_std_dev[370]), .feature_accum(feature_accums[370]));
  accum_calculator ac371(.scan_win(scan_win371), .rectangle1_x(rectangle1_xs[371]), .rectangle1_y(rectangle1_ys[371]), .rectangle1_width(rectangle1_widths[371]), .rectangle1_height(rectangle1_heights[371]), .rectangle1_weight(rectangle1_weights[371]), .rectangle2_x(rectangle2_xs[371]), .rectangle2_y(rectangle2_ys[371]), .rectangle2_width(rectangle2_widths[371]), .rectangle2_height(rectangle2_heights[371]), .rectangle2_weight(rectangle2_weights[371]), .rectangle3_x(rectangle3_xs[371]), .rectangle3_y(rectangle3_ys[371]), .rectangle3_width(rectangle3_widths[371]), .rectangle3_height(rectangle3_heights[371]), .rectangle3_weight(rectangle3_weights[371]), .feature_threshold(feature_thresholds[371]), .feature_above(feature_aboves[371]), .feature_below(feature_belows[371]), .scan_win_std_dev(scan_win_std_dev[371]), .feature_accum(feature_accums[371]));
  accum_calculator ac372(.scan_win(scan_win372), .rectangle1_x(rectangle1_xs[372]), .rectangle1_y(rectangle1_ys[372]), .rectangle1_width(rectangle1_widths[372]), .rectangle1_height(rectangle1_heights[372]), .rectangle1_weight(rectangle1_weights[372]), .rectangle2_x(rectangle2_xs[372]), .rectangle2_y(rectangle2_ys[372]), .rectangle2_width(rectangle2_widths[372]), .rectangle2_height(rectangle2_heights[372]), .rectangle2_weight(rectangle2_weights[372]), .rectangle3_x(rectangle3_xs[372]), .rectangle3_y(rectangle3_ys[372]), .rectangle3_width(rectangle3_widths[372]), .rectangle3_height(rectangle3_heights[372]), .rectangle3_weight(rectangle3_weights[372]), .feature_threshold(feature_thresholds[372]), .feature_above(feature_aboves[372]), .feature_below(feature_belows[372]), .scan_win_std_dev(scan_win_std_dev[372]), .feature_accum(feature_accums[372]));
  accum_calculator ac373(.scan_win(scan_win373), .rectangle1_x(rectangle1_xs[373]), .rectangle1_y(rectangle1_ys[373]), .rectangle1_width(rectangle1_widths[373]), .rectangle1_height(rectangle1_heights[373]), .rectangle1_weight(rectangle1_weights[373]), .rectangle2_x(rectangle2_xs[373]), .rectangle2_y(rectangle2_ys[373]), .rectangle2_width(rectangle2_widths[373]), .rectangle2_height(rectangle2_heights[373]), .rectangle2_weight(rectangle2_weights[373]), .rectangle3_x(rectangle3_xs[373]), .rectangle3_y(rectangle3_ys[373]), .rectangle3_width(rectangle3_widths[373]), .rectangle3_height(rectangle3_heights[373]), .rectangle3_weight(rectangle3_weights[373]), .feature_threshold(feature_thresholds[373]), .feature_above(feature_aboves[373]), .feature_below(feature_belows[373]), .scan_win_std_dev(scan_win_std_dev[373]), .feature_accum(feature_accums[373]));
  accum_calculator ac374(.scan_win(scan_win374), .rectangle1_x(rectangle1_xs[374]), .rectangle1_y(rectangle1_ys[374]), .rectangle1_width(rectangle1_widths[374]), .rectangle1_height(rectangle1_heights[374]), .rectangle1_weight(rectangle1_weights[374]), .rectangle2_x(rectangle2_xs[374]), .rectangle2_y(rectangle2_ys[374]), .rectangle2_width(rectangle2_widths[374]), .rectangle2_height(rectangle2_heights[374]), .rectangle2_weight(rectangle2_weights[374]), .rectangle3_x(rectangle3_xs[374]), .rectangle3_y(rectangle3_ys[374]), .rectangle3_width(rectangle3_widths[374]), .rectangle3_height(rectangle3_heights[374]), .rectangle3_weight(rectangle3_weights[374]), .feature_threshold(feature_thresholds[374]), .feature_above(feature_aboves[374]), .feature_below(feature_belows[374]), .scan_win_std_dev(scan_win_std_dev[374]), .feature_accum(feature_accums[374]));
  accum_calculator ac375(.scan_win(scan_win375), .rectangle1_x(rectangle1_xs[375]), .rectangle1_y(rectangle1_ys[375]), .rectangle1_width(rectangle1_widths[375]), .rectangle1_height(rectangle1_heights[375]), .rectangle1_weight(rectangle1_weights[375]), .rectangle2_x(rectangle2_xs[375]), .rectangle2_y(rectangle2_ys[375]), .rectangle2_width(rectangle2_widths[375]), .rectangle2_height(rectangle2_heights[375]), .rectangle2_weight(rectangle2_weights[375]), .rectangle3_x(rectangle3_xs[375]), .rectangle3_y(rectangle3_ys[375]), .rectangle3_width(rectangle3_widths[375]), .rectangle3_height(rectangle3_heights[375]), .rectangle3_weight(rectangle3_weights[375]), .feature_threshold(feature_thresholds[375]), .feature_above(feature_aboves[375]), .feature_below(feature_belows[375]), .scan_win_std_dev(scan_win_std_dev[375]), .feature_accum(feature_accums[375]));
  accum_calculator ac376(.scan_win(scan_win376), .rectangle1_x(rectangle1_xs[376]), .rectangle1_y(rectangle1_ys[376]), .rectangle1_width(rectangle1_widths[376]), .rectangle1_height(rectangle1_heights[376]), .rectangle1_weight(rectangle1_weights[376]), .rectangle2_x(rectangle2_xs[376]), .rectangle2_y(rectangle2_ys[376]), .rectangle2_width(rectangle2_widths[376]), .rectangle2_height(rectangle2_heights[376]), .rectangle2_weight(rectangle2_weights[376]), .rectangle3_x(rectangle3_xs[376]), .rectangle3_y(rectangle3_ys[376]), .rectangle3_width(rectangle3_widths[376]), .rectangle3_height(rectangle3_heights[376]), .rectangle3_weight(rectangle3_weights[376]), .feature_threshold(feature_thresholds[376]), .feature_above(feature_aboves[376]), .feature_below(feature_belows[376]), .scan_win_std_dev(scan_win_std_dev[376]), .feature_accum(feature_accums[376]));
  accum_calculator ac377(.scan_win(scan_win377), .rectangle1_x(rectangle1_xs[377]), .rectangle1_y(rectangle1_ys[377]), .rectangle1_width(rectangle1_widths[377]), .rectangle1_height(rectangle1_heights[377]), .rectangle1_weight(rectangle1_weights[377]), .rectangle2_x(rectangle2_xs[377]), .rectangle2_y(rectangle2_ys[377]), .rectangle2_width(rectangle2_widths[377]), .rectangle2_height(rectangle2_heights[377]), .rectangle2_weight(rectangle2_weights[377]), .rectangle3_x(rectangle3_xs[377]), .rectangle3_y(rectangle3_ys[377]), .rectangle3_width(rectangle3_widths[377]), .rectangle3_height(rectangle3_heights[377]), .rectangle3_weight(rectangle3_weights[377]), .feature_threshold(feature_thresholds[377]), .feature_above(feature_aboves[377]), .feature_below(feature_belows[377]), .scan_win_std_dev(scan_win_std_dev[377]), .feature_accum(feature_accums[377]));
  accum_calculator ac378(.scan_win(scan_win378), .rectangle1_x(rectangle1_xs[378]), .rectangle1_y(rectangle1_ys[378]), .rectangle1_width(rectangle1_widths[378]), .rectangle1_height(rectangle1_heights[378]), .rectangle1_weight(rectangle1_weights[378]), .rectangle2_x(rectangle2_xs[378]), .rectangle2_y(rectangle2_ys[378]), .rectangle2_width(rectangle2_widths[378]), .rectangle2_height(rectangle2_heights[378]), .rectangle2_weight(rectangle2_weights[378]), .rectangle3_x(rectangle3_xs[378]), .rectangle3_y(rectangle3_ys[378]), .rectangle3_width(rectangle3_widths[378]), .rectangle3_height(rectangle3_heights[378]), .rectangle3_weight(rectangle3_weights[378]), .feature_threshold(feature_thresholds[378]), .feature_above(feature_aboves[378]), .feature_below(feature_belows[378]), .scan_win_std_dev(scan_win_std_dev[378]), .feature_accum(feature_accums[378]));
  accum_calculator ac379(.scan_win(scan_win379), .rectangle1_x(rectangle1_xs[379]), .rectangle1_y(rectangle1_ys[379]), .rectangle1_width(rectangle1_widths[379]), .rectangle1_height(rectangle1_heights[379]), .rectangle1_weight(rectangle1_weights[379]), .rectangle2_x(rectangle2_xs[379]), .rectangle2_y(rectangle2_ys[379]), .rectangle2_width(rectangle2_widths[379]), .rectangle2_height(rectangle2_heights[379]), .rectangle2_weight(rectangle2_weights[379]), .rectangle3_x(rectangle3_xs[379]), .rectangle3_y(rectangle3_ys[379]), .rectangle3_width(rectangle3_widths[379]), .rectangle3_height(rectangle3_heights[379]), .rectangle3_weight(rectangle3_weights[379]), .feature_threshold(feature_thresholds[379]), .feature_above(feature_aboves[379]), .feature_below(feature_belows[379]), .scan_win_std_dev(scan_win_std_dev[379]), .feature_accum(feature_accums[379]));
  accum_calculator ac380(.scan_win(scan_win380), .rectangle1_x(rectangle1_xs[380]), .rectangle1_y(rectangle1_ys[380]), .rectangle1_width(rectangle1_widths[380]), .rectangle1_height(rectangle1_heights[380]), .rectangle1_weight(rectangle1_weights[380]), .rectangle2_x(rectangle2_xs[380]), .rectangle2_y(rectangle2_ys[380]), .rectangle2_width(rectangle2_widths[380]), .rectangle2_height(rectangle2_heights[380]), .rectangle2_weight(rectangle2_weights[380]), .rectangle3_x(rectangle3_xs[380]), .rectangle3_y(rectangle3_ys[380]), .rectangle3_width(rectangle3_widths[380]), .rectangle3_height(rectangle3_heights[380]), .rectangle3_weight(rectangle3_weights[380]), .feature_threshold(feature_thresholds[380]), .feature_above(feature_aboves[380]), .feature_below(feature_belows[380]), .scan_win_std_dev(scan_win_std_dev[380]), .feature_accum(feature_accums[380]));
  accum_calculator ac381(.scan_win(scan_win381), .rectangle1_x(rectangle1_xs[381]), .rectangle1_y(rectangle1_ys[381]), .rectangle1_width(rectangle1_widths[381]), .rectangle1_height(rectangle1_heights[381]), .rectangle1_weight(rectangle1_weights[381]), .rectangle2_x(rectangle2_xs[381]), .rectangle2_y(rectangle2_ys[381]), .rectangle2_width(rectangle2_widths[381]), .rectangle2_height(rectangle2_heights[381]), .rectangle2_weight(rectangle2_weights[381]), .rectangle3_x(rectangle3_xs[381]), .rectangle3_y(rectangle3_ys[381]), .rectangle3_width(rectangle3_widths[381]), .rectangle3_height(rectangle3_heights[381]), .rectangle3_weight(rectangle3_weights[381]), .feature_threshold(feature_thresholds[381]), .feature_above(feature_aboves[381]), .feature_below(feature_belows[381]), .scan_win_std_dev(scan_win_std_dev[381]), .feature_accum(feature_accums[381]));
  accum_calculator ac382(.scan_win(scan_win382), .rectangle1_x(rectangle1_xs[382]), .rectangle1_y(rectangle1_ys[382]), .rectangle1_width(rectangle1_widths[382]), .rectangle1_height(rectangle1_heights[382]), .rectangle1_weight(rectangle1_weights[382]), .rectangle2_x(rectangle2_xs[382]), .rectangle2_y(rectangle2_ys[382]), .rectangle2_width(rectangle2_widths[382]), .rectangle2_height(rectangle2_heights[382]), .rectangle2_weight(rectangle2_weights[382]), .rectangle3_x(rectangle3_xs[382]), .rectangle3_y(rectangle3_ys[382]), .rectangle3_width(rectangle3_widths[382]), .rectangle3_height(rectangle3_heights[382]), .rectangle3_weight(rectangle3_weights[382]), .feature_threshold(feature_thresholds[382]), .feature_above(feature_aboves[382]), .feature_below(feature_belows[382]), .scan_win_std_dev(scan_win_std_dev[382]), .feature_accum(feature_accums[382]));
  accum_calculator ac383(.scan_win(scan_win383), .rectangle1_x(rectangle1_xs[383]), .rectangle1_y(rectangle1_ys[383]), .rectangle1_width(rectangle1_widths[383]), .rectangle1_height(rectangle1_heights[383]), .rectangle1_weight(rectangle1_weights[383]), .rectangle2_x(rectangle2_xs[383]), .rectangle2_y(rectangle2_ys[383]), .rectangle2_width(rectangle2_widths[383]), .rectangle2_height(rectangle2_heights[383]), .rectangle2_weight(rectangle2_weights[383]), .rectangle3_x(rectangle3_xs[383]), .rectangle3_y(rectangle3_ys[383]), .rectangle3_width(rectangle3_widths[383]), .rectangle3_height(rectangle3_heights[383]), .rectangle3_weight(rectangle3_weights[383]), .feature_threshold(feature_thresholds[383]), .feature_above(feature_aboves[383]), .feature_below(feature_belows[383]), .scan_win_std_dev(scan_win_std_dev[383]), .feature_accum(feature_accums[383]));
  accum_calculator ac384(.scan_win(scan_win384), .rectangle1_x(rectangle1_xs[384]), .rectangle1_y(rectangle1_ys[384]), .rectangle1_width(rectangle1_widths[384]), .rectangle1_height(rectangle1_heights[384]), .rectangle1_weight(rectangle1_weights[384]), .rectangle2_x(rectangle2_xs[384]), .rectangle2_y(rectangle2_ys[384]), .rectangle2_width(rectangle2_widths[384]), .rectangle2_height(rectangle2_heights[384]), .rectangle2_weight(rectangle2_weights[384]), .rectangle3_x(rectangle3_xs[384]), .rectangle3_y(rectangle3_ys[384]), .rectangle3_width(rectangle3_widths[384]), .rectangle3_height(rectangle3_heights[384]), .rectangle3_weight(rectangle3_weights[384]), .feature_threshold(feature_thresholds[384]), .feature_above(feature_aboves[384]), .feature_below(feature_belows[384]), .scan_win_std_dev(scan_win_std_dev[384]), .feature_accum(feature_accums[384]));
  accum_calculator ac385(.scan_win(scan_win385), .rectangle1_x(rectangle1_xs[385]), .rectangle1_y(rectangle1_ys[385]), .rectangle1_width(rectangle1_widths[385]), .rectangle1_height(rectangle1_heights[385]), .rectangle1_weight(rectangle1_weights[385]), .rectangle2_x(rectangle2_xs[385]), .rectangle2_y(rectangle2_ys[385]), .rectangle2_width(rectangle2_widths[385]), .rectangle2_height(rectangle2_heights[385]), .rectangle2_weight(rectangle2_weights[385]), .rectangle3_x(rectangle3_xs[385]), .rectangle3_y(rectangle3_ys[385]), .rectangle3_width(rectangle3_widths[385]), .rectangle3_height(rectangle3_heights[385]), .rectangle3_weight(rectangle3_weights[385]), .feature_threshold(feature_thresholds[385]), .feature_above(feature_aboves[385]), .feature_below(feature_belows[385]), .scan_win_std_dev(scan_win_std_dev[385]), .feature_accum(feature_accums[385]));
  accum_calculator ac386(.scan_win(scan_win386), .rectangle1_x(rectangle1_xs[386]), .rectangle1_y(rectangle1_ys[386]), .rectangle1_width(rectangle1_widths[386]), .rectangle1_height(rectangle1_heights[386]), .rectangle1_weight(rectangle1_weights[386]), .rectangle2_x(rectangle2_xs[386]), .rectangle2_y(rectangle2_ys[386]), .rectangle2_width(rectangle2_widths[386]), .rectangle2_height(rectangle2_heights[386]), .rectangle2_weight(rectangle2_weights[386]), .rectangle3_x(rectangle3_xs[386]), .rectangle3_y(rectangle3_ys[386]), .rectangle3_width(rectangle3_widths[386]), .rectangle3_height(rectangle3_heights[386]), .rectangle3_weight(rectangle3_weights[386]), .feature_threshold(feature_thresholds[386]), .feature_above(feature_aboves[386]), .feature_below(feature_belows[386]), .scan_win_std_dev(scan_win_std_dev[386]), .feature_accum(feature_accums[386]));
  accum_calculator ac387(.scan_win(scan_win387), .rectangle1_x(rectangle1_xs[387]), .rectangle1_y(rectangle1_ys[387]), .rectangle1_width(rectangle1_widths[387]), .rectangle1_height(rectangle1_heights[387]), .rectangle1_weight(rectangle1_weights[387]), .rectangle2_x(rectangle2_xs[387]), .rectangle2_y(rectangle2_ys[387]), .rectangle2_width(rectangle2_widths[387]), .rectangle2_height(rectangle2_heights[387]), .rectangle2_weight(rectangle2_weights[387]), .rectangle3_x(rectangle3_xs[387]), .rectangle3_y(rectangle3_ys[387]), .rectangle3_width(rectangle3_widths[387]), .rectangle3_height(rectangle3_heights[387]), .rectangle3_weight(rectangle3_weights[387]), .feature_threshold(feature_thresholds[387]), .feature_above(feature_aboves[387]), .feature_below(feature_belows[387]), .scan_win_std_dev(scan_win_std_dev[387]), .feature_accum(feature_accums[387]));
  accum_calculator ac388(.scan_win(scan_win388), .rectangle1_x(rectangle1_xs[388]), .rectangle1_y(rectangle1_ys[388]), .rectangle1_width(rectangle1_widths[388]), .rectangle1_height(rectangle1_heights[388]), .rectangle1_weight(rectangle1_weights[388]), .rectangle2_x(rectangle2_xs[388]), .rectangle2_y(rectangle2_ys[388]), .rectangle2_width(rectangle2_widths[388]), .rectangle2_height(rectangle2_heights[388]), .rectangle2_weight(rectangle2_weights[388]), .rectangle3_x(rectangle3_xs[388]), .rectangle3_y(rectangle3_ys[388]), .rectangle3_width(rectangle3_widths[388]), .rectangle3_height(rectangle3_heights[388]), .rectangle3_weight(rectangle3_weights[388]), .feature_threshold(feature_thresholds[388]), .feature_above(feature_aboves[388]), .feature_below(feature_belows[388]), .scan_win_std_dev(scan_win_std_dev[388]), .feature_accum(feature_accums[388]));
  accum_calculator ac389(.scan_win(scan_win389), .rectangle1_x(rectangle1_xs[389]), .rectangle1_y(rectangle1_ys[389]), .rectangle1_width(rectangle1_widths[389]), .rectangle1_height(rectangle1_heights[389]), .rectangle1_weight(rectangle1_weights[389]), .rectangle2_x(rectangle2_xs[389]), .rectangle2_y(rectangle2_ys[389]), .rectangle2_width(rectangle2_widths[389]), .rectangle2_height(rectangle2_heights[389]), .rectangle2_weight(rectangle2_weights[389]), .rectangle3_x(rectangle3_xs[389]), .rectangle3_y(rectangle3_ys[389]), .rectangle3_width(rectangle3_widths[389]), .rectangle3_height(rectangle3_heights[389]), .rectangle3_weight(rectangle3_weights[389]), .feature_threshold(feature_thresholds[389]), .feature_above(feature_aboves[389]), .feature_below(feature_belows[389]), .scan_win_std_dev(scan_win_std_dev[389]), .feature_accum(feature_accums[389]));
  accum_calculator ac390(.scan_win(scan_win390), .rectangle1_x(rectangle1_xs[390]), .rectangle1_y(rectangle1_ys[390]), .rectangle1_width(rectangle1_widths[390]), .rectangle1_height(rectangle1_heights[390]), .rectangle1_weight(rectangle1_weights[390]), .rectangle2_x(rectangle2_xs[390]), .rectangle2_y(rectangle2_ys[390]), .rectangle2_width(rectangle2_widths[390]), .rectangle2_height(rectangle2_heights[390]), .rectangle2_weight(rectangle2_weights[390]), .rectangle3_x(rectangle3_xs[390]), .rectangle3_y(rectangle3_ys[390]), .rectangle3_width(rectangle3_widths[390]), .rectangle3_height(rectangle3_heights[390]), .rectangle3_weight(rectangle3_weights[390]), .feature_threshold(feature_thresholds[390]), .feature_above(feature_aboves[390]), .feature_below(feature_belows[390]), .scan_win_std_dev(scan_win_std_dev[390]), .feature_accum(feature_accums[390]));
  accum_calculator ac391(.scan_win(scan_win391), .rectangle1_x(rectangle1_xs[391]), .rectangle1_y(rectangle1_ys[391]), .rectangle1_width(rectangle1_widths[391]), .rectangle1_height(rectangle1_heights[391]), .rectangle1_weight(rectangle1_weights[391]), .rectangle2_x(rectangle2_xs[391]), .rectangle2_y(rectangle2_ys[391]), .rectangle2_width(rectangle2_widths[391]), .rectangle2_height(rectangle2_heights[391]), .rectangle2_weight(rectangle2_weights[391]), .rectangle3_x(rectangle3_xs[391]), .rectangle3_y(rectangle3_ys[391]), .rectangle3_width(rectangle3_widths[391]), .rectangle3_height(rectangle3_heights[391]), .rectangle3_weight(rectangle3_weights[391]), .feature_threshold(feature_thresholds[391]), .feature_above(feature_aboves[391]), .feature_below(feature_belows[391]), .scan_win_std_dev(scan_win_std_dev[391]), .feature_accum(feature_accums[391]));
  accum_calculator ac392(.scan_win(scan_win392), .rectangle1_x(rectangle1_xs[392]), .rectangle1_y(rectangle1_ys[392]), .rectangle1_width(rectangle1_widths[392]), .rectangle1_height(rectangle1_heights[392]), .rectangle1_weight(rectangle1_weights[392]), .rectangle2_x(rectangle2_xs[392]), .rectangle2_y(rectangle2_ys[392]), .rectangle2_width(rectangle2_widths[392]), .rectangle2_height(rectangle2_heights[392]), .rectangle2_weight(rectangle2_weights[392]), .rectangle3_x(rectangle3_xs[392]), .rectangle3_y(rectangle3_ys[392]), .rectangle3_width(rectangle3_widths[392]), .rectangle3_height(rectangle3_heights[392]), .rectangle3_weight(rectangle3_weights[392]), .feature_threshold(feature_thresholds[392]), .feature_above(feature_aboves[392]), .feature_below(feature_belows[392]), .scan_win_std_dev(scan_win_std_dev[392]), .feature_accum(feature_accums[392]));
  accum_calculator ac393(.scan_win(scan_win393), .rectangle1_x(rectangle1_xs[393]), .rectangle1_y(rectangle1_ys[393]), .rectangle1_width(rectangle1_widths[393]), .rectangle1_height(rectangle1_heights[393]), .rectangle1_weight(rectangle1_weights[393]), .rectangle2_x(rectangle2_xs[393]), .rectangle2_y(rectangle2_ys[393]), .rectangle2_width(rectangle2_widths[393]), .rectangle2_height(rectangle2_heights[393]), .rectangle2_weight(rectangle2_weights[393]), .rectangle3_x(rectangle3_xs[393]), .rectangle3_y(rectangle3_ys[393]), .rectangle3_width(rectangle3_widths[393]), .rectangle3_height(rectangle3_heights[393]), .rectangle3_weight(rectangle3_weights[393]), .feature_threshold(feature_thresholds[393]), .feature_above(feature_aboves[393]), .feature_below(feature_belows[393]), .scan_win_std_dev(scan_win_std_dev[393]), .feature_accum(feature_accums[393]));
  accum_calculator ac394(.scan_win(scan_win394), .rectangle1_x(rectangle1_xs[394]), .rectangle1_y(rectangle1_ys[394]), .rectangle1_width(rectangle1_widths[394]), .rectangle1_height(rectangle1_heights[394]), .rectangle1_weight(rectangle1_weights[394]), .rectangle2_x(rectangle2_xs[394]), .rectangle2_y(rectangle2_ys[394]), .rectangle2_width(rectangle2_widths[394]), .rectangle2_height(rectangle2_heights[394]), .rectangle2_weight(rectangle2_weights[394]), .rectangle3_x(rectangle3_xs[394]), .rectangle3_y(rectangle3_ys[394]), .rectangle3_width(rectangle3_widths[394]), .rectangle3_height(rectangle3_heights[394]), .rectangle3_weight(rectangle3_weights[394]), .feature_threshold(feature_thresholds[394]), .feature_above(feature_aboves[394]), .feature_below(feature_belows[394]), .scan_win_std_dev(scan_win_std_dev[394]), .feature_accum(feature_accums[394]));
  accum_calculator ac395(.scan_win(scan_win395), .rectangle1_x(rectangle1_xs[395]), .rectangle1_y(rectangle1_ys[395]), .rectangle1_width(rectangle1_widths[395]), .rectangle1_height(rectangle1_heights[395]), .rectangle1_weight(rectangle1_weights[395]), .rectangle2_x(rectangle2_xs[395]), .rectangle2_y(rectangle2_ys[395]), .rectangle2_width(rectangle2_widths[395]), .rectangle2_height(rectangle2_heights[395]), .rectangle2_weight(rectangle2_weights[395]), .rectangle3_x(rectangle3_xs[395]), .rectangle3_y(rectangle3_ys[395]), .rectangle3_width(rectangle3_widths[395]), .rectangle3_height(rectangle3_heights[395]), .rectangle3_weight(rectangle3_weights[395]), .feature_threshold(feature_thresholds[395]), .feature_above(feature_aboves[395]), .feature_below(feature_belows[395]), .scan_win_std_dev(scan_win_std_dev[395]), .feature_accum(feature_accums[395]));
  accum_calculator ac396(.scan_win(scan_win396), .rectangle1_x(rectangle1_xs[396]), .rectangle1_y(rectangle1_ys[396]), .rectangle1_width(rectangle1_widths[396]), .rectangle1_height(rectangle1_heights[396]), .rectangle1_weight(rectangle1_weights[396]), .rectangle2_x(rectangle2_xs[396]), .rectangle2_y(rectangle2_ys[396]), .rectangle2_width(rectangle2_widths[396]), .rectangle2_height(rectangle2_heights[396]), .rectangle2_weight(rectangle2_weights[396]), .rectangle3_x(rectangle3_xs[396]), .rectangle3_y(rectangle3_ys[396]), .rectangle3_width(rectangle3_widths[396]), .rectangle3_height(rectangle3_heights[396]), .rectangle3_weight(rectangle3_weights[396]), .feature_threshold(feature_thresholds[396]), .feature_above(feature_aboves[396]), .feature_below(feature_belows[396]), .scan_win_std_dev(scan_win_std_dev[396]), .feature_accum(feature_accums[396]));
  accum_calculator ac397(.scan_win(scan_win397), .rectangle1_x(rectangle1_xs[397]), .rectangle1_y(rectangle1_ys[397]), .rectangle1_width(rectangle1_widths[397]), .rectangle1_height(rectangle1_heights[397]), .rectangle1_weight(rectangle1_weights[397]), .rectangle2_x(rectangle2_xs[397]), .rectangle2_y(rectangle2_ys[397]), .rectangle2_width(rectangle2_widths[397]), .rectangle2_height(rectangle2_heights[397]), .rectangle2_weight(rectangle2_weights[397]), .rectangle3_x(rectangle3_xs[397]), .rectangle3_y(rectangle3_ys[397]), .rectangle3_width(rectangle3_widths[397]), .rectangle3_height(rectangle3_heights[397]), .rectangle3_weight(rectangle3_weights[397]), .feature_threshold(feature_thresholds[397]), .feature_above(feature_aboves[397]), .feature_below(feature_belows[397]), .scan_win_std_dev(scan_win_std_dev[397]), .feature_accum(feature_accums[397]));
  accum_calculator ac398(.scan_win(scan_win398), .rectangle1_x(rectangle1_xs[398]), .rectangle1_y(rectangle1_ys[398]), .rectangle1_width(rectangle1_widths[398]), .rectangle1_height(rectangle1_heights[398]), .rectangle1_weight(rectangle1_weights[398]), .rectangle2_x(rectangle2_xs[398]), .rectangle2_y(rectangle2_ys[398]), .rectangle2_width(rectangle2_widths[398]), .rectangle2_height(rectangle2_heights[398]), .rectangle2_weight(rectangle2_weights[398]), .rectangle3_x(rectangle3_xs[398]), .rectangle3_y(rectangle3_ys[398]), .rectangle3_width(rectangle3_widths[398]), .rectangle3_height(rectangle3_heights[398]), .rectangle3_weight(rectangle3_weights[398]), .feature_threshold(feature_thresholds[398]), .feature_above(feature_aboves[398]), .feature_below(feature_belows[398]), .scan_win_std_dev(scan_win_std_dev[398]), .feature_accum(feature_accums[398]));
  accum_calculator ac399(.scan_win(scan_win399), .rectangle1_x(rectangle1_xs[399]), .rectangle1_y(rectangle1_ys[399]), .rectangle1_width(rectangle1_widths[399]), .rectangle1_height(rectangle1_heights[399]), .rectangle1_weight(rectangle1_weights[399]), .rectangle2_x(rectangle2_xs[399]), .rectangle2_y(rectangle2_ys[399]), .rectangle2_width(rectangle2_widths[399]), .rectangle2_height(rectangle2_heights[399]), .rectangle2_weight(rectangle2_weights[399]), .rectangle3_x(rectangle3_xs[399]), .rectangle3_y(rectangle3_ys[399]), .rectangle3_width(rectangle3_widths[399]), .rectangle3_height(rectangle3_heights[399]), .rectangle3_weight(rectangle3_weights[399]), .feature_threshold(feature_thresholds[399]), .feature_above(feature_aboves[399]), .feature_below(feature_belows[399]), .scan_win_std_dev(scan_win_std_dev[399]), .feature_accum(feature_accums[399]));
  accum_calculator ac400(.scan_win(scan_win400), .rectangle1_x(rectangle1_xs[400]), .rectangle1_y(rectangle1_ys[400]), .rectangle1_width(rectangle1_widths[400]), .rectangle1_height(rectangle1_heights[400]), .rectangle1_weight(rectangle1_weights[400]), .rectangle2_x(rectangle2_xs[400]), .rectangle2_y(rectangle2_ys[400]), .rectangle2_width(rectangle2_widths[400]), .rectangle2_height(rectangle2_heights[400]), .rectangle2_weight(rectangle2_weights[400]), .rectangle3_x(rectangle3_xs[400]), .rectangle3_y(rectangle3_ys[400]), .rectangle3_width(rectangle3_widths[400]), .rectangle3_height(rectangle3_heights[400]), .rectangle3_weight(rectangle3_weights[400]), .feature_threshold(feature_thresholds[400]), .feature_above(feature_aboves[400]), .feature_below(feature_belows[400]), .scan_win_std_dev(scan_win_std_dev[400]), .feature_accum(feature_accums[400]));
  accum_calculator ac401(.scan_win(scan_win401), .rectangle1_x(rectangle1_xs[401]), .rectangle1_y(rectangle1_ys[401]), .rectangle1_width(rectangle1_widths[401]), .rectangle1_height(rectangle1_heights[401]), .rectangle1_weight(rectangle1_weights[401]), .rectangle2_x(rectangle2_xs[401]), .rectangle2_y(rectangle2_ys[401]), .rectangle2_width(rectangle2_widths[401]), .rectangle2_height(rectangle2_heights[401]), .rectangle2_weight(rectangle2_weights[401]), .rectangle3_x(rectangle3_xs[401]), .rectangle3_y(rectangle3_ys[401]), .rectangle3_width(rectangle3_widths[401]), .rectangle3_height(rectangle3_heights[401]), .rectangle3_weight(rectangle3_weights[401]), .feature_threshold(feature_thresholds[401]), .feature_above(feature_aboves[401]), .feature_below(feature_belows[401]), .scan_win_std_dev(scan_win_std_dev[401]), .feature_accum(feature_accums[401]));
  accum_calculator ac402(.scan_win(scan_win402), .rectangle1_x(rectangle1_xs[402]), .rectangle1_y(rectangle1_ys[402]), .rectangle1_width(rectangle1_widths[402]), .rectangle1_height(rectangle1_heights[402]), .rectangle1_weight(rectangle1_weights[402]), .rectangle2_x(rectangle2_xs[402]), .rectangle2_y(rectangle2_ys[402]), .rectangle2_width(rectangle2_widths[402]), .rectangle2_height(rectangle2_heights[402]), .rectangle2_weight(rectangle2_weights[402]), .rectangle3_x(rectangle3_xs[402]), .rectangle3_y(rectangle3_ys[402]), .rectangle3_width(rectangle3_widths[402]), .rectangle3_height(rectangle3_heights[402]), .rectangle3_weight(rectangle3_weights[402]), .feature_threshold(feature_thresholds[402]), .feature_above(feature_aboves[402]), .feature_below(feature_belows[402]), .scan_win_std_dev(scan_win_std_dev[402]), .feature_accum(feature_accums[402]));
  accum_calculator ac403(.scan_win(scan_win403), .rectangle1_x(rectangle1_xs[403]), .rectangle1_y(rectangle1_ys[403]), .rectangle1_width(rectangle1_widths[403]), .rectangle1_height(rectangle1_heights[403]), .rectangle1_weight(rectangle1_weights[403]), .rectangle2_x(rectangle2_xs[403]), .rectangle2_y(rectangle2_ys[403]), .rectangle2_width(rectangle2_widths[403]), .rectangle2_height(rectangle2_heights[403]), .rectangle2_weight(rectangle2_weights[403]), .rectangle3_x(rectangle3_xs[403]), .rectangle3_y(rectangle3_ys[403]), .rectangle3_width(rectangle3_widths[403]), .rectangle3_height(rectangle3_heights[403]), .rectangle3_weight(rectangle3_weights[403]), .feature_threshold(feature_thresholds[403]), .feature_above(feature_aboves[403]), .feature_below(feature_belows[403]), .scan_win_std_dev(scan_win_std_dev[403]), .feature_accum(feature_accums[403]));
  accum_calculator ac404(.scan_win(scan_win404), .rectangle1_x(rectangle1_xs[404]), .rectangle1_y(rectangle1_ys[404]), .rectangle1_width(rectangle1_widths[404]), .rectangle1_height(rectangle1_heights[404]), .rectangle1_weight(rectangle1_weights[404]), .rectangle2_x(rectangle2_xs[404]), .rectangle2_y(rectangle2_ys[404]), .rectangle2_width(rectangle2_widths[404]), .rectangle2_height(rectangle2_heights[404]), .rectangle2_weight(rectangle2_weights[404]), .rectangle3_x(rectangle3_xs[404]), .rectangle3_y(rectangle3_ys[404]), .rectangle3_width(rectangle3_widths[404]), .rectangle3_height(rectangle3_heights[404]), .rectangle3_weight(rectangle3_weights[404]), .feature_threshold(feature_thresholds[404]), .feature_above(feature_aboves[404]), .feature_below(feature_belows[404]), .scan_win_std_dev(scan_win_std_dev[404]), .feature_accum(feature_accums[404]));
  accum_calculator ac405(.scan_win(scan_win405), .rectangle1_x(rectangle1_xs[405]), .rectangle1_y(rectangle1_ys[405]), .rectangle1_width(rectangle1_widths[405]), .rectangle1_height(rectangle1_heights[405]), .rectangle1_weight(rectangle1_weights[405]), .rectangle2_x(rectangle2_xs[405]), .rectangle2_y(rectangle2_ys[405]), .rectangle2_width(rectangle2_widths[405]), .rectangle2_height(rectangle2_heights[405]), .rectangle2_weight(rectangle2_weights[405]), .rectangle3_x(rectangle3_xs[405]), .rectangle3_y(rectangle3_ys[405]), .rectangle3_width(rectangle3_widths[405]), .rectangle3_height(rectangle3_heights[405]), .rectangle3_weight(rectangle3_weights[405]), .feature_threshold(feature_thresholds[405]), .feature_above(feature_aboves[405]), .feature_below(feature_belows[405]), .scan_win_std_dev(scan_win_std_dev[405]), .feature_accum(feature_accums[405]));
  accum_calculator ac406(.scan_win(scan_win406), .rectangle1_x(rectangle1_xs[406]), .rectangle1_y(rectangle1_ys[406]), .rectangle1_width(rectangle1_widths[406]), .rectangle1_height(rectangle1_heights[406]), .rectangle1_weight(rectangle1_weights[406]), .rectangle2_x(rectangle2_xs[406]), .rectangle2_y(rectangle2_ys[406]), .rectangle2_width(rectangle2_widths[406]), .rectangle2_height(rectangle2_heights[406]), .rectangle2_weight(rectangle2_weights[406]), .rectangle3_x(rectangle3_xs[406]), .rectangle3_y(rectangle3_ys[406]), .rectangle3_width(rectangle3_widths[406]), .rectangle3_height(rectangle3_heights[406]), .rectangle3_weight(rectangle3_weights[406]), .feature_threshold(feature_thresholds[406]), .feature_above(feature_aboves[406]), .feature_below(feature_belows[406]), .scan_win_std_dev(scan_win_std_dev[406]), .feature_accum(feature_accums[406]));
  accum_calculator ac407(.scan_win(scan_win407), .rectangle1_x(rectangle1_xs[407]), .rectangle1_y(rectangle1_ys[407]), .rectangle1_width(rectangle1_widths[407]), .rectangle1_height(rectangle1_heights[407]), .rectangle1_weight(rectangle1_weights[407]), .rectangle2_x(rectangle2_xs[407]), .rectangle2_y(rectangle2_ys[407]), .rectangle2_width(rectangle2_widths[407]), .rectangle2_height(rectangle2_heights[407]), .rectangle2_weight(rectangle2_weights[407]), .rectangle3_x(rectangle3_xs[407]), .rectangle3_y(rectangle3_ys[407]), .rectangle3_width(rectangle3_widths[407]), .rectangle3_height(rectangle3_heights[407]), .rectangle3_weight(rectangle3_weights[407]), .feature_threshold(feature_thresholds[407]), .feature_above(feature_aboves[407]), .feature_below(feature_belows[407]), .scan_win_std_dev(scan_win_std_dev[407]), .feature_accum(feature_accums[407]));
  accum_calculator ac408(.scan_win(scan_win408), .rectangle1_x(rectangle1_xs[408]), .rectangle1_y(rectangle1_ys[408]), .rectangle1_width(rectangle1_widths[408]), .rectangle1_height(rectangle1_heights[408]), .rectangle1_weight(rectangle1_weights[408]), .rectangle2_x(rectangle2_xs[408]), .rectangle2_y(rectangle2_ys[408]), .rectangle2_width(rectangle2_widths[408]), .rectangle2_height(rectangle2_heights[408]), .rectangle2_weight(rectangle2_weights[408]), .rectangle3_x(rectangle3_xs[408]), .rectangle3_y(rectangle3_ys[408]), .rectangle3_width(rectangle3_widths[408]), .rectangle3_height(rectangle3_heights[408]), .rectangle3_weight(rectangle3_weights[408]), .feature_threshold(feature_thresholds[408]), .feature_above(feature_aboves[408]), .feature_below(feature_belows[408]), .scan_win_std_dev(scan_win_std_dev[408]), .feature_accum(feature_accums[408]));
  accum_calculator ac409(.scan_win(scan_win409), .rectangle1_x(rectangle1_xs[409]), .rectangle1_y(rectangle1_ys[409]), .rectangle1_width(rectangle1_widths[409]), .rectangle1_height(rectangle1_heights[409]), .rectangle1_weight(rectangle1_weights[409]), .rectangle2_x(rectangle2_xs[409]), .rectangle2_y(rectangle2_ys[409]), .rectangle2_width(rectangle2_widths[409]), .rectangle2_height(rectangle2_heights[409]), .rectangle2_weight(rectangle2_weights[409]), .rectangle3_x(rectangle3_xs[409]), .rectangle3_y(rectangle3_ys[409]), .rectangle3_width(rectangle3_widths[409]), .rectangle3_height(rectangle3_heights[409]), .rectangle3_weight(rectangle3_weights[409]), .feature_threshold(feature_thresholds[409]), .feature_above(feature_aboves[409]), .feature_below(feature_belows[409]), .scan_win_std_dev(scan_win_std_dev[409]), .feature_accum(feature_accums[409]));
  accum_calculator ac410(.scan_win(scan_win410), .rectangle1_x(rectangle1_xs[410]), .rectangle1_y(rectangle1_ys[410]), .rectangle1_width(rectangle1_widths[410]), .rectangle1_height(rectangle1_heights[410]), .rectangle1_weight(rectangle1_weights[410]), .rectangle2_x(rectangle2_xs[410]), .rectangle2_y(rectangle2_ys[410]), .rectangle2_width(rectangle2_widths[410]), .rectangle2_height(rectangle2_heights[410]), .rectangle2_weight(rectangle2_weights[410]), .rectangle3_x(rectangle3_xs[410]), .rectangle3_y(rectangle3_ys[410]), .rectangle3_width(rectangle3_widths[410]), .rectangle3_height(rectangle3_heights[410]), .rectangle3_weight(rectangle3_weights[410]), .feature_threshold(feature_thresholds[410]), .feature_above(feature_aboves[410]), .feature_below(feature_belows[410]), .scan_win_std_dev(scan_win_std_dev[410]), .feature_accum(feature_accums[410]));
  accum_calculator ac411(.scan_win(scan_win411), .rectangle1_x(rectangle1_xs[411]), .rectangle1_y(rectangle1_ys[411]), .rectangle1_width(rectangle1_widths[411]), .rectangle1_height(rectangle1_heights[411]), .rectangle1_weight(rectangle1_weights[411]), .rectangle2_x(rectangle2_xs[411]), .rectangle2_y(rectangle2_ys[411]), .rectangle2_width(rectangle2_widths[411]), .rectangle2_height(rectangle2_heights[411]), .rectangle2_weight(rectangle2_weights[411]), .rectangle3_x(rectangle3_xs[411]), .rectangle3_y(rectangle3_ys[411]), .rectangle3_width(rectangle3_widths[411]), .rectangle3_height(rectangle3_heights[411]), .rectangle3_weight(rectangle3_weights[411]), .feature_threshold(feature_thresholds[411]), .feature_above(feature_aboves[411]), .feature_below(feature_belows[411]), .scan_win_std_dev(scan_win_std_dev[411]), .feature_accum(feature_accums[411]));
  accum_calculator ac412(.scan_win(scan_win412), .rectangle1_x(rectangle1_xs[412]), .rectangle1_y(rectangle1_ys[412]), .rectangle1_width(rectangle1_widths[412]), .rectangle1_height(rectangle1_heights[412]), .rectangle1_weight(rectangle1_weights[412]), .rectangle2_x(rectangle2_xs[412]), .rectangle2_y(rectangle2_ys[412]), .rectangle2_width(rectangle2_widths[412]), .rectangle2_height(rectangle2_heights[412]), .rectangle2_weight(rectangle2_weights[412]), .rectangle3_x(rectangle3_xs[412]), .rectangle3_y(rectangle3_ys[412]), .rectangle3_width(rectangle3_widths[412]), .rectangle3_height(rectangle3_heights[412]), .rectangle3_weight(rectangle3_weights[412]), .feature_threshold(feature_thresholds[412]), .feature_above(feature_aboves[412]), .feature_below(feature_belows[412]), .scan_win_std_dev(scan_win_std_dev[412]), .feature_accum(feature_accums[412]));
  accum_calculator ac413(.scan_win(scan_win413), .rectangle1_x(rectangle1_xs[413]), .rectangle1_y(rectangle1_ys[413]), .rectangle1_width(rectangle1_widths[413]), .rectangle1_height(rectangle1_heights[413]), .rectangle1_weight(rectangle1_weights[413]), .rectangle2_x(rectangle2_xs[413]), .rectangle2_y(rectangle2_ys[413]), .rectangle2_width(rectangle2_widths[413]), .rectangle2_height(rectangle2_heights[413]), .rectangle2_weight(rectangle2_weights[413]), .rectangle3_x(rectangle3_xs[413]), .rectangle3_y(rectangle3_ys[413]), .rectangle3_width(rectangle3_widths[413]), .rectangle3_height(rectangle3_heights[413]), .rectangle3_weight(rectangle3_weights[413]), .feature_threshold(feature_thresholds[413]), .feature_above(feature_aboves[413]), .feature_below(feature_belows[413]), .scan_win_std_dev(scan_win_std_dev[413]), .feature_accum(feature_accums[413]));
  accum_calculator ac414(.scan_win(scan_win414), .rectangle1_x(rectangle1_xs[414]), .rectangle1_y(rectangle1_ys[414]), .rectangle1_width(rectangle1_widths[414]), .rectangle1_height(rectangle1_heights[414]), .rectangle1_weight(rectangle1_weights[414]), .rectangle2_x(rectangle2_xs[414]), .rectangle2_y(rectangle2_ys[414]), .rectangle2_width(rectangle2_widths[414]), .rectangle2_height(rectangle2_heights[414]), .rectangle2_weight(rectangle2_weights[414]), .rectangle3_x(rectangle3_xs[414]), .rectangle3_y(rectangle3_ys[414]), .rectangle3_width(rectangle3_widths[414]), .rectangle3_height(rectangle3_heights[414]), .rectangle3_weight(rectangle3_weights[414]), .feature_threshold(feature_thresholds[414]), .feature_above(feature_aboves[414]), .feature_below(feature_belows[414]), .scan_win_std_dev(scan_win_std_dev[414]), .feature_accum(feature_accums[414]));
  accum_calculator ac415(.scan_win(scan_win415), .rectangle1_x(rectangle1_xs[415]), .rectangle1_y(rectangle1_ys[415]), .rectangle1_width(rectangle1_widths[415]), .rectangle1_height(rectangle1_heights[415]), .rectangle1_weight(rectangle1_weights[415]), .rectangle2_x(rectangle2_xs[415]), .rectangle2_y(rectangle2_ys[415]), .rectangle2_width(rectangle2_widths[415]), .rectangle2_height(rectangle2_heights[415]), .rectangle2_weight(rectangle2_weights[415]), .rectangle3_x(rectangle3_xs[415]), .rectangle3_y(rectangle3_ys[415]), .rectangle3_width(rectangle3_widths[415]), .rectangle3_height(rectangle3_heights[415]), .rectangle3_weight(rectangle3_weights[415]), .feature_threshold(feature_thresholds[415]), .feature_above(feature_aboves[415]), .feature_below(feature_belows[415]), .scan_win_std_dev(scan_win_std_dev[415]), .feature_accum(feature_accums[415]));
  accum_calculator ac416(.scan_win(scan_win416), .rectangle1_x(rectangle1_xs[416]), .rectangle1_y(rectangle1_ys[416]), .rectangle1_width(rectangle1_widths[416]), .rectangle1_height(rectangle1_heights[416]), .rectangle1_weight(rectangle1_weights[416]), .rectangle2_x(rectangle2_xs[416]), .rectangle2_y(rectangle2_ys[416]), .rectangle2_width(rectangle2_widths[416]), .rectangle2_height(rectangle2_heights[416]), .rectangle2_weight(rectangle2_weights[416]), .rectangle3_x(rectangle3_xs[416]), .rectangle3_y(rectangle3_ys[416]), .rectangle3_width(rectangle3_widths[416]), .rectangle3_height(rectangle3_heights[416]), .rectangle3_weight(rectangle3_weights[416]), .feature_threshold(feature_thresholds[416]), .feature_above(feature_aboves[416]), .feature_below(feature_belows[416]), .scan_win_std_dev(scan_win_std_dev[416]), .feature_accum(feature_accums[416]));
  accum_calculator ac417(.scan_win(scan_win417), .rectangle1_x(rectangle1_xs[417]), .rectangle1_y(rectangle1_ys[417]), .rectangle1_width(rectangle1_widths[417]), .rectangle1_height(rectangle1_heights[417]), .rectangle1_weight(rectangle1_weights[417]), .rectangle2_x(rectangle2_xs[417]), .rectangle2_y(rectangle2_ys[417]), .rectangle2_width(rectangle2_widths[417]), .rectangle2_height(rectangle2_heights[417]), .rectangle2_weight(rectangle2_weights[417]), .rectangle3_x(rectangle3_xs[417]), .rectangle3_y(rectangle3_ys[417]), .rectangle3_width(rectangle3_widths[417]), .rectangle3_height(rectangle3_heights[417]), .rectangle3_weight(rectangle3_weights[417]), .feature_threshold(feature_thresholds[417]), .feature_above(feature_aboves[417]), .feature_below(feature_belows[417]), .scan_win_std_dev(scan_win_std_dev[417]), .feature_accum(feature_accums[417]));
  accum_calculator ac418(.scan_win(scan_win418), .rectangle1_x(rectangle1_xs[418]), .rectangle1_y(rectangle1_ys[418]), .rectangle1_width(rectangle1_widths[418]), .rectangle1_height(rectangle1_heights[418]), .rectangle1_weight(rectangle1_weights[418]), .rectangle2_x(rectangle2_xs[418]), .rectangle2_y(rectangle2_ys[418]), .rectangle2_width(rectangle2_widths[418]), .rectangle2_height(rectangle2_heights[418]), .rectangle2_weight(rectangle2_weights[418]), .rectangle3_x(rectangle3_xs[418]), .rectangle3_y(rectangle3_ys[418]), .rectangle3_width(rectangle3_widths[418]), .rectangle3_height(rectangle3_heights[418]), .rectangle3_weight(rectangle3_weights[418]), .feature_threshold(feature_thresholds[418]), .feature_above(feature_aboves[418]), .feature_below(feature_belows[418]), .scan_win_std_dev(scan_win_std_dev[418]), .feature_accum(feature_accums[418]));
  accum_calculator ac419(.scan_win(scan_win419), .rectangle1_x(rectangle1_xs[419]), .rectangle1_y(rectangle1_ys[419]), .rectangle1_width(rectangle1_widths[419]), .rectangle1_height(rectangle1_heights[419]), .rectangle1_weight(rectangle1_weights[419]), .rectangle2_x(rectangle2_xs[419]), .rectangle2_y(rectangle2_ys[419]), .rectangle2_width(rectangle2_widths[419]), .rectangle2_height(rectangle2_heights[419]), .rectangle2_weight(rectangle2_weights[419]), .rectangle3_x(rectangle3_xs[419]), .rectangle3_y(rectangle3_ys[419]), .rectangle3_width(rectangle3_widths[419]), .rectangle3_height(rectangle3_heights[419]), .rectangle3_weight(rectangle3_weights[419]), .feature_threshold(feature_thresholds[419]), .feature_above(feature_aboves[419]), .feature_below(feature_belows[419]), .scan_win_std_dev(scan_win_std_dev[419]), .feature_accum(feature_accums[419]));
  accum_calculator ac420(.scan_win(scan_win420), .rectangle1_x(rectangle1_xs[420]), .rectangle1_y(rectangle1_ys[420]), .rectangle1_width(rectangle1_widths[420]), .rectangle1_height(rectangle1_heights[420]), .rectangle1_weight(rectangle1_weights[420]), .rectangle2_x(rectangle2_xs[420]), .rectangle2_y(rectangle2_ys[420]), .rectangle2_width(rectangle2_widths[420]), .rectangle2_height(rectangle2_heights[420]), .rectangle2_weight(rectangle2_weights[420]), .rectangle3_x(rectangle3_xs[420]), .rectangle3_y(rectangle3_ys[420]), .rectangle3_width(rectangle3_widths[420]), .rectangle3_height(rectangle3_heights[420]), .rectangle3_weight(rectangle3_weights[420]), .feature_threshold(feature_thresholds[420]), .feature_above(feature_aboves[420]), .feature_below(feature_belows[420]), .scan_win_std_dev(scan_win_std_dev[420]), .feature_accum(feature_accums[420]));
  accum_calculator ac421(.scan_win(scan_win421), .rectangle1_x(rectangle1_xs[421]), .rectangle1_y(rectangle1_ys[421]), .rectangle1_width(rectangle1_widths[421]), .rectangle1_height(rectangle1_heights[421]), .rectangle1_weight(rectangle1_weights[421]), .rectangle2_x(rectangle2_xs[421]), .rectangle2_y(rectangle2_ys[421]), .rectangle2_width(rectangle2_widths[421]), .rectangle2_height(rectangle2_heights[421]), .rectangle2_weight(rectangle2_weights[421]), .rectangle3_x(rectangle3_xs[421]), .rectangle3_y(rectangle3_ys[421]), .rectangle3_width(rectangle3_widths[421]), .rectangle3_height(rectangle3_heights[421]), .rectangle3_weight(rectangle3_weights[421]), .feature_threshold(feature_thresholds[421]), .feature_above(feature_aboves[421]), .feature_below(feature_belows[421]), .scan_win_std_dev(scan_win_std_dev[421]), .feature_accum(feature_accums[421]));
  accum_calculator ac422(.scan_win(scan_win422), .rectangle1_x(rectangle1_xs[422]), .rectangle1_y(rectangle1_ys[422]), .rectangle1_width(rectangle1_widths[422]), .rectangle1_height(rectangle1_heights[422]), .rectangle1_weight(rectangle1_weights[422]), .rectangle2_x(rectangle2_xs[422]), .rectangle2_y(rectangle2_ys[422]), .rectangle2_width(rectangle2_widths[422]), .rectangle2_height(rectangle2_heights[422]), .rectangle2_weight(rectangle2_weights[422]), .rectangle3_x(rectangle3_xs[422]), .rectangle3_y(rectangle3_ys[422]), .rectangle3_width(rectangle3_widths[422]), .rectangle3_height(rectangle3_heights[422]), .rectangle3_weight(rectangle3_weights[422]), .feature_threshold(feature_thresholds[422]), .feature_above(feature_aboves[422]), .feature_below(feature_belows[422]), .scan_win_std_dev(scan_win_std_dev[422]), .feature_accum(feature_accums[422]));
  accum_calculator ac423(.scan_win(scan_win423), .rectangle1_x(rectangle1_xs[423]), .rectangle1_y(rectangle1_ys[423]), .rectangle1_width(rectangle1_widths[423]), .rectangle1_height(rectangle1_heights[423]), .rectangle1_weight(rectangle1_weights[423]), .rectangle2_x(rectangle2_xs[423]), .rectangle2_y(rectangle2_ys[423]), .rectangle2_width(rectangle2_widths[423]), .rectangle2_height(rectangle2_heights[423]), .rectangle2_weight(rectangle2_weights[423]), .rectangle3_x(rectangle3_xs[423]), .rectangle3_y(rectangle3_ys[423]), .rectangle3_width(rectangle3_widths[423]), .rectangle3_height(rectangle3_heights[423]), .rectangle3_weight(rectangle3_weights[423]), .feature_threshold(feature_thresholds[423]), .feature_above(feature_aboves[423]), .feature_below(feature_belows[423]), .scan_win_std_dev(scan_win_std_dev[423]), .feature_accum(feature_accums[423]));
  accum_calculator ac424(.scan_win(scan_win424), .rectangle1_x(rectangle1_xs[424]), .rectangle1_y(rectangle1_ys[424]), .rectangle1_width(rectangle1_widths[424]), .rectangle1_height(rectangle1_heights[424]), .rectangle1_weight(rectangle1_weights[424]), .rectangle2_x(rectangle2_xs[424]), .rectangle2_y(rectangle2_ys[424]), .rectangle2_width(rectangle2_widths[424]), .rectangle2_height(rectangle2_heights[424]), .rectangle2_weight(rectangle2_weights[424]), .rectangle3_x(rectangle3_xs[424]), .rectangle3_y(rectangle3_ys[424]), .rectangle3_width(rectangle3_widths[424]), .rectangle3_height(rectangle3_heights[424]), .rectangle3_weight(rectangle3_weights[424]), .feature_threshold(feature_thresholds[424]), .feature_above(feature_aboves[424]), .feature_below(feature_belows[424]), .scan_win_std_dev(scan_win_std_dev[424]), .feature_accum(feature_accums[424]));
  accum_calculator ac425(.scan_win(scan_win425), .rectangle1_x(rectangle1_xs[425]), .rectangle1_y(rectangle1_ys[425]), .rectangle1_width(rectangle1_widths[425]), .rectangle1_height(rectangle1_heights[425]), .rectangle1_weight(rectangle1_weights[425]), .rectangle2_x(rectangle2_xs[425]), .rectangle2_y(rectangle2_ys[425]), .rectangle2_width(rectangle2_widths[425]), .rectangle2_height(rectangle2_heights[425]), .rectangle2_weight(rectangle2_weights[425]), .rectangle3_x(rectangle3_xs[425]), .rectangle3_y(rectangle3_ys[425]), .rectangle3_width(rectangle3_widths[425]), .rectangle3_height(rectangle3_heights[425]), .rectangle3_weight(rectangle3_weights[425]), .feature_threshold(feature_thresholds[425]), .feature_above(feature_aboves[425]), .feature_below(feature_belows[425]), .scan_win_std_dev(scan_win_std_dev[425]), .feature_accum(feature_accums[425]));
  accum_calculator ac426(.scan_win(scan_win426), .rectangle1_x(rectangle1_xs[426]), .rectangle1_y(rectangle1_ys[426]), .rectangle1_width(rectangle1_widths[426]), .rectangle1_height(rectangle1_heights[426]), .rectangle1_weight(rectangle1_weights[426]), .rectangle2_x(rectangle2_xs[426]), .rectangle2_y(rectangle2_ys[426]), .rectangle2_width(rectangle2_widths[426]), .rectangle2_height(rectangle2_heights[426]), .rectangle2_weight(rectangle2_weights[426]), .rectangle3_x(rectangle3_xs[426]), .rectangle3_y(rectangle3_ys[426]), .rectangle3_width(rectangle3_widths[426]), .rectangle3_height(rectangle3_heights[426]), .rectangle3_weight(rectangle3_weights[426]), .feature_threshold(feature_thresholds[426]), .feature_above(feature_aboves[426]), .feature_below(feature_belows[426]), .scan_win_std_dev(scan_win_std_dev[426]), .feature_accum(feature_accums[426]));
  accum_calculator ac427(.scan_win(scan_win427), .rectangle1_x(rectangle1_xs[427]), .rectangle1_y(rectangle1_ys[427]), .rectangle1_width(rectangle1_widths[427]), .rectangle1_height(rectangle1_heights[427]), .rectangle1_weight(rectangle1_weights[427]), .rectangle2_x(rectangle2_xs[427]), .rectangle2_y(rectangle2_ys[427]), .rectangle2_width(rectangle2_widths[427]), .rectangle2_height(rectangle2_heights[427]), .rectangle2_weight(rectangle2_weights[427]), .rectangle3_x(rectangle3_xs[427]), .rectangle3_y(rectangle3_ys[427]), .rectangle3_width(rectangle3_widths[427]), .rectangle3_height(rectangle3_heights[427]), .rectangle3_weight(rectangle3_weights[427]), .feature_threshold(feature_thresholds[427]), .feature_above(feature_aboves[427]), .feature_below(feature_belows[427]), .scan_win_std_dev(scan_win_std_dev[427]), .feature_accum(feature_accums[427]));
  accum_calculator ac428(.scan_win(scan_win428), .rectangle1_x(rectangle1_xs[428]), .rectangle1_y(rectangle1_ys[428]), .rectangle1_width(rectangle1_widths[428]), .rectangle1_height(rectangle1_heights[428]), .rectangle1_weight(rectangle1_weights[428]), .rectangle2_x(rectangle2_xs[428]), .rectangle2_y(rectangle2_ys[428]), .rectangle2_width(rectangle2_widths[428]), .rectangle2_height(rectangle2_heights[428]), .rectangle2_weight(rectangle2_weights[428]), .rectangle3_x(rectangle3_xs[428]), .rectangle3_y(rectangle3_ys[428]), .rectangle3_width(rectangle3_widths[428]), .rectangle3_height(rectangle3_heights[428]), .rectangle3_weight(rectangle3_weights[428]), .feature_threshold(feature_thresholds[428]), .feature_above(feature_aboves[428]), .feature_below(feature_belows[428]), .scan_win_std_dev(scan_win_std_dev[428]), .feature_accum(feature_accums[428]));
  accum_calculator ac429(.scan_win(scan_win429), .rectangle1_x(rectangle1_xs[429]), .rectangle1_y(rectangle1_ys[429]), .rectangle1_width(rectangle1_widths[429]), .rectangle1_height(rectangle1_heights[429]), .rectangle1_weight(rectangle1_weights[429]), .rectangle2_x(rectangle2_xs[429]), .rectangle2_y(rectangle2_ys[429]), .rectangle2_width(rectangle2_widths[429]), .rectangle2_height(rectangle2_heights[429]), .rectangle2_weight(rectangle2_weights[429]), .rectangle3_x(rectangle3_xs[429]), .rectangle3_y(rectangle3_ys[429]), .rectangle3_width(rectangle3_widths[429]), .rectangle3_height(rectangle3_heights[429]), .rectangle3_weight(rectangle3_weights[429]), .feature_threshold(feature_thresholds[429]), .feature_above(feature_aboves[429]), .feature_below(feature_belows[429]), .scan_win_std_dev(scan_win_std_dev[429]), .feature_accum(feature_accums[429]));
  accum_calculator ac430(.scan_win(scan_win430), .rectangle1_x(rectangle1_xs[430]), .rectangle1_y(rectangle1_ys[430]), .rectangle1_width(rectangle1_widths[430]), .rectangle1_height(rectangle1_heights[430]), .rectangle1_weight(rectangle1_weights[430]), .rectangle2_x(rectangle2_xs[430]), .rectangle2_y(rectangle2_ys[430]), .rectangle2_width(rectangle2_widths[430]), .rectangle2_height(rectangle2_heights[430]), .rectangle2_weight(rectangle2_weights[430]), .rectangle3_x(rectangle3_xs[430]), .rectangle3_y(rectangle3_ys[430]), .rectangle3_width(rectangle3_widths[430]), .rectangle3_height(rectangle3_heights[430]), .rectangle3_weight(rectangle3_weights[430]), .feature_threshold(feature_thresholds[430]), .feature_above(feature_aboves[430]), .feature_below(feature_belows[430]), .scan_win_std_dev(scan_win_std_dev[430]), .feature_accum(feature_accums[430]));
  accum_calculator ac431(.scan_win(scan_win431), .rectangle1_x(rectangle1_xs[431]), .rectangle1_y(rectangle1_ys[431]), .rectangle1_width(rectangle1_widths[431]), .rectangle1_height(rectangle1_heights[431]), .rectangle1_weight(rectangle1_weights[431]), .rectangle2_x(rectangle2_xs[431]), .rectangle2_y(rectangle2_ys[431]), .rectangle2_width(rectangle2_widths[431]), .rectangle2_height(rectangle2_heights[431]), .rectangle2_weight(rectangle2_weights[431]), .rectangle3_x(rectangle3_xs[431]), .rectangle3_y(rectangle3_ys[431]), .rectangle3_width(rectangle3_widths[431]), .rectangle3_height(rectangle3_heights[431]), .rectangle3_weight(rectangle3_weights[431]), .feature_threshold(feature_thresholds[431]), .feature_above(feature_aboves[431]), .feature_below(feature_belows[431]), .scan_win_std_dev(scan_win_std_dev[431]), .feature_accum(feature_accums[431]));
  accum_calculator ac432(.scan_win(scan_win432), .rectangle1_x(rectangle1_xs[432]), .rectangle1_y(rectangle1_ys[432]), .rectangle1_width(rectangle1_widths[432]), .rectangle1_height(rectangle1_heights[432]), .rectangle1_weight(rectangle1_weights[432]), .rectangle2_x(rectangle2_xs[432]), .rectangle2_y(rectangle2_ys[432]), .rectangle2_width(rectangle2_widths[432]), .rectangle2_height(rectangle2_heights[432]), .rectangle2_weight(rectangle2_weights[432]), .rectangle3_x(rectangle3_xs[432]), .rectangle3_y(rectangle3_ys[432]), .rectangle3_width(rectangle3_widths[432]), .rectangle3_height(rectangle3_heights[432]), .rectangle3_weight(rectangle3_weights[432]), .feature_threshold(feature_thresholds[432]), .feature_above(feature_aboves[432]), .feature_below(feature_belows[432]), .scan_win_std_dev(scan_win_std_dev[432]), .feature_accum(feature_accums[432]));
  accum_calculator ac433(.scan_win(scan_win433), .rectangle1_x(rectangle1_xs[433]), .rectangle1_y(rectangle1_ys[433]), .rectangle1_width(rectangle1_widths[433]), .rectangle1_height(rectangle1_heights[433]), .rectangle1_weight(rectangle1_weights[433]), .rectangle2_x(rectangle2_xs[433]), .rectangle2_y(rectangle2_ys[433]), .rectangle2_width(rectangle2_widths[433]), .rectangle2_height(rectangle2_heights[433]), .rectangle2_weight(rectangle2_weights[433]), .rectangle3_x(rectangle3_xs[433]), .rectangle3_y(rectangle3_ys[433]), .rectangle3_width(rectangle3_widths[433]), .rectangle3_height(rectangle3_heights[433]), .rectangle3_weight(rectangle3_weights[433]), .feature_threshold(feature_thresholds[433]), .feature_above(feature_aboves[433]), .feature_below(feature_belows[433]), .scan_win_std_dev(scan_win_std_dev[433]), .feature_accum(feature_accums[433]));
  accum_calculator ac434(.scan_win(scan_win434), .rectangle1_x(rectangle1_xs[434]), .rectangle1_y(rectangle1_ys[434]), .rectangle1_width(rectangle1_widths[434]), .rectangle1_height(rectangle1_heights[434]), .rectangle1_weight(rectangle1_weights[434]), .rectangle2_x(rectangle2_xs[434]), .rectangle2_y(rectangle2_ys[434]), .rectangle2_width(rectangle2_widths[434]), .rectangle2_height(rectangle2_heights[434]), .rectangle2_weight(rectangle2_weights[434]), .rectangle3_x(rectangle3_xs[434]), .rectangle3_y(rectangle3_ys[434]), .rectangle3_width(rectangle3_widths[434]), .rectangle3_height(rectangle3_heights[434]), .rectangle3_weight(rectangle3_weights[434]), .feature_threshold(feature_thresholds[434]), .feature_above(feature_aboves[434]), .feature_below(feature_belows[434]), .scan_win_std_dev(scan_win_std_dev[434]), .feature_accum(feature_accums[434]));
  accum_calculator ac435(.scan_win(scan_win435), .rectangle1_x(rectangle1_xs[435]), .rectangle1_y(rectangle1_ys[435]), .rectangle1_width(rectangle1_widths[435]), .rectangle1_height(rectangle1_heights[435]), .rectangle1_weight(rectangle1_weights[435]), .rectangle2_x(rectangle2_xs[435]), .rectangle2_y(rectangle2_ys[435]), .rectangle2_width(rectangle2_widths[435]), .rectangle2_height(rectangle2_heights[435]), .rectangle2_weight(rectangle2_weights[435]), .rectangle3_x(rectangle3_xs[435]), .rectangle3_y(rectangle3_ys[435]), .rectangle3_width(rectangle3_widths[435]), .rectangle3_height(rectangle3_heights[435]), .rectangle3_weight(rectangle3_weights[435]), .feature_threshold(feature_thresholds[435]), .feature_above(feature_aboves[435]), .feature_below(feature_belows[435]), .scan_win_std_dev(scan_win_std_dev[435]), .feature_accum(feature_accums[435]));
  accum_calculator ac436(.scan_win(scan_win436), .rectangle1_x(rectangle1_xs[436]), .rectangle1_y(rectangle1_ys[436]), .rectangle1_width(rectangle1_widths[436]), .rectangle1_height(rectangle1_heights[436]), .rectangle1_weight(rectangle1_weights[436]), .rectangle2_x(rectangle2_xs[436]), .rectangle2_y(rectangle2_ys[436]), .rectangle2_width(rectangle2_widths[436]), .rectangle2_height(rectangle2_heights[436]), .rectangle2_weight(rectangle2_weights[436]), .rectangle3_x(rectangle3_xs[436]), .rectangle3_y(rectangle3_ys[436]), .rectangle3_width(rectangle3_widths[436]), .rectangle3_height(rectangle3_heights[436]), .rectangle3_weight(rectangle3_weights[436]), .feature_threshold(feature_thresholds[436]), .feature_above(feature_aboves[436]), .feature_below(feature_belows[436]), .scan_win_std_dev(scan_win_std_dev[436]), .feature_accum(feature_accums[436]));
  accum_calculator ac437(.scan_win(scan_win437), .rectangle1_x(rectangle1_xs[437]), .rectangle1_y(rectangle1_ys[437]), .rectangle1_width(rectangle1_widths[437]), .rectangle1_height(rectangle1_heights[437]), .rectangle1_weight(rectangle1_weights[437]), .rectangle2_x(rectangle2_xs[437]), .rectangle2_y(rectangle2_ys[437]), .rectangle2_width(rectangle2_widths[437]), .rectangle2_height(rectangle2_heights[437]), .rectangle2_weight(rectangle2_weights[437]), .rectangle3_x(rectangle3_xs[437]), .rectangle3_y(rectangle3_ys[437]), .rectangle3_width(rectangle3_widths[437]), .rectangle3_height(rectangle3_heights[437]), .rectangle3_weight(rectangle3_weights[437]), .feature_threshold(feature_thresholds[437]), .feature_above(feature_aboves[437]), .feature_below(feature_belows[437]), .scan_win_std_dev(scan_win_std_dev[437]), .feature_accum(feature_accums[437]));
  accum_calculator ac438(.scan_win(scan_win438), .rectangle1_x(rectangle1_xs[438]), .rectangle1_y(rectangle1_ys[438]), .rectangle1_width(rectangle1_widths[438]), .rectangle1_height(rectangle1_heights[438]), .rectangle1_weight(rectangle1_weights[438]), .rectangle2_x(rectangle2_xs[438]), .rectangle2_y(rectangle2_ys[438]), .rectangle2_width(rectangle2_widths[438]), .rectangle2_height(rectangle2_heights[438]), .rectangle2_weight(rectangle2_weights[438]), .rectangle3_x(rectangle3_xs[438]), .rectangle3_y(rectangle3_ys[438]), .rectangle3_width(rectangle3_widths[438]), .rectangle3_height(rectangle3_heights[438]), .rectangle3_weight(rectangle3_weights[438]), .feature_threshold(feature_thresholds[438]), .feature_above(feature_aboves[438]), .feature_below(feature_belows[438]), .scan_win_std_dev(scan_win_std_dev[438]), .feature_accum(feature_accums[438]));
  accum_calculator ac439(.scan_win(scan_win439), .rectangle1_x(rectangle1_xs[439]), .rectangle1_y(rectangle1_ys[439]), .rectangle1_width(rectangle1_widths[439]), .rectangle1_height(rectangle1_heights[439]), .rectangle1_weight(rectangle1_weights[439]), .rectangle2_x(rectangle2_xs[439]), .rectangle2_y(rectangle2_ys[439]), .rectangle2_width(rectangle2_widths[439]), .rectangle2_height(rectangle2_heights[439]), .rectangle2_weight(rectangle2_weights[439]), .rectangle3_x(rectangle3_xs[439]), .rectangle3_y(rectangle3_ys[439]), .rectangle3_width(rectangle3_widths[439]), .rectangle3_height(rectangle3_heights[439]), .rectangle3_weight(rectangle3_weights[439]), .feature_threshold(feature_thresholds[439]), .feature_above(feature_aboves[439]), .feature_below(feature_belows[439]), .scan_win_std_dev(scan_win_std_dev[439]), .feature_accum(feature_accums[439]));
  accum_calculator ac440(.scan_win(scan_win440), .rectangle1_x(rectangle1_xs[440]), .rectangle1_y(rectangle1_ys[440]), .rectangle1_width(rectangle1_widths[440]), .rectangle1_height(rectangle1_heights[440]), .rectangle1_weight(rectangle1_weights[440]), .rectangle2_x(rectangle2_xs[440]), .rectangle2_y(rectangle2_ys[440]), .rectangle2_width(rectangle2_widths[440]), .rectangle2_height(rectangle2_heights[440]), .rectangle2_weight(rectangle2_weights[440]), .rectangle3_x(rectangle3_xs[440]), .rectangle3_y(rectangle3_ys[440]), .rectangle3_width(rectangle3_widths[440]), .rectangle3_height(rectangle3_heights[440]), .rectangle3_weight(rectangle3_weights[440]), .feature_threshold(feature_thresholds[440]), .feature_above(feature_aboves[440]), .feature_below(feature_belows[440]), .scan_win_std_dev(scan_win_std_dev[440]), .feature_accum(feature_accums[440]));
  accum_calculator ac441(.scan_win(scan_win441), .rectangle1_x(rectangle1_xs[441]), .rectangle1_y(rectangle1_ys[441]), .rectangle1_width(rectangle1_widths[441]), .rectangle1_height(rectangle1_heights[441]), .rectangle1_weight(rectangle1_weights[441]), .rectangle2_x(rectangle2_xs[441]), .rectangle2_y(rectangle2_ys[441]), .rectangle2_width(rectangle2_widths[441]), .rectangle2_height(rectangle2_heights[441]), .rectangle2_weight(rectangle2_weights[441]), .rectangle3_x(rectangle3_xs[441]), .rectangle3_y(rectangle3_ys[441]), .rectangle3_width(rectangle3_widths[441]), .rectangle3_height(rectangle3_heights[441]), .rectangle3_weight(rectangle3_weights[441]), .feature_threshold(feature_thresholds[441]), .feature_above(feature_aboves[441]), .feature_below(feature_belows[441]), .scan_win_std_dev(scan_win_std_dev[441]), .feature_accum(feature_accums[441]));
  accum_calculator ac442(.scan_win(scan_win442), .rectangle1_x(rectangle1_xs[442]), .rectangle1_y(rectangle1_ys[442]), .rectangle1_width(rectangle1_widths[442]), .rectangle1_height(rectangle1_heights[442]), .rectangle1_weight(rectangle1_weights[442]), .rectangle2_x(rectangle2_xs[442]), .rectangle2_y(rectangle2_ys[442]), .rectangle2_width(rectangle2_widths[442]), .rectangle2_height(rectangle2_heights[442]), .rectangle2_weight(rectangle2_weights[442]), .rectangle3_x(rectangle3_xs[442]), .rectangle3_y(rectangle3_ys[442]), .rectangle3_width(rectangle3_widths[442]), .rectangle3_height(rectangle3_heights[442]), .rectangle3_weight(rectangle3_weights[442]), .feature_threshold(feature_thresholds[442]), .feature_above(feature_aboves[442]), .feature_below(feature_belows[442]), .scan_win_std_dev(scan_win_std_dev[442]), .feature_accum(feature_accums[442]));
  accum_calculator ac443(.scan_win(scan_win443), .rectangle1_x(rectangle1_xs[443]), .rectangle1_y(rectangle1_ys[443]), .rectangle1_width(rectangle1_widths[443]), .rectangle1_height(rectangle1_heights[443]), .rectangle1_weight(rectangle1_weights[443]), .rectangle2_x(rectangle2_xs[443]), .rectangle2_y(rectangle2_ys[443]), .rectangle2_width(rectangle2_widths[443]), .rectangle2_height(rectangle2_heights[443]), .rectangle2_weight(rectangle2_weights[443]), .rectangle3_x(rectangle3_xs[443]), .rectangle3_y(rectangle3_ys[443]), .rectangle3_width(rectangle3_widths[443]), .rectangle3_height(rectangle3_heights[443]), .rectangle3_weight(rectangle3_weights[443]), .feature_threshold(feature_thresholds[443]), .feature_above(feature_aboves[443]), .feature_below(feature_belows[443]), .scan_win_std_dev(scan_win_std_dev[443]), .feature_accum(feature_accums[443]));
  accum_calculator ac444(.scan_win(scan_win444), .rectangle1_x(rectangle1_xs[444]), .rectangle1_y(rectangle1_ys[444]), .rectangle1_width(rectangle1_widths[444]), .rectangle1_height(rectangle1_heights[444]), .rectangle1_weight(rectangle1_weights[444]), .rectangle2_x(rectangle2_xs[444]), .rectangle2_y(rectangle2_ys[444]), .rectangle2_width(rectangle2_widths[444]), .rectangle2_height(rectangle2_heights[444]), .rectangle2_weight(rectangle2_weights[444]), .rectangle3_x(rectangle3_xs[444]), .rectangle3_y(rectangle3_ys[444]), .rectangle3_width(rectangle3_widths[444]), .rectangle3_height(rectangle3_heights[444]), .rectangle3_weight(rectangle3_weights[444]), .feature_threshold(feature_thresholds[444]), .feature_above(feature_aboves[444]), .feature_below(feature_belows[444]), .scan_win_std_dev(scan_win_std_dev[444]), .feature_accum(feature_accums[444]));
  accum_calculator ac445(.scan_win(scan_win445), .rectangle1_x(rectangle1_xs[445]), .rectangle1_y(rectangle1_ys[445]), .rectangle1_width(rectangle1_widths[445]), .rectangle1_height(rectangle1_heights[445]), .rectangle1_weight(rectangle1_weights[445]), .rectangle2_x(rectangle2_xs[445]), .rectangle2_y(rectangle2_ys[445]), .rectangle2_width(rectangle2_widths[445]), .rectangle2_height(rectangle2_heights[445]), .rectangle2_weight(rectangle2_weights[445]), .rectangle3_x(rectangle3_xs[445]), .rectangle3_y(rectangle3_ys[445]), .rectangle3_width(rectangle3_widths[445]), .rectangle3_height(rectangle3_heights[445]), .rectangle3_weight(rectangle3_weights[445]), .feature_threshold(feature_thresholds[445]), .feature_above(feature_aboves[445]), .feature_below(feature_belows[445]), .scan_win_std_dev(scan_win_std_dev[445]), .feature_accum(feature_accums[445]));
  accum_calculator ac446(.scan_win(scan_win446), .rectangle1_x(rectangle1_xs[446]), .rectangle1_y(rectangle1_ys[446]), .rectangle1_width(rectangle1_widths[446]), .rectangle1_height(rectangle1_heights[446]), .rectangle1_weight(rectangle1_weights[446]), .rectangle2_x(rectangle2_xs[446]), .rectangle2_y(rectangle2_ys[446]), .rectangle2_width(rectangle2_widths[446]), .rectangle2_height(rectangle2_heights[446]), .rectangle2_weight(rectangle2_weights[446]), .rectangle3_x(rectangle3_xs[446]), .rectangle3_y(rectangle3_ys[446]), .rectangle3_width(rectangle3_widths[446]), .rectangle3_height(rectangle3_heights[446]), .rectangle3_weight(rectangle3_weights[446]), .feature_threshold(feature_thresholds[446]), .feature_above(feature_aboves[446]), .feature_below(feature_belows[446]), .scan_win_std_dev(scan_win_std_dev[446]), .feature_accum(feature_accums[446]));
  accum_calculator ac447(.scan_win(scan_win447), .rectangle1_x(rectangle1_xs[447]), .rectangle1_y(rectangle1_ys[447]), .rectangle1_width(rectangle1_widths[447]), .rectangle1_height(rectangle1_heights[447]), .rectangle1_weight(rectangle1_weights[447]), .rectangle2_x(rectangle2_xs[447]), .rectangle2_y(rectangle2_ys[447]), .rectangle2_width(rectangle2_widths[447]), .rectangle2_height(rectangle2_heights[447]), .rectangle2_weight(rectangle2_weights[447]), .rectangle3_x(rectangle3_xs[447]), .rectangle3_y(rectangle3_ys[447]), .rectangle3_width(rectangle3_widths[447]), .rectangle3_height(rectangle3_heights[447]), .rectangle3_weight(rectangle3_weights[447]), .feature_threshold(feature_thresholds[447]), .feature_above(feature_aboves[447]), .feature_below(feature_belows[447]), .scan_win_std_dev(scan_win_std_dev[447]), .feature_accum(feature_accums[447]));
  accum_calculator ac448(.scan_win(scan_win448), .rectangle1_x(rectangle1_xs[448]), .rectangle1_y(rectangle1_ys[448]), .rectangle1_width(rectangle1_widths[448]), .rectangle1_height(rectangle1_heights[448]), .rectangle1_weight(rectangle1_weights[448]), .rectangle2_x(rectangle2_xs[448]), .rectangle2_y(rectangle2_ys[448]), .rectangle2_width(rectangle2_widths[448]), .rectangle2_height(rectangle2_heights[448]), .rectangle2_weight(rectangle2_weights[448]), .rectangle3_x(rectangle3_xs[448]), .rectangle3_y(rectangle3_ys[448]), .rectangle3_width(rectangle3_widths[448]), .rectangle3_height(rectangle3_heights[448]), .rectangle3_weight(rectangle3_weights[448]), .feature_threshold(feature_thresholds[448]), .feature_above(feature_aboves[448]), .feature_below(feature_belows[448]), .scan_win_std_dev(scan_win_std_dev[448]), .feature_accum(feature_accums[448]));
  accum_calculator ac449(.scan_win(scan_win449), .rectangle1_x(rectangle1_xs[449]), .rectangle1_y(rectangle1_ys[449]), .rectangle1_width(rectangle1_widths[449]), .rectangle1_height(rectangle1_heights[449]), .rectangle1_weight(rectangle1_weights[449]), .rectangle2_x(rectangle2_xs[449]), .rectangle2_y(rectangle2_ys[449]), .rectangle2_width(rectangle2_widths[449]), .rectangle2_height(rectangle2_heights[449]), .rectangle2_weight(rectangle2_weights[449]), .rectangle3_x(rectangle3_xs[449]), .rectangle3_y(rectangle3_ys[449]), .rectangle3_width(rectangle3_widths[449]), .rectangle3_height(rectangle3_heights[449]), .rectangle3_weight(rectangle3_weights[449]), .feature_threshold(feature_thresholds[449]), .feature_above(feature_aboves[449]), .feature_below(feature_belows[449]), .scan_win_std_dev(scan_win_std_dev[449]), .feature_accum(feature_accums[449]));
  accum_calculator ac450(.scan_win(scan_win450), .rectangle1_x(rectangle1_xs[450]), .rectangle1_y(rectangle1_ys[450]), .rectangle1_width(rectangle1_widths[450]), .rectangle1_height(rectangle1_heights[450]), .rectangle1_weight(rectangle1_weights[450]), .rectangle2_x(rectangle2_xs[450]), .rectangle2_y(rectangle2_ys[450]), .rectangle2_width(rectangle2_widths[450]), .rectangle2_height(rectangle2_heights[450]), .rectangle2_weight(rectangle2_weights[450]), .rectangle3_x(rectangle3_xs[450]), .rectangle3_y(rectangle3_ys[450]), .rectangle3_width(rectangle3_widths[450]), .rectangle3_height(rectangle3_heights[450]), .rectangle3_weight(rectangle3_weights[450]), .feature_threshold(feature_thresholds[450]), .feature_above(feature_aboves[450]), .feature_below(feature_belows[450]), .scan_win_std_dev(scan_win_std_dev[450]), .feature_accum(feature_accums[450]));
  accum_calculator ac451(.scan_win(scan_win451), .rectangle1_x(rectangle1_xs[451]), .rectangle1_y(rectangle1_ys[451]), .rectangle1_width(rectangle1_widths[451]), .rectangle1_height(rectangle1_heights[451]), .rectangle1_weight(rectangle1_weights[451]), .rectangle2_x(rectangle2_xs[451]), .rectangle2_y(rectangle2_ys[451]), .rectangle2_width(rectangle2_widths[451]), .rectangle2_height(rectangle2_heights[451]), .rectangle2_weight(rectangle2_weights[451]), .rectangle3_x(rectangle3_xs[451]), .rectangle3_y(rectangle3_ys[451]), .rectangle3_width(rectangle3_widths[451]), .rectangle3_height(rectangle3_heights[451]), .rectangle3_weight(rectangle3_weights[451]), .feature_threshold(feature_thresholds[451]), .feature_above(feature_aboves[451]), .feature_below(feature_belows[451]), .scan_win_std_dev(scan_win_std_dev[451]), .feature_accum(feature_accums[451]));
  accum_calculator ac452(.scan_win(scan_win452), .rectangle1_x(rectangle1_xs[452]), .rectangle1_y(rectangle1_ys[452]), .rectangle1_width(rectangle1_widths[452]), .rectangle1_height(rectangle1_heights[452]), .rectangle1_weight(rectangle1_weights[452]), .rectangle2_x(rectangle2_xs[452]), .rectangle2_y(rectangle2_ys[452]), .rectangle2_width(rectangle2_widths[452]), .rectangle2_height(rectangle2_heights[452]), .rectangle2_weight(rectangle2_weights[452]), .rectangle3_x(rectangle3_xs[452]), .rectangle3_y(rectangle3_ys[452]), .rectangle3_width(rectangle3_widths[452]), .rectangle3_height(rectangle3_heights[452]), .rectangle3_weight(rectangle3_weights[452]), .feature_threshold(feature_thresholds[452]), .feature_above(feature_aboves[452]), .feature_below(feature_belows[452]), .scan_win_std_dev(scan_win_std_dev[452]), .feature_accum(feature_accums[452]));
  accum_calculator ac453(.scan_win(scan_win453), .rectangle1_x(rectangle1_xs[453]), .rectangle1_y(rectangle1_ys[453]), .rectangle1_width(rectangle1_widths[453]), .rectangle1_height(rectangle1_heights[453]), .rectangle1_weight(rectangle1_weights[453]), .rectangle2_x(rectangle2_xs[453]), .rectangle2_y(rectangle2_ys[453]), .rectangle2_width(rectangle2_widths[453]), .rectangle2_height(rectangle2_heights[453]), .rectangle2_weight(rectangle2_weights[453]), .rectangle3_x(rectangle3_xs[453]), .rectangle3_y(rectangle3_ys[453]), .rectangle3_width(rectangle3_widths[453]), .rectangle3_height(rectangle3_heights[453]), .rectangle3_weight(rectangle3_weights[453]), .feature_threshold(feature_thresholds[453]), .feature_above(feature_aboves[453]), .feature_below(feature_belows[453]), .scan_win_std_dev(scan_win_std_dev[453]), .feature_accum(feature_accums[453]));
  accum_calculator ac454(.scan_win(scan_win454), .rectangle1_x(rectangle1_xs[454]), .rectangle1_y(rectangle1_ys[454]), .rectangle1_width(rectangle1_widths[454]), .rectangle1_height(rectangle1_heights[454]), .rectangle1_weight(rectangle1_weights[454]), .rectangle2_x(rectangle2_xs[454]), .rectangle2_y(rectangle2_ys[454]), .rectangle2_width(rectangle2_widths[454]), .rectangle2_height(rectangle2_heights[454]), .rectangle2_weight(rectangle2_weights[454]), .rectangle3_x(rectangle3_xs[454]), .rectangle3_y(rectangle3_ys[454]), .rectangle3_width(rectangle3_widths[454]), .rectangle3_height(rectangle3_heights[454]), .rectangle3_weight(rectangle3_weights[454]), .feature_threshold(feature_thresholds[454]), .feature_above(feature_aboves[454]), .feature_below(feature_belows[454]), .scan_win_std_dev(scan_win_std_dev[454]), .feature_accum(feature_accums[454]));
  accum_calculator ac455(.scan_win(scan_win455), .rectangle1_x(rectangle1_xs[455]), .rectangle1_y(rectangle1_ys[455]), .rectangle1_width(rectangle1_widths[455]), .rectangle1_height(rectangle1_heights[455]), .rectangle1_weight(rectangle1_weights[455]), .rectangle2_x(rectangle2_xs[455]), .rectangle2_y(rectangle2_ys[455]), .rectangle2_width(rectangle2_widths[455]), .rectangle2_height(rectangle2_heights[455]), .rectangle2_weight(rectangle2_weights[455]), .rectangle3_x(rectangle3_xs[455]), .rectangle3_y(rectangle3_ys[455]), .rectangle3_width(rectangle3_widths[455]), .rectangle3_height(rectangle3_heights[455]), .rectangle3_weight(rectangle3_weights[455]), .feature_threshold(feature_thresholds[455]), .feature_above(feature_aboves[455]), .feature_below(feature_belows[455]), .scan_win_std_dev(scan_win_std_dev[455]), .feature_accum(feature_accums[455]));
  accum_calculator ac456(.scan_win(scan_win456), .rectangle1_x(rectangle1_xs[456]), .rectangle1_y(rectangle1_ys[456]), .rectangle1_width(rectangle1_widths[456]), .rectangle1_height(rectangle1_heights[456]), .rectangle1_weight(rectangle1_weights[456]), .rectangle2_x(rectangle2_xs[456]), .rectangle2_y(rectangle2_ys[456]), .rectangle2_width(rectangle2_widths[456]), .rectangle2_height(rectangle2_heights[456]), .rectangle2_weight(rectangle2_weights[456]), .rectangle3_x(rectangle3_xs[456]), .rectangle3_y(rectangle3_ys[456]), .rectangle3_width(rectangle3_widths[456]), .rectangle3_height(rectangle3_heights[456]), .rectangle3_weight(rectangle3_weights[456]), .feature_threshold(feature_thresholds[456]), .feature_above(feature_aboves[456]), .feature_below(feature_belows[456]), .scan_win_std_dev(scan_win_std_dev[456]), .feature_accum(feature_accums[456]));
  accum_calculator ac457(.scan_win(scan_win457), .rectangle1_x(rectangle1_xs[457]), .rectangle1_y(rectangle1_ys[457]), .rectangle1_width(rectangle1_widths[457]), .rectangle1_height(rectangle1_heights[457]), .rectangle1_weight(rectangle1_weights[457]), .rectangle2_x(rectangle2_xs[457]), .rectangle2_y(rectangle2_ys[457]), .rectangle2_width(rectangle2_widths[457]), .rectangle2_height(rectangle2_heights[457]), .rectangle2_weight(rectangle2_weights[457]), .rectangle3_x(rectangle3_xs[457]), .rectangle3_y(rectangle3_ys[457]), .rectangle3_width(rectangle3_widths[457]), .rectangle3_height(rectangle3_heights[457]), .rectangle3_weight(rectangle3_weights[457]), .feature_threshold(feature_thresholds[457]), .feature_above(feature_aboves[457]), .feature_below(feature_belows[457]), .scan_win_std_dev(scan_win_std_dev[457]), .feature_accum(feature_accums[457]));
  accum_calculator ac458(.scan_win(scan_win458), .rectangle1_x(rectangle1_xs[458]), .rectangle1_y(rectangle1_ys[458]), .rectangle1_width(rectangle1_widths[458]), .rectangle1_height(rectangle1_heights[458]), .rectangle1_weight(rectangle1_weights[458]), .rectangle2_x(rectangle2_xs[458]), .rectangle2_y(rectangle2_ys[458]), .rectangle2_width(rectangle2_widths[458]), .rectangle2_height(rectangle2_heights[458]), .rectangle2_weight(rectangle2_weights[458]), .rectangle3_x(rectangle3_xs[458]), .rectangle3_y(rectangle3_ys[458]), .rectangle3_width(rectangle3_widths[458]), .rectangle3_height(rectangle3_heights[458]), .rectangle3_weight(rectangle3_weights[458]), .feature_threshold(feature_thresholds[458]), .feature_above(feature_aboves[458]), .feature_below(feature_belows[458]), .scan_win_std_dev(scan_win_std_dev[458]), .feature_accum(feature_accums[458]));
  accum_calculator ac459(.scan_win(scan_win459), .rectangle1_x(rectangle1_xs[459]), .rectangle1_y(rectangle1_ys[459]), .rectangle1_width(rectangle1_widths[459]), .rectangle1_height(rectangle1_heights[459]), .rectangle1_weight(rectangle1_weights[459]), .rectangle2_x(rectangle2_xs[459]), .rectangle2_y(rectangle2_ys[459]), .rectangle2_width(rectangle2_widths[459]), .rectangle2_height(rectangle2_heights[459]), .rectangle2_weight(rectangle2_weights[459]), .rectangle3_x(rectangle3_xs[459]), .rectangle3_y(rectangle3_ys[459]), .rectangle3_width(rectangle3_widths[459]), .rectangle3_height(rectangle3_heights[459]), .rectangle3_weight(rectangle3_weights[459]), .feature_threshold(feature_thresholds[459]), .feature_above(feature_aboves[459]), .feature_below(feature_belows[459]), .scan_win_std_dev(scan_win_std_dev[459]), .feature_accum(feature_accums[459]));
  accum_calculator ac460(.scan_win(scan_win460), .rectangle1_x(rectangle1_xs[460]), .rectangle1_y(rectangle1_ys[460]), .rectangle1_width(rectangle1_widths[460]), .rectangle1_height(rectangle1_heights[460]), .rectangle1_weight(rectangle1_weights[460]), .rectangle2_x(rectangle2_xs[460]), .rectangle2_y(rectangle2_ys[460]), .rectangle2_width(rectangle2_widths[460]), .rectangle2_height(rectangle2_heights[460]), .rectangle2_weight(rectangle2_weights[460]), .rectangle3_x(rectangle3_xs[460]), .rectangle3_y(rectangle3_ys[460]), .rectangle3_width(rectangle3_widths[460]), .rectangle3_height(rectangle3_heights[460]), .rectangle3_weight(rectangle3_weights[460]), .feature_threshold(feature_thresholds[460]), .feature_above(feature_aboves[460]), .feature_below(feature_belows[460]), .scan_win_std_dev(scan_win_std_dev[460]), .feature_accum(feature_accums[460]));
  accum_calculator ac461(.scan_win(scan_win461), .rectangle1_x(rectangle1_xs[461]), .rectangle1_y(rectangle1_ys[461]), .rectangle1_width(rectangle1_widths[461]), .rectangle1_height(rectangle1_heights[461]), .rectangle1_weight(rectangle1_weights[461]), .rectangle2_x(rectangle2_xs[461]), .rectangle2_y(rectangle2_ys[461]), .rectangle2_width(rectangle2_widths[461]), .rectangle2_height(rectangle2_heights[461]), .rectangle2_weight(rectangle2_weights[461]), .rectangle3_x(rectangle3_xs[461]), .rectangle3_y(rectangle3_ys[461]), .rectangle3_width(rectangle3_widths[461]), .rectangle3_height(rectangle3_heights[461]), .rectangle3_weight(rectangle3_weights[461]), .feature_threshold(feature_thresholds[461]), .feature_above(feature_aboves[461]), .feature_below(feature_belows[461]), .scan_win_std_dev(scan_win_std_dev[461]), .feature_accum(feature_accums[461]));
  accum_calculator ac462(.scan_win(scan_win462), .rectangle1_x(rectangle1_xs[462]), .rectangle1_y(rectangle1_ys[462]), .rectangle1_width(rectangle1_widths[462]), .rectangle1_height(rectangle1_heights[462]), .rectangle1_weight(rectangle1_weights[462]), .rectangle2_x(rectangle2_xs[462]), .rectangle2_y(rectangle2_ys[462]), .rectangle2_width(rectangle2_widths[462]), .rectangle2_height(rectangle2_heights[462]), .rectangle2_weight(rectangle2_weights[462]), .rectangle3_x(rectangle3_xs[462]), .rectangle3_y(rectangle3_ys[462]), .rectangle3_width(rectangle3_widths[462]), .rectangle3_height(rectangle3_heights[462]), .rectangle3_weight(rectangle3_weights[462]), .feature_threshold(feature_thresholds[462]), .feature_above(feature_aboves[462]), .feature_below(feature_belows[462]), .scan_win_std_dev(scan_win_std_dev[462]), .feature_accum(feature_accums[462]));
  accum_calculator ac463(.scan_win(scan_win463), .rectangle1_x(rectangle1_xs[463]), .rectangle1_y(rectangle1_ys[463]), .rectangle1_width(rectangle1_widths[463]), .rectangle1_height(rectangle1_heights[463]), .rectangle1_weight(rectangle1_weights[463]), .rectangle2_x(rectangle2_xs[463]), .rectangle2_y(rectangle2_ys[463]), .rectangle2_width(rectangle2_widths[463]), .rectangle2_height(rectangle2_heights[463]), .rectangle2_weight(rectangle2_weights[463]), .rectangle3_x(rectangle3_xs[463]), .rectangle3_y(rectangle3_ys[463]), .rectangle3_width(rectangle3_widths[463]), .rectangle3_height(rectangle3_heights[463]), .rectangle3_weight(rectangle3_weights[463]), .feature_threshold(feature_thresholds[463]), .feature_above(feature_aboves[463]), .feature_below(feature_belows[463]), .scan_win_std_dev(scan_win_std_dev[463]), .feature_accum(feature_accums[463]));
  accum_calculator ac464(.scan_win(scan_win464), .rectangle1_x(rectangle1_xs[464]), .rectangle1_y(rectangle1_ys[464]), .rectangle1_width(rectangle1_widths[464]), .rectangle1_height(rectangle1_heights[464]), .rectangle1_weight(rectangle1_weights[464]), .rectangle2_x(rectangle2_xs[464]), .rectangle2_y(rectangle2_ys[464]), .rectangle2_width(rectangle2_widths[464]), .rectangle2_height(rectangle2_heights[464]), .rectangle2_weight(rectangle2_weights[464]), .rectangle3_x(rectangle3_xs[464]), .rectangle3_y(rectangle3_ys[464]), .rectangle3_width(rectangle3_widths[464]), .rectangle3_height(rectangle3_heights[464]), .rectangle3_weight(rectangle3_weights[464]), .feature_threshold(feature_thresholds[464]), .feature_above(feature_aboves[464]), .feature_below(feature_belows[464]), .scan_win_std_dev(scan_win_std_dev[464]), .feature_accum(feature_accums[464]));
  accum_calculator ac465(.scan_win(scan_win465), .rectangle1_x(rectangle1_xs[465]), .rectangle1_y(rectangle1_ys[465]), .rectangle1_width(rectangle1_widths[465]), .rectangle1_height(rectangle1_heights[465]), .rectangle1_weight(rectangle1_weights[465]), .rectangle2_x(rectangle2_xs[465]), .rectangle2_y(rectangle2_ys[465]), .rectangle2_width(rectangle2_widths[465]), .rectangle2_height(rectangle2_heights[465]), .rectangle2_weight(rectangle2_weights[465]), .rectangle3_x(rectangle3_xs[465]), .rectangle3_y(rectangle3_ys[465]), .rectangle3_width(rectangle3_widths[465]), .rectangle3_height(rectangle3_heights[465]), .rectangle3_weight(rectangle3_weights[465]), .feature_threshold(feature_thresholds[465]), .feature_above(feature_aboves[465]), .feature_below(feature_belows[465]), .scan_win_std_dev(scan_win_std_dev[465]), .feature_accum(feature_accums[465]));
  accum_calculator ac466(.scan_win(scan_win466), .rectangle1_x(rectangle1_xs[466]), .rectangle1_y(rectangle1_ys[466]), .rectangle1_width(rectangle1_widths[466]), .rectangle1_height(rectangle1_heights[466]), .rectangle1_weight(rectangle1_weights[466]), .rectangle2_x(rectangle2_xs[466]), .rectangle2_y(rectangle2_ys[466]), .rectangle2_width(rectangle2_widths[466]), .rectangle2_height(rectangle2_heights[466]), .rectangle2_weight(rectangle2_weights[466]), .rectangle3_x(rectangle3_xs[466]), .rectangle3_y(rectangle3_ys[466]), .rectangle3_width(rectangle3_widths[466]), .rectangle3_height(rectangle3_heights[466]), .rectangle3_weight(rectangle3_weights[466]), .feature_threshold(feature_thresholds[466]), .feature_above(feature_aboves[466]), .feature_below(feature_belows[466]), .scan_win_std_dev(scan_win_std_dev[466]), .feature_accum(feature_accums[466]));
  accum_calculator ac467(.scan_win(scan_win467), .rectangle1_x(rectangle1_xs[467]), .rectangle1_y(rectangle1_ys[467]), .rectangle1_width(rectangle1_widths[467]), .rectangle1_height(rectangle1_heights[467]), .rectangle1_weight(rectangle1_weights[467]), .rectangle2_x(rectangle2_xs[467]), .rectangle2_y(rectangle2_ys[467]), .rectangle2_width(rectangle2_widths[467]), .rectangle2_height(rectangle2_heights[467]), .rectangle2_weight(rectangle2_weights[467]), .rectangle3_x(rectangle3_xs[467]), .rectangle3_y(rectangle3_ys[467]), .rectangle3_width(rectangle3_widths[467]), .rectangle3_height(rectangle3_heights[467]), .rectangle3_weight(rectangle3_weights[467]), .feature_threshold(feature_thresholds[467]), .feature_above(feature_aboves[467]), .feature_below(feature_belows[467]), .scan_win_std_dev(scan_win_std_dev[467]), .feature_accum(feature_accums[467]));
  accum_calculator ac468(.scan_win(scan_win468), .rectangle1_x(rectangle1_xs[468]), .rectangle1_y(rectangle1_ys[468]), .rectangle1_width(rectangle1_widths[468]), .rectangle1_height(rectangle1_heights[468]), .rectangle1_weight(rectangle1_weights[468]), .rectangle2_x(rectangle2_xs[468]), .rectangle2_y(rectangle2_ys[468]), .rectangle2_width(rectangle2_widths[468]), .rectangle2_height(rectangle2_heights[468]), .rectangle2_weight(rectangle2_weights[468]), .rectangle3_x(rectangle3_xs[468]), .rectangle3_y(rectangle3_ys[468]), .rectangle3_width(rectangle3_widths[468]), .rectangle3_height(rectangle3_heights[468]), .rectangle3_weight(rectangle3_weights[468]), .feature_threshold(feature_thresholds[468]), .feature_above(feature_aboves[468]), .feature_below(feature_belows[468]), .scan_win_std_dev(scan_win_std_dev[468]), .feature_accum(feature_accums[468]));
  accum_calculator ac469(.scan_win(scan_win469), .rectangle1_x(rectangle1_xs[469]), .rectangle1_y(rectangle1_ys[469]), .rectangle1_width(rectangle1_widths[469]), .rectangle1_height(rectangle1_heights[469]), .rectangle1_weight(rectangle1_weights[469]), .rectangle2_x(rectangle2_xs[469]), .rectangle2_y(rectangle2_ys[469]), .rectangle2_width(rectangle2_widths[469]), .rectangle2_height(rectangle2_heights[469]), .rectangle2_weight(rectangle2_weights[469]), .rectangle3_x(rectangle3_xs[469]), .rectangle3_y(rectangle3_ys[469]), .rectangle3_width(rectangle3_widths[469]), .rectangle3_height(rectangle3_heights[469]), .rectangle3_weight(rectangle3_weights[469]), .feature_threshold(feature_thresholds[469]), .feature_above(feature_aboves[469]), .feature_below(feature_belows[469]), .scan_win_std_dev(scan_win_std_dev[469]), .feature_accum(feature_accums[469]));
  accum_calculator ac470(.scan_win(scan_win470), .rectangle1_x(rectangle1_xs[470]), .rectangle1_y(rectangle1_ys[470]), .rectangle1_width(rectangle1_widths[470]), .rectangle1_height(rectangle1_heights[470]), .rectangle1_weight(rectangle1_weights[470]), .rectangle2_x(rectangle2_xs[470]), .rectangle2_y(rectangle2_ys[470]), .rectangle2_width(rectangle2_widths[470]), .rectangle2_height(rectangle2_heights[470]), .rectangle2_weight(rectangle2_weights[470]), .rectangle3_x(rectangle3_xs[470]), .rectangle3_y(rectangle3_ys[470]), .rectangle3_width(rectangle3_widths[470]), .rectangle3_height(rectangle3_heights[470]), .rectangle3_weight(rectangle3_weights[470]), .feature_threshold(feature_thresholds[470]), .feature_above(feature_aboves[470]), .feature_below(feature_belows[470]), .scan_win_std_dev(scan_win_std_dev[470]), .feature_accum(feature_accums[470]));
  accum_calculator ac471(.scan_win(scan_win471), .rectangle1_x(rectangle1_xs[471]), .rectangle1_y(rectangle1_ys[471]), .rectangle1_width(rectangle1_widths[471]), .rectangle1_height(rectangle1_heights[471]), .rectangle1_weight(rectangle1_weights[471]), .rectangle2_x(rectangle2_xs[471]), .rectangle2_y(rectangle2_ys[471]), .rectangle2_width(rectangle2_widths[471]), .rectangle2_height(rectangle2_heights[471]), .rectangle2_weight(rectangle2_weights[471]), .rectangle3_x(rectangle3_xs[471]), .rectangle3_y(rectangle3_ys[471]), .rectangle3_width(rectangle3_widths[471]), .rectangle3_height(rectangle3_heights[471]), .rectangle3_weight(rectangle3_weights[471]), .feature_threshold(feature_thresholds[471]), .feature_above(feature_aboves[471]), .feature_below(feature_belows[471]), .scan_win_std_dev(scan_win_std_dev[471]), .feature_accum(feature_accums[471]));
  accum_calculator ac472(.scan_win(scan_win472), .rectangle1_x(rectangle1_xs[472]), .rectangle1_y(rectangle1_ys[472]), .rectangle1_width(rectangle1_widths[472]), .rectangle1_height(rectangle1_heights[472]), .rectangle1_weight(rectangle1_weights[472]), .rectangle2_x(rectangle2_xs[472]), .rectangle2_y(rectangle2_ys[472]), .rectangle2_width(rectangle2_widths[472]), .rectangle2_height(rectangle2_heights[472]), .rectangle2_weight(rectangle2_weights[472]), .rectangle3_x(rectangle3_xs[472]), .rectangle3_y(rectangle3_ys[472]), .rectangle3_width(rectangle3_widths[472]), .rectangle3_height(rectangle3_heights[472]), .rectangle3_weight(rectangle3_weights[472]), .feature_threshold(feature_thresholds[472]), .feature_above(feature_aboves[472]), .feature_below(feature_belows[472]), .scan_win_std_dev(scan_win_std_dev[472]), .feature_accum(feature_accums[472]));
  accum_calculator ac473(.scan_win(scan_win473), .rectangle1_x(rectangle1_xs[473]), .rectangle1_y(rectangle1_ys[473]), .rectangle1_width(rectangle1_widths[473]), .rectangle1_height(rectangle1_heights[473]), .rectangle1_weight(rectangle1_weights[473]), .rectangle2_x(rectangle2_xs[473]), .rectangle2_y(rectangle2_ys[473]), .rectangle2_width(rectangle2_widths[473]), .rectangle2_height(rectangle2_heights[473]), .rectangle2_weight(rectangle2_weights[473]), .rectangle3_x(rectangle3_xs[473]), .rectangle3_y(rectangle3_ys[473]), .rectangle3_width(rectangle3_widths[473]), .rectangle3_height(rectangle3_heights[473]), .rectangle3_weight(rectangle3_weights[473]), .feature_threshold(feature_thresholds[473]), .feature_above(feature_aboves[473]), .feature_below(feature_belows[473]), .scan_win_std_dev(scan_win_std_dev[473]), .feature_accum(feature_accums[473]));
  accum_calculator ac474(.scan_win(scan_win474), .rectangle1_x(rectangle1_xs[474]), .rectangle1_y(rectangle1_ys[474]), .rectangle1_width(rectangle1_widths[474]), .rectangle1_height(rectangle1_heights[474]), .rectangle1_weight(rectangle1_weights[474]), .rectangle2_x(rectangle2_xs[474]), .rectangle2_y(rectangle2_ys[474]), .rectangle2_width(rectangle2_widths[474]), .rectangle2_height(rectangle2_heights[474]), .rectangle2_weight(rectangle2_weights[474]), .rectangle3_x(rectangle3_xs[474]), .rectangle3_y(rectangle3_ys[474]), .rectangle3_width(rectangle3_widths[474]), .rectangle3_height(rectangle3_heights[474]), .rectangle3_weight(rectangle3_weights[474]), .feature_threshold(feature_thresholds[474]), .feature_above(feature_aboves[474]), .feature_below(feature_belows[474]), .scan_win_std_dev(scan_win_std_dev[474]), .feature_accum(feature_accums[474]));
  accum_calculator ac475(.scan_win(scan_win475), .rectangle1_x(rectangle1_xs[475]), .rectangle1_y(rectangle1_ys[475]), .rectangle1_width(rectangle1_widths[475]), .rectangle1_height(rectangle1_heights[475]), .rectangle1_weight(rectangle1_weights[475]), .rectangle2_x(rectangle2_xs[475]), .rectangle2_y(rectangle2_ys[475]), .rectangle2_width(rectangle2_widths[475]), .rectangle2_height(rectangle2_heights[475]), .rectangle2_weight(rectangle2_weights[475]), .rectangle3_x(rectangle3_xs[475]), .rectangle3_y(rectangle3_ys[475]), .rectangle3_width(rectangle3_widths[475]), .rectangle3_height(rectangle3_heights[475]), .rectangle3_weight(rectangle3_weights[475]), .feature_threshold(feature_thresholds[475]), .feature_above(feature_aboves[475]), .feature_below(feature_belows[475]), .scan_win_std_dev(scan_win_std_dev[475]), .feature_accum(feature_accums[475]));
  accum_calculator ac476(.scan_win(scan_win476), .rectangle1_x(rectangle1_xs[476]), .rectangle1_y(rectangle1_ys[476]), .rectangle1_width(rectangle1_widths[476]), .rectangle1_height(rectangle1_heights[476]), .rectangle1_weight(rectangle1_weights[476]), .rectangle2_x(rectangle2_xs[476]), .rectangle2_y(rectangle2_ys[476]), .rectangle2_width(rectangle2_widths[476]), .rectangle2_height(rectangle2_heights[476]), .rectangle2_weight(rectangle2_weights[476]), .rectangle3_x(rectangle3_xs[476]), .rectangle3_y(rectangle3_ys[476]), .rectangle3_width(rectangle3_widths[476]), .rectangle3_height(rectangle3_heights[476]), .rectangle3_weight(rectangle3_weights[476]), .feature_threshold(feature_thresholds[476]), .feature_above(feature_aboves[476]), .feature_below(feature_belows[476]), .scan_win_std_dev(scan_win_std_dev[476]), .feature_accum(feature_accums[476]));
  accum_calculator ac477(.scan_win(scan_win477), .rectangle1_x(rectangle1_xs[477]), .rectangle1_y(rectangle1_ys[477]), .rectangle1_width(rectangle1_widths[477]), .rectangle1_height(rectangle1_heights[477]), .rectangle1_weight(rectangle1_weights[477]), .rectangle2_x(rectangle2_xs[477]), .rectangle2_y(rectangle2_ys[477]), .rectangle2_width(rectangle2_widths[477]), .rectangle2_height(rectangle2_heights[477]), .rectangle2_weight(rectangle2_weights[477]), .rectangle3_x(rectangle3_xs[477]), .rectangle3_y(rectangle3_ys[477]), .rectangle3_width(rectangle3_widths[477]), .rectangle3_height(rectangle3_heights[477]), .rectangle3_weight(rectangle3_weights[477]), .feature_threshold(feature_thresholds[477]), .feature_above(feature_aboves[477]), .feature_below(feature_belows[477]), .scan_win_std_dev(scan_win_std_dev[477]), .feature_accum(feature_accums[477]));
  accum_calculator ac478(.scan_win(scan_win478), .rectangle1_x(rectangle1_xs[478]), .rectangle1_y(rectangle1_ys[478]), .rectangle1_width(rectangle1_widths[478]), .rectangle1_height(rectangle1_heights[478]), .rectangle1_weight(rectangle1_weights[478]), .rectangle2_x(rectangle2_xs[478]), .rectangle2_y(rectangle2_ys[478]), .rectangle2_width(rectangle2_widths[478]), .rectangle2_height(rectangle2_heights[478]), .rectangle2_weight(rectangle2_weights[478]), .rectangle3_x(rectangle3_xs[478]), .rectangle3_y(rectangle3_ys[478]), .rectangle3_width(rectangle3_widths[478]), .rectangle3_height(rectangle3_heights[478]), .rectangle3_weight(rectangle3_weights[478]), .feature_threshold(feature_thresholds[478]), .feature_above(feature_aboves[478]), .feature_below(feature_belows[478]), .scan_win_std_dev(scan_win_std_dev[478]), .feature_accum(feature_accums[478]));
  accum_calculator ac479(.scan_win(scan_win479), .rectangle1_x(rectangle1_xs[479]), .rectangle1_y(rectangle1_ys[479]), .rectangle1_width(rectangle1_widths[479]), .rectangle1_height(rectangle1_heights[479]), .rectangle1_weight(rectangle1_weights[479]), .rectangle2_x(rectangle2_xs[479]), .rectangle2_y(rectangle2_ys[479]), .rectangle2_width(rectangle2_widths[479]), .rectangle2_height(rectangle2_heights[479]), .rectangle2_weight(rectangle2_weights[479]), .rectangle3_x(rectangle3_xs[479]), .rectangle3_y(rectangle3_ys[479]), .rectangle3_width(rectangle3_widths[479]), .rectangle3_height(rectangle3_heights[479]), .rectangle3_weight(rectangle3_weights[479]), .feature_threshold(feature_thresholds[479]), .feature_above(feature_aboves[479]), .feature_below(feature_belows[479]), .scan_win_std_dev(scan_win_std_dev[479]), .feature_accum(feature_accums[479]));
  accum_calculator ac480(.scan_win(scan_win480), .rectangle1_x(rectangle1_xs[480]), .rectangle1_y(rectangle1_ys[480]), .rectangle1_width(rectangle1_widths[480]), .rectangle1_height(rectangle1_heights[480]), .rectangle1_weight(rectangle1_weights[480]), .rectangle2_x(rectangle2_xs[480]), .rectangle2_y(rectangle2_ys[480]), .rectangle2_width(rectangle2_widths[480]), .rectangle2_height(rectangle2_heights[480]), .rectangle2_weight(rectangle2_weights[480]), .rectangle3_x(rectangle3_xs[480]), .rectangle3_y(rectangle3_ys[480]), .rectangle3_width(rectangle3_widths[480]), .rectangle3_height(rectangle3_heights[480]), .rectangle3_weight(rectangle3_weights[480]), .feature_threshold(feature_thresholds[480]), .feature_above(feature_aboves[480]), .feature_below(feature_belows[480]), .scan_win_std_dev(scan_win_std_dev[480]), .feature_accum(feature_accums[480]));
  accum_calculator ac481(.scan_win(scan_win481), .rectangle1_x(rectangle1_xs[481]), .rectangle1_y(rectangle1_ys[481]), .rectangle1_width(rectangle1_widths[481]), .rectangle1_height(rectangle1_heights[481]), .rectangle1_weight(rectangle1_weights[481]), .rectangle2_x(rectangle2_xs[481]), .rectangle2_y(rectangle2_ys[481]), .rectangle2_width(rectangle2_widths[481]), .rectangle2_height(rectangle2_heights[481]), .rectangle2_weight(rectangle2_weights[481]), .rectangle3_x(rectangle3_xs[481]), .rectangle3_y(rectangle3_ys[481]), .rectangle3_width(rectangle3_widths[481]), .rectangle3_height(rectangle3_heights[481]), .rectangle3_weight(rectangle3_weights[481]), .feature_threshold(feature_thresholds[481]), .feature_above(feature_aboves[481]), .feature_below(feature_belows[481]), .scan_win_std_dev(scan_win_std_dev[481]), .feature_accum(feature_accums[481]));
  accum_calculator ac482(.scan_win(scan_win482), .rectangle1_x(rectangle1_xs[482]), .rectangle1_y(rectangle1_ys[482]), .rectangle1_width(rectangle1_widths[482]), .rectangle1_height(rectangle1_heights[482]), .rectangle1_weight(rectangle1_weights[482]), .rectangle2_x(rectangle2_xs[482]), .rectangle2_y(rectangle2_ys[482]), .rectangle2_width(rectangle2_widths[482]), .rectangle2_height(rectangle2_heights[482]), .rectangle2_weight(rectangle2_weights[482]), .rectangle3_x(rectangle3_xs[482]), .rectangle3_y(rectangle3_ys[482]), .rectangle3_width(rectangle3_widths[482]), .rectangle3_height(rectangle3_heights[482]), .rectangle3_weight(rectangle3_weights[482]), .feature_threshold(feature_thresholds[482]), .feature_above(feature_aboves[482]), .feature_below(feature_belows[482]), .scan_win_std_dev(scan_win_std_dev[482]), .feature_accum(feature_accums[482]));
  accum_calculator ac483(.scan_win(scan_win483), .rectangle1_x(rectangle1_xs[483]), .rectangle1_y(rectangle1_ys[483]), .rectangle1_width(rectangle1_widths[483]), .rectangle1_height(rectangle1_heights[483]), .rectangle1_weight(rectangle1_weights[483]), .rectangle2_x(rectangle2_xs[483]), .rectangle2_y(rectangle2_ys[483]), .rectangle2_width(rectangle2_widths[483]), .rectangle2_height(rectangle2_heights[483]), .rectangle2_weight(rectangle2_weights[483]), .rectangle3_x(rectangle3_xs[483]), .rectangle3_y(rectangle3_ys[483]), .rectangle3_width(rectangle3_widths[483]), .rectangle3_height(rectangle3_heights[483]), .rectangle3_weight(rectangle3_weights[483]), .feature_threshold(feature_thresholds[483]), .feature_above(feature_aboves[483]), .feature_below(feature_belows[483]), .scan_win_std_dev(scan_win_std_dev[483]), .feature_accum(feature_accums[483]));
  accum_calculator ac484(.scan_win(scan_win484), .rectangle1_x(rectangle1_xs[484]), .rectangle1_y(rectangle1_ys[484]), .rectangle1_width(rectangle1_widths[484]), .rectangle1_height(rectangle1_heights[484]), .rectangle1_weight(rectangle1_weights[484]), .rectangle2_x(rectangle2_xs[484]), .rectangle2_y(rectangle2_ys[484]), .rectangle2_width(rectangle2_widths[484]), .rectangle2_height(rectangle2_heights[484]), .rectangle2_weight(rectangle2_weights[484]), .rectangle3_x(rectangle3_xs[484]), .rectangle3_y(rectangle3_ys[484]), .rectangle3_width(rectangle3_widths[484]), .rectangle3_height(rectangle3_heights[484]), .rectangle3_weight(rectangle3_weights[484]), .feature_threshold(feature_thresholds[484]), .feature_above(feature_aboves[484]), .feature_below(feature_belows[484]), .scan_win_std_dev(scan_win_std_dev[484]), .feature_accum(feature_accums[484]));
  accum_calculator ac485(.scan_win(scan_win485), .rectangle1_x(rectangle1_xs[485]), .rectangle1_y(rectangle1_ys[485]), .rectangle1_width(rectangle1_widths[485]), .rectangle1_height(rectangle1_heights[485]), .rectangle1_weight(rectangle1_weights[485]), .rectangle2_x(rectangle2_xs[485]), .rectangle2_y(rectangle2_ys[485]), .rectangle2_width(rectangle2_widths[485]), .rectangle2_height(rectangle2_heights[485]), .rectangle2_weight(rectangle2_weights[485]), .rectangle3_x(rectangle3_xs[485]), .rectangle3_y(rectangle3_ys[485]), .rectangle3_width(rectangle3_widths[485]), .rectangle3_height(rectangle3_heights[485]), .rectangle3_weight(rectangle3_weights[485]), .feature_threshold(feature_thresholds[485]), .feature_above(feature_aboves[485]), .feature_below(feature_belows[485]), .scan_win_std_dev(scan_win_std_dev[485]), .feature_accum(feature_accums[485]));
  accum_calculator ac486(.scan_win(scan_win486), .rectangle1_x(rectangle1_xs[486]), .rectangle1_y(rectangle1_ys[486]), .rectangle1_width(rectangle1_widths[486]), .rectangle1_height(rectangle1_heights[486]), .rectangle1_weight(rectangle1_weights[486]), .rectangle2_x(rectangle2_xs[486]), .rectangle2_y(rectangle2_ys[486]), .rectangle2_width(rectangle2_widths[486]), .rectangle2_height(rectangle2_heights[486]), .rectangle2_weight(rectangle2_weights[486]), .rectangle3_x(rectangle3_xs[486]), .rectangle3_y(rectangle3_ys[486]), .rectangle3_width(rectangle3_widths[486]), .rectangle3_height(rectangle3_heights[486]), .rectangle3_weight(rectangle3_weights[486]), .feature_threshold(feature_thresholds[486]), .feature_above(feature_aboves[486]), .feature_below(feature_belows[486]), .scan_win_std_dev(scan_win_std_dev[486]), .feature_accum(feature_accums[486]));
  accum_calculator ac487(.scan_win(scan_win487), .rectangle1_x(rectangle1_xs[487]), .rectangle1_y(rectangle1_ys[487]), .rectangle1_width(rectangle1_widths[487]), .rectangle1_height(rectangle1_heights[487]), .rectangle1_weight(rectangle1_weights[487]), .rectangle2_x(rectangle2_xs[487]), .rectangle2_y(rectangle2_ys[487]), .rectangle2_width(rectangle2_widths[487]), .rectangle2_height(rectangle2_heights[487]), .rectangle2_weight(rectangle2_weights[487]), .rectangle3_x(rectangle3_xs[487]), .rectangle3_y(rectangle3_ys[487]), .rectangle3_width(rectangle3_widths[487]), .rectangle3_height(rectangle3_heights[487]), .rectangle3_weight(rectangle3_weights[487]), .feature_threshold(feature_thresholds[487]), .feature_above(feature_aboves[487]), .feature_below(feature_belows[487]), .scan_win_std_dev(scan_win_std_dev[487]), .feature_accum(feature_accums[487]));
  accum_calculator ac488(.scan_win(scan_win488), .rectangle1_x(rectangle1_xs[488]), .rectangle1_y(rectangle1_ys[488]), .rectangle1_width(rectangle1_widths[488]), .rectangle1_height(rectangle1_heights[488]), .rectangle1_weight(rectangle1_weights[488]), .rectangle2_x(rectangle2_xs[488]), .rectangle2_y(rectangle2_ys[488]), .rectangle2_width(rectangle2_widths[488]), .rectangle2_height(rectangle2_heights[488]), .rectangle2_weight(rectangle2_weights[488]), .rectangle3_x(rectangle3_xs[488]), .rectangle3_y(rectangle3_ys[488]), .rectangle3_width(rectangle3_widths[488]), .rectangle3_height(rectangle3_heights[488]), .rectangle3_weight(rectangle3_weights[488]), .feature_threshold(feature_thresholds[488]), .feature_above(feature_aboves[488]), .feature_below(feature_belows[488]), .scan_win_std_dev(scan_win_std_dev[488]), .feature_accum(feature_accums[488]));
  accum_calculator ac489(.scan_win(scan_win489), .rectangle1_x(rectangle1_xs[489]), .rectangle1_y(rectangle1_ys[489]), .rectangle1_width(rectangle1_widths[489]), .rectangle1_height(rectangle1_heights[489]), .rectangle1_weight(rectangle1_weights[489]), .rectangle2_x(rectangle2_xs[489]), .rectangle2_y(rectangle2_ys[489]), .rectangle2_width(rectangle2_widths[489]), .rectangle2_height(rectangle2_heights[489]), .rectangle2_weight(rectangle2_weights[489]), .rectangle3_x(rectangle3_xs[489]), .rectangle3_y(rectangle3_ys[489]), .rectangle3_width(rectangle3_widths[489]), .rectangle3_height(rectangle3_heights[489]), .rectangle3_weight(rectangle3_weights[489]), .feature_threshold(feature_thresholds[489]), .feature_above(feature_aboves[489]), .feature_below(feature_belows[489]), .scan_win_std_dev(scan_win_std_dev[489]), .feature_accum(feature_accums[489]));
  accum_calculator ac490(.scan_win(scan_win490), .rectangle1_x(rectangle1_xs[490]), .rectangle1_y(rectangle1_ys[490]), .rectangle1_width(rectangle1_widths[490]), .rectangle1_height(rectangle1_heights[490]), .rectangle1_weight(rectangle1_weights[490]), .rectangle2_x(rectangle2_xs[490]), .rectangle2_y(rectangle2_ys[490]), .rectangle2_width(rectangle2_widths[490]), .rectangle2_height(rectangle2_heights[490]), .rectangle2_weight(rectangle2_weights[490]), .rectangle3_x(rectangle3_xs[490]), .rectangle3_y(rectangle3_ys[490]), .rectangle3_width(rectangle3_widths[490]), .rectangle3_height(rectangle3_heights[490]), .rectangle3_weight(rectangle3_weights[490]), .feature_threshold(feature_thresholds[490]), .feature_above(feature_aboves[490]), .feature_below(feature_belows[490]), .scan_win_std_dev(scan_win_std_dev[490]), .feature_accum(feature_accums[490]));
  accum_calculator ac491(.scan_win(scan_win491), .rectangle1_x(rectangle1_xs[491]), .rectangle1_y(rectangle1_ys[491]), .rectangle1_width(rectangle1_widths[491]), .rectangle1_height(rectangle1_heights[491]), .rectangle1_weight(rectangle1_weights[491]), .rectangle2_x(rectangle2_xs[491]), .rectangle2_y(rectangle2_ys[491]), .rectangle2_width(rectangle2_widths[491]), .rectangle2_height(rectangle2_heights[491]), .rectangle2_weight(rectangle2_weights[491]), .rectangle3_x(rectangle3_xs[491]), .rectangle3_y(rectangle3_ys[491]), .rectangle3_width(rectangle3_widths[491]), .rectangle3_height(rectangle3_heights[491]), .rectangle3_weight(rectangle3_weights[491]), .feature_threshold(feature_thresholds[491]), .feature_above(feature_aboves[491]), .feature_below(feature_belows[491]), .scan_win_std_dev(scan_win_std_dev[491]), .feature_accum(feature_accums[491]));
  accum_calculator ac492(.scan_win(scan_win492), .rectangle1_x(rectangle1_xs[492]), .rectangle1_y(rectangle1_ys[492]), .rectangle1_width(rectangle1_widths[492]), .rectangle1_height(rectangle1_heights[492]), .rectangle1_weight(rectangle1_weights[492]), .rectangle2_x(rectangle2_xs[492]), .rectangle2_y(rectangle2_ys[492]), .rectangle2_width(rectangle2_widths[492]), .rectangle2_height(rectangle2_heights[492]), .rectangle2_weight(rectangle2_weights[492]), .rectangle3_x(rectangle3_xs[492]), .rectangle3_y(rectangle3_ys[492]), .rectangle3_width(rectangle3_widths[492]), .rectangle3_height(rectangle3_heights[492]), .rectangle3_weight(rectangle3_weights[492]), .feature_threshold(feature_thresholds[492]), .feature_above(feature_aboves[492]), .feature_below(feature_belows[492]), .scan_win_std_dev(scan_win_std_dev[492]), .feature_accum(feature_accums[492]));
  accum_calculator ac493(.scan_win(scan_win493), .rectangle1_x(rectangle1_xs[493]), .rectangle1_y(rectangle1_ys[493]), .rectangle1_width(rectangle1_widths[493]), .rectangle1_height(rectangle1_heights[493]), .rectangle1_weight(rectangle1_weights[493]), .rectangle2_x(rectangle2_xs[493]), .rectangle2_y(rectangle2_ys[493]), .rectangle2_width(rectangle2_widths[493]), .rectangle2_height(rectangle2_heights[493]), .rectangle2_weight(rectangle2_weights[493]), .rectangle3_x(rectangle3_xs[493]), .rectangle3_y(rectangle3_ys[493]), .rectangle3_width(rectangle3_widths[493]), .rectangle3_height(rectangle3_heights[493]), .rectangle3_weight(rectangle3_weights[493]), .feature_threshold(feature_thresholds[493]), .feature_above(feature_aboves[493]), .feature_below(feature_belows[493]), .scan_win_std_dev(scan_win_std_dev[493]), .feature_accum(feature_accums[493]));
  accum_calculator ac494(.scan_win(scan_win494), .rectangle1_x(rectangle1_xs[494]), .rectangle1_y(rectangle1_ys[494]), .rectangle1_width(rectangle1_widths[494]), .rectangle1_height(rectangle1_heights[494]), .rectangle1_weight(rectangle1_weights[494]), .rectangle2_x(rectangle2_xs[494]), .rectangle2_y(rectangle2_ys[494]), .rectangle2_width(rectangle2_widths[494]), .rectangle2_height(rectangle2_heights[494]), .rectangle2_weight(rectangle2_weights[494]), .rectangle3_x(rectangle3_xs[494]), .rectangle3_y(rectangle3_ys[494]), .rectangle3_width(rectangle3_widths[494]), .rectangle3_height(rectangle3_heights[494]), .rectangle3_weight(rectangle3_weights[494]), .feature_threshold(feature_thresholds[494]), .feature_above(feature_aboves[494]), .feature_below(feature_belows[494]), .scan_win_std_dev(scan_win_std_dev[494]), .feature_accum(feature_accums[494]));
  accum_calculator ac495(.scan_win(scan_win495), .rectangle1_x(rectangle1_xs[495]), .rectangle1_y(rectangle1_ys[495]), .rectangle1_width(rectangle1_widths[495]), .rectangle1_height(rectangle1_heights[495]), .rectangle1_weight(rectangle1_weights[495]), .rectangle2_x(rectangle2_xs[495]), .rectangle2_y(rectangle2_ys[495]), .rectangle2_width(rectangle2_widths[495]), .rectangle2_height(rectangle2_heights[495]), .rectangle2_weight(rectangle2_weights[495]), .rectangle3_x(rectangle3_xs[495]), .rectangle3_y(rectangle3_ys[495]), .rectangle3_width(rectangle3_widths[495]), .rectangle3_height(rectangle3_heights[495]), .rectangle3_weight(rectangle3_weights[495]), .feature_threshold(feature_thresholds[495]), .feature_above(feature_aboves[495]), .feature_below(feature_belows[495]), .scan_win_std_dev(scan_win_std_dev[495]), .feature_accum(feature_accums[495]));
  accum_calculator ac496(.scan_win(scan_win496), .rectangle1_x(rectangle1_xs[496]), .rectangle1_y(rectangle1_ys[496]), .rectangle1_width(rectangle1_widths[496]), .rectangle1_height(rectangle1_heights[496]), .rectangle1_weight(rectangle1_weights[496]), .rectangle2_x(rectangle2_xs[496]), .rectangle2_y(rectangle2_ys[496]), .rectangle2_width(rectangle2_widths[496]), .rectangle2_height(rectangle2_heights[496]), .rectangle2_weight(rectangle2_weights[496]), .rectangle3_x(rectangle3_xs[496]), .rectangle3_y(rectangle3_ys[496]), .rectangle3_width(rectangle3_widths[496]), .rectangle3_height(rectangle3_heights[496]), .rectangle3_weight(rectangle3_weights[496]), .feature_threshold(feature_thresholds[496]), .feature_above(feature_aboves[496]), .feature_below(feature_belows[496]), .scan_win_std_dev(scan_win_std_dev[496]), .feature_accum(feature_accums[496]));
  accum_calculator ac497(.scan_win(scan_win497), .rectangle1_x(rectangle1_xs[497]), .rectangle1_y(rectangle1_ys[497]), .rectangle1_width(rectangle1_widths[497]), .rectangle1_height(rectangle1_heights[497]), .rectangle1_weight(rectangle1_weights[497]), .rectangle2_x(rectangle2_xs[497]), .rectangle2_y(rectangle2_ys[497]), .rectangle2_width(rectangle2_widths[497]), .rectangle2_height(rectangle2_heights[497]), .rectangle2_weight(rectangle2_weights[497]), .rectangle3_x(rectangle3_xs[497]), .rectangle3_y(rectangle3_ys[497]), .rectangle3_width(rectangle3_widths[497]), .rectangle3_height(rectangle3_heights[497]), .rectangle3_weight(rectangle3_weights[497]), .feature_threshold(feature_thresholds[497]), .feature_above(feature_aboves[497]), .feature_below(feature_belows[497]), .scan_win_std_dev(scan_win_std_dev[497]), .feature_accum(feature_accums[497]));
  accum_calculator ac498(.scan_win(scan_win498), .rectangle1_x(rectangle1_xs[498]), .rectangle1_y(rectangle1_ys[498]), .rectangle1_width(rectangle1_widths[498]), .rectangle1_height(rectangle1_heights[498]), .rectangle1_weight(rectangle1_weights[498]), .rectangle2_x(rectangle2_xs[498]), .rectangle2_y(rectangle2_ys[498]), .rectangle2_width(rectangle2_widths[498]), .rectangle2_height(rectangle2_heights[498]), .rectangle2_weight(rectangle2_weights[498]), .rectangle3_x(rectangle3_xs[498]), .rectangle3_y(rectangle3_ys[498]), .rectangle3_width(rectangle3_widths[498]), .rectangle3_height(rectangle3_heights[498]), .rectangle3_weight(rectangle3_weights[498]), .feature_threshold(feature_thresholds[498]), .feature_above(feature_aboves[498]), .feature_below(feature_belows[498]), .scan_win_std_dev(scan_win_std_dev[498]), .feature_accum(feature_accums[498]));
  accum_calculator ac499(.scan_win(scan_win499), .rectangle1_x(rectangle1_xs[499]), .rectangle1_y(rectangle1_ys[499]), .rectangle1_width(rectangle1_widths[499]), .rectangle1_height(rectangle1_heights[499]), .rectangle1_weight(rectangle1_weights[499]), .rectangle2_x(rectangle2_xs[499]), .rectangle2_y(rectangle2_ys[499]), .rectangle2_width(rectangle2_widths[499]), .rectangle2_height(rectangle2_heights[499]), .rectangle2_weight(rectangle2_weights[499]), .rectangle3_x(rectangle3_xs[499]), .rectangle3_y(rectangle3_ys[499]), .rectangle3_width(rectangle3_widths[499]), .rectangle3_height(rectangle3_heights[499]), .rectangle3_weight(rectangle3_weights[499]), .feature_threshold(feature_thresholds[499]), .feature_above(feature_aboves[499]), .feature_below(feature_belows[499]), .scan_win_std_dev(scan_win_std_dev[499]), .feature_accum(feature_accums[499]));
  accum_calculator ac500(.scan_win(scan_win500), .rectangle1_x(rectangle1_xs[500]), .rectangle1_y(rectangle1_ys[500]), .rectangle1_width(rectangle1_widths[500]), .rectangle1_height(rectangle1_heights[500]), .rectangle1_weight(rectangle1_weights[500]), .rectangle2_x(rectangle2_xs[500]), .rectangle2_y(rectangle2_ys[500]), .rectangle2_width(rectangle2_widths[500]), .rectangle2_height(rectangle2_heights[500]), .rectangle2_weight(rectangle2_weights[500]), .rectangle3_x(rectangle3_xs[500]), .rectangle3_y(rectangle3_ys[500]), .rectangle3_width(rectangle3_widths[500]), .rectangle3_height(rectangle3_heights[500]), .rectangle3_weight(rectangle3_weights[500]), .feature_threshold(feature_thresholds[500]), .feature_above(feature_aboves[500]), .feature_below(feature_belows[500]), .scan_win_std_dev(scan_win_std_dev[500]), .feature_accum(feature_accums[500]));
  accum_calculator ac501(.scan_win(scan_win501), .rectangle1_x(rectangle1_xs[501]), .rectangle1_y(rectangle1_ys[501]), .rectangle1_width(rectangle1_widths[501]), .rectangle1_height(rectangle1_heights[501]), .rectangle1_weight(rectangle1_weights[501]), .rectangle2_x(rectangle2_xs[501]), .rectangle2_y(rectangle2_ys[501]), .rectangle2_width(rectangle2_widths[501]), .rectangle2_height(rectangle2_heights[501]), .rectangle2_weight(rectangle2_weights[501]), .rectangle3_x(rectangle3_xs[501]), .rectangle3_y(rectangle3_ys[501]), .rectangle3_width(rectangle3_widths[501]), .rectangle3_height(rectangle3_heights[501]), .rectangle3_weight(rectangle3_weights[501]), .feature_threshold(feature_thresholds[501]), .feature_above(feature_aboves[501]), .feature_below(feature_belows[501]), .scan_win_std_dev(scan_win_std_dev[501]), .feature_accum(feature_accums[501]));
  accum_calculator ac502(.scan_win(scan_win502), .rectangle1_x(rectangle1_xs[502]), .rectangle1_y(rectangle1_ys[502]), .rectangle1_width(rectangle1_widths[502]), .rectangle1_height(rectangle1_heights[502]), .rectangle1_weight(rectangle1_weights[502]), .rectangle2_x(rectangle2_xs[502]), .rectangle2_y(rectangle2_ys[502]), .rectangle2_width(rectangle2_widths[502]), .rectangle2_height(rectangle2_heights[502]), .rectangle2_weight(rectangle2_weights[502]), .rectangle3_x(rectangle3_xs[502]), .rectangle3_y(rectangle3_ys[502]), .rectangle3_width(rectangle3_widths[502]), .rectangle3_height(rectangle3_heights[502]), .rectangle3_weight(rectangle3_weights[502]), .feature_threshold(feature_thresholds[502]), .feature_above(feature_aboves[502]), .feature_below(feature_belows[502]), .scan_win_std_dev(scan_win_std_dev[502]), .feature_accum(feature_accums[502]));
  accum_calculator ac503(.scan_win(scan_win503), .rectangle1_x(rectangle1_xs[503]), .rectangle1_y(rectangle1_ys[503]), .rectangle1_width(rectangle1_widths[503]), .rectangle1_height(rectangle1_heights[503]), .rectangle1_weight(rectangle1_weights[503]), .rectangle2_x(rectangle2_xs[503]), .rectangle2_y(rectangle2_ys[503]), .rectangle2_width(rectangle2_widths[503]), .rectangle2_height(rectangle2_heights[503]), .rectangle2_weight(rectangle2_weights[503]), .rectangle3_x(rectangle3_xs[503]), .rectangle3_y(rectangle3_ys[503]), .rectangle3_width(rectangle3_widths[503]), .rectangle3_height(rectangle3_heights[503]), .rectangle3_weight(rectangle3_weights[503]), .feature_threshold(feature_thresholds[503]), .feature_above(feature_aboves[503]), .feature_below(feature_belows[503]), .scan_win_std_dev(scan_win_std_dev[503]), .feature_accum(feature_accums[503]));
  accum_calculator ac504(.scan_win(scan_win504), .rectangle1_x(rectangle1_xs[504]), .rectangle1_y(rectangle1_ys[504]), .rectangle1_width(rectangle1_widths[504]), .rectangle1_height(rectangle1_heights[504]), .rectangle1_weight(rectangle1_weights[504]), .rectangle2_x(rectangle2_xs[504]), .rectangle2_y(rectangle2_ys[504]), .rectangle2_width(rectangle2_widths[504]), .rectangle2_height(rectangle2_heights[504]), .rectangle2_weight(rectangle2_weights[504]), .rectangle3_x(rectangle3_xs[504]), .rectangle3_y(rectangle3_ys[504]), .rectangle3_width(rectangle3_widths[504]), .rectangle3_height(rectangle3_heights[504]), .rectangle3_weight(rectangle3_weights[504]), .feature_threshold(feature_thresholds[504]), .feature_above(feature_aboves[504]), .feature_below(feature_belows[504]), .scan_win_std_dev(scan_win_std_dev[504]), .feature_accum(feature_accums[504]));
  accum_calculator ac505(.scan_win(scan_win505), .rectangle1_x(rectangle1_xs[505]), .rectangle1_y(rectangle1_ys[505]), .rectangle1_width(rectangle1_widths[505]), .rectangle1_height(rectangle1_heights[505]), .rectangle1_weight(rectangle1_weights[505]), .rectangle2_x(rectangle2_xs[505]), .rectangle2_y(rectangle2_ys[505]), .rectangle2_width(rectangle2_widths[505]), .rectangle2_height(rectangle2_heights[505]), .rectangle2_weight(rectangle2_weights[505]), .rectangle3_x(rectangle3_xs[505]), .rectangle3_y(rectangle3_ys[505]), .rectangle3_width(rectangle3_widths[505]), .rectangle3_height(rectangle3_heights[505]), .rectangle3_weight(rectangle3_weights[505]), .feature_threshold(feature_thresholds[505]), .feature_above(feature_aboves[505]), .feature_below(feature_belows[505]), .scan_win_std_dev(scan_win_std_dev[505]), .feature_accum(feature_accums[505]));
  accum_calculator ac506(.scan_win(scan_win506), .rectangle1_x(rectangle1_xs[506]), .rectangle1_y(rectangle1_ys[506]), .rectangle1_width(rectangle1_widths[506]), .rectangle1_height(rectangle1_heights[506]), .rectangle1_weight(rectangle1_weights[506]), .rectangle2_x(rectangle2_xs[506]), .rectangle2_y(rectangle2_ys[506]), .rectangle2_width(rectangle2_widths[506]), .rectangle2_height(rectangle2_heights[506]), .rectangle2_weight(rectangle2_weights[506]), .rectangle3_x(rectangle3_xs[506]), .rectangle3_y(rectangle3_ys[506]), .rectangle3_width(rectangle3_widths[506]), .rectangle3_height(rectangle3_heights[506]), .rectangle3_weight(rectangle3_weights[506]), .feature_threshold(feature_thresholds[506]), .feature_above(feature_aboves[506]), .feature_below(feature_belows[506]), .scan_win_std_dev(scan_win_std_dev[506]), .feature_accum(feature_accums[506]));
  accum_calculator ac507(.scan_win(scan_win507), .rectangle1_x(rectangle1_xs[507]), .rectangle1_y(rectangle1_ys[507]), .rectangle1_width(rectangle1_widths[507]), .rectangle1_height(rectangle1_heights[507]), .rectangle1_weight(rectangle1_weights[507]), .rectangle2_x(rectangle2_xs[507]), .rectangle2_y(rectangle2_ys[507]), .rectangle2_width(rectangle2_widths[507]), .rectangle2_height(rectangle2_heights[507]), .rectangle2_weight(rectangle2_weights[507]), .rectangle3_x(rectangle3_xs[507]), .rectangle3_y(rectangle3_ys[507]), .rectangle3_width(rectangle3_widths[507]), .rectangle3_height(rectangle3_heights[507]), .rectangle3_weight(rectangle3_weights[507]), .feature_threshold(feature_thresholds[507]), .feature_above(feature_aboves[507]), .feature_below(feature_belows[507]), .scan_win_std_dev(scan_win_std_dev[507]), .feature_accum(feature_accums[507]));
  accum_calculator ac508(.scan_win(scan_win508), .rectangle1_x(rectangle1_xs[508]), .rectangle1_y(rectangle1_ys[508]), .rectangle1_width(rectangle1_widths[508]), .rectangle1_height(rectangle1_heights[508]), .rectangle1_weight(rectangle1_weights[508]), .rectangle2_x(rectangle2_xs[508]), .rectangle2_y(rectangle2_ys[508]), .rectangle2_width(rectangle2_widths[508]), .rectangle2_height(rectangle2_heights[508]), .rectangle2_weight(rectangle2_weights[508]), .rectangle3_x(rectangle3_xs[508]), .rectangle3_y(rectangle3_ys[508]), .rectangle3_width(rectangle3_widths[508]), .rectangle3_height(rectangle3_heights[508]), .rectangle3_weight(rectangle3_weights[508]), .feature_threshold(feature_thresholds[508]), .feature_above(feature_aboves[508]), .feature_below(feature_belows[508]), .scan_win_std_dev(scan_win_std_dev[508]), .feature_accum(feature_accums[508]));
  accum_calculator ac509(.scan_win(scan_win509), .rectangle1_x(rectangle1_xs[509]), .rectangle1_y(rectangle1_ys[509]), .rectangle1_width(rectangle1_widths[509]), .rectangle1_height(rectangle1_heights[509]), .rectangle1_weight(rectangle1_weights[509]), .rectangle2_x(rectangle2_xs[509]), .rectangle2_y(rectangle2_ys[509]), .rectangle2_width(rectangle2_widths[509]), .rectangle2_height(rectangle2_heights[509]), .rectangle2_weight(rectangle2_weights[509]), .rectangle3_x(rectangle3_xs[509]), .rectangle3_y(rectangle3_ys[509]), .rectangle3_width(rectangle3_widths[509]), .rectangle3_height(rectangle3_heights[509]), .rectangle3_weight(rectangle3_weights[509]), .feature_threshold(feature_thresholds[509]), .feature_above(feature_aboves[509]), .feature_below(feature_belows[509]), .scan_win_std_dev(scan_win_std_dev[509]), .feature_accum(feature_accums[509]));
  accum_calculator ac510(.scan_win(scan_win510), .rectangle1_x(rectangle1_xs[510]), .rectangle1_y(rectangle1_ys[510]), .rectangle1_width(rectangle1_widths[510]), .rectangle1_height(rectangle1_heights[510]), .rectangle1_weight(rectangle1_weights[510]), .rectangle2_x(rectangle2_xs[510]), .rectangle2_y(rectangle2_ys[510]), .rectangle2_width(rectangle2_widths[510]), .rectangle2_height(rectangle2_heights[510]), .rectangle2_weight(rectangle2_weights[510]), .rectangle3_x(rectangle3_xs[510]), .rectangle3_y(rectangle3_ys[510]), .rectangle3_width(rectangle3_widths[510]), .rectangle3_height(rectangle3_heights[510]), .rectangle3_weight(rectangle3_weights[510]), .feature_threshold(feature_thresholds[510]), .feature_above(feature_aboves[510]), .feature_below(feature_belows[510]), .scan_win_std_dev(scan_win_std_dev[510]), .feature_accum(feature_accums[510]));
  accum_calculator ac511(.scan_win(scan_win511), .rectangle1_x(rectangle1_xs[511]), .rectangle1_y(rectangle1_ys[511]), .rectangle1_width(rectangle1_widths[511]), .rectangle1_height(rectangle1_heights[511]), .rectangle1_weight(rectangle1_weights[511]), .rectangle2_x(rectangle2_xs[511]), .rectangle2_y(rectangle2_ys[511]), .rectangle2_width(rectangle2_widths[511]), .rectangle2_height(rectangle2_heights[511]), .rectangle2_weight(rectangle2_weights[511]), .rectangle3_x(rectangle3_xs[511]), .rectangle3_y(rectangle3_ys[511]), .rectangle3_width(rectangle3_widths[511]), .rectangle3_height(rectangle3_heights[511]), .rectangle3_weight(rectangle3_weights[511]), .feature_threshold(feature_thresholds[511]), .feature_above(feature_aboves[511]), .feature_below(feature_belows[511]), .scan_win_std_dev(scan_win_std_dev[511]), .feature_accum(feature_accums[511]));
  accum_calculator ac512(.scan_win(scan_win512), .rectangle1_x(rectangle1_xs[512]), .rectangle1_y(rectangle1_ys[512]), .rectangle1_width(rectangle1_widths[512]), .rectangle1_height(rectangle1_heights[512]), .rectangle1_weight(rectangle1_weights[512]), .rectangle2_x(rectangle2_xs[512]), .rectangle2_y(rectangle2_ys[512]), .rectangle2_width(rectangle2_widths[512]), .rectangle2_height(rectangle2_heights[512]), .rectangle2_weight(rectangle2_weights[512]), .rectangle3_x(rectangle3_xs[512]), .rectangle3_y(rectangle3_ys[512]), .rectangle3_width(rectangle3_widths[512]), .rectangle3_height(rectangle3_heights[512]), .rectangle3_weight(rectangle3_weights[512]), .feature_threshold(feature_thresholds[512]), .feature_above(feature_aboves[512]), .feature_below(feature_belows[512]), .scan_win_std_dev(scan_win_std_dev[512]), .feature_accum(feature_accums[512]));
  accum_calculator ac513(.scan_win(scan_win513), .rectangle1_x(rectangle1_xs[513]), .rectangle1_y(rectangle1_ys[513]), .rectangle1_width(rectangle1_widths[513]), .rectangle1_height(rectangle1_heights[513]), .rectangle1_weight(rectangle1_weights[513]), .rectangle2_x(rectangle2_xs[513]), .rectangle2_y(rectangle2_ys[513]), .rectangle2_width(rectangle2_widths[513]), .rectangle2_height(rectangle2_heights[513]), .rectangle2_weight(rectangle2_weights[513]), .rectangle3_x(rectangle3_xs[513]), .rectangle3_y(rectangle3_ys[513]), .rectangle3_width(rectangle3_widths[513]), .rectangle3_height(rectangle3_heights[513]), .rectangle3_weight(rectangle3_weights[513]), .feature_threshold(feature_thresholds[513]), .feature_above(feature_aboves[513]), .feature_below(feature_belows[513]), .scan_win_std_dev(scan_win_std_dev[513]), .feature_accum(feature_accums[513]));
  accum_calculator ac514(.scan_win(scan_win514), .rectangle1_x(rectangle1_xs[514]), .rectangle1_y(rectangle1_ys[514]), .rectangle1_width(rectangle1_widths[514]), .rectangle1_height(rectangle1_heights[514]), .rectangle1_weight(rectangle1_weights[514]), .rectangle2_x(rectangle2_xs[514]), .rectangle2_y(rectangle2_ys[514]), .rectangle2_width(rectangle2_widths[514]), .rectangle2_height(rectangle2_heights[514]), .rectangle2_weight(rectangle2_weights[514]), .rectangle3_x(rectangle3_xs[514]), .rectangle3_y(rectangle3_ys[514]), .rectangle3_width(rectangle3_widths[514]), .rectangle3_height(rectangle3_heights[514]), .rectangle3_weight(rectangle3_weights[514]), .feature_threshold(feature_thresholds[514]), .feature_above(feature_aboves[514]), .feature_below(feature_belows[514]), .scan_win_std_dev(scan_win_std_dev[514]), .feature_accum(feature_accums[514]));
  accum_calculator ac515(.scan_win(scan_win515), .rectangle1_x(rectangle1_xs[515]), .rectangle1_y(rectangle1_ys[515]), .rectangle1_width(rectangle1_widths[515]), .rectangle1_height(rectangle1_heights[515]), .rectangle1_weight(rectangle1_weights[515]), .rectangle2_x(rectangle2_xs[515]), .rectangle2_y(rectangle2_ys[515]), .rectangle2_width(rectangle2_widths[515]), .rectangle2_height(rectangle2_heights[515]), .rectangle2_weight(rectangle2_weights[515]), .rectangle3_x(rectangle3_xs[515]), .rectangle3_y(rectangle3_ys[515]), .rectangle3_width(rectangle3_widths[515]), .rectangle3_height(rectangle3_heights[515]), .rectangle3_weight(rectangle3_weights[515]), .feature_threshold(feature_thresholds[515]), .feature_above(feature_aboves[515]), .feature_below(feature_belows[515]), .scan_win_std_dev(scan_win_std_dev[515]), .feature_accum(feature_accums[515]));
  accum_calculator ac516(.scan_win(scan_win516), .rectangle1_x(rectangle1_xs[516]), .rectangle1_y(rectangle1_ys[516]), .rectangle1_width(rectangle1_widths[516]), .rectangle1_height(rectangle1_heights[516]), .rectangle1_weight(rectangle1_weights[516]), .rectangle2_x(rectangle2_xs[516]), .rectangle2_y(rectangle2_ys[516]), .rectangle2_width(rectangle2_widths[516]), .rectangle2_height(rectangle2_heights[516]), .rectangle2_weight(rectangle2_weights[516]), .rectangle3_x(rectangle3_xs[516]), .rectangle3_y(rectangle3_ys[516]), .rectangle3_width(rectangle3_widths[516]), .rectangle3_height(rectangle3_heights[516]), .rectangle3_weight(rectangle3_weights[516]), .feature_threshold(feature_thresholds[516]), .feature_above(feature_aboves[516]), .feature_below(feature_belows[516]), .scan_win_std_dev(scan_win_std_dev[516]), .feature_accum(feature_accums[516]));
  accum_calculator ac517(.scan_win(scan_win517), .rectangle1_x(rectangle1_xs[517]), .rectangle1_y(rectangle1_ys[517]), .rectangle1_width(rectangle1_widths[517]), .rectangle1_height(rectangle1_heights[517]), .rectangle1_weight(rectangle1_weights[517]), .rectangle2_x(rectangle2_xs[517]), .rectangle2_y(rectangle2_ys[517]), .rectangle2_width(rectangle2_widths[517]), .rectangle2_height(rectangle2_heights[517]), .rectangle2_weight(rectangle2_weights[517]), .rectangle3_x(rectangle3_xs[517]), .rectangle3_y(rectangle3_ys[517]), .rectangle3_width(rectangle3_widths[517]), .rectangle3_height(rectangle3_heights[517]), .rectangle3_weight(rectangle3_weights[517]), .feature_threshold(feature_thresholds[517]), .feature_above(feature_aboves[517]), .feature_below(feature_belows[517]), .scan_win_std_dev(scan_win_std_dev[517]), .feature_accum(feature_accums[517]));
  accum_calculator ac518(.scan_win(scan_win518), .rectangle1_x(rectangle1_xs[518]), .rectangle1_y(rectangle1_ys[518]), .rectangle1_width(rectangle1_widths[518]), .rectangle1_height(rectangle1_heights[518]), .rectangle1_weight(rectangle1_weights[518]), .rectangle2_x(rectangle2_xs[518]), .rectangle2_y(rectangle2_ys[518]), .rectangle2_width(rectangle2_widths[518]), .rectangle2_height(rectangle2_heights[518]), .rectangle2_weight(rectangle2_weights[518]), .rectangle3_x(rectangle3_xs[518]), .rectangle3_y(rectangle3_ys[518]), .rectangle3_width(rectangle3_widths[518]), .rectangle3_height(rectangle3_heights[518]), .rectangle3_weight(rectangle3_weights[518]), .feature_threshold(feature_thresholds[518]), .feature_above(feature_aboves[518]), .feature_below(feature_belows[518]), .scan_win_std_dev(scan_win_std_dev[518]), .feature_accum(feature_accums[518]));
  accum_calculator ac519(.scan_win(scan_win519), .rectangle1_x(rectangle1_xs[519]), .rectangle1_y(rectangle1_ys[519]), .rectangle1_width(rectangle1_widths[519]), .rectangle1_height(rectangle1_heights[519]), .rectangle1_weight(rectangle1_weights[519]), .rectangle2_x(rectangle2_xs[519]), .rectangle2_y(rectangle2_ys[519]), .rectangle2_width(rectangle2_widths[519]), .rectangle2_height(rectangle2_heights[519]), .rectangle2_weight(rectangle2_weights[519]), .rectangle3_x(rectangle3_xs[519]), .rectangle3_y(rectangle3_ys[519]), .rectangle3_width(rectangle3_widths[519]), .rectangle3_height(rectangle3_heights[519]), .rectangle3_weight(rectangle3_weights[519]), .feature_threshold(feature_thresholds[519]), .feature_above(feature_aboves[519]), .feature_below(feature_belows[519]), .scan_win_std_dev(scan_win_std_dev[519]), .feature_accum(feature_accums[519]));
  accum_calculator ac520(.scan_win(scan_win520), .rectangle1_x(rectangle1_xs[520]), .rectangle1_y(rectangle1_ys[520]), .rectangle1_width(rectangle1_widths[520]), .rectangle1_height(rectangle1_heights[520]), .rectangle1_weight(rectangle1_weights[520]), .rectangle2_x(rectangle2_xs[520]), .rectangle2_y(rectangle2_ys[520]), .rectangle2_width(rectangle2_widths[520]), .rectangle2_height(rectangle2_heights[520]), .rectangle2_weight(rectangle2_weights[520]), .rectangle3_x(rectangle3_xs[520]), .rectangle3_y(rectangle3_ys[520]), .rectangle3_width(rectangle3_widths[520]), .rectangle3_height(rectangle3_heights[520]), .rectangle3_weight(rectangle3_weights[520]), .feature_threshold(feature_thresholds[520]), .feature_above(feature_aboves[520]), .feature_below(feature_belows[520]), .scan_win_std_dev(scan_win_std_dev[520]), .feature_accum(feature_accums[520]));
  accum_calculator ac521(.scan_win(scan_win521), .rectangle1_x(rectangle1_xs[521]), .rectangle1_y(rectangle1_ys[521]), .rectangle1_width(rectangle1_widths[521]), .rectangle1_height(rectangle1_heights[521]), .rectangle1_weight(rectangle1_weights[521]), .rectangle2_x(rectangle2_xs[521]), .rectangle2_y(rectangle2_ys[521]), .rectangle2_width(rectangle2_widths[521]), .rectangle2_height(rectangle2_heights[521]), .rectangle2_weight(rectangle2_weights[521]), .rectangle3_x(rectangle3_xs[521]), .rectangle3_y(rectangle3_ys[521]), .rectangle3_width(rectangle3_widths[521]), .rectangle3_height(rectangle3_heights[521]), .rectangle3_weight(rectangle3_weights[521]), .feature_threshold(feature_thresholds[521]), .feature_above(feature_aboves[521]), .feature_below(feature_belows[521]), .scan_win_std_dev(scan_win_std_dev[521]), .feature_accum(feature_accums[521]));
  accum_calculator ac522(.scan_win(scan_win522), .rectangle1_x(rectangle1_xs[522]), .rectangle1_y(rectangle1_ys[522]), .rectangle1_width(rectangle1_widths[522]), .rectangle1_height(rectangle1_heights[522]), .rectangle1_weight(rectangle1_weights[522]), .rectangle2_x(rectangle2_xs[522]), .rectangle2_y(rectangle2_ys[522]), .rectangle2_width(rectangle2_widths[522]), .rectangle2_height(rectangle2_heights[522]), .rectangle2_weight(rectangle2_weights[522]), .rectangle3_x(rectangle3_xs[522]), .rectangle3_y(rectangle3_ys[522]), .rectangle3_width(rectangle3_widths[522]), .rectangle3_height(rectangle3_heights[522]), .rectangle3_weight(rectangle3_weights[522]), .feature_threshold(feature_thresholds[522]), .feature_above(feature_aboves[522]), .feature_below(feature_belows[522]), .scan_win_std_dev(scan_win_std_dev[522]), .feature_accum(feature_accums[522]));
  accum_calculator ac523(.scan_win(scan_win523), .rectangle1_x(rectangle1_xs[523]), .rectangle1_y(rectangle1_ys[523]), .rectangle1_width(rectangle1_widths[523]), .rectangle1_height(rectangle1_heights[523]), .rectangle1_weight(rectangle1_weights[523]), .rectangle2_x(rectangle2_xs[523]), .rectangle2_y(rectangle2_ys[523]), .rectangle2_width(rectangle2_widths[523]), .rectangle2_height(rectangle2_heights[523]), .rectangle2_weight(rectangle2_weights[523]), .rectangle3_x(rectangle3_xs[523]), .rectangle3_y(rectangle3_ys[523]), .rectangle3_width(rectangle3_widths[523]), .rectangle3_height(rectangle3_heights[523]), .rectangle3_weight(rectangle3_weights[523]), .feature_threshold(feature_thresholds[523]), .feature_above(feature_aboves[523]), .feature_below(feature_belows[523]), .scan_win_std_dev(scan_win_std_dev[523]), .feature_accum(feature_accums[523]));
  accum_calculator ac524(.scan_win(scan_win524), .rectangle1_x(rectangle1_xs[524]), .rectangle1_y(rectangle1_ys[524]), .rectangle1_width(rectangle1_widths[524]), .rectangle1_height(rectangle1_heights[524]), .rectangle1_weight(rectangle1_weights[524]), .rectangle2_x(rectangle2_xs[524]), .rectangle2_y(rectangle2_ys[524]), .rectangle2_width(rectangle2_widths[524]), .rectangle2_height(rectangle2_heights[524]), .rectangle2_weight(rectangle2_weights[524]), .rectangle3_x(rectangle3_xs[524]), .rectangle3_y(rectangle3_ys[524]), .rectangle3_width(rectangle3_widths[524]), .rectangle3_height(rectangle3_heights[524]), .rectangle3_weight(rectangle3_weights[524]), .feature_threshold(feature_thresholds[524]), .feature_above(feature_aboves[524]), .feature_below(feature_belows[524]), .scan_win_std_dev(scan_win_std_dev[524]), .feature_accum(feature_accums[524]));
  accum_calculator ac525(.scan_win(scan_win525), .rectangle1_x(rectangle1_xs[525]), .rectangle1_y(rectangle1_ys[525]), .rectangle1_width(rectangle1_widths[525]), .rectangle1_height(rectangle1_heights[525]), .rectangle1_weight(rectangle1_weights[525]), .rectangle2_x(rectangle2_xs[525]), .rectangle2_y(rectangle2_ys[525]), .rectangle2_width(rectangle2_widths[525]), .rectangle2_height(rectangle2_heights[525]), .rectangle2_weight(rectangle2_weights[525]), .rectangle3_x(rectangle3_xs[525]), .rectangle3_y(rectangle3_ys[525]), .rectangle3_width(rectangle3_widths[525]), .rectangle3_height(rectangle3_heights[525]), .rectangle3_weight(rectangle3_weights[525]), .feature_threshold(feature_thresholds[525]), .feature_above(feature_aboves[525]), .feature_below(feature_belows[525]), .scan_win_std_dev(scan_win_std_dev[525]), .feature_accum(feature_accums[525]));
  accum_calculator ac526(.scan_win(scan_win526), .rectangle1_x(rectangle1_xs[526]), .rectangle1_y(rectangle1_ys[526]), .rectangle1_width(rectangle1_widths[526]), .rectangle1_height(rectangle1_heights[526]), .rectangle1_weight(rectangle1_weights[526]), .rectangle2_x(rectangle2_xs[526]), .rectangle2_y(rectangle2_ys[526]), .rectangle2_width(rectangle2_widths[526]), .rectangle2_height(rectangle2_heights[526]), .rectangle2_weight(rectangle2_weights[526]), .rectangle3_x(rectangle3_xs[526]), .rectangle3_y(rectangle3_ys[526]), .rectangle3_width(rectangle3_widths[526]), .rectangle3_height(rectangle3_heights[526]), .rectangle3_weight(rectangle3_weights[526]), .feature_threshold(feature_thresholds[526]), .feature_above(feature_aboves[526]), .feature_below(feature_belows[526]), .scan_win_std_dev(scan_win_std_dev[526]), .feature_accum(feature_accums[526]));
  accum_calculator ac527(.scan_win(scan_win527), .rectangle1_x(rectangle1_xs[527]), .rectangle1_y(rectangle1_ys[527]), .rectangle1_width(rectangle1_widths[527]), .rectangle1_height(rectangle1_heights[527]), .rectangle1_weight(rectangle1_weights[527]), .rectangle2_x(rectangle2_xs[527]), .rectangle2_y(rectangle2_ys[527]), .rectangle2_width(rectangle2_widths[527]), .rectangle2_height(rectangle2_heights[527]), .rectangle2_weight(rectangle2_weights[527]), .rectangle3_x(rectangle3_xs[527]), .rectangle3_y(rectangle3_ys[527]), .rectangle3_width(rectangle3_widths[527]), .rectangle3_height(rectangle3_heights[527]), .rectangle3_weight(rectangle3_weights[527]), .feature_threshold(feature_thresholds[527]), .feature_above(feature_aboves[527]), .feature_below(feature_belows[527]), .scan_win_std_dev(scan_win_std_dev[527]), .feature_accum(feature_accums[527]));
  accum_calculator ac528(.scan_win(scan_win528), .rectangle1_x(rectangle1_xs[528]), .rectangle1_y(rectangle1_ys[528]), .rectangle1_width(rectangle1_widths[528]), .rectangle1_height(rectangle1_heights[528]), .rectangle1_weight(rectangle1_weights[528]), .rectangle2_x(rectangle2_xs[528]), .rectangle2_y(rectangle2_ys[528]), .rectangle2_width(rectangle2_widths[528]), .rectangle2_height(rectangle2_heights[528]), .rectangle2_weight(rectangle2_weights[528]), .rectangle3_x(rectangle3_xs[528]), .rectangle3_y(rectangle3_ys[528]), .rectangle3_width(rectangle3_widths[528]), .rectangle3_height(rectangle3_heights[528]), .rectangle3_weight(rectangle3_weights[528]), .feature_threshold(feature_thresholds[528]), .feature_above(feature_aboves[528]), .feature_below(feature_belows[528]), .scan_win_std_dev(scan_win_std_dev[528]), .feature_accum(feature_accums[528]));
  accum_calculator ac529(.scan_win(scan_win529), .rectangle1_x(rectangle1_xs[529]), .rectangle1_y(rectangle1_ys[529]), .rectangle1_width(rectangle1_widths[529]), .rectangle1_height(rectangle1_heights[529]), .rectangle1_weight(rectangle1_weights[529]), .rectangle2_x(rectangle2_xs[529]), .rectangle2_y(rectangle2_ys[529]), .rectangle2_width(rectangle2_widths[529]), .rectangle2_height(rectangle2_heights[529]), .rectangle2_weight(rectangle2_weights[529]), .rectangle3_x(rectangle3_xs[529]), .rectangle3_y(rectangle3_ys[529]), .rectangle3_width(rectangle3_widths[529]), .rectangle3_height(rectangle3_heights[529]), .rectangle3_weight(rectangle3_weights[529]), .feature_threshold(feature_thresholds[529]), .feature_above(feature_aboves[529]), .feature_below(feature_belows[529]), .scan_win_std_dev(scan_win_std_dev[529]), .feature_accum(feature_accums[529]));
  accum_calculator ac530(.scan_win(scan_win530), .rectangle1_x(rectangle1_xs[530]), .rectangle1_y(rectangle1_ys[530]), .rectangle1_width(rectangle1_widths[530]), .rectangle1_height(rectangle1_heights[530]), .rectangle1_weight(rectangle1_weights[530]), .rectangle2_x(rectangle2_xs[530]), .rectangle2_y(rectangle2_ys[530]), .rectangle2_width(rectangle2_widths[530]), .rectangle2_height(rectangle2_heights[530]), .rectangle2_weight(rectangle2_weights[530]), .rectangle3_x(rectangle3_xs[530]), .rectangle3_y(rectangle3_ys[530]), .rectangle3_width(rectangle3_widths[530]), .rectangle3_height(rectangle3_heights[530]), .rectangle3_weight(rectangle3_weights[530]), .feature_threshold(feature_thresholds[530]), .feature_above(feature_aboves[530]), .feature_below(feature_belows[530]), .scan_win_std_dev(scan_win_std_dev[530]), .feature_accum(feature_accums[530]));
  accum_calculator ac531(.scan_win(scan_win531), .rectangle1_x(rectangle1_xs[531]), .rectangle1_y(rectangle1_ys[531]), .rectangle1_width(rectangle1_widths[531]), .rectangle1_height(rectangle1_heights[531]), .rectangle1_weight(rectangle1_weights[531]), .rectangle2_x(rectangle2_xs[531]), .rectangle2_y(rectangle2_ys[531]), .rectangle2_width(rectangle2_widths[531]), .rectangle2_height(rectangle2_heights[531]), .rectangle2_weight(rectangle2_weights[531]), .rectangle3_x(rectangle3_xs[531]), .rectangle3_y(rectangle3_ys[531]), .rectangle3_width(rectangle3_widths[531]), .rectangle3_height(rectangle3_heights[531]), .rectangle3_weight(rectangle3_weights[531]), .feature_threshold(feature_thresholds[531]), .feature_above(feature_aboves[531]), .feature_below(feature_belows[531]), .scan_win_std_dev(scan_win_std_dev[531]), .feature_accum(feature_accums[531]));
  accum_calculator ac532(.scan_win(scan_win532), .rectangle1_x(rectangle1_xs[532]), .rectangle1_y(rectangle1_ys[532]), .rectangle1_width(rectangle1_widths[532]), .rectangle1_height(rectangle1_heights[532]), .rectangle1_weight(rectangle1_weights[532]), .rectangle2_x(rectangle2_xs[532]), .rectangle2_y(rectangle2_ys[532]), .rectangle2_width(rectangle2_widths[532]), .rectangle2_height(rectangle2_heights[532]), .rectangle2_weight(rectangle2_weights[532]), .rectangle3_x(rectangle3_xs[532]), .rectangle3_y(rectangle3_ys[532]), .rectangle3_width(rectangle3_widths[532]), .rectangle3_height(rectangle3_heights[532]), .rectangle3_weight(rectangle3_weights[532]), .feature_threshold(feature_thresholds[532]), .feature_above(feature_aboves[532]), .feature_below(feature_belows[532]), .scan_win_std_dev(scan_win_std_dev[532]), .feature_accum(feature_accums[532]));
  accum_calculator ac533(.scan_win(scan_win533), .rectangle1_x(rectangle1_xs[533]), .rectangle1_y(rectangle1_ys[533]), .rectangle1_width(rectangle1_widths[533]), .rectangle1_height(rectangle1_heights[533]), .rectangle1_weight(rectangle1_weights[533]), .rectangle2_x(rectangle2_xs[533]), .rectangle2_y(rectangle2_ys[533]), .rectangle2_width(rectangle2_widths[533]), .rectangle2_height(rectangle2_heights[533]), .rectangle2_weight(rectangle2_weights[533]), .rectangle3_x(rectangle3_xs[533]), .rectangle3_y(rectangle3_ys[533]), .rectangle3_width(rectangle3_widths[533]), .rectangle3_height(rectangle3_heights[533]), .rectangle3_weight(rectangle3_weights[533]), .feature_threshold(feature_thresholds[533]), .feature_above(feature_aboves[533]), .feature_below(feature_belows[533]), .scan_win_std_dev(scan_win_std_dev[533]), .feature_accum(feature_accums[533]));
  accum_calculator ac534(.scan_win(scan_win534), .rectangle1_x(rectangle1_xs[534]), .rectangle1_y(rectangle1_ys[534]), .rectangle1_width(rectangle1_widths[534]), .rectangle1_height(rectangle1_heights[534]), .rectangle1_weight(rectangle1_weights[534]), .rectangle2_x(rectangle2_xs[534]), .rectangle2_y(rectangle2_ys[534]), .rectangle2_width(rectangle2_widths[534]), .rectangle2_height(rectangle2_heights[534]), .rectangle2_weight(rectangle2_weights[534]), .rectangle3_x(rectangle3_xs[534]), .rectangle3_y(rectangle3_ys[534]), .rectangle3_width(rectangle3_widths[534]), .rectangle3_height(rectangle3_heights[534]), .rectangle3_weight(rectangle3_weights[534]), .feature_threshold(feature_thresholds[534]), .feature_above(feature_aboves[534]), .feature_below(feature_belows[534]), .scan_win_std_dev(scan_win_std_dev[534]), .feature_accum(feature_accums[534]));
  accum_calculator ac535(.scan_win(scan_win535), .rectangle1_x(rectangle1_xs[535]), .rectangle1_y(rectangle1_ys[535]), .rectangle1_width(rectangle1_widths[535]), .rectangle1_height(rectangle1_heights[535]), .rectangle1_weight(rectangle1_weights[535]), .rectangle2_x(rectangle2_xs[535]), .rectangle2_y(rectangle2_ys[535]), .rectangle2_width(rectangle2_widths[535]), .rectangle2_height(rectangle2_heights[535]), .rectangle2_weight(rectangle2_weights[535]), .rectangle3_x(rectangle3_xs[535]), .rectangle3_y(rectangle3_ys[535]), .rectangle3_width(rectangle3_widths[535]), .rectangle3_height(rectangle3_heights[535]), .rectangle3_weight(rectangle3_weights[535]), .feature_threshold(feature_thresholds[535]), .feature_above(feature_aboves[535]), .feature_below(feature_belows[535]), .scan_win_std_dev(scan_win_std_dev[535]), .feature_accum(feature_accums[535]));
  accum_calculator ac536(.scan_win(scan_win536), .rectangle1_x(rectangle1_xs[536]), .rectangle1_y(rectangle1_ys[536]), .rectangle1_width(rectangle1_widths[536]), .rectangle1_height(rectangle1_heights[536]), .rectangle1_weight(rectangle1_weights[536]), .rectangle2_x(rectangle2_xs[536]), .rectangle2_y(rectangle2_ys[536]), .rectangle2_width(rectangle2_widths[536]), .rectangle2_height(rectangle2_heights[536]), .rectangle2_weight(rectangle2_weights[536]), .rectangle3_x(rectangle3_xs[536]), .rectangle3_y(rectangle3_ys[536]), .rectangle3_width(rectangle3_widths[536]), .rectangle3_height(rectangle3_heights[536]), .rectangle3_weight(rectangle3_weights[536]), .feature_threshold(feature_thresholds[536]), .feature_above(feature_aboves[536]), .feature_below(feature_belows[536]), .scan_win_std_dev(scan_win_std_dev[536]), .feature_accum(feature_accums[536]));
  accum_calculator ac537(.scan_win(scan_win537), .rectangle1_x(rectangle1_xs[537]), .rectangle1_y(rectangle1_ys[537]), .rectangle1_width(rectangle1_widths[537]), .rectangle1_height(rectangle1_heights[537]), .rectangle1_weight(rectangle1_weights[537]), .rectangle2_x(rectangle2_xs[537]), .rectangle2_y(rectangle2_ys[537]), .rectangle2_width(rectangle2_widths[537]), .rectangle2_height(rectangle2_heights[537]), .rectangle2_weight(rectangle2_weights[537]), .rectangle3_x(rectangle3_xs[537]), .rectangle3_y(rectangle3_ys[537]), .rectangle3_width(rectangle3_widths[537]), .rectangle3_height(rectangle3_heights[537]), .rectangle3_weight(rectangle3_weights[537]), .feature_threshold(feature_thresholds[537]), .feature_above(feature_aboves[537]), .feature_below(feature_belows[537]), .scan_win_std_dev(scan_win_std_dev[537]), .feature_accum(feature_accums[537]));
  accum_calculator ac538(.scan_win(scan_win538), .rectangle1_x(rectangle1_xs[538]), .rectangle1_y(rectangle1_ys[538]), .rectangle1_width(rectangle1_widths[538]), .rectangle1_height(rectangle1_heights[538]), .rectangle1_weight(rectangle1_weights[538]), .rectangle2_x(rectangle2_xs[538]), .rectangle2_y(rectangle2_ys[538]), .rectangle2_width(rectangle2_widths[538]), .rectangle2_height(rectangle2_heights[538]), .rectangle2_weight(rectangle2_weights[538]), .rectangle3_x(rectangle3_xs[538]), .rectangle3_y(rectangle3_ys[538]), .rectangle3_width(rectangle3_widths[538]), .rectangle3_height(rectangle3_heights[538]), .rectangle3_weight(rectangle3_weights[538]), .feature_threshold(feature_thresholds[538]), .feature_above(feature_aboves[538]), .feature_below(feature_belows[538]), .scan_win_std_dev(scan_win_std_dev[538]), .feature_accum(feature_accums[538]));
  accum_calculator ac539(.scan_win(scan_win539), .rectangle1_x(rectangle1_xs[539]), .rectangle1_y(rectangle1_ys[539]), .rectangle1_width(rectangle1_widths[539]), .rectangle1_height(rectangle1_heights[539]), .rectangle1_weight(rectangle1_weights[539]), .rectangle2_x(rectangle2_xs[539]), .rectangle2_y(rectangle2_ys[539]), .rectangle2_width(rectangle2_widths[539]), .rectangle2_height(rectangle2_heights[539]), .rectangle2_weight(rectangle2_weights[539]), .rectangle3_x(rectangle3_xs[539]), .rectangle3_y(rectangle3_ys[539]), .rectangle3_width(rectangle3_widths[539]), .rectangle3_height(rectangle3_heights[539]), .rectangle3_weight(rectangle3_weights[539]), .feature_threshold(feature_thresholds[539]), .feature_above(feature_aboves[539]), .feature_below(feature_belows[539]), .scan_win_std_dev(scan_win_std_dev[539]), .feature_accum(feature_accums[539]));
  accum_calculator ac540(.scan_win(scan_win540), .rectangle1_x(rectangle1_xs[540]), .rectangle1_y(rectangle1_ys[540]), .rectangle1_width(rectangle1_widths[540]), .rectangle1_height(rectangle1_heights[540]), .rectangle1_weight(rectangle1_weights[540]), .rectangle2_x(rectangle2_xs[540]), .rectangle2_y(rectangle2_ys[540]), .rectangle2_width(rectangle2_widths[540]), .rectangle2_height(rectangle2_heights[540]), .rectangle2_weight(rectangle2_weights[540]), .rectangle3_x(rectangle3_xs[540]), .rectangle3_y(rectangle3_ys[540]), .rectangle3_width(rectangle3_widths[540]), .rectangle3_height(rectangle3_heights[540]), .rectangle3_weight(rectangle3_weights[540]), .feature_threshold(feature_thresholds[540]), .feature_above(feature_aboves[540]), .feature_below(feature_belows[540]), .scan_win_std_dev(scan_win_std_dev[540]), .feature_accum(feature_accums[540]));
  accum_calculator ac541(.scan_win(scan_win541), .rectangle1_x(rectangle1_xs[541]), .rectangle1_y(rectangle1_ys[541]), .rectangle1_width(rectangle1_widths[541]), .rectangle1_height(rectangle1_heights[541]), .rectangle1_weight(rectangle1_weights[541]), .rectangle2_x(rectangle2_xs[541]), .rectangle2_y(rectangle2_ys[541]), .rectangle2_width(rectangle2_widths[541]), .rectangle2_height(rectangle2_heights[541]), .rectangle2_weight(rectangle2_weights[541]), .rectangle3_x(rectangle3_xs[541]), .rectangle3_y(rectangle3_ys[541]), .rectangle3_width(rectangle3_widths[541]), .rectangle3_height(rectangle3_heights[541]), .rectangle3_weight(rectangle3_weights[541]), .feature_threshold(feature_thresholds[541]), .feature_above(feature_aboves[541]), .feature_below(feature_belows[541]), .scan_win_std_dev(scan_win_std_dev[541]), .feature_accum(feature_accums[541]));
  accum_calculator ac542(.scan_win(scan_win542), .rectangle1_x(rectangle1_xs[542]), .rectangle1_y(rectangle1_ys[542]), .rectangle1_width(rectangle1_widths[542]), .rectangle1_height(rectangle1_heights[542]), .rectangle1_weight(rectangle1_weights[542]), .rectangle2_x(rectangle2_xs[542]), .rectangle2_y(rectangle2_ys[542]), .rectangle2_width(rectangle2_widths[542]), .rectangle2_height(rectangle2_heights[542]), .rectangle2_weight(rectangle2_weights[542]), .rectangle3_x(rectangle3_xs[542]), .rectangle3_y(rectangle3_ys[542]), .rectangle3_width(rectangle3_widths[542]), .rectangle3_height(rectangle3_heights[542]), .rectangle3_weight(rectangle3_weights[542]), .feature_threshold(feature_thresholds[542]), .feature_above(feature_aboves[542]), .feature_below(feature_belows[542]), .scan_win_std_dev(scan_win_std_dev[542]), .feature_accum(feature_accums[542]));
  accum_calculator ac543(.scan_win(scan_win543), .rectangle1_x(rectangle1_xs[543]), .rectangle1_y(rectangle1_ys[543]), .rectangle1_width(rectangle1_widths[543]), .rectangle1_height(rectangle1_heights[543]), .rectangle1_weight(rectangle1_weights[543]), .rectangle2_x(rectangle2_xs[543]), .rectangle2_y(rectangle2_ys[543]), .rectangle2_width(rectangle2_widths[543]), .rectangle2_height(rectangle2_heights[543]), .rectangle2_weight(rectangle2_weights[543]), .rectangle3_x(rectangle3_xs[543]), .rectangle3_y(rectangle3_ys[543]), .rectangle3_width(rectangle3_widths[543]), .rectangle3_height(rectangle3_heights[543]), .rectangle3_weight(rectangle3_weights[543]), .feature_threshold(feature_thresholds[543]), .feature_above(feature_aboves[543]), .feature_below(feature_belows[543]), .scan_win_std_dev(scan_win_std_dev[543]), .feature_accum(feature_accums[543]));
  accum_calculator ac544(.scan_win(scan_win544), .rectangle1_x(rectangle1_xs[544]), .rectangle1_y(rectangle1_ys[544]), .rectangle1_width(rectangle1_widths[544]), .rectangle1_height(rectangle1_heights[544]), .rectangle1_weight(rectangle1_weights[544]), .rectangle2_x(rectangle2_xs[544]), .rectangle2_y(rectangle2_ys[544]), .rectangle2_width(rectangle2_widths[544]), .rectangle2_height(rectangle2_heights[544]), .rectangle2_weight(rectangle2_weights[544]), .rectangle3_x(rectangle3_xs[544]), .rectangle3_y(rectangle3_ys[544]), .rectangle3_width(rectangle3_widths[544]), .rectangle3_height(rectangle3_heights[544]), .rectangle3_weight(rectangle3_weights[544]), .feature_threshold(feature_thresholds[544]), .feature_above(feature_aboves[544]), .feature_below(feature_belows[544]), .scan_win_std_dev(scan_win_std_dev[544]), .feature_accum(feature_accums[544]));
  accum_calculator ac545(.scan_win(scan_win545), .rectangle1_x(rectangle1_xs[545]), .rectangle1_y(rectangle1_ys[545]), .rectangle1_width(rectangle1_widths[545]), .rectangle1_height(rectangle1_heights[545]), .rectangle1_weight(rectangle1_weights[545]), .rectangle2_x(rectangle2_xs[545]), .rectangle2_y(rectangle2_ys[545]), .rectangle2_width(rectangle2_widths[545]), .rectangle2_height(rectangle2_heights[545]), .rectangle2_weight(rectangle2_weights[545]), .rectangle3_x(rectangle3_xs[545]), .rectangle3_y(rectangle3_ys[545]), .rectangle3_width(rectangle3_widths[545]), .rectangle3_height(rectangle3_heights[545]), .rectangle3_weight(rectangle3_weights[545]), .feature_threshold(feature_thresholds[545]), .feature_above(feature_aboves[545]), .feature_below(feature_belows[545]), .scan_win_std_dev(scan_win_std_dev[545]), .feature_accum(feature_accums[545]));
  accum_calculator ac546(.scan_win(scan_win546), .rectangle1_x(rectangle1_xs[546]), .rectangle1_y(rectangle1_ys[546]), .rectangle1_width(rectangle1_widths[546]), .rectangle1_height(rectangle1_heights[546]), .rectangle1_weight(rectangle1_weights[546]), .rectangle2_x(rectangle2_xs[546]), .rectangle2_y(rectangle2_ys[546]), .rectangle2_width(rectangle2_widths[546]), .rectangle2_height(rectangle2_heights[546]), .rectangle2_weight(rectangle2_weights[546]), .rectangle3_x(rectangle3_xs[546]), .rectangle3_y(rectangle3_ys[546]), .rectangle3_width(rectangle3_widths[546]), .rectangle3_height(rectangle3_heights[546]), .rectangle3_weight(rectangle3_weights[546]), .feature_threshold(feature_thresholds[546]), .feature_above(feature_aboves[546]), .feature_below(feature_belows[546]), .scan_win_std_dev(scan_win_std_dev[546]), .feature_accum(feature_accums[546]));
  accum_calculator ac547(.scan_win(scan_win547), .rectangle1_x(rectangle1_xs[547]), .rectangle1_y(rectangle1_ys[547]), .rectangle1_width(rectangle1_widths[547]), .rectangle1_height(rectangle1_heights[547]), .rectangle1_weight(rectangle1_weights[547]), .rectangle2_x(rectangle2_xs[547]), .rectangle2_y(rectangle2_ys[547]), .rectangle2_width(rectangle2_widths[547]), .rectangle2_height(rectangle2_heights[547]), .rectangle2_weight(rectangle2_weights[547]), .rectangle3_x(rectangle3_xs[547]), .rectangle3_y(rectangle3_ys[547]), .rectangle3_width(rectangle3_widths[547]), .rectangle3_height(rectangle3_heights[547]), .rectangle3_weight(rectangle3_weights[547]), .feature_threshold(feature_thresholds[547]), .feature_above(feature_aboves[547]), .feature_below(feature_belows[547]), .scan_win_std_dev(scan_win_std_dev[547]), .feature_accum(feature_accums[547]));
  accum_calculator ac548(.scan_win(scan_win548), .rectangle1_x(rectangle1_xs[548]), .rectangle1_y(rectangle1_ys[548]), .rectangle1_width(rectangle1_widths[548]), .rectangle1_height(rectangle1_heights[548]), .rectangle1_weight(rectangle1_weights[548]), .rectangle2_x(rectangle2_xs[548]), .rectangle2_y(rectangle2_ys[548]), .rectangle2_width(rectangle2_widths[548]), .rectangle2_height(rectangle2_heights[548]), .rectangle2_weight(rectangle2_weights[548]), .rectangle3_x(rectangle3_xs[548]), .rectangle3_y(rectangle3_ys[548]), .rectangle3_width(rectangle3_widths[548]), .rectangle3_height(rectangle3_heights[548]), .rectangle3_weight(rectangle3_weights[548]), .feature_threshold(feature_thresholds[548]), .feature_above(feature_aboves[548]), .feature_below(feature_belows[548]), .scan_win_std_dev(scan_win_std_dev[548]), .feature_accum(feature_accums[548]));
  accum_calculator ac549(.scan_win(scan_win549), .rectangle1_x(rectangle1_xs[549]), .rectangle1_y(rectangle1_ys[549]), .rectangle1_width(rectangle1_widths[549]), .rectangle1_height(rectangle1_heights[549]), .rectangle1_weight(rectangle1_weights[549]), .rectangle2_x(rectangle2_xs[549]), .rectangle2_y(rectangle2_ys[549]), .rectangle2_width(rectangle2_widths[549]), .rectangle2_height(rectangle2_heights[549]), .rectangle2_weight(rectangle2_weights[549]), .rectangle3_x(rectangle3_xs[549]), .rectangle3_y(rectangle3_ys[549]), .rectangle3_width(rectangle3_widths[549]), .rectangle3_height(rectangle3_heights[549]), .rectangle3_weight(rectangle3_weights[549]), .feature_threshold(feature_thresholds[549]), .feature_above(feature_aboves[549]), .feature_below(feature_belows[549]), .scan_win_std_dev(scan_win_std_dev[549]), .feature_accum(feature_accums[549]));
  accum_calculator ac550(.scan_win(scan_win550), .rectangle1_x(rectangle1_xs[550]), .rectangle1_y(rectangle1_ys[550]), .rectangle1_width(rectangle1_widths[550]), .rectangle1_height(rectangle1_heights[550]), .rectangle1_weight(rectangle1_weights[550]), .rectangle2_x(rectangle2_xs[550]), .rectangle2_y(rectangle2_ys[550]), .rectangle2_width(rectangle2_widths[550]), .rectangle2_height(rectangle2_heights[550]), .rectangle2_weight(rectangle2_weights[550]), .rectangle3_x(rectangle3_xs[550]), .rectangle3_y(rectangle3_ys[550]), .rectangle3_width(rectangle3_widths[550]), .rectangle3_height(rectangle3_heights[550]), .rectangle3_weight(rectangle3_weights[550]), .feature_threshold(feature_thresholds[550]), .feature_above(feature_aboves[550]), .feature_below(feature_belows[550]), .scan_win_std_dev(scan_win_std_dev[550]), .feature_accum(feature_accums[550]));
  accum_calculator ac551(.scan_win(scan_win551), .rectangle1_x(rectangle1_xs[551]), .rectangle1_y(rectangle1_ys[551]), .rectangle1_width(rectangle1_widths[551]), .rectangle1_height(rectangle1_heights[551]), .rectangle1_weight(rectangle1_weights[551]), .rectangle2_x(rectangle2_xs[551]), .rectangle2_y(rectangle2_ys[551]), .rectangle2_width(rectangle2_widths[551]), .rectangle2_height(rectangle2_heights[551]), .rectangle2_weight(rectangle2_weights[551]), .rectangle3_x(rectangle3_xs[551]), .rectangle3_y(rectangle3_ys[551]), .rectangle3_width(rectangle3_widths[551]), .rectangle3_height(rectangle3_heights[551]), .rectangle3_weight(rectangle3_weights[551]), .feature_threshold(feature_thresholds[551]), .feature_above(feature_aboves[551]), .feature_below(feature_belows[551]), .scan_win_std_dev(scan_win_std_dev[551]), .feature_accum(feature_accums[551]));
  accum_calculator ac552(.scan_win(scan_win552), .rectangle1_x(rectangle1_xs[552]), .rectangle1_y(rectangle1_ys[552]), .rectangle1_width(rectangle1_widths[552]), .rectangle1_height(rectangle1_heights[552]), .rectangle1_weight(rectangle1_weights[552]), .rectangle2_x(rectangle2_xs[552]), .rectangle2_y(rectangle2_ys[552]), .rectangle2_width(rectangle2_widths[552]), .rectangle2_height(rectangle2_heights[552]), .rectangle2_weight(rectangle2_weights[552]), .rectangle3_x(rectangle3_xs[552]), .rectangle3_y(rectangle3_ys[552]), .rectangle3_width(rectangle3_widths[552]), .rectangle3_height(rectangle3_heights[552]), .rectangle3_weight(rectangle3_weights[552]), .feature_threshold(feature_thresholds[552]), .feature_above(feature_aboves[552]), .feature_below(feature_belows[552]), .scan_win_std_dev(scan_win_std_dev[552]), .feature_accum(feature_accums[552]));
  accum_calculator ac553(.scan_win(scan_win553), .rectangle1_x(rectangle1_xs[553]), .rectangle1_y(rectangle1_ys[553]), .rectangle1_width(rectangle1_widths[553]), .rectangle1_height(rectangle1_heights[553]), .rectangle1_weight(rectangle1_weights[553]), .rectangle2_x(rectangle2_xs[553]), .rectangle2_y(rectangle2_ys[553]), .rectangle2_width(rectangle2_widths[553]), .rectangle2_height(rectangle2_heights[553]), .rectangle2_weight(rectangle2_weights[553]), .rectangle3_x(rectangle3_xs[553]), .rectangle3_y(rectangle3_ys[553]), .rectangle3_width(rectangle3_widths[553]), .rectangle3_height(rectangle3_heights[553]), .rectangle3_weight(rectangle3_weights[553]), .feature_threshold(feature_thresholds[553]), .feature_above(feature_aboves[553]), .feature_below(feature_belows[553]), .scan_win_std_dev(scan_win_std_dev[553]), .feature_accum(feature_accums[553]));
  accum_calculator ac554(.scan_win(scan_win554), .rectangle1_x(rectangle1_xs[554]), .rectangle1_y(rectangle1_ys[554]), .rectangle1_width(rectangle1_widths[554]), .rectangle1_height(rectangle1_heights[554]), .rectangle1_weight(rectangle1_weights[554]), .rectangle2_x(rectangle2_xs[554]), .rectangle2_y(rectangle2_ys[554]), .rectangle2_width(rectangle2_widths[554]), .rectangle2_height(rectangle2_heights[554]), .rectangle2_weight(rectangle2_weights[554]), .rectangle3_x(rectangle3_xs[554]), .rectangle3_y(rectangle3_ys[554]), .rectangle3_width(rectangle3_widths[554]), .rectangle3_height(rectangle3_heights[554]), .rectangle3_weight(rectangle3_weights[554]), .feature_threshold(feature_thresholds[554]), .feature_above(feature_aboves[554]), .feature_below(feature_belows[554]), .scan_win_std_dev(scan_win_std_dev[554]), .feature_accum(feature_accums[554]));
  accum_calculator ac555(.scan_win(scan_win555), .rectangle1_x(rectangle1_xs[555]), .rectangle1_y(rectangle1_ys[555]), .rectangle1_width(rectangle1_widths[555]), .rectangle1_height(rectangle1_heights[555]), .rectangle1_weight(rectangle1_weights[555]), .rectangle2_x(rectangle2_xs[555]), .rectangle2_y(rectangle2_ys[555]), .rectangle2_width(rectangle2_widths[555]), .rectangle2_height(rectangle2_heights[555]), .rectangle2_weight(rectangle2_weights[555]), .rectangle3_x(rectangle3_xs[555]), .rectangle3_y(rectangle3_ys[555]), .rectangle3_width(rectangle3_widths[555]), .rectangle3_height(rectangle3_heights[555]), .rectangle3_weight(rectangle3_weights[555]), .feature_threshold(feature_thresholds[555]), .feature_above(feature_aboves[555]), .feature_below(feature_belows[555]), .scan_win_std_dev(scan_win_std_dev[555]), .feature_accum(feature_accums[555]));
  accum_calculator ac556(.scan_win(scan_win556), .rectangle1_x(rectangle1_xs[556]), .rectangle1_y(rectangle1_ys[556]), .rectangle1_width(rectangle1_widths[556]), .rectangle1_height(rectangle1_heights[556]), .rectangle1_weight(rectangle1_weights[556]), .rectangle2_x(rectangle2_xs[556]), .rectangle2_y(rectangle2_ys[556]), .rectangle2_width(rectangle2_widths[556]), .rectangle2_height(rectangle2_heights[556]), .rectangle2_weight(rectangle2_weights[556]), .rectangle3_x(rectangle3_xs[556]), .rectangle3_y(rectangle3_ys[556]), .rectangle3_width(rectangle3_widths[556]), .rectangle3_height(rectangle3_heights[556]), .rectangle3_weight(rectangle3_weights[556]), .feature_threshold(feature_thresholds[556]), .feature_above(feature_aboves[556]), .feature_below(feature_belows[556]), .scan_win_std_dev(scan_win_std_dev[556]), .feature_accum(feature_accums[556]));
  accum_calculator ac557(.scan_win(scan_win557), .rectangle1_x(rectangle1_xs[557]), .rectangle1_y(rectangle1_ys[557]), .rectangle1_width(rectangle1_widths[557]), .rectangle1_height(rectangle1_heights[557]), .rectangle1_weight(rectangle1_weights[557]), .rectangle2_x(rectangle2_xs[557]), .rectangle2_y(rectangle2_ys[557]), .rectangle2_width(rectangle2_widths[557]), .rectangle2_height(rectangle2_heights[557]), .rectangle2_weight(rectangle2_weights[557]), .rectangle3_x(rectangle3_xs[557]), .rectangle3_y(rectangle3_ys[557]), .rectangle3_width(rectangle3_widths[557]), .rectangle3_height(rectangle3_heights[557]), .rectangle3_weight(rectangle3_weights[557]), .feature_threshold(feature_thresholds[557]), .feature_above(feature_aboves[557]), .feature_below(feature_belows[557]), .scan_win_std_dev(scan_win_std_dev[557]), .feature_accum(feature_accums[557]));
  accum_calculator ac558(.scan_win(scan_win558), .rectangle1_x(rectangle1_xs[558]), .rectangle1_y(rectangle1_ys[558]), .rectangle1_width(rectangle1_widths[558]), .rectangle1_height(rectangle1_heights[558]), .rectangle1_weight(rectangle1_weights[558]), .rectangle2_x(rectangle2_xs[558]), .rectangle2_y(rectangle2_ys[558]), .rectangle2_width(rectangle2_widths[558]), .rectangle2_height(rectangle2_heights[558]), .rectangle2_weight(rectangle2_weights[558]), .rectangle3_x(rectangle3_xs[558]), .rectangle3_y(rectangle3_ys[558]), .rectangle3_width(rectangle3_widths[558]), .rectangle3_height(rectangle3_heights[558]), .rectangle3_weight(rectangle3_weights[558]), .feature_threshold(feature_thresholds[558]), .feature_above(feature_aboves[558]), .feature_below(feature_belows[558]), .scan_win_std_dev(scan_win_std_dev[558]), .feature_accum(feature_accums[558]));
  accum_calculator ac559(.scan_win(scan_win559), .rectangle1_x(rectangle1_xs[559]), .rectangle1_y(rectangle1_ys[559]), .rectangle1_width(rectangle1_widths[559]), .rectangle1_height(rectangle1_heights[559]), .rectangle1_weight(rectangle1_weights[559]), .rectangle2_x(rectangle2_xs[559]), .rectangle2_y(rectangle2_ys[559]), .rectangle2_width(rectangle2_widths[559]), .rectangle2_height(rectangle2_heights[559]), .rectangle2_weight(rectangle2_weights[559]), .rectangle3_x(rectangle3_xs[559]), .rectangle3_y(rectangle3_ys[559]), .rectangle3_width(rectangle3_widths[559]), .rectangle3_height(rectangle3_heights[559]), .rectangle3_weight(rectangle3_weights[559]), .feature_threshold(feature_thresholds[559]), .feature_above(feature_aboves[559]), .feature_below(feature_belows[559]), .scan_win_std_dev(scan_win_std_dev[559]), .feature_accum(feature_accums[559]));
  accum_calculator ac560(.scan_win(scan_win560), .rectangle1_x(rectangle1_xs[560]), .rectangle1_y(rectangle1_ys[560]), .rectangle1_width(rectangle1_widths[560]), .rectangle1_height(rectangle1_heights[560]), .rectangle1_weight(rectangle1_weights[560]), .rectangle2_x(rectangle2_xs[560]), .rectangle2_y(rectangle2_ys[560]), .rectangle2_width(rectangle2_widths[560]), .rectangle2_height(rectangle2_heights[560]), .rectangle2_weight(rectangle2_weights[560]), .rectangle3_x(rectangle3_xs[560]), .rectangle3_y(rectangle3_ys[560]), .rectangle3_width(rectangle3_widths[560]), .rectangle3_height(rectangle3_heights[560]), .rectangle3_weight(rectangle3_weights[560]), .feature_threshold(feature_thresholds[560]), .feature_above(feature_aboves[560]), .feature_below(feature_belows[560]), .scan_win_std_dev(scan_win_std_dev[560]), .feature_accum(feature_accums[560]));
  accum_calculator ac561(.scan_win(scan_win561), .rectangle1_x(rectangle1_xs[561]), .rectangle1_y(rectangle1_ys[561]), .rectangle1_width(rectangle1_widths[561]), .rectangle1_height(rectangle1_heights[561]), .rectangle1_weight(rectangle1_weights[561]), .rectangle2_x(rectangle2_xs[561]), .rectangle2_y(rectangle2_ys[561]), .rectangle2_width(rectangle2_widths[561]), .rectangle2_height(rectangle2_heights[561]), .rectangle2_weight(rectangle2_weights[561]), .rectangle3_x(rectangle3_xs[561]), .rectangle3_y(rectangle3_ys[561]), .rectangle3_width(rectangle3_widths[561]), .rectangle3_height(rectangle3_heights[561]), .rectangle3_weight(rectangle3_weights[561]), .feature_threshold(feature_thresholds[561]), .feature_above(feature_aboves[561]), .feature_below(feature_belows[561]), .scan_win_std_dev(scan_win_std_dev[561]), .feature_accum(feature_accums[561]));
  accum_calculator ac562(.scan_win(scan_win562), .rectangle1_x(rectangle1_xs[562]), .rectangle1_y(rectangle1_ys[562]), .rectangle1_width(rectangle1_widths[562]), .rectangle1_height(rectangle1_heights[562]), .rectangle1_weight(rectangle1_weights[562]), .rectangle2_x(rectangle2_xs[562]), .rectangle2_y(rectangle2_ys[562]), .rectangle2_width(rectangle2_widths[562]), .rectangle2_height(rectangle2_heights[562]), .rectangle2_weight(rectangle2_weights[562]), .rectangle3_x(rectangle3_xs[562]), .rectangle3_y(rectangle3_ys[562]), .rectangle3_width(rectangle3_widths[562]), .rectangle3_height(rectangle3_heights[562]), .rectangle3_weight(rectangle3_weights[562]), .feature_threshold(feature_thresholds[562]), .feature_above(feature_aboves[562]), .feature_below(feature_belows[562]), .scan_win_std_dev(scan_win_std_dev[562]), .feature_accum(feature_accums[562]));
  accum_calculator ac563(.scan_win(scan_win563), .rectangle1_x(rectangle1_xs[563]), .rectangle1_y(rectangle1_ys[563]), .rectangle1_width(rectangle1_widths[563]), .rectangle1_height(rectangle1_heights[563]), .rectangle1_weight(rectangle1_weights[563]), .rectangle2_x(rectangle2_xs[563]), .rectangle2_y(rectangle2_ys[563]), .rectangle2_width(rectangle2_widths[563]), .rectangle2_height(rectangle2_heights[563]), .rectangle2_weight(rectangle2_weights[563]), .rectangle3_x(rectangle3_xs[563]), .rectangle3_y(rectangle3_ys[563]), .rectangle3_width(rectangle3_widths[563]), .rectangle3_height(rectangle3_heights[563]), .rectangle3_weight(rectangle3_weights[563]), .feature_threshold(feature_thresholds[563]), .feature_above(feature_aboves[563]), .feature_below(feature_belows[563]), .scan_win_std_dev(scan_win_std_dev[563]), .feature_accum(feature_accums[563]));
  accum_calculator ac564(.scan_win(scan_win564), .rectangle1_x(rectangle1_xs[564]), .rectangle1_y(rectangle1_ys[564]), .rectangle1_width(rectangle1_widths[564]), .rectangle1_height(rectangle1_heights[564]), .rectangle1_weight(rectangle1_weights[564]), .rectangle2_x(rectangle2_xs[564]), .rectangle2_y(rectangle2_ys[564]), .rectangle2_width(rectangle2_widths[564]), .rectangle2_height(rectangle2_heights[564]), .rectangle2_weight(rectangle2_weights[564]), .rectangle3_x(rectangle3_xs[564]), .rectangle3_y(rectangle3_ys[564]), .rectangle3_width(rectangle3_widths[564]), .rectangle3_height(rectangle3_heights[564]), .rectangle3_weight(rectangle3_weights[564]), .feature_threshold(feature_thresholds[564]), .feature_above(feature_aboves[564]), .feature_below(feature_belows[564]), .scan_win_std_dev(scan_win_std_dev[564]), .feature_accum(feature_accums[564]));
  accum_calculator ac565(.scan_win(scan_win565), .rectangle1_x(rectangle1_xs[565]), .rectangle1_y(rectangle1_ys[565]), .rectangle1_width(rectangle1_widths[565]), .rectangle1_height(rectangle1_heights[565]), .rectangle1_weight(rectangle1_weights[565]), .rectangle2_x(rectangle2_xs[565]), .rectangle2_y(rectangle2_ys[565]), .rectangle2_width(rectangle2_widths[565]), .rectangle2_height(rectangle2_heights[565]), .rectangle2_weight(rectangle2_weights[565]), .rectangle3_x(rectangle3_xs[565]), .rectangle3_y(rectangle3_ys[565]), .rectangle3_width(rectangle3_widths[565]), .rectangle3_height(rectangle3_heights[565]), .rectangle3_weight(rectangle3_weights[565]), .feature_threshold(feature_thresholds[565]), .feature_above(feature_aboves[565]), .feature_below(feature_belows[565]), .scan_win_std_dev(scan_win_std_dev[565]), .feature_accum(feature_accums[565]));
  accum_calculator ac566(.scan_win(scan_win566), .rectangle1_x(rectangle1_xs[566]), .rectangle1_y(rectangle1_ys[566]), .rectangle1_width(rectangle1_widths[566]), .rectangle1_height(rectangle1_heights[566]), .rectangle1_weight(rectangle1_weights[566]), .rectangle2_x(rectangle2_xs[566]), .rectangle2_y(rectangle2_ys[566]), .rectangle2_width(rectangle2_widths[566]), .rectangle2_height(rectangle2_heights[566]), .rectangle2_weight(rectangle2_weights[566]), .rectangle3_x(rectangle3_xs[566]), .rectangle3_y(rectangle3_ys[566]), .rectangle3_width(rectangle3_widths[566]), .rectangle3_height(rectangle3_heights[566]), .rectangle3_weight(rectangle3_weights[566]), .feature_threshold(feature_thresholds[566]), .feature_above(feature_aboves[566]), .feature_below(feature_belows[566]), .scan_win_std_dev(scan_win_std_dev[566]), .feature_accum(feature_accums[566]));
  accum_calculator ac567(.scan_win(scan_win567), .rectangle1_x(rectangle1_xs[567]), .rectangle1_y(rectangle1_ys[567]), .rectangle1_width(rectangle1_widths[567]), .rectangle1_height(rectangle1_heights[567]), .rectangle1_weight(rectangle1_weights[567]), .rectangle2_x(rectangle2_xs[567]), .rectangle2_y(rectangle2_ys[567]), .rectangle2_width(rectangle2_widths[567]), .rectangle2_height(rectangle2_heights[567]), .rectangle2_weight(rectangle2_weights[567]), .rectangle3_x(rectangle3_xs[567]), .rectangle3_y(rectangle3_ys[567]), .rectangle3_width(rectangle3_widths[567]), .rectangle3_height(rectangle3_heights[567]), .rectangle3_weight(rectangle3_weights[567]), .feature_threshold(feature_thresholds[567]), .feature_above(feature_aboves[567]), .feature_below(feature_belows[567]), .scan_win_std_dev(scan_win_std_dev[567]), .feature_accum(feature_accums[567]));
  accum_calculator ac568(.scan_win(scan_win568), .rectangle1_x(rectangle1_xs[568]), .rectangle1_y(rectangle1_ys[568]), .rectangle1_width(rectangle1_widths[568]), .rectangle1_height(rectangle1_heights[568]), .rectangle1_weight(rectangle1_weights[568]), .rectangle2_x(rectangle2_xs[568]), .rectangle2_y(rectangle2_ys[568]), .rectangle2_width(rectangle2_widths[568]), .rectangle2_height(rectangle2_heights[568]), .rectangle2_weight(rectangle2_weights[568]), .rectangle3_x(rectangle3_xs[568]), .rectangle3_y(rectangle3_ys[568]), .rectangle3_width(rectangle3_widths[568]), .rectangle3_height(rectangle3_heights[568]), .rectangle3_weight(rectangle3_weights[568]), .feature_threshold(feature_thresholds[568]), .feature_above(feature_aboves[568]), .feature_below(feature_belows[568]), .scan_win_std_dev(scan_win_std_dev[568]), .feature_accum(feature_accums[568]));
  accum_calculator ac569(.scan_win(scan_win569), .rectangle1_x(rectangle1_xs[569]), .rectangle1_y(rectangle1_ys[569]), .rectangle1_width(rectangle1_widths[569]), .rectangle1_height(rectangle1_heights[569]), .rectangle1_weight(rectangle1_weights[569]), .rectangle2_x(rectangle2_xs[569]), .rectangle2_y(rectangle2_ys[569]), .rectangle2_width(rectangle2_widths[569]), .rectangle2_height(rectangle2_heights[569]), .rectangle2_weight(rectangle2_weights[569]), .rectangle3_x(rectangle3_xs[569]), .rectangle3_y(rectangle3_ys[569]), .rectangle3_width(rectangle3_widths[569]), .rectangle3_height(rectangle3_heights[569]), .rectangle3_weight(rectangle3_weights[569]), .feature_threshold(feature_thresholds[569]), .feature_above(feature_aboves[569]), .feature_below(feature_belows[569]), .scan_win_std_dev(scan_win_std_dev[569]), .feature_accum(feature_accums[569]));
  accum_calculator ac570(.scan_win(scan_win570), .rectangle1_x(rectangle1_xs[570]), .rectangle1_y(rectangle1_ys[570]), .rectangle1_width(rectangle1_widths[570]), .rectangle1_height(rectangle1_heights[570]), .rectangle1_weight(rectangle1_weights[570]), .rectangle2_x(rectangle2_xs[570]), .rectangle2_y(rectangle2_ys[570]), .rectangle2_width(rectangle2_widths[570]), .rectangle2_height(rectangle2_heights[570]), .rectangle2_weight(rectangle2_weights[570]), .rectangle3_x(rectangle3_xs[570]), .rectangle3_y(rectangle3_ys[570]), .rectangle3_width(rectangle3_widths[570]), .rectangle3_height(rectangle3_heights[570]), .rectangle3_weight(rectangle3_weights[570]), .feature_threshold(feature_thresholds[570]), .feature_above(feature_aboves[570]), .feature_below(feature_belows[570]), .scan_win_std_dev(scan_win_std_dev[570]), .feature_accum(feature_accums[570]));
  accum_calculator ac571(.scan_win(scan_win571), .rectangle1_x(rectangle1_xs[571]), .rectangle1_y(rectangle1_ys[571]), .rectangle1_width(rectangle1_widths[571]), .rectangle1_height(rectangle1_heights[571]), .rectangle1_weight(rectangle1_weights[571]), .rectangle2_x(rectangle2_xs[571]), .rectangle2_y(rectangle2_ys[571]), .rectangle2_width(rectangle2_widths[571]), .rectangle2_height(rectangle2_heights[571]), .rectangle2_weight(rectangle2_weights[571]), .rectangle3_x(rectangle3_xs[571]), .rectangle3_y(rectangle3_ys[571]), .rectangle3_width(rectangle3_widths[571]), .rectangle3_height(rectangle3_heights[571]), .rectangle3_weight(rectangle3_weights[571]), .feature_threshold(feature_thresholds[571]), .feature_above(feature_aboves[571]), .feature_below(feature_belows[571]), .scan_win_std_dev(scan_win_std_dev[571]), .feature_accum(feature_accums[571]));
  accum_calculator ac572(.scan_win(scan_win572), .rectangle1_x(rectangle1_xs[572]), .rectangle1_y(rectangle1_ys[572]), .rectangle1_width(rectangle1_widths[572]), .rectangle1_height(rectangle1_heights[572]), .rectangle1_weight(rectangle1_weights[572]), .rectangle2_x(rectangle2_xs[572]), .rectangle2_y(rectangle2_ys[572]), .rectangle2_width(rectangle2_widths[572]), .rectangle2_height(rectangle2_heights[572]), .rectangle2_weight(rectangle2_weights[572]), .rectangle3_x(rectangle3_xs[572]), .rectangle3_y(rectangle3_ys[572]), .rectangle3_width(rectangle3_widths[572]), .rectangle3_height(rectangle3_heights[572]), .rectangle3_weight(rectangle3_weights[572]), .feature_threshold(feature_thresholds[572]), .feature_above(feature_aboves[572]), .feature_below(feature_belows[572]), .scan_win_std_dev(scan_win_std_dev[572]), .feature_accum(feature_accums[572]));
  accum_calculator ac573(.scan_win(scan_win573), .rectangle1_x(rectangle1_xs[573]), .rectangle1_y(rectangle1_ys[573]), .rectangle1_width(rectangle1_widths[573]), .rectangle1_height(rectangle1_heights[573]), .rectangle1_weight(rectangle1_weights[573]), .rectangle2_x(rectangle2_xs[573]), .rectangle2_y(rectangle2_ys[573]), .rectangle2_width(rectangle2_widths[573]), .rectangle2_height(rectangle2_heights[573]), .rectangle2_weight(rectangle2_weights[573]), .rectangle3_x(rectangle3_xs[573]), .rectangle3_y(rectangle3_ys[573]), .rectangle3_width(rectangle3_widths[573]), .rectangle3_height(rectangle3_heights[573]), .rectangle3_weight(rectangle3_weights[573]), .feature_threshold(feature_thresholds[573]), .feature_above(feature_aboves[573]), .feature_below(feature_belows[573]), .scan_win_std_dev(scan_win_std_dev[573]), .feature_accum(feature_accums[573]));
  accum_calculator ac574(.scan_win(scan_win574), .rectangle1_x(rectangle1_xs[574]), .rectangle1_y(rectangle1_ys[574]), .rectangle1_width(rectangle1_widths[574]), .rectangle1_height(rectangle1_heights[574]), .rectangle1_weight(rectangle1_weights[574]), .rectangle2_x(rectangle2_xs[574]), .rectangle2_y(rectangle2_ys[574]), .rectangle2_width(rectangle2_widths[574]), .rectangle2_height(rectangle2_heights[574]), .rectangle2_weight(rectangle2_weights[574]), .rectangle3_x(rectangle3_xs[574]), .rectangle3_y(rectangle3_ys[574]), .rectangle3_width(rectangle3_widths[574]), .rectangle3_height(rectangle3_heights[574]), .rectangle3_weight(rectangle3_weights[574]), .feature_threshold(feature_thresholds[574]), .feature_above(feature_aboves[574]), .feature_below(feature_belows[574]), .scan_win_std_dev(scan_win_std_dev[574]), .feature_accum(feature_accums[574]));
  accum_calculator ac575(.scan_win(scan_win575), .rectangle1_x(rectangle1_xs[575]), .rectangle1_y(rectangle1_ys[575]), .rectangle1_width(rectangle1_widths[575]), .rectangle1_height(rectangle1_heights[575]), .rectangle1_weight(rectangle1_weights[575]), .rectangle2_x(rectangle2_xs[575]), .rectangle2_y(rectangle2_ys[575]), .rectangle2_width(rectangle2_widths[575]), .rectangle2_height(rectangle2_heights[575]), .rectangle2_weight(rectangle2_weights[575]), .rectangle3_x(rectangle3_xs[575]), .rectangle3_y(rectangle3_ys[575]), .rectangle3_width(rectangle3_widths[575]), .rectangle3_height(rectangle3_heights[575]), .rectangle3_weight(rectangle3_weights[575]), .feature_threshold(feature_thresholds[575]), .feature_above(feature_aboves[575]), .feature_below(feature_belows[575]), .scan_win_std_dev(scan_win_std_dev[575]), .feature_accum(feature_accums[575]));
  accum_calculator ac576(.scan_win(scan_win576), .rectangle1_x(rectangle1_xs[576]), .rectangle1_y(rectangle1_ys[576]), .rectangle1_width(rectangle1_widths[576]), .rectangle1_height(rectangle1_heights[576]), .rectangle1_weight(rectangle1_weights[576]), .rectangle2_x(rectangle2_xs[576]), .rectangle2_y(rectangle2_ys[576]), .rectangle2_width(rectangle2_widths[576]), .rectangle2_height(rectangle2_heights[576]), .rectangle2_weight(rectangle2_weights[576]), .rectangle3_x(rectangle3_xs[576]), .rectangle3_y(rectangle3_ys[576]), .rectangle3_width(rectangle3_widths[576]), .rectangle3_height(rectangle3_heights[576]), .rectangle3_weight(rectangle3_weights[576]), .feature_threshold(feature_thresholds[576]), .feature_above(feature_aboves[576]), .feature_below(feature_belows[576]), .scan_win_std_dev(scan_win_std_dev[576]), .feature_accum(feature_accums[576]));
  accum_calculator ac577(.scan_win(scan_win577), .rectangle1_x(rectangle1_xs[577]), .rectangle1_y(rectangle1_ys[577]), .rectangle1_width(rectangle1_widths[577]), .rectangle1_height(rectangle1_heights[577]), .rectangle1_weight(rectangle1_weights[577]), .rectangle2_x(rectangle2_xs[577]), .rectangle2_y(rectangle2_ys[577]), .rectangle2_width(rectangle2_widths[577]), .rectangle2_height(rectangle2_heights[577]), .rectangle2_weight(rectangle2_weights[577]), .rectangle3_x(rectangle3_xs[577]), .rectangle3_y(rectangle3_ys[577]), .rectangle3_width(rectangle3_widths[577]), .rectangle3_height(rectangle3_heights[577]), .rectangle3_weight(rectangle3_weights[577]), .feature_threshold(feature_thresholds[577]), .feature_above(feature_aboves[577]), .feature_below(feature_belows[577]), .scan_win_std_dev(scan_win_std_dev[577]), .feature_accum(feature_accums[577]));
  accum_calculator ac578(.scan_win(scan_win578), .rectangle1_x(rectangle1_xs[578]), .rectangle1_y(rectangle1_ys[578]), .rectangle1_width(rectangle1_widths[578]), .rectangle1_height(rectangle1_heights[578]), .rectangle1_weight(rectangle1_weights[578]), .rectangle2_x(rectangle2_xs[578]), .rectangle2_y(rectangle2_ys[578]), .rectangle2_width(rectangle2_widths[578]), .rectangle2_height(rectangle2_heights[578]), .rectangle2_weight(rectangle2_weights[578]), .rectangle3_x(rectangle3_xs[578]), .rectangle3_y(rectangle3_ys[578]), .rectangle3_width(rectangle3_widths[578]), .rectangle3_height(rectangle3_heights[578]), .rectangle3_weight(rectangle3_weights[578]), .feature_threshold(feature_thresholds[578]), .feature_above(feature_aboves[578]), .feature_below(feature_belows[578]), .scan_win_std_dev(scan_win_std_dev[578]), .feature_accum(feature_accums[578]));
  accum_calculator ac579(.scan_win(scan_win579), .rectangle1_x(rectangle1_xs[579]), .rectangle1_y(rectangle1_ys[579]), .rectangle1_width(rectangle1_widths[579]), .rectangle1_height(rectangle1_heights[579]), .rectangle1_weight(rectangle1_weights[579]), .rectangle2_x(rectangle2_xs[579]), .rectangle2_y(rectangle2_ys[579]), .rectangle2_width(rectangle2_widths[579]), .rectangle2_height(rectangle2_heights[579]), .rectangle2_weight(rectangle2_weights[579]), .rectangle3_x(rectangle3_xs[579]), .rectangle3_y(rectangle3_ys[579]), .rectangle3_width(rectangle3_widths[579]), .rectangle3_height(rectangle3_heights[579]), .rectangle3_weight(rectangle3_weights[579]), .feature_threshold(feature_thresholds[579]), .feature_above(feature_aboves[579]), .feature_below(feature_belows[579]), .scan_win_std_dev(scan_win_std_dev[579]), .feature_accum(feature_accums[579]));
  accum_calculator ac580(.scan_win(scan_win580), .rectangle1_x(rectangle1_xs[580]), .rectangle1_y(rectangle1_ys[580]), .rectangle1_width(rectangle1_widths[580]), .rectangle1_height(rectangle1_heights[580]), .rectangle1_weight(rectangle1_weights[580]), .rectangle2_x(rectangle2_xs[580]), .rectangle2_y(rectangle2_ys[580]), .rectangle2_width(rectangle2_widths[580]), .rectangle2_height(rectangle2_heights[580]), .rectangle2_weight(rectangle2_weights[580]), .rectangle3_x(rectangle3_xs[580]), .rectangle3_y(rectangle3_ys[580]), .rectangle3_width(rectangle3_widths[580]), .rectangle3_height(rectangle3_heights[580]), .rectangle3_weight(rectangle3_weights[580]), .feature_threshold(feature_thresholds[580]), .feature_above(feature_aboves[580]), .feature_below(feature_belows[580]), .scan_win_std_dev(scan_win_std_dev[580]), .feature_accum(feature_accums[580]));
  accum_calculator ac581(.scan_win(scan_win581), .rectangle1_x(rectangle1_xs[581]), .rectangle1_y(rectangle1_ys[581]), .rectangle1_width(rectangle1_widths[581]), .rectangle1_height(rectangle1_heights[581]), .rectangle1_weight(rectangle1_weights[581]), .rectangle2_x(rectangle2_xs[581]), .rectangle2_y(rectangle2_ys[581]), .rectangle2_width(rectangle2_widths[581]), .rectangle2_height(rectangle2_heights[581]), .rectangle2_weight(rectangle2_weights[581]), .rectangle3_x(rectangle3_xs[581]), .rectangle3_y(rectangle3_ys[581]), .rectangle3_width(rectangle3_widths[581]), .rectangle3_height(rectangle3_heights[581]), .rectangle3_weight(rectangle3_weights[581]), .feature_threshold(feature_thresholds[581]), .feature_above(feature_aboves[581]), .feature_below(feature_belows[581]), .scan_win_std_dev(scan_win_std_dev[581]), .feature_accum(feature_accums[581]));
  accum_calculator ac582(.scan_win(scan_win582), .rectangle1_x(rectangle1_xs[582]), .rectangle1_y(rectangle1_ys[582]), .rectangle1_width(rectangle1_widths[582]), .rectangle1_height(rectangle1_heights[582]), .rectangle1_weight(rectangle1_weights[582]), .rectangle2_x(rectangle2_xs[582]), .rectangle2_y(rectangle2_ys[582]), .rectangle2_width(rectangle2_widths[582]), .rectangle2_height(rectangle2_heights[582]), .rectangle2_weight(rectangle2_weights[582]), .rectangle3_x(rectangle3_xs[582]), .rectangle3_y(rectangle3_ys[582]), .rectangle3_width(rectangle3_widths[582]), .rectangle3_height(rectangle3_heights[582]), .rectangle3_weight(rectangle3_weights[582]), .feature_threshold(feature_thresholds[582]), .feature_above(feature_aboves[582]), .feature_below(feature_belows[582]), .scan_win_std_dev(scan_win_std_dev[582]), .feature_accum(feature_accums[582]));
  accum_calculator ac583(.scan_win(scan_win583), .rectangle1_x(rectangle1_xs[583]), .rectangle1_y(rectangle1_ys[583]), .rectangle1_width(rectangle1_widths[583]), .rectangle1_height(rectangle1_heights[583]), .rectangle1_weight(rectangle1_weights[583]), .rectangle2_x(rectangle2_xs[583]), .rectangle2_y(rectangle2_ys[583]), .rectangle2_width(rectangle2_widths[583]), .rectangle2_height(rectangle2_heights[583]), .rectangle2_weight(rectangle2_weights[583]), .rectangle3_x(rectangle3_xs[583]), .rectangle3_y(rectangle3_ys[583]), .rectangle3_width(rectangle3_widths[583]), .rectangle3_height(rectangle3_heights[583]), .rectangle3_weight(rectangle3_weights[583]), .feature_threshold(feature_thresholds[583]), .feature_above(feature_aboves[583]), .feature_below(feature_belows[583]), .scan_win_std_dev(scan_win_std_dev[583]), .feature_accum(feature_accums[583]));
  accum_calculator ac584(.scan_win(scan_win584), .rectangle1_x(rectangle1_xs[584]), .rectangle1_y(rectangle1_ys[584]), .rectangle1_width(rectangle1_widths[584]), .rectangle1_height(rectangle1_heights[584]), .rectangle1_weight(rectangle1_weights[584]), .rectangle2_x(rectangle2_xs[584]), .rectangle2_y(rectangle2_ys[584]), .rectangle2_width(rectangle2_widths[584]), .rectangle2_height(rectangle2_heights[584]), .rectangle2_weight(rectangle2_weights[584]), .rectangle3_x(rectangle3_xs[584]), .rectangle3_y(rectangle3_ys[584]), .rectangle3_width(rectangle3_widths[584]), .rectangle3_height(rectangle3_heights[584]), .rectangle3_weight(rectangle3_weights[584]), .feature_threshold(feature_thresholds[584]), .feature_above(feature_aboves[584]), .feature_below(feature_belows[584]), .scan_win_std_dev(scan_win_std_dev[584]), .feature_accum(feature_accums[584]));
  accum_calculator ac585(.scan_win(scan_win585), .rectangle1_x(rectangle1_xs[585]), .rectangle1_y(rectangle1_ys[585]), .rectangle1_width(rectangle1_widths[585]), .rectangle1_height(rectangle1_heights[585]), .rectangle1_weight(rectangle1_weights[585]), .rectangle2_x(rectangle2_xs[585]), .rectangle2_y(rectangle2_ys[585]), .rectangle2_width(rectangle2_widths[585]), .rectangle2_height(rectangle2_heights[585]), .rectangle2_weight(rectangle2_weights[585]), .rectangle3_x(rectangle3_xs[585]), .rectangle3_y(rectangle3_ys[585]), .rectangle3_width(rectangle3_widths[585]), .rectangle3_height(rectangle3_heights[585]), .rectangle3_weight(rectangle3_weights[585]), .feature_threshold(feature_thresholds[585]), .feature_above(feature_aboves[585]), .feature_below(feature_belows[585]), .scan_win_std_dev(scan_win_std_dev[585]), .feature_accum(feature_accums[585]));
  accum_calculator ac586(.scan_win(scan_win586), .rectangle1_x(rectangle1_xs[586]), .rectangle1_y(rectangle1_ys[586]), .rectangle1_width(rectangle1_widths[586]), .rectangle1_height(rectangle1_heights[586]), .rectangle1_weight(rectangle1_weights[586]), .rectangle2_x(rectangle2_xs[586]), .rectangle2_y(rectangle2_ys[586]), .rectangle2_width(rectangle2_widths[586]), .rectangle2_height(rectangle2_heights[586]), .rectangle2_weight(rectangle2_weights[586]), .rectangle3_x(rectangle3_xs[586]), .rectangle3_y(rectangle3_ys[586]), .rectangle3_width(rectangle3_widths[586]), .rectangle3_height(rectangle3_heights[586]), .rectangle3_weight(rectangle3_weights[586]), .feature_threshold(feature_thresholds[586]), .feature_above(feature_aboves[586]), .feature_below(feature_belows[586]), .scan_win_std_dev(scan_win_std_dev[586]), .feature_accum(feature_accums[586]));
  accum_calculator ac587(.scan_win(scan_win587), .rectangle1_x(rectangle1_xs[587]), .rectangle1_y(rectangle1_ys[587]), .rectangle1_width(rectangle1_widths[587]), .rectangle1_height(rectangle1_heights[587]), .rectangle1_weight(rectangle1_weights[587]), .rectangle2_x(rectangle2_xs[587]), .rectangle2_y(rectangle2_ys[587]), .rectangle2_width(rectangle2_widths[587]), .rectangle2_height(rectangle2_heights[587]), .rectangle2_weight(rectangle2_weights[587]), .rectangle3_x(rectangle3_xs[587]), .rectangle3_y(rectangle3_ys[587]), .rectangle3_width(rectangle3_widths[587]), .rectangle3_height(rectangle3_heights[587]), .rectangle3_weight(rectangle3_weights[587]), .feature_threshold(feature_thresholds[587]), .feature_above(feature_aboves[587]), .feature_below(feature_belows[587]), .scan_win_std_dev(scan_win_std_dev[587]), .feature_accum(feature_accums[587]));
  accum_calculator ac588(.scan_win(scan_win588), .rectangle1_x(rectangle1_xs[588]), .rectangle1_y(rectangle1_ys[588]), .rectangle1_width(rectangle1_widths[588]), .rectangle1_height(rectangle1_heights[588]), .rectangle1_weight(rectangle1_weights[588]), .rectangle2_x(rectangle2_xs[588]), .rectangle2_y(rectangle2_ys[588]), .rectangle2_width(rectangle2_widths[588]), .rectangle2_height(rectangle2_heights[588]), .rectangle2_weight(rectangle2_weights[588]), .rectangle3_x(rectangle3_xs[588]), .rectangle3_y(rectangle3_ys[588]), .rectangle3_width(rectangle3_widths[588]), .rectangle3_height(rectangle3_heights[588]), .rectangle3_weight(rectangle3_weights[588]), .feature_threshold(feature_thresholds[588]), .feature_above(feature_aboves[588]), .feature_below(feature_belows[588]), .scan_win_std_dev(scan_win_std_dev[588]), .feature_accum(feature_accums[588]));
  accum_calculator ac589(.scan_win(scan_win589), .rectangle1_x(rectangle1_xs[589]), .rectangle1_y(rectangle1_ys[589]), .rectangle1_width(rectangle1_widths[589]), .rectangle1_height(rectangle1_heights[589]), .rectangle1_weight(rectangle1_weights[589]), .rectangle2_x(rectangle2_xs[589]), .rectangle2_y(rectangle2_ys[589]), .rectangle2_width(rectangle2_widths[589]), .rectangle2_height(rectangle2_heights[589]), .rectangle2_weight(rectangle2_weights[589]), .rectangle3_x(rectangle3_xs[589]), .rectangle3_y(rectangle3_ys[589]), .rectangle3_width(rectangle3_widths[589]), .rectangle3_height(rectangle3_heights[589]), .rectangle3_weight(rectangle3_weights[589]), .feature_threshold(feature_thresholds[589]), .feature_above(feature_aboves[589]), .feature_below(feature_belows[589]), .scan_win_std_dev(scan_win_std_dev[589]), .feature_accum(feature_accums[589]));
  accum_calculator ac590(.scan_win(scan_win590), .rectangle1_x(rectangle1_xs[590]), .rectangle1_y(rectangle1_ys[590]), .rectangle1_width(rectangle1_widths[590]), .rectangle1_height(rectangle1_heights[590]), .rectangle1_weight(rectangle1_weights[590]), .rectangle2_x(rectangle2_xs[590]), .rectangle2_y(rectangle2_ys[590]), .rectangle2_width(rectangle2_widths[590]), .rectangle2_height(rectangle2_heights[590]), .rectangle2_weight(rectangle2_weights[590]), .rectangle3_x(rectangle3_xs[590]), .rectangle3_y(rectangle3_ys[590]), .rectangle3_width(rectangle3_widths[590]), .rectangle3_height(rectangle3_heights[590]), .rectangle3_weight(rectangle3_weights[590]), .feature_threshold(feature_thresholds[590]), .feature_above(feature_aboves[590]), .feature_below(feature_belows[590]), .scan_win_std_dev(scan_win_std_dev[590]), .feature_accum(feature_accums[590]));
  accum_calculator ac591(.scan_win(scan_win591), .rectangle1_x(rectangle1_xs[591]), .rectangle1_y(rectangle1_ys[591]), .rectangle1_width(rectangle1_widths[591]), .rectangle1_height(rectangle1_heights[591]), .rectangle1_weight(rectangle1_weights[591]), .rectangle2_x(rectangle2_xs[591]), .rectangle2_y(rectangle2_ys[591]), .rectangle2_width(rectangle2_widths[591]), .rectangle2_height(rectangle2_heights[591]), .rectangle2_weight(rectangle2_weights[591]), .rectangle3_x(rectangle3_xs[591]), .rectangle3_y(rectangle3_ys[591]), .rectangle3_width(rectangle3_widths[591]), .rectangle3_height(rectangle3_heights[591]), .rectangle3_weight(rectangle3_weights[591]), .feature_threshold(feature_thresholds[591]), .feature_above(feature_aboves[591]), .feature_below(feature_belows[591]), .scan_win_std_dev(scan_win_std_dev[591]), .feature_accum(feature_accums[591]));
  accum_calculator ac592(.scan_win(scan_win592), .rectangle1_x(rectangle1_xs[592]), .rectangle1_y(rectangle1_ys[592]), .rectangle1_width(rectangle1_widths[592]), .rectangle1_height(rectangle1_heights[592]), .rectangle1_weight(rectangle1_weights[592]), .rectangle2_x(rectangle2_xs[592]), .rectangle2_y(rectangle2_ys[592]), .rectangle2_width(rectangle2_widths[592]), .rectangle2_height(rectangle2_heights[592]), .rectangle2_weight(rectangle2_weights[592]), .rectangle3_x(rectangle3_xs[592]), .rectangle3_y(rectangle3_ys[592]), .rectangle3_width(rectangle3_widths[592]), .rectangle3_height(rectangle3_heights[592]), .rectangle3_weight(rectangle3_weights[592]), .feature_threshold(feature_thresholds[592]), .feature_above(feature_aboves[592]), .feature_below(feature_belows[592]), .scan_win_std_dev(scan_win_std_dev[592]), .feature_accum(feature_accums[592]));
  accum_calculator ac593(.scan_win(scan_win593), .rectangle1_x(rectangle1_xs[593]), .rectangle1_y(rectangle1_ys[593]), .rectangle1_width(rectangle1_widths[593]), .rectangle1_height(rectangle1_heights[593]), .rectangle1_weight(rectangle1_weights[593]), .rectangle2_x(rectangle2_xs[593]), .rectangle2_y(rectangle2_ys[593]), .rectangle2_width(rectangle2_widths[593]), .rectangle2_height(rectangle2_heights[593]), .rectangle2_weight(rectangle2_weights[593]), .rectangle3_x(rectangle3_xs[593]), .rectangle3_y(rectangle3_ys[593]), .rectangle3_width(rectangle3_widths[593]), .rectangle3_height(rectangle3_heights[593]), .rectangle3_weight(rectangle3_weights[593]), .feature_threshold(feature_thresholds[593]), .feature_above(feature_aboves[593]), .feature_below(feature_belows[593]), .scan_win_std_dev(scan_win_std_dev[593]), .feature_accum(feature_accums[593]));
  accum_calculator ac594(.scan_win(scan_win594), .rectangle1_x(rectangle1_xs[594]), .rectangle1_y(rectangle1_ys[594]), .rectangle1_width(rectangle1_widths[594]), .rectangle1_height(rectangle1_heights[594]), .rectangle1_weight(rectangle1_weights[594]), .rectangle2_x(rectangle2_xs[594]), .rectangle2_y(rectangle2_ys[594]), .rectangle2_width(rectangle2_widths[594]), .rectangle2_height(rectangle2_heights[594]), .rectangle2_weight(rectangle2_weights[594]), .rectangle3_x(rectangle3_xs[594]), .rectangle3_y(rectangle3_ys[594]), .rectangle3_width(rectangle3_widths[594]), .rectangle3_height(rectangle3_heights[594]), .rectangle3_weight(rectangle3_weights[594]), .feature_threshold(feature_thresholds[594]), .feature_above(feature_aboves[594]), .feature_below(feature_belows[594]), .scan_win_std_dev(scan_win_std_dev[594]), .feature_accum(feature_accums[594]));
  accum_calculator ac595(.scan_win(scan_win595), .rectangle1_x(rectangle1_xs[595]), .rectangle1_y(rectangle1_ys[595]), .rectangle1_width(rectangle1_widths[595]), .rectangle1_height(rectangle1_heights[595]), .rectangle1_weight(rectangle1_weights[595]), .rectangle2_x(rectangle2_xs[595]), .rectangle2_y(rectangle2_ys[595]), .rectangle2_width(rectangle2_widths[595]), .rectangle2_height(rectangle2_heights[595]), .rectangle2_weight(rectangle2_weights[595]), .rectangle3_x(rectangle3_xs[595]), .rectangle3_y(rectangle3_ys[595]), .rectangle3_width(rectangle3_widths[595]), .rectangle3_height(rectangle3_heights[595]), .rectangle3_weight(rectangle3_weights[595]), .feature_threshold(feature_thresholds[595]), .feature_above(feature_aboves[595]), .feature_below(feature_belows[595]), .scan_win_std_dev(scan_win_std_dev[595]), .feature_accum(feature_accums[595]));
  accum_calculator ac596(.scan_win(scan_win596), .rectangle1_x(rectangle1_xs[596]), .rectangle1_y(rectangle1_ys[596]), .rectangle1_width(rectangle1_widths[596]), .rectangle1_height(rectangle1_heights[596]), .rectangle1_weight(rectangle1_weights[596]), .rectangle2_x(rectangle2_xs[596]), .rectangle2_y(rectangle2_ys[596]), .rectangle2_width(rectangle2_widths[596]), .rectangle2_height(rectangle2_heights[596]), .rectangle2_weight(rectangle2_weights[596]), .rectangle3_x(rectangle3_xs[596]), .rectangle3_y(rectangle3_ys[596]), .rectangle3_width(rectangle3_widths[596]), .rectangle3_height(rectangle3_heights[596]), .rectangle3_weight(rectangle3_weights[596]), .feature_threshold(feature_thresholds[596]), .feature_above(feature_aboves[596]), .feature_below(feature_belows[596]), .scan_win_std_dev(scan_win_std_dev[596]), .feature_accum(feature_accums[596]));
  accum_calculator ac597(.scan_win(scan_win597), .rectangle1_x(rectangle1_xs[597]), .rectangle1_y(rectangle1_ys[597]), .rectangle1_width(rectangle1_widths[597]), .rectangle1_height(rectangle1_heights[597]), .rectangle1_weight(rectangle1_weights[597]), .rectangle2_x(rectangle2_xs[597]), .rectangle2_y(rectangle2_ys[597]), .rectangle2_width(rectangle2_widths[597]), .rectangle2_height(rectangle2_heights[597]), .rectangle2_weight(rectangle2_weights[597]), .rectangle3_x(rectangle3_xs[597]), .rectangle3_y(rectangle3_ys[597]), .rectangle3_width(rectangle3_widths[597]), .rectangle3_height(rectangle3_heights[597]), .rectangle3_weight(rectangle3_weights[597]), .feature_threshold(feature_thresholds[597]), .feature_above(feature_aboves[597]), .feature_below(feature_belows[597]), .scan_win_std_dev(scan_win_std_dev[597]), .feature_accum(feature_accums[597]));
  accum_calculator ac598(.scan_win(scan_win598), .rectangle1_x(rectangle1_xs[598]), .rectangle1_y(rectangle1_ys[598]), .rectangle1_width(rectangle1_widths[598]), .rectangle1_height(rectangle1_heights[598]), .rectangle1_weight(rectangle1_weights[598]), .rectangle2_x(rectangle2_xs[598]), .rectangle2_y(rectangle2_ys[598]), .rectangle2_width(rectangle2_widths[598]), .rectangle2_height(rectangle2_heights[598]), .rectangle2_weight(rectangle2_weights[598]), .rectangle3_x(rectangle3_xs[598]), .rectangle3_y(rectangle3_ys[598]), .rectangle3_width(rectangle3_widths[598]), .rectangle3_height(rectangle3_heights[598]), .rectangle3_weight(rectangle3_weights[598]), .feature_threshold(feature_thresholds[598]), .feature_above(feature_aboves[598]), .feature_below(feature_belows[598]), .scan_win_std_dev(scan_win_std_dev[598]), .feature_accum(feature_accums[598]));
  accum_calculator ac599(.scan_win(scan_win599), .rectangle1_x(rectangle1_xs[599]), .rectangle1_y(rectangle1_ys[599]), .rectangle1_width(rectangle1_widths[599]), .rectangle1_height(rectangle1_heights[599]), .rectangle1_weight(rectangle1_weights[599]), .rectangle2_x(rectangle2_xs[599]), .rectangle2_y(rectangle2_ys[599]), .rectangle2_width(rectangle2_widths[599]), .rectangle2_height(rectangle2_heights[599]), .rectangle2_weight(rectangle2_weights[599]), .rectangle3_x(rectangle3_xs[599]), .rectangle3_y(rectangle3_ys[599]), .rectangle3_width(rectangle3_widths[599]), .rectangle3_height(rectangle3_heights[599]), .rectangle3_weight(rectangle3_weights[599]), .feature_threshold(feature_thresholds[599]), .feature_above(feature_aboves[599]), .feature_below(feature_belows[599]), .scan_win_std_dev(scan_win_std_dev[599]), .feature_accum(feature_accums[599]));
  accum_calculator ac600(.scan_win(scan_win600), .rectangle1_x(rectangle1_xs[600]), .rectangle1_y(rectangle1_ys[600]), .rectangle1_width(rectangle1_widths[600]), .rectangle1_height(rectangle1_heights[600]), .rectangle1_weight(rectangle1_weights[600]), .rectangle2_x(rectangle2_xs[600]), .rectangle2_y(rectangle2_ys[600]), .rectangle2_width(rectangle2_widths[600]), .rectangle2_height(rectangle2_heights[600]), .rectangle2_weight(rectangle2_weights[600]), .rectangle3_x(rectangle3_xs[600]), .rectangle3_y(rectangle3_ys[600]), .rectangle3_width(rectangle3_widths[600]), .rectangle3_height(rectangle3_heights[600]), .rectangle3_weight(rectangle3_weights[600]), .feature_threshold(feature_thresholds[600]), .feature_above(feature_aboves[600]), .feature_below(feature_belows[600]), .scan_win_std_dev(scan_win_std_dev[600]), .feature_accum(feature_accums[600]));
  accum_calculator ac601(.scan_win(scan_win601), .rectangle1_x(rectangle1_xs[601]), .rectangle1_y(rectangle1_ys[601]), .rectangle1_width(rectangle1_widths[601]), .rectangle1_height(rectangle1_heights[601]), .rectangle1_weight(rectangle1_weights[601]), .rectangle2_x(rectangle2_xs[601]), .rectangle2_y(rectangle2_ys[601]), .rectangle2_width(rectangle2_widths[601]), .rectangle2_height(rectangle2_heights[601]), .rectangle2_weight(rectangle2_weights[601]), .rectangle3_x(rectangle3_xs[601]), .rectangle3_y(rectangle3_ys[601]), .rectangle3_width(rectangle3_widths[601]), .rectangle3_height(rectangle3_heights[601]), .rectangle3_weight(rectangle3_weights[601]), .feature_threshold(feature_thresholds[601]), .feature_above(feature_aboves[601]), .feature_below(feature_belows[601]), .scan_win_std_dev(scan_win_std_dev[601]), .feature_accum(feature_accums[601]));
  accum_calculator ac602(.scan_win(scan_win602), .rectangle1_x(rectangle1_xs[602]), .rectangle1_y(rectangle1_ys[602]), .rectangle1_width(rectangle1_widths[602]), .rectangle1_height(rectangle1_heights[602]), .rectangle1_weight(rectangle1_weights[602]), .rectangle2_x(rectangle2_xs[602]), .rectangle2_y(rectangle2_ys[602]), .rectangle2_width(rectangle2_widths[602]), .rectangle2_height(rectangle2_heights[602]), .rectangle2_weight(rectangle2_weights[602]), .rectangle3_x(rectangle3_xs[602]), .rectangle3_y(rectangle3_ys[602]), .rectangle3_width(rectangle3_widths[602]), .rectangle3_height(rectangle3_heights[602]), .rectangle3_weight(rectangle3_weights[602]), .feature_threshold(feature_thresholds[602]), .feature_above(feature_aboves[602]), .feature_below(feature_belows[602]), .scan_win_std_dev(scan_win_std_dev[602]), .feature_accum(feature_accums[602]));
  accum_calculator ac603(.scan_win(scan_win603), .rectangle1_x(rectangle1_xs[603]), .rectangle1_y(rectangle1_ys[603]), .rectangle1_width(rectangle1_widths[603]), .rectangle1_height(rectangle1_heights[603]), .rectangle1_weight(rectangle1_weights[603]), .rectangle2_x(rectangle2_xs[603]), .rectangle2_y(rectangle2_ys[603]), .rectangle2_width(rectangle2_widths[603]), .rectangle2_height(rectangle2_heights[603]), .rectangle2_weight(rectangle2_weights[603]), .rectangle3_x(rectangle3_xs[603]), .rectangle3_y(rectangle3_ys[603]), .rectangle3_width(rectangle3_widths[603]), .rectangle3_height(rectangle3_heights[603]), .rectangle3_weight(rectangle3_weights[603]), .feature_threshold(feature_thresholds[603]), .feature_above(feature_aboves[603]), .feature_below(feature_belows[603]), .scan_win_std_dev(scan_win_std_dev[603]), .feature_accum(feature_accums[603]));
  accum_calculator ac604(.scan_win(scan_win604), .rectangle1_x(rectangle1_xs[604]), .rectangle1_y(rectangle1_ys[604]), .rectangle1_width(rectangle1_widths[604]), .rectangle1_height(rectangle1_heights[604]), .rectangle1_weight(rectangle1_weights[604]), .rectangle2_x(rectangle2_xs[604]), .rectangle2_y(rectangle2_ys[604]), .rectangle2_width(rectangle2_widths[604]), .rectangle2_height(rectangle2_heights[604]), .rectangle2_weight(rectangle2_weights[604]), .rectangle3_x(rectangle3_xs[604]), .rectangle3_y(rectangle3_ys[604]), .rectangle3_width(rectangle3_widths[604]), .rectangle3_height(rectangle3_heights[604]), .rectangle3_weight(rectangle3_weights[604]), .feature_threshold(feature_thresholds[604]), .feature_above(feature_aboves[604]), .feature_below(feature_belows[604]), .scan_win_std_dev(scan_win_std_dev[604]), .feature_accum(feature_accums[604]));
  accum_calculator ac605(.scan_win(scan_win605), .rectangle1_x(rectangle1_xs[605]), .rectangle1_y(rectangle1_ys[605]), .rectangle1_width(rectangle1_widths[605]), .rectangle1_height(rectangle1_heights[605]), .rectangle1_weight(rectangle1_weights[605]), .rectangle2_x(rectangle2_xs[605]), .rectangle2_y(rectangle2_ys[605]), .rectangle2_width(rectangle2_widths[605]), .rectangle2_height(rectangle2_heights[605]), .rectangle2_weight(rectangle2_weights[605]), .rectangle3_x(rectangle3_xs[605]), .rectangle3_y(rectangle3_ys[605]), .rectangle3_width(rectangle3_widths[605]), .rectangle3_height(rectangle3_heights[605]), .rectangle3_weight(rectangle3_weights[605]), .feature_threshold(feature_thresholds[605]), .feature_above(feature_aboves[605]), .feature_below(feature_belows[605]), .scan_win_std_dev(scan_win_std_dev[605]), .feature_accum(feature_accums[605]));
  accum_calculator ac606(.scan_win(scan_win606), .rectangle1_x(rectangle1_xs[606]), .rectangle1_y(rectangle1_ys[606]), .rectangle1_width(rectangle1_widths[606]), .rectangle1_height(rectangle1_heights[606]), .rectangle1_weight(rectangle1_weights[606]), .rectangle2_x(rectangle2_xs[606]), .rectangle2_y(rectangle2_ys[606]), .rectangle2_width(rectangle2_widths[606]), .rectangle2_height(rectangle2_heights[606]), .rectangle2_weight(rectangle2_weights[606]), .rectangle3_x(rectangle3_xs[606]), .rectangle3_y(rectangle3_ys[606]), .rectangle3_width(rectangle3_widths[606]), .rectangle3_height(rectangle3_heights[606]), .rectangle3_weight(rectangle3_weights[606]), .feature_threshold(feature_thresholds[606]), .feature_above(feature_aboves[606]), .feature_below(feature_belows[606]), .scan_win_std_dev(scan_win_std_dev[606]), .feature_accum(feature_accums[606]));
  accum_calculator ac607(.scan_win(scan_win607), .rectangle1_x(rectangle1_xs[607]), .rectangle1_y(rectangle1_ys[607]), .rectangle1_width(rectangle1_widths[607]), .rectangle1_height(rectangle1_heights[607]), .rectangle1_weight(rectangle1_weights[607]), .rectangle2_x(rectangle2_xs[607]), .rectangle2_y(rectangle2_ys[607]), .rectangle2_width(rectangle2_widths[607]), .rectangle2_height(rectangle2_heights[607]), .rectangle2_weight(rectangle2_weights[607]), .rectangle3_x(rectangle3_xs[607]), .rectangle3_y(rectangle3_ys[607]), .rectangle3_width(rectangle3_widths[607]), .rectangle3_height(rectangle3_heights[607]), .rectangle3_weight(rectangle3_weights[607]), .feature_threshold(feature_thresholds[607]), .feature_above(feature_aboves[607]), .feature_below(feature_belows[607]), .scan_win_std_dev(scan_win_std_dev[607]), .feature_accum(feature_accums[607]));
  accum_calculator ac608(.scan_win(scan_win608), .rectangle1_x(rectangle1_xs[608]), .rectangle1_y(rectangle1_ys[608]), .rectangle1_width(rectangle1_widths[608]), .rectangle1_height(rectangle1_heights[608]), .rectangle1_weight(rectangle1_weights[608]), .rectangle2_x(rectangle2_xs[608]), .rectangle2_y(rectangle2_ys[608]), .rectangle2_width(rectangle2_widths[608]), .rectangle2_height(rectangle2_heights[608]), .rectangle2_weight(rectangle2_weights[608]), .rectangle3_x(rectangle3_xs[608]), .rectangle3_y(rectangle3_ys[608]), .rectangle3_width(rectangle3_widths[608]), .rectangle3_height(rectangle3_heights[608]), .rectangle3_weight(rectangle3_weights[608]), .feature_threshold(feature_thresholds[608]), .feature_above(feature_aboves[608]), .feature_below(feature_belows[608]), .scan_win_std_dev(scan_win_std_dev[608]), .feature_accum(feature_accums[608]));
  accum_calculator ac609(.scan_win(scan_win609), .rectangle1_x(rectangle1_xs[609]), .rectangle1_y(rectangle1_ys[609]), .rectangle1_width(rectangle1_widths[609]), .rectangle1_height(rectangle1_heights[609]), .rectangle1_weight(rectangle1_weights[609]), .rectangle2_x(rectangle2_xs[609]), .rectangle2_y(rectangle2_ys[609]), .rectangle2_width(rectangle2_widths[609]), .rectangle2_height(rectangle2_heights[609]), .rectangle2_weight(rectangle2_weights[609]), .rectangle3_x(rectangle3_xs[609]), .rectangle3_y(rectangle3_ys[609]), .rectangle3_width(rectangle3_widths[609]), .rectangle3_height(rectangle3_heights[609]), .rectangle3_weight(rectangle3_weights[609]), .feature_threshold(feature_thresholds[609]), .feature_above(feature_aboves[609]), .feature_below(feature_belows[609]), .scan_win_std_dev(scan_win_std_dev[609]), .feature_accum(feature_accums[609]));
  accum_calculator ac610(.scan_win(scan_win610), .rectangle1_x(rectangle1_xs[610]), .rectangle1_y(rectangle1_ys[610]), .rectangle1_width(rectangle1_widths[610]), .rectangle1_height(rectangle1_heights[610]), .rectangle1_weight(rectangle1_weights[610]), .rectangle2_x(rectangle2_xs[610]), .rectangle2_y(rectangle2_ys[610]), .rectangle2_width(rectangle2_widths[610]), .rectangle2_height(rectangle2_heights[610]), .rectangle2_weight(rectangle2_weights[610]), .rectangle3_x(rectangle3_xs[610]), .rectangle3_y(rectangle3_ys[610]), .rectangle3_width(rectangle3_widths[610]), .rectangle3_height(rectangle3_heights[610]), .rectangle3_weight(rectangle3_weights[610]), .feature_threshold(feature_thresholds[610]), .feature_above(feature_aboves[610]), .feature_below(feature_belows[610]), .scan_win_std_dev(scan_win_std_dev[610]), .feature_accum(feature_accums[610]));
  accum_calculator ac611(.scan_win(scan_win611), .rectangle1_x(rectangle1_xs[611]), .rectangle1_y(rectangle1_ys[611]), .rectangle1_width(rectangle1_widths[611]), .rectangle1_height(rectangle1_heights[611]), .rectangle1_weight(rectangle1_weights[611]), .rectangle2_x(rectangle2_xs[611]), .rectangle2_y(rectangle2_ys[611]), .rectangle2_width(rectangle2_widths[611]), .rectangle2_height(rectangle2_heights[611]), .rectangle2_weight(rectangle2_weights[611]), .rectangle3_x(rectangle3_xs[611]), .rectangle3_y(rectangle3_ys[611]), .rectangle3_width(rectangle3_widths[611]), .rectangle3_height(rectangle3_heights[611]), .rectangle3_weight(rectangle3_weights[611]), .feature_threshold(feature_thresholds[611]), .feature_above(feature_aboves[611]), .feature_below(feature_belows[611]), .scan_win_std_dev(scan_win_std_dev[611]), .feature_accum(feature_accums[611]));
  accum_calculator ac612(.scan_win(scan_win612), .rectangle1_x(rectangle1_xs[612]), .rectangle1_y(rectangle1_ys[612]), .rectangle1_width(rectangle1_widths[612]), .rectangle1_height(rectangle1_heights[612]), .rectangle1_weight(rectangle1_weights[612]), .rectangle2_x(rectangle2_xs[612]), .rectangle2_y(rectangle2_ys[612]), .rectangle2_width(rectangle2_widths[612]), .rectangle2_height(rectangle2_heights[612]), .rectangle2_weight(rectangle2_weights[612]), .rectangle3_x(rectangle3_xs[612]), .rectangle3_y(rectangle3_ys[612]), .rectangle3_width(rectangle3_widths[612]), .rectangle3_height(rectangle3_heights[612]), .rectangle3_weight(rectangle3_weights[612]), .feature_threshold(feature_thresholds[612]), .feature_above(feature_aboves[612]), .feature_below(feature_belows[612]), .scan_win_std_dev(scan_win_std_dev[612]), .feature_accum(feature_accums[612]));
  accum_calculator ac613(.scan_win(scan_win613), .rectangle1_x(rectangle1_xs[613]), .rectangle1_y(rectangle1_ys[613]), .rectangle1_width(rectangle1_widths[613]), .rectangle1_height(rectangle1_heights[613]), .rectangle1_weight(rectangle1_weights[613]), .rectangle2_x(rectangle2_xs[613]), .rectangle2_y(rectangle2_ys[613]), .rectangle2_width(rectangle2_widths[613]), .rectangle2_height(rectangle2_heights[613]), .rectangle2_weight(rectangle2_weights[613]), .rectangle3_x(rectangle3_xs[613]), .rectangle3_y(rectangle3_ys[613]), .rectangle3_width(rectangle3_widths[613]), .rectangle3_height(rectangle3_heights[613]), .rectangle3_weight(rectangle3_weights[613]), .feature_threshold(feature_thresholds[613]), .feature_above(feature_aboves[613]), .feature_below(feature_belows[613]), .scan_win_std_dev(scan_win_std_dev[613]), .feature_accum(feature_accums[613]));
  accum_calculator ac614(.scan_win(scan_win614), .rectangle1_x(rectangle1_xs[614]), .rectangle1_y(rectangle1_ys[614]), .rectangle1_width(rectangle1_widths[614]), .rectangle1_height(rectangle1_heights[614]), .rectangle1_weight(rectangle1_weights[614]), .rectangle2_x(rectangle2_xs[614]), .rectangle2_y(rectangle2_ys[614]), .rectangle2_width(rectangle2_widths[614]), .rectangle2_height(rectangle2_heights[614]), .rectangle2_weight(rectangle2_weights[614]), .rectangle3_x(rectangle3_xs[614]), .rectangle3_y(rectangle3_ys[614]), .rectangle3_width(rectangle3_widths[614]), .rectangle3_height(rectangle3_heights[614]), .rectangle3_weight(rectangle3_weights[614]), .feature_threshold(feature_thresholds[614]), .feature_above(feature_aboves[614]), .feature_below(feature_belows[614]), .scan_win_std_dev(scan_win_std_dev[614]), .feature_accum(feature_accums[614]));
  accum_calculator ac615(.scan_win(scan_win615), .rectangle1_x(rectangle1_xs[615]), .rectangle1_y(rectangle1_ys[615]), .rectangle1_width(rectangle1_widths[615]), .rectangle1_height(rectangle1_heights[615]), .rectangle1_weight(rectangle1_weights[615]), .rectangle2_x(rectangle2_xs[615]), .rectangle2_y(rectangle2_ys[615]), .rectangle2_width(rectangle2_widths[615]), .rectangle2_height(rectangle2_heights[615]), .rectangle2_weight(rectangle2_weights[615]), .rectangle3_x(rectangle3_xs[615]), .rectangle3_y(rectangle3_ys[615]), .rectangle3_width(rectangle3_widths[615]), .rectangle3_height(rectangle3_heights[615]), .rectangle3_weight(rectangle3_weights[615]), .feature_threshold(feature_thresholds[615]), .feature_above(feature_aboves[615]), .feature_below(feature_belows[615]), .scan_win_std_dev(scan_win_std_dev[615]), .feature_accum(feature_accums[615]));
  accum_calculator ac616(.scan_win(scan_win616), .rectangle1_x(rectangle1_xs[616]), .rectangle1_y(rectangle1_ys[616]), .rectangle1_width(rectangle1_widths[616]), .rectangle1_height(rectangle1_heights[616]), .rectangle1_weight(rectangle1_weights[616]), .rectangle2_x(rectangle2_xs[616]), .rectangle2_y(rectangle2_ys[616]), .rectangle2_width(rectangle2_widths[616]), .rectangle2_height(rectangle2_heights[616]), .rectangle2_weight(rectangle2_weights[616]), .rectangle3_x(rectangle3_xs[616]), .rectangle3_y(rectangle3_ys[616]), .rectangle3_width(rectangle3_widths[616]), .rectangle3_height(rectangle3_heights[616]), .rectangle3_weight(rectangle3_weights[616]), .feature_threshold(feature_thresholds[616]), .feature_above(feature_aboves[616]), .feature_below(feature_belows[616]), .scan_win_std_dev(scan_win_std_dev[616]), .feature_accum(feature_accums[616]));
  accum_calculator ac617(.scan_win(scan_win617), .rectangle1_x(rectangle1_xs[617]), .rectangle1_y(rectangle1_ys[617]), .rectangle1_width(rectangle1_widths[617]), .rectangle1_height(rectangle1_heights[617]), .rectangle1_weight(rectangle1_weights[617]), .rectangle2_x(rectangle2_xs[617]), .rectangle2_y(rectangle2_ys[617]), .rectangle2_width(rectangle2_widths[617]), .rectangle2_height(rectangle2_heights[617]), .rectangle2_weight(rectangle2_weights[617]), .rectangle3_x(rectangle3_xs[617]), .rectangle3_y(rectangle3_ys[617]), .rectangle3_width(rectangle3_widths[617]), .rectangle3_height(rectangle3_heights[617]), .rectangle3_weight(rectangle3_weights[617]), .feature_threshold(feature_thresholds[617]), .feature_above(feature_aboves[617]), .feature_below(feature_belows[617]), .scan_win_std_dev(scan_win_std_dev[617]), .feature_accum(feature_accums[617]));
  accum_calculator ac618(.scan_win(scan_win618), .rectangle1_x(rectangle1_xs[618]), .rectangle1_y(rectangle1_ys[618]), .rectangle1_width(rectangle1_widths[618]), .rectangle1_height(rectangle1_heights[618]), .rectangle1_weight(rectangle1_weights[618]), .rectangle2_x(rectangle2_xs[618]), .rectangle2_y(rectangle2_ys[618]), .rectangle2_width(rectangle2_widths[618]), .rectangle2_height(rectangle2_heights[618]), .rectangle2_weight(rectangle2_weights[618]), .rectangle3_x(rectangle3_xs[618]), .rectangle3_y(rectangle3_ys[618]), .rectangle3_width(rectangle3_widths[618]), .rectangle3_height(rectangle3_heights[618]), .rectangle3_weight(rectangle3_weights[618]), .feature_threshold(feature_thresholds[618]), .feature_above(feature_aboves[618]), .feature_below(feature_belows[618]), .scan_win_std_dev(scan_win_std_dev[618]), .feature_accum(feature_accums[618]));
  accum_calculator ac619(.scan_win(scan_win619), .rectangle1_x(rectangle1_xs[619]), .rectangle1_y(rectangle1_ys[619]), .rectangle1_width(rectangle1_widths[619]), .rectangle1_height(rectangle1_heights[619]), .rectangle1_weight(rectangle1_weights[619]), .rectangle2_x(rectangle2_xs[619]), .rectangle2_y(rectangle2_ys[619]), .rectangle2_width(rectangle2_widths[619]), .rectangle2_height(rectangle2_heights[619]), .rectangle2_weight(rectangle2_weights[619]), .rectangle3_x(rectangle3_xs[619]), .rectangle3_y(rectangle3_ys[619]), .rectangle3_width(rectangle3_widths[619]), .rectangle3_height(rectangle3_heights[619]), .rectangle3_weight(rectangle3_weights[619]), .feature_threshold(feature_thresholds[619]), .feature_above(feature_aboves[619]), .feature_below(feature_belows[619]), .scan_win_std_dev(scan_win_std_dev[619]), .feature_accum(feature_accums[619]));
  accum_calculator ac620(.scan_win(scan_win620), .rectangle1_x(rectangle1_xs[620]), .rectangle1_y(rectangle1_ys[620]), .rectangle1_width(rectangle1_widths[620]), .rectangle1_height(rectangle1_heights[620]), .rectangle1_weight(rectangle1_weights[620]), .rectangle2_x(rectangle2_xs[620]), .rectangle2_y(rectangle2_ys[620]), .rectangle2_width(rectangle2_widths[620]), .rectangle2_height(rectangle2_heights[620]), .rectangle2_weight(rectangle2_weights[620]), .rectangle3_x(rectangle3_xs[620]), .rectangle3_y(rectangle3_ys[620]), .rectangle3_width(rectangle3_widths[620]), .rectangle3_height(rectangle3_heights[620]), .rectangle3_weight(rectangle3_weights[620]), .feature_threshold(feature_thresholds[620]), .feature_above(feature_aboves[620]), .feature_below(feature_belows[620]), .scan_win_std_dev(scan_win_std_dev[620]), .feature_accum(feature_accums[620]));
  accum_calculator ac621(.scan_win(scan_win621), .rectangle1_x(rectangle1_xs[621]), .rectangle1_y(rectangle1_ys[621]), .rectangle1_width(rectangle1_widths[621]), .rectangle1_height(rectangle1_heights[621]), .rectangle1_weight(rectangle1_weights[621]), .rectangle2_x(rectangle2_xs[621]), .rectangle2_y(rectangle2_ys[621]), .rectangle2_width(rectangle2_widths[621]), .rectangle2_height(rectangle2_heights[621]), .rectangle2_weight(rectangle2_weights[621]), .rectangle3_x(rectangle3_xs[621]), .rectangle3_y(rectangle3_ys[621]), .rectangle3_width(rectangle3_widths[621]), .rectangle3_height(rectangle3_heights[621]), .rectangle3_weight(rectangle3_weights[621]), .feature_threshold(feature_thresholds[621]), .feature_above(feature_aboves[621]), .feature_below(feature_belows[621]), .scan_win_std_dev(scan_win_std_dev[621]), .feature_accum(feature_accums[621]));
  accum_calculator ac622(.scan_win(scan_win622), .rectangle1_x(rectangle1_xs[622]), .rectangle1_y(rectangle1_ys[622]), .rectangle1_width(rectangle1_widths[622]), .rectangle1_height(rectangle1_heights[622]), .rectangle1_weight(rectangle1_weights[622]), .rectangle2_x(rectangle2_xs[622]), .rectangle2_y(rectangle2_ys[622]), .rectangle2_width(rectangle2_widths[622]), .rectangle2_height(rectangle2_heights[622]), .rectangle2_weight(rectangle2_weights[622]), .rectangle3_x(rectangle3_xs[622]), .rectangle3_y(rectangle3_ys[622]), .rectangle3_width(rectangle3_widths[622]), .rectangle3_height(rectangle3_heights[622]), .rectangle3_weight(rectangle3_weights[622]), .feature_threshold(feature_thresholds[622]), .feature_above(feature_aboves[622]), .feature_below(feature_belows[622]), .scan_win_std_dev(scan_win_std_dev[622]), .feature_accum(feature_accums[622]));
  accum_calculator ac623(.scan_win(scan_win623), .rectangle1_x(rectangle1_xs[623]), .rectangle1_y(rectangle1_ys[623]), .rectangle1_width(rectangle1_widths[623]), .rectangle1_height(rectangle1_heights[623]), .rectangle1_weight(rectangle1_weights[623]), .rectangle2_x(rectangle2_xs[623]), .rectangle2_y(rectangle2_ys[623]), .rectangle2_width(rectangle2_widths[623]), .rectangle2_height(rectangle2_heights[623]), .rectangle2_weight(rectangle2_weights[623]), .rectangle3_x(rectangle3_xs[623]), .rectangle3_y(rectangle3_ys[623]), .rectangle3_width(rectangle3_widths[623]), .rectangle3_height(rectangle3_heights[623]), .rectangle3_weight(rectangle3_weights[623]), .feature_threshold(feature_thresholds[623]), .feature_above(feature_aboves[623]), .feature_below(feature_belows[623]), .scan_win_std_dev(scan_win_std_dev[623]), .feature_accum(feature_accums[623]));
  accum_calculator ac624(.scan_win(scan_win624), .rectangle1_x(rectangle1_xs[624]), .rectangle1_y(rectangle1_ys[624]), .rectangle1_width(rectangle1_widths[624]), .rectangle1_height(rectangle1_heights[624]), .rectangle1_weight(rectangle1_weights[624]), .rectangle2_x(rectangle2_xs[624]), .rectangle2_y(rectangle2_ys[624]), .rectangle2_width(rectangle2_widths[624]), .rectangle2_height(rectangle2_heights[624]), .rectangle2_weight(rectangle2_weights[624]), .rectangle3_x(rectangle3_xs[624]), .rectangle3_y(rectangle3_ys[624]), .rectangle3_width(rectangle3_widths[624]), .rectangle3_height(rectangle3_heights[624]), .rectangle3_weight(rectangle3_weights[624]), .feature_threshold(feature_thresholds[624]), .feature_above(feature_aboves[624]), .feature_below(feature_belows[624]), .scan_win_std_dev(scan_win_std_dev[624]), .feature_accum(feature_accums[624]));
  accum_calculator ac625(.scan_win(scan_win625), .rectangle1_x(rectangle1_xs[625]), .rectangle1_y(rectangle1_ys[625]), .rectangle1_width(rectangle1_widths[625]), .rectangle1_height(rectangle1_heights[625]), .rectangle1_weight(rectangle1_weights[625]), .rectangle2_x(rectangle2_xs[625]), .rectangle2_y(rectangle2_ys[625]), .rectangle2_width(rectangle2_widths[625]), .rectangle2_height(rectangle2_heights[625]), .rectangle2_weight(rectangle2_weights[625]), .rectangle3_x(rectangle3_xs[625]), .rectangle3_y(rectangle3_ys[625]), .rectangle3_width(rectangle3_widths[625]), .rectangle3_height(rectangle3_heights[625]), .rectangle3_weight(rectangle3_weights[625]), .feature_threshold(feature_thresholds[625]), .feature_above(feature_aboves[625]), .feature_below(feature_belows[625]), .scan_win_std_dev(scan_win_std_dev[625]), .feature_accum(feature_accums[625]));
  accum_calculator ac626(.scan_win(scan_win626), .rectangle1_x(rectangle1_xs[626]), .rectangle1_y(rectangle1_ys[626]), .rectangle1_width(rectangle1_widths[626]), .rectangle1_height(rectangle1_heights[626]), .rectangle1_weight(rectangle1_weights[626]), .rectangle2_x(rectangle2_xs[626]), .rectangle2_y(rectangle2_ys[626]), .rectangle2_width(rectangle2_widths[626]), .rectangle2_height(rectangle2_heights[626]), .rectangle2_weight(rectangle2_weights[626]), .rectangle3_x(rectangle3_xs[626]), .rectangle3_y(rectangle3_ys[626]), .rectangle3_width(rectangle3_widths[626]), .rectangle3_height(rectangle3_heights[626]), .rectangle3_weight(rectangle3_weights[626]), .feature_threshold(feature_thresholds[626]), .feature_above(feature_aboves[626]), .feature_below(feature_belows[626]), .scan_win_std_dev(scan_win_std_dev[626]), .feature_accum(feature_accums[626]));
  accum_calculator ac627(.scan_win(scan_win627), .rectangle1_x(rectangle1_xs[627]), .rectangle1_y(rectangle1_ys[627]), .rectangle1_width(rectangle1_widths[627]), .rectangle1_height(rectangle1_heights[627]), .rectangle1_weight(rectangle1_weights[627]), .rectangle2_x(rectangle2_xs[627]), .rectangle2_y(rectangle2_ys[627]), .rectangle2_width(rectangle2_widths[627]), .rectangle2_height(rectangle2_heights[627]), .rectangle2_weight(rectangle2_weights[627]), .rectangle3_x(rectangle3_xs[627]), .rectangle3_y(rectangle3_ys[627]), .rectangle3_width(rectangle3_widths[627]), .rectangle3_height(rectangle3_heights[627]), .rectangle3_weight(rectangle3_weights[627]), .feature_threshold(feature_thresholds[627]), .feature_above(feature_aboves[627]), .feature_below(feature_belows[627]), .scan_win_std_dev(scan_win_std_dev[627]), .feature_accum(feature_accums[627]));
  accum_calculator ac628(.scan_win(scan_win628), .rectangle1_x(rectangle1_xs[628]), .rectangle1_y(rectangle1_ys[628]), .rectangle1_width(rectangle1_widths[628]), .rectangle1_height(rectangle1_heights[628]), .rectangle1_weight(rectangle1_weights[628]), .rectangle2_x(rectangle2_xs[628]), .rectangle2_y(rectangle2_ys[628]), .rectangle2_width(rectangle2_widths[628]), .rectangle2_height(rectangle2_heights[628]), .rectangle2_weight(rectangle2_weights[628]), .rectangle3_x(rectangle3_xs[628]), .rectangle3_y(rectangle3_ys[628]), .rectangle3_width(rectangle3_widths[628]), .rectangle3_height(rectangle3_heights[628]), .rectangle3_weight(rectangle3_weights[628]), .feature_threshold(feature_thresholds[628]), .feature_above(feature_aboves[628]), .feature_below(feature_belows[628]), .scan_win_std_dev(scan_win_std_dev[628]), .feature_accum(feature_accums[628]));
  accum_calculator ac629(.scan_win(scan_win629), .rectangle1_x(rectangle1_xs[629]), .rectangle1_y(rectangle1_ys[629]), .rectangle1_width(rectangle1_widths[629]), .rectangle1_height(rectangle1_heights[629]), .rectangle1_weight(rectangle1_weights[629]), .rectangle2_x(rectangle2_xs[629]), .rectangle2_y(rectangle2_ys[629]), .rectangle2_width(rectangle2_widths[629]), .rectangle2_height(rectangle2_heights[629]), .rectangle2_weight(rectangle2_weights[629]), .rectangle3_x(rectangle3_xs[629]), .rectangle3_y(rectangle3_ys[629]), .rectangle3_width(rectangle3_widths[629]), .rectangle3_height(rectangle3_heights[629]), .rectangle3_weight(rectangle3_weights[629]), .feature_threshold(feature_thresholds[629]), .feature_above(feature_aboves[629]), .feature_below(feature_belows[629]), .scan_win_std_dev(scan_win_std_dev[629]), .feature_accum(feature_accums[629]));
  accum_calculator ac630(.scan_win(scan_win630), .rectangle1_x(rectangle1_xs[630]), .rectangle1_y(rectangle1_ys[630]), .rectangle1_width(rectangle1_widths[630]), .rectangle1_height(rectangle1_heights[630]), .rectangle1_weight(rectangle1_weights[630]), .rectangle2_x(rectangle2_xs[630]), .rectangle2_y(rectangle2_ys[630]), .rectangle2_width(rectangle2_widths[630]), .rectangle2_height(rectangle2_heights[630]), .rectangle2_weight(rectangle2_weights[630]), .rectangle3_x(rectangle3_xs[630]), .rectangle3_y(rectangle3_ys[630]), .rectangle3_width(rectangle3_widths[630]), .rectangle3_height(rectangle3_heights[630]), .rectangle3_weight(rectangle3_weights[630]), .feature_threshold(feature_thresholds[630]), .feature_above(feature_aboves[630]), .feature_below(feature_belows[630]), .scan_win_std_dev(scan_win_std_dev[630]), .feature_accum(feature_accums[630]));
  accum_calculator ac631(.scan_win(scan_win631), .rectangle1_x(rectangle1_xs[631]), .rectangle1_y(rectangle1_ys[631]), .rectangle1_width(rectangle1_widths[631]), .rectangle1_height(rectangle1_heights[631]), .rectangle1_weight(rectangle1_weights[631]), .rectangle2_x(rectangle2_xs[631]), .rectangle2_y(rectangle2_ys[631]), .rectangle2_width(rectangle2_widths[631]), .rectangle2_height(rectangle2_heights[631]), .rectangle2_weight(rectangle2_weights[631]), .rectangle3_x(rectangle3_xs[631]), .rectangle3_y(rectangle3_ys[631]), .rectangle3_width(rectangle3_widths[631]), .rectangle3_height(rectangle3_heights[631]), .rectangle3_weight(rectangle3_weights[631]), .feature_threshold(feature_thresholds[631]), .feature_above(feature_aboves[631]), .feature_below(feature_belows[631]), .scan_win_std_dev(scan_win_std_dev[631]), .feature_accum(feature_accums[631]));
  accum_calculator ac632(.scan_win(scan_win632), .rectangle1_x(rectangle1_xs[632]), .rectangle1_y(rectangle1_ys[632]), .rectangle1_width(rectangle1_widths[632]), .rectangle1_height(rectangle1_heights[632]), .rectangle1_weight(rectangle1_weights[632]), .rectangle2_x(rectangle2_xs[632]), .rectangle2_y(rectangle2_ys[632]), .rectangle2_width(rectangle2_widths[632]), .rectangle2_height(rectangle2_heights[632]), .rectangle2_weight(rectangle2_weights[632]), .rectangle3_x(rectangle3_xs[632]), .rectangle3_y(rectangle3_ys[632]), .rectangle3_width(rectangle3_widths[632]), .rectangle3_height(rectangle3_heights[632]), .rectangle3_weight(rectangle3_weights[632]), .feature_threshold(feature_thresholds[632]), .feature_above(feature_aboves[632]), .feature_below(feature_belows[632]), .scan_win_std_dev(scan_win_std_dev[632]), .feature_accum(feature_accums[632]));
  accum_calculator ac633(.scan_win(scan_win633), .rectangle1_x(rectangle1_xs[633]), .rectangle1_y(rectangle1_ys[633]), .rectangle1_width(rectangle1_widths[633]), .rectangle1_height(rectangle1_heights[633]), .rectangle1_weight(rectangle1_weights[633]), .rectangle2_x(rectangle2_xs[633]), .rectangle2_y(rectangle2_ys[633]), .rectangle2_width(rectangle2_widths[633]), .rectangle2_height(rectangle2_heights[633]), .rectangle2_weight(rectangle2_weights[633]), .rectangle3_x(rectangle3_xs[633]), .rectangle3_y(rectangle3_ys[633]), .rectangle3_width(rectangle3_widths[633]), .rectangle3_height(rectangle3_heights[633]), .rectangle3_weight(rectangle3_weights[633]), .feature_threshold(feature_thresholds[633]), .feature_above(feature_aboves[633]), .feature_below(feature_belows[633]), .scan_win_std_dev(scan_win_std_dev[633]), .feature_accum(feature_accums[633]));
  accum_calculator ac634(.scan_win(scan_win634), .rectangle1_x(rectangle1_xs[634]), .rectangle1_y(rectangle1_ys[634]), .rectangle1_width(rectangle1_widths[634]), .rectangle1_height(rectangle1_heights[634]), .rectangle1_weight(rectangle1_weights[634]), .rectangle2_x(rectangle2_xs[634]), .rectangle2_y(rectangle2_ys[634]), .rectangle2_width(rectangle2_widths[634]), .rectangle2_height(rectangle2_heights[634]), .rectangle2_weight(rectangle2_weights[634]), .rectangle3_x(rectangle3_xs[634]), .rectangle3_y(rectangle3_ys[634]), .rectangle3_width(rectangle3_widths[634]), .rectangle3_height(rectangle3_heights[634]), .rectangle3_weight(rectangle3_weights[634]), .feature_threshold(feature_thresholds[634]), .feature_above(feature_aboves[634]), .feature_below(feature_belows[634]), .scan_win_std_dev(scan_win_std_dev[634]), .feature_accum(feature_accums[634]));
  accum_calculator ac635(.scan_win(scan_win635), .rectangle1_x(rectangle1_xs[635]), .rectangle1_y(rectangle1_ys[635]), .rectangle1_width(rectangle1_widths[635]), .rectangle1_height(rectangle1_heights[635]), .rectangle1_weight(rectangle1_weights[635]), .rectangle2_x(rectangle2_xs[635]), .rectangle2_y(rectangle2_ys[635]), .rectangle2_width(rectangle2_widths[635]), .rectangle2_height(rectangle2_heights[635]), .rectangle2_weight(rectangle2_weights[635]), .rectangle3_x(rectangle3_xs[635]), .rectangle3_y(rectangle3_ys[635]), .rectangle3_width(rectangle3_widths[635]), .rectangle3_height(rectangle3_heights[635]), .rectangle3_weight(rectangle3_weights[635]), .feature_threshold(feature_thresholds[635]), .feature_above(feature_aboves[635]), .feature_below(feature_belows[635]), .scan_win_std_dev(scan_win_std_dev[635]), .feature_accum(feature_accums[635]));
  accum_calculator ac636(.scan_win(scan_win636), .rectangle1_x(rectangle1_xs[636]), .rectangle1_y(rectangle1_ys[636]), .rectangle1_width(rectangle1_widths[636]), .rectangle1_height(rectangle1_heights[636]), .rectangle1_weight(rectangle1_weights[636]), .rectangle2_x(rectangle2_xs[636]), .rectangle2_y(rectangle2_ys[636]), .rectangle2_width(rectangle2_widths[636]), .rectangle2_height(rectangle2_heights[636]), .rectangle2_weight(rectangle2_weights[636]), .rectangle3_x(rectangle3_xs[636]), .rectangle3_y(rectangle3_ys[636]), .rectangle3_width(rectangle3_widths[636]), .rectangle3_height(rectangle3_heights[636]), .rectangle3_weight(rectangle3_weights[636]), .feature_threshold(feature_thresholds[636]), .feature_above(feature_aboves[636]), .feature_below(feature_belows[636]), .scan_win_std_dev(scan_win_std_dev[636]), .feature_accum(feature_accums[636]));
  accum_calculator ac637(.scan_win(scan_win637), .rectangle1_x(rectangle1_xs[637]), .rectangle1_y(rectangle1_ys[637]), .rectangle1_width(rectangle1_widths[637]), .rectangle1_height(rectangle1_heights[637]), .rectangle1_weight(rectangle1_weights[637]), .rectangle2_x(rectangle2_xs[637]), .rectangle2_y(rectangle2_ys[637]), .rectangle2_width(rectangle2_widths[637]), .rectangle2_height(rectangle2_heights[637]), .rectangle2_weight(rectangle2_weights[637]), .rectangle3_x(rectangle3_xs[637]), .rectangle3_y(rectangle3_ys[637]), .rectangle3_width(rectangle3_widths[637]), .rectangle3_height(rectangle3_heights[637]), .rectangle3_weight(rectangle3_weights[637]), .feature_threshold(feature_thresholds[637]), .feature_above(feature_aboves[637]), .feature_below(feature_belows[637]), .scan_win_std_dev(scan_win_std_dev[637]), .feature_accum(feature_accums[637]));
  accum_calculator ac638(.scan_win(scan_win638), .rectangle1_x(rectangle1_xs[638]), .rectangle1_y(rectangle1_ys[638]), .rectangle1_width(rectangle1_widths[638]), .rectangle1_height(rectangle1_heights[638]), .rectangle1_weight(rectangle1_weights[638]), .rectangle2_x(rectangle2_xs[638]), .rectangle2_y(rectangle2_ys[638]), .rectangle2_width(rectangle2_widths[638]), .rectangle2_height(rectangle2_heights[638]), .rectangle2_weight(rectangle2_weights[638]), .rectangle3_x(rectangle3_xs[638]), .rectangle3_y(rectangle3_ys[638]), .rectangle3_width(rectangle3_widths[638]), .rectangle3_height(rectangle3_heights[638]), .rectangle3_weight(rectangle3_weights[638]), .feature_threshold(feature_thresholds[638]), .feature_above(feature_aboves[638]), .feature_below(feature_belows[638]), .scan_win_std_dev(scan_win_std_dev[638]), .feature_accum(feature_accums[638]));
  accum_calculator ac639(.scan_win(scan_win639), .rectangle1_x(rectangle1_xs[639]), .rectangle1_y(rectangle1_ys[639]), .rectangle1_width(rectangle1_widths[639]), .rectangle1_height(rectangle1_heights[639]), .rectangle1_weight(rectangle1_weights[639]), .rectangle2_x(rectangle2_xs[639]), .rectangle2_y(rectangle2_ys[639]), .rectangle2_width(rectangle2_widths[639]), .rectangle2_height(rectangle2_heights[639]), .rectangle2_weight(rectangle2_weights[639]), .rectangle3_x(rectangle3_xs[639]), .rectangle3_y(rectangle3_ys[639]), .rectangle3_width(rectangle3_widths[639]), .rectangle3_height(rectangle3_heights[639]), .rectangle3_weight(rectangle3_weights[639]), .feature_threshold(feature_thresholds[639]), .feature_above(feature_aboves[639]), .feature_below(feature_belows[639]), .scan_win_std_dev(scan_win_std_dev[639]), .feature_accum(feature_accums[639]));
  accum_calculator ac640(.scan_win(scan_win640), .rectangle1_x(rectangle1_xs[640]), .rectangle1_y(rectangle1_ys[640]), .rectangle1_width(rectangle1_widths[640]), .rectangle1_height(rectangle1_heights[640]), .rectangle1_weight(rectangle1_weights[640]), .rectangle2_x(rectangle2_xs[640]), .rectangle2_y(rectangle2_ys[640]), .rectangle2_width(rectangle2_widths[640]), .rectangle2_height(rectangle2_heights[640]), .rectangle2_weight(rectangle2_weights[640]), .rectangle3_x(rectangle3_xs[640]), .rectangle3_y(rectangle3_ys[640]), .rectangle3_width(rectangle3_widths[640]), .rectangle3_height(rectangle3_heights[640]), .rectangle3_weight(rectangle3_weights[640]), .feature_threshold(feature_thresholds[640]), .feature_above(feature_aboves[640]), .feature_below(feature_belows[640]), .scan_win_std_dev(scan_win_std_dev[640]), .feature_accum(feature_accums[640]));
  accum_calculator ac641(.scan_win(scan_win641), .rectangle1_x(rectangle1_xs[641]), .rectangle1_y(rectangle1_ys[641]), .rectangle1_width(rectangle1_widths[641]), .rectangle1_height(rectangle1_heights[641]), .rectangle1_weight(rectangle1_weights[641]), .rectangle2_x(rectangle2_xs[641]), .rectangle2_y(rectangle2_ys[641]), .rectangle2_width(rectangle2_widths[641]), .rectangle2_height(rectangle2_heights[641]), .rectangle2_weight(rectangle2_weights[641]), .rectangle3_x(rectangle3_xs[641]), .rectangle3_y(rectangle3_ys[641]), .rectangle3_width(rectangle3_widths[641]), .rectangle3_height(rectangle3_heights[641]), .rectangle3_weight(rectangle3_weights[641]), .feature_threshold(feature_thresholds[641]), .feature_above(feature_aboves[641]), .feature_below(feature_belows[641]), .scan_win_std_dev(scan_win_std_dev[641]), .feature_accum(feature_accums[641]));
  accum_calculator ac642(.scan_win(scan_win642), .rectangle1_x(rectangle1_xs[642]), .rectangle1_y(rectangle1_ys[642]), .rectangle1_width(rectangle1_widths[642]), .rectangle1_height(rectangle1_heights[642]), .rectangle1_weight(rectangle1_weights[642]), .rectangle2_x(rectangle2_xs[642]), .rectangle2_y(rectangle2_ys[642]), .rectangle2_width(rectangle2_widths[642]), .rectangle2_height(rectangle2_heights[642]), .rectangle2_weight(rectangle2_weights[642]), .rectangle3_x(rectangle3_xs[642]), .rectangle3_y(rectangle3_ys[642]), .rectangle3_width(rectangle3_widths[642]), .rectangle3_height(rectangle3_heights[642]), .rectangle3_weight(rectangle3_weights[642]), .feature_threshold(feature_thresholds[642]), .feature_above(feature_aboves[642]), .feature_below(feature_belows[642]), .scan_win_std_dev(scan_win_std_dev[642]), .feature_accum(feature_accums[642]));
  accum_calculator ac643(.scan_win(scan_win643), .rectangle1_x(rectangle1_xs[643]), .rectangle1_y(rectangle1_ys[643]), .rectangle1_width(rectangle1_widths[643]), .rectangle1_height(rectangle1_heights[643]), .rectangle1_weight(rectangle1_weights[643]), .rectangle2_x(rectangle2_xs[643]), .rectangle2_y(rectangle2_ys[643]), .rectangle2_width(rectangle2_widths[643]), .rectangle2_height(rectangle2_heights[643]), .rectangle2_weight(rectangle2_weights[643]), .rectangle3_x(rectangle3_xs[643]), .rectangle3_y(rectangle3_ys[643]), .rectangle3_width(rectangle3_widths[643]), .rectangle3_height(rectangle3_heights[643]), .rectangle3_weight(rectangle3_weights[643]), .feature_threshold(feature_thresholds[643]), .feature_above(feature_aboves[643]), .feature_below(feature_belows[643]), .scan_win_std_dev(scan_win_std_dev[643]), .feature_accum(feature_accums[643]));
  accum_calculator ac644(.scan_win(scan_win644), .rectangle1_x(rectangle1_xs[644]), .rectangle1_y(rectangle1_ys[644]), .rectangle1_width(rectangle1_widths[644]), .rectangle1_height(rectangle1_heights[644]), .rectangle1_weight(rectangle1_weights[644]), .rectangle2_x(rectangle2_xs[644]), .rectangle2_y(rectangle2_ys[644]), .rectangle2_width(rectangle2_widths[644]), .rectangle2_height(rectangle2_heights[644]), .rectangle2_weight(rectangle2_weights[644]), .rectangle3_x(rectangle3_xs[644]), .rectangle3_y(rectangle3_ys[644]), .rectangle3_width(rectangle3_widths[644]), .rectangle3_height(rectangle3_heights[644]), .rectangle3_weight(rectangle3_weights[644]), .feature_threshold(feature_thresholds[644]), .feature_above(feature_aboves[644]), .feature_below(feature_belows[644]), .scan_win_std_dev(scan_win_std_dev[644]), .feature_accum(feature_accums[644]));
  accum_calculator ac645(.scan_win(scan_win645), .rectangle1_x(rectangle1_xs[645]), .rectangle1_y(rectangle1_ys[645]), .rectangle1_width(rectangle1_widths[645]), .rectangle1_height(rectangle1_heights[645]), .rectangle1_weight(rectangle1_weights[645]), .rectangle2_x(rectangle2_xs[645]), .rectangle2_y(rectangle2_ys[645]), .rectangle2_width(rectangle2_widths[645]), .rectangle2_height(rectangle2_heights[645]), .rectangle2_weight(rectangle2_weights[645]), .rectangle3_x(rectangle3_xs[645]), .rectangle3_y(rectangle3_ys[645]), .rectangle3_width(rectangle3_widths[645]), .rectangle3_height(rectangle3_heights[645]), .rectangle3_weight(rectangle3_weights[645]), .feature_threshold(feature_thresholds[645]), .feature_above(feature_aboves[645]), .feature_below(feature_belows[645]), .scan_win_std_dev(scan_win_std_dev[645]), .feature_accum(feature_accums[645]));
  accum_calculator ac646(.scan_win(scan_win646), .rectangle1_x(rectangle1_xs[646]), .rectangle1_y(rectangle1_ys[646]), .rectangle1_width(rectangle1_widths[646]), .rectangle1_height(rectangle1_heights[646]), .rectangle1_weight(rectangle1_weights[646]), .rectangle2_x(rectangle2_xs[646]), .rectangle2_y(rectangle2_ys[646]), .rectangle2_width(rectangle2_widths[646]), .rectangle2_height(rectangle2_heights[646]), .rectangle2_weight(rectangle2_weights[646]), .rectangle3_x(rectangle3_xs[646]), .rectangle3_y(rectangle3_ys[646]), .rectangle3_width(rectangle3_widths[646]), .rectangle3_height(rectangle3_heights[646]), .rectangle3_weight(rectangle3_weights[646]), .feature_threshold(feature_thresholds[646]), .feature_above(feature_aboves[646]), .feature_below(feature_belows[646]), .scan_win_std_dev(scan_win_std_dev[646]), .feature_accum(feature_accums[646]));
  accum_calculator ac647(.scan_win(scan_win647), .rectangle1_x(rectangle1_xs[647]), .rectangle1_y(rectangle1_ys[647]), .rectangle1_width(rectangle1_widths[647]), .rectangle1_height(rectangle1_heights[647]), .rectangle1_weight(rectangle1_weights[647]), .rectangle2_x(rectangle2_xs[647]), .rectangle2_y(rectangle2_ys[647]), .rectangle2_width(rectangle2_widths[647]), .rectangle2_height(rectangle2_heights[647]), .rectangle2_weight(rectangle2_weights[647]), .rectangle3_x(rectangle3_xs[647]), .rectangle3_y(rectangle3_ys[647]), .rectangle3_width(rectangle3_widths[647]), .rectangle3_height(rectangle3_heights[647]), .rectangle3_weight(rectangle3_weights[647]), .feature_threshold(feature_thresholds[647]), .feature_above(feature_aboves[647]), .feature_below(feature_belows[647]), .scan_win_std_dev(scan_win_std_dev[647]), .feature_accum(feature_accums[647]));
  accum_calculator ac648(.scan_win(scan_win648), .rectangle1_x(rectangle1_xs[648]), .rectangle1_y(rectangle1_ys[648]), .rectangle1_width(rectangle1_widths[648]), .rectangle1_height(rectangle1_heights[648]), .rectangle1_weight(rectangle1_weights[648]), .rectangle2_x(rectangle2_xs[648]), .rectangle2_y(rectangle2_ys[648]), .rectangle2_width(rectangle2_widths[648]), .rectangle2_height(rectangle2_heights[648]), .rectangle2_weight(rectangle2_weights[648]), .rectangle3_x(rectangle3_xs[648]), .rectangle3_y(rectangle3_ys[648]), .rectangle3_width(rectangle3_widths[648]), .rectangle3_height(rectangle3_heights[648]), .rectangle3_weight(rectangle3_weights[648]), .feature_threshold(feature_thresholds[648]), .feature_above(feature_aboves[648]), .feature_below(feature_belows[648]), .scan_win_std_dev(scan_win_std_dev[648]), .feature_accum(feature_accums[648]));
  accum_calculator ac649(.scan_win(scan_win649), .rectangle1_x(rectangle1_xs[649]), .rectangle1_y(rectangle1_ys[649]), .rectangle1_width(rectangle1_widths[649]), .rectangle1_height(rectangle1_heights[649]), .rectangle1_weight(rectangle1_weights[649]), .rectangle2_x(rectangle2_xs[649]), .rectangle2_y(rectangle2_ys[649]), .rectangle2_width(rectangle2_widths[649]), .rectangle2_height(rectangle2_heights[649]), .rectangle2_weight(rectangle2_weights[649]), .rectangle3_x(rectangle3_xs[649]), .rectangle3_y(rectangle3_ys[649]), .rectangle3_width(rectangle3_widths[649]), .rectangle3_height(rectangle3_heights[649]), .rectangle3_weight(rectangle3_weights[649]), .feature_threshold(feature_thresholds[649]), .feature_above(feature_aboves[649]), .feature_below(feature_belows[649]), .scan_win_std_dev(scan_win_std_dev[649]), .feature_accum(feature_accums[649]));
  accum_calculator ac650(.scan_win(scan_win650), .rectangle1_x(rectangle1_xs[650]), .rectangle1_y(rectangle1_ys[650]), .rectangle1_width(rectangle1_widths[650]), .rectangle1_height(rectangle1_heights[650]), .rectangle1_weight(rectangle1_weights[650]), .rectangle2_x(rectangle2_xs[650]), .rectangle2_y(rectangle2_ys[650]), .rectangle2_width(rectangle2_widths[650]), .rectangle2_height(rectangle2_heights[650]), .rectangle2_weight(rectangle2_weights[650]), .rectangle3_x(rectangle3_xs[650]), .rectangle3_y(rectangle3_ys[650]), .rectangle3_width(rectangle3_widths[650]), .rectangle3_height(rectangle3_heights[650]), .rectangle3_weight(rectangle3_weights[650]), .feature_threshold(feature_thresholds[650]), .feature_above(feature_aboves[650]), .feature_below(feature_belows[650]), .scan_win_std_dev(scan_win_std_dev[650]), .feature_accum(feature_accums[650]));
  accum_calculator ac651(.scan_win(scan_win651), .rectangle1_x(rectangle1_xs[651]), .rectangle1_y(rectangle1_ys[651]), .rectangle1_width(rectangle1_widths[651]), .rectangle1_height(rectangle1_heights[651]), .rectangle1_weight(rectangle1_weights[651]), .rectangle2_x(rectangle2_xs[651]), .rectangle2_y(rectangle2_ys[651]), .rectangle2_width(rectangle2_widths[651]), .rectangle2_height(rectangle2_heights[651]), .rectangle2_weight(rectangle2_weights[651]), .rectangle3_x(rectangle3_xs[651]), .rectangle3_y(rectangle3_ys[651]), .rectangle3_width(rectangle3_widths[651]), .rectangle3_height(rectangle3_heights[651]), .rectangle3_weight(rectangle3_weights[651]), .feature_threshold(feature_thresholds[651]), .feature_above(feature_aboves[651]), .feature_below(feature_belows[651]), .scan_win_std_dev(scan_win_std_dev[651]), .feature_accum(feature_accums[651]));
  accum_calculator ac652(.scan_win(scan_win652), .rectangle1_x(rectangle1_xs[652]), .rectangle1_y(rectangle1_ys[652]), .rectangle1_width(rectangle1_widths[652]), .rectangle1_height(rectangle1_heights[652]), .rectangle1_weight(rectangle1_weights[652]), .rectangle2_x(rectangle2_xs[652]), .rectangle2_y(rectangle2_ys[652]), .rectangle2_width(rectangle2_widths[652]), .rectangle2_height(rectangle2_heights[652]), .rectangle2_weight(rectangle2_weights[652]), .rectangle3_x(rectangle3_xs[652]), .rectangle3_y(rectangle3_ys[652]), .rectangle3_width(rectangle3_widths[652]), .rectangle3_height(rectangle3_heights[652]), .rectangle3_weight(rectangle3_weights[652]), .feature_threshold(feature_thresholds[652]), .feature_above(feature_aboves[652]), .feature_below(feature_belows[652]), .scan_win_std_dev(scan_win_std_dev[652]), .feature_accum(feature_accums[652]));
  accum_calculator ac653(.scan_win(scan_win653), .rectangle1_x(rectangle1_xs[653]), .rectangle1_y(rectangle1_ys[653]), .rectangle1_width(rectangle1_widths[653]), .rectangle1_height(rectangle1_heights[653]), .rectangle1_weight(rectangle1_weights[653]), .rectangle2_x(rectangle2_xs[653]), .rectangle2_y(rectangle2_ys[653]), .rectangle2_width(rectangle2_widths[653]), .rectangle2_height(rectangle2_heights[653]), .rectangle2_weight(rectangle2_weights[653]), .rectangle3_x(rectangle3_xs[653]), .rectangle3_y(rectangle3_ys[653]), .rectangle3_width(rectangle3_widths[653]), .rectangle3_height(rectangle3_heights[653]), .rectangle3_weight(rectangle3_weights[653]), .feature_threshold(feature_thresholds[653]), .feature_above(feature_aboves[653]), .feature_below(feature_belows[653]), .scan_win_std_dev(scan_win_std_dev[653]), .feature_accum(feature_accums[653]));
  accum_calculator ac654(.scan_win(scan_win654), .rectangle1_x(rectangle1_xs[654]), .rectangle1_y(rectangle1_ys[654]), .rectangle1_width(rectangle1_widths[654]), .rectangle1_height(rectangle1_heights[654]), .rectangle1_weight(rectangle1_weights[654]), .rectangle2_x(rectangle2_xs[654]), .rectangle2_y(rectangle2_ys[654]), .rectangle2_width(rectangle2_widths[654]), .rectangle2_height(rectangle2_heights[654]), .rectangle2_weight(rectangle2_weights[654]), .rectangle3_x(rectangle3_xs[654]), .rectangle3_y(rectangle3_ys[654]), .rectangle3_width(rectangle3_widths[654]), .rectangle3_height(rectangle3_heights[654]), .rectangle3_weight(rectangle3_weights[654]), .feature_threshold(feature_thresholds[654]), .feature_above(feature_aboves[654]), .feature_below(feature_belows[654]), .scan_win_std_dev(scan_win_std_dev[654]), .feature_accum(feature_accums[654]));
  accum_calculator ac655(.scan_win(scan_win655), .rectangle1_x(rectangle1_xs[655]), .rectangle1_y(rectangle1_ys[655]), .rectangle1_width(rectangle1_widths[655]), .rectangle1_height(rectangle1_heights[655]), .rectangle1_weight(rectangle1_weights[655]), .rectangle2_x(rectangle2_xs[655]), .rectangle2_y(rectangle2_ys[655]), .rectangle2_width(rectangle2_widths[655]), .rectangle2_height(rectangle2_heights[655]), .rectangle2_weight(rectangle2_weights[655]), .rectangle3_x(rectangle3_xs[655]), .rectangle3_y(rectangle3_ys[655]), .rectangle3_width(rectangle3_widths[655]), .rectangle3_height(rectangle3_heights[655]), .rectangle3_weight(rectangle3_weights[655]), .feature_threshold(feature_thresholds[655]), .feature_above(feature_aboves[655]), .feature_below(feature_belows[655]), .scan_win_std_dev(scan_win_std_dev[655]), .feature_accum(feature_accums[655]));
  accum_calculator ac656(.scan_win(scan_win656), .rectangle1_x(rectangle1_xs[656]), .rectangle1_y(rectangle1_ys[656]), .rectangle1_width(rectangle1_widths[656]), .rectangle1_height(rectangle1_heights[656]), .rectangle1_weight(rectangle1_weights[656]), .rectangle2_x(rectangle2_xs[656]), .rectangle2_y(rectangle2_ys[656]), .rectangle2_width(rectangle2_widths[656]), .rectangle2_height(rectangle2_heights[656]), .rectangle2_weight(rectangle2_weights[656]), .rectangle3_x(rectangle3_xs[656]), .rectangle3_y(rectangle3_ys[656]), .rectangle3_width(rectangle3_widths[656]), .rectangle3_height(rectangle3_heights[656]), .rectangle3_weight(rectangle3_weights[656]), .feature_threshold(feature_thresholds[656]), .feature_above(feature_aboves[656]), .feature_below(feature_belows[656]), .scan_win_std_dev(scan_win_std_dev[656]), .feature_accum(feature_accums[656]));
  accum_calculator ac657(.scan_win(scan_win657), .rectangle1_x(rectangle1_xs[657]), .rectangle1_y(rectangle1_ys[657]), .rectangle1_width(rectangle1_widths[657]), .rectangle1_height(rectangle1_heights[657]), .rectangle1_weight(rectangle1_weights[657]), .rectangle2_x(rectangle2_xs[657]), .rectangle2_y(rectangle2_ys[657]), .rectangle2_width(rectangle2_widths[657]), .rectangle2_height(rectangle2_heights[657]), .rectangle2_weight(rectangle2_weights[657]), .rectangle3_x(rectangle3_xs[657]), .rectangle3_y(rectangle3_ys[657]), .rectangle3_width(rectangle3_widths[657]), .rectangle3_height(rectangle3_heights[657]), .rectangle3_weight(rectangle3_weights[657]), .feature_threshold(feature_thresholds[657]), .feature_above(feature_aboves[657]), .feature_below(feature_belows[657]), .scan_win_std_dev(scan_win_std_dev[657]), .feature_accum(feature_accums[657]));
  accum_calculator ac658(.scan_win(scan_win658), .rectangle1_x(rectangle1_xs[658]), .rectangle1_y(rectangle1_ys[658]), .rectangle1_width(rectangle1_widths[658]), .rectangle1_height(rectangle1_heights[658]), .rectangle1_weight(rectangle1_weights[658]), .rectangle2_x(rectangle2_xs[658]), .rectangle2_y(rectangle2_ys[658]), .rectangle2_width(rectangle2_widths[658]), .rectangle2_height(rectangle2_heights[658]), .rectangle2_weight(rectangle2_weights[658]), .rectangle3_x(rectangle3_xs[658]), .rectangle3_y(rectangle3_ys[658]), .rectangle3_width(rectangle3_widths[658]), .rectangle3_height(rectangle3_heights[658]), .rectangle3_weight(rectangle3_weights[658]), .feature_threshold(feature_thresholds[658]), .feature_above(feature_aboves[658]), .feature_below(feature_belows[658]), .scan_win_std_dev(scan_win_std_dev[658]), .feature_accum(feature_accums[658]));
  accum_calculator ac659(.scan_win(scan_win659), .rectangle1_x(rectangle1_xs[659]), .rectangle1_y(rectangle1_ys[659]), .rectangle1_width(rectangle1_widths[659]), .rectangle1_height(rectangle1_heights[659]), .rectangle1_weight(rectangle1_weights[659]), .rectangle2_x(rectangle2_xs[659]), .rectangle2_y(rectangle2_ys[659]), .rectangle2_width(rectangle2_widths[659]), .rectangle2_height(rectangle2_heights[659]), .rectangle2_weight(rectangle2_weights[659]), .rectangle3_x(rectangle3_xs[659]), .rectangle3_y(rectangle3_ys[659]), .rectangle3_width(rectangle3_widths[659]), .rectangle3_height(rectangle3_heights[659]), .rectangle3_weight(rectangle3_weights[659]), .feature_threshold(feature_thresholds[659]), .feature_above(feature_aboves[659]), .feature_below(feature_belows[659]), .scan_win_std_dev(scan_win_std_dev[659]), .feature_accum(feature_accums[659]));
  accum_calculator ac660(.scan_win(scan_win660), .rectangle1_x(rectangle1_xs[660]), .rectangle1_y(rectangle1_ys[660]), .rectangle1_width(rectangle1_widths[660]), .rectangle1_height(rectangle1_heights[660]), .rectangle1_weight(rectangle1_weights[660]), .rectangle2_x(rectangle2_xs[660]), .rectangle2_y(rectangle2_ys[660]), .rectangle2_width(rectangle2_widths[660]), .rectangle2_height(rectangle2_heights[660]), .rectangle2_weight(rectangle2_weights[660]), .rectangle3_x(rectangle3_xs[660]), .rectangle3_y(rectangle3_ys[660]), .rectangle3_width(rectangle3_widths[660]), .rectangle3_height(rectangle3_heights[660]), .rectangle3_weight(rectangle3_weights[660]), .feature_threshold(feature_thresholds[660]), .feature_above(feature_aboves[660]), .feature_below(feature_belows[660]), .scan_win_std_dev(scan_win_std_dev[660]), .feature_accum(feature_accums[660]));
  accum_calculator ac661(.scan_win(scan_win661), .rectangle1_x(rectangle1_xs[661]), .rectangle1_y(rectangle1_ys[661]), .rectangle1_width(rectangle1_widths[661]), .rectangle1_height(rectangle1_heights[661]), .rectangle1_weight(rectangle1_weights[661]), .rectangle2_x(rectangle2_xs[661]), .rectangle2_y(rectangle2_ys[661]), .rectangle2_width(rectangle2_widths[661]), .rectangle2_height(rectangle2_heights[661]), .rectangle2_weight(rectangle2_weights[661]), .rectangle3_x(rectangle3_xs[661]), .rectangle3_y(rectangle3_ys[661]), .rectangle3_width(rectangle3_widths[661]), .rectangle3_height(rectangle3_heights[661]), .rectangle3_weight(rectangle3_weights[661]), .feature_threshold(feature_thresholds[661]), .feature_above(feature_aboves[661]), .feature_below(feature_belows[661]), .scan_win_std_dev(scan_win_std_dev[661]), .feature_accum(feature_accums[661]));
  accum_calculator ac662(.scan_win(scan_win662), .rectangle1_x(rectangle1_xs[662]), .rectangle1_y(rectangle1_ys[662]), .rectangle1_width(rectangle1_widths[662]), .rectangle1_height(rectangle1_heights[662]), .rectangle1_weight(rectangle1_weights[662]), .rectangle2_x(rectangle2_xs[662]), .rectangle2_y(rectangle2_ys[662]), .rectangle2_width(rectangle2_widths[662]), .rectangle2_height(rectangle2_heights[662]), .rectangle2_weight(rectangle2_weights[662]), .rectangle3_x(rectangle3_xs[662]), .rectangle3_y(rectangle3_ys[662]), .rectangle3_width(rectangle3_widths[662]), .rectangle3_height(rectangle3_heights[662]), .rectangle3_weight(rectangle3_weights[662]), .feature_threshold(feature_thresholds[662]), .feature_above(feature_aboves[662]), .feature_below(feature_belows[662]), .scan_win_std_dev(scan_win_std_dev[662]), .feature_accum(feature_accums[662]));
  accum_calculator ac663(.scan_win(scan_win663), .rectangle1_x(rectangle1_xs[663]), .rectangle1_y(rectangle1_ys[663]), .rectangle1_width(rectangle1_widths[663]), .rectangle1_height(rectangle1_heights[663]), .rectangle1_weight(rectangle1_weights[663]), .rectangle2_x(rectangle2_xs[663]), .rectangle2_y(rectangle2_ys[663]), .rectangle2_width(rectangle2_widths[663]), .rectangle2_height(rectangle2_heights[663]), .rectangle2_weight(rectangle2_weights[663]), .rectangle3_x(rectangle3_xs[663]), .rectangle3_y(rectangle3_ys[663]), .rectangle3_width(rectangle3_widths[663]), .rectangle3_height(rectangle3_heights[663]), .rectangle3_weight(rectangle3_weights[663]), .feature_threshold(feature_thresholds[663]), .feature_above(feature_aboves[663]), .feature_below(feature_belows[663]), .scan_win_std_dev(scan_win_std_dev[663]), .feature_accum(feature_accums[663]));
  accum_calculator ac664(.scan_win(scan_win664), .rectangle1_x(rectangle1_xs[664]), .rectangle1_y(rectangle1_ys[664]), .rectangle1_width(rectangle1_widths[664]), .rectangle1_height(rectangle1_heights[664]), .rectangle1_weight(rectangle1_weights[664]), .rectangle2_x(rectangle2_xs[664]), .rectangle2_y(rectangle2_ys[664]), .rectangle2_width(rectangle2_widths[664]), .rectangle2_height(rectangle2_heights[664]), .rectangle2_weight(rectangle2_weights[664]), .rectangle3_x(rectangle3_xs[664]), .rectangle3_y(rectangle3_ys[664]), .rectangle3_width(rectangle3_widths[664]), .rectangle3_height(rectangle3_heights[664]), .rectangle3_weight(rectangle3_weights[664]), .feature_threshold(feature_thresholds[664]), .feature_above(feature_aboves[664]), .feature_below(feature_belows[664]), .scan_win_std_dev(scan_win_std_dev[664]), .feature_accum(feature_accums[664]));
  accum_calculator ac665(.scan_win(scan_win665), .rectangle1_x(rectangle1_xs[665]), .rectangle1_y(rectangle1_ys[665]), .rectangle1_width(rectangle1_widths[665]), .rectangle1_height(rectangle1_heights[665]), .rectangle1_weight(rectangle1_weights[665]), .rectangle2_x(rectangle2_xs[665]), .rectangle2_y(rectangle2_ys[665]), .rectangle2_width(rectangle2_widths[665]), .rectangle2_height(rectangle2_heights[665]), .rectangle2_weight(rectangle2_weights[665]), .rectangle3_x(rectangle3_xs[665]), .rectangle3_y(rectangle3_ys[665]), .rectangle3_width(rectangle3_widths[665]), .rectangle3_height(rectangle3_heights[665]), .rectangle3_weight(rectangle3_weights[665]), .feature_threshold(feature_thresholds[665]), .feature_above(feature_aboves[665]), .feature_below(feature_belows[665]), .scan_win_std_dev(scan_win_std_dev[665]), .feature_accum(feature_accums[665]));
  accum_calculator ac666(.scan_win(scan_win666), .rectangle1_x(rectangle1_xs[666]), .rectangle1_y(rectangle1_ys[666]), .rectangle1_width(rectangle1_widths[666]), .rectangle1_height(rectangle1_heights[666]), .rectangle1_weight(rectangle1_weights[666]), .rectangle2_x(rectangle2_xs[666]), .rectangle2_y(rectangle2_ys[666]), .rectangle2_width(rectangle2_widths[666]), .rectangle2_height(rectangle2_heights[666]), .rectangle2_weight(rectangle2_weights[666]), .rectangle3_x(rectangle3_xs[666]), .rectangle3_y(rectangle3_ys[666]), .rectangle3_width(rectangle3_widths[666]), .rectangle3_height(rectangle3_heights[666]), .rectangle3_weight(rectangle3_weights[666]), .feature_threshold(feature_thresholds[666]), .feature_above(feature_aboves[666]), .feature_below(feature_belows[666]), .scan_win_std_dev(scan_win_std_dev[666]), .feature_accum(feature_accums[666]));
  accum_calculator ac667(.scan_win(scan_win667), .rectangle1_x(rectangle1_xs[667]), .rectangle1_y(rectangle1_ys[667]), .rectangle1_width(rectangle1_widths[667]), .rectangle1_height(rectangle1_heights[667]), .rectangle1_weight(rectangle1_weights[667]), .rectangle2_x(rectangle2_xs[667]), .rectangle2_y(rectangle2_ys[667]), .rectangle2_width(rectangle2_widths[667]), .rectangle2_height(rectangle2_heights[667]), .rectangle2_weight(rectangle2_weights[667]), .rectangle3_x(rectangle3_xs[667]), .rectangle3_y(rectangle3_ys[667]), .rectangle3_width(rectangle3_widths[667]), .rectangle3_height(rectangle3_heights[667]), .rectangle3_weight(rectangle3_weights[667]), .feature_threshold(feature_thresholds[667]), .feature_above(feature_aboves[667]), .feature_below(feature_belows[667]), .scan_win_std_dev(scan_win_std_dev[667]), .feature_accum(feature_accums[667]));
  accum_calculator ac668(.scan_win(scan_win668), .rectangle1_x(rectangle1_xs[668]), .rectangle1_y(rectangle1_ys[668]), .rectangle1_width(rectangle1_widths[668]), .rectangle1_height(rectangle1_heights[668]), .rectangle1_weight(rectangle1_weights[668]), .rectangle2_x(rectangle2_xs[668]), .rectangle2_y(rectangle2_ys[668]), .rectangle2_width(rectangle2_widths[668]), .rectangle2_height(rectangle2_heights[668]), .rectangle2_weight(rectangle2_weights[668]), .rectangle3_x(rectangle3_xs[668]), .rectangle3_y(rectangle3_ys[668]), .rectangle3_width(rectangle3_widths[668]), .rectangle3_height(rectangle3_heights[668]), .rectangle3_weight(rectangle3_weights[668]), .feature_threshold(feature_thresholds[668]), .feature_above(feature_aboves[668]), .feature_below(feature_belows[668]), .scan_win_std_dev(scan_win_std_dev[668]), .feature_accum(feature_accums[668]));
  accum_calculator ac669(.scan_win(scan_win669), .rectangle1_x(rectangle1_xs[669]), .rectangle1_y(rectangle1_ys[669]), .rectangle1_width(rectangle1_widths[669]), .rectangle1_height(rectangle1_heights[669]), .rectangle1_weight(rectangle1_weights[669]), .rectangle2_x(rectangle2_xs[669]), .rectangle2_y(rectangle2_ys[669]), .rectangle2_width(rectangle2_widths[669]), .rectangle2_height(rectangle2_heights[669]), .rectangle2_weight(rectangle2_weights[669]), .rectangle3_x(rectangle3_xs[669]), .rectangle3_y(rectangle3_ys[669]), .rectangle3_width(rectangle3_widths[669]), .rectangle3_height(rectangle3_heights[669]), .rectangle3_weight(rectangle3_weights[669]), .feature_threshold(feature_thresholds[669]), .feature_above(feature_aboves[669]), .feature_below(feature_belows[669]), .scan_win_std_dev(scan_win_std_dev[669]), .feature_accum(feature_accums[669]));
  accum_calculator ac670(.scan_win(scan_win670), .rectangle1_x(rectangle1_xs[670]), .rectangle1_y(rectangle1_ys[670]), .rectangle1_width(rectangle1_widths[670]), .rectangle1_height(rectangle1_heights[670]), .rectangle1_weight(rectangle1_weights[670]), .rectangle2_x(rectangle2_xs[670]), .rectangle2_y(rectangle2_ys[670]), .rectangle2_width(rectangle2_widths[670]), .rectangle2_height(rectangle2_heights[670]), .rectangle2_weight(rectangle2_weights[670]), .rectangle3_x(rectangle3_xs[670]), .rectangle3_y(rectangle3_ys[670]), .rectangle3_width(rectangle3_widths[670]), .rectangle3_height(rectangle3_heights[670]), .rectangle3_weight(rectangle3_weights[670]), .feature_threshold(feature_thresholds[670]), .feature_above(feature_aboves[670]), .feature_below(feature_belows[670]), .scan_win_std_dev(scan_win_std_dev[670]), .feature_accum(feature_accums[670]));
  accum_calculator ac671(.scan_win(scan_win671), .rectangle1_x(rectangle1_xs[671]), .rectangle1_y(rectangle1_ys[671]), .rectangle1_width(rectangle1_widths[671]), .rectangle1_height(rectangle1_heights[671]), .rectangle1_weight(rectangle1_weights[671]), .rectangle2_x(rectangle2_xs[671]), .rectangle2_y(rectangle2_ys[671]), .rectangle2_width(rectangle2_widths[671]), .rectangle2_height(rectangle2_heights[671]), .rectangle2_weight(rectangle2_weights[671]), .rectangle3_x(rectangle3_xs[671]), .rectangle3_y(rectangle3_ys[671]), .rectangle3_width(rectangle3_widths[671]), .rectangle3_height(rectangle3_heights[671]), .rectangle3_weight(rectangle3_weights[671]), .feature_threshold(feature_thresholds[671]), .feature_above(feature_aboves[671]), .feature_below(feature_belows[671]), .scan_win_std_dev(scan_win_std_dev[671]), .feature_accum(feature_accums[671]));
  accum_calculator ac672(.scan_win(scan_win672), .rectangle1_x(rectangle1_xs[672]), .rectangle1_y(rectangle1_ys[672]), .rectangle1_width(rectangle1_widths[672]), .rectangle1_height(rectangle1_heights[672]), .rectangle1_weight(rectangle1_weights[672]), .rectangle2_x(rectangle2_xs[672]), .rectangle2_y(rectangle2_ys[672]), .rectangle2_width(rectangle2_widths[672]), .rectangle2_height(rectangle2_heights[672]), .rectangle2_weight(rectangle2_weights[672]), .rectangle3_x(rectangle3_xs[672]), .rectangle3_y(rectangle3_ys[672]), .rectangle3_width(rectangle3_widths[672]), .rectangle3_height(rectangle3_heights[672]), .rectangle3_weight(rectangle3_weights[672]), .feature_threshold(feature_thresholds[672]), .feature_above(feature_aboves[672]), .feature_below(feature_belows[672]), .scan_win_std_dev(scan_win_std_dev[672]), .feature_accum(feature_accums[672]));
  accum_calculator ac673(.scan_win(scan_win673), .rectangle1_x(rectangle1_xs[673]), .rectangle1_y(rectangle1_ys[673]), .rectangle1_width(rectangle1_widths[673]), .rectangle1_height(rectangle1_heights[673]), .rectangle1_weight(rectangle1_weights[673]), .rectangle2_x(rectangle2_xs[673]), .rectangle2_y(rectangle2_ys[673]), .rectangle2_width(rectangle2_widths[673]), .rectangle2_height(rectangle2_heights[673]), .rectangle2_weight(rectangle2_weights[673]), .rectangle3_x(rectangle3_xs[673]), .rectangle3_y(rectangle3_ys[673]), .rectangle3_width(rectangle3_widths[673]), .rectangle3_height(rectangle3_heights[673]), .rectangle3_weight(rectangle3_weights[673]), .feature_threshold(feature_thresholds[673]), .feature_above(feature_aboves[673]), .feature_below(feature_belows[673]), .scan_win_std_dev(scan_win_std_dev[673]), .feature_accum(feature_accums[673]));
  accum_calculator ac674(.scan_win(scan_win674), .rectangle1_x(rectangle1_xs[674]), .rectangle1_y(rectangle1_ys[674]), .rectangle1_width(rectangle1_widths[674]), .rectangle1_height(rectangle1_heights[674]), .rectangle1_weight(rectangle1_weights[674]), .rectangle2_x(rectangle2_xs[674]), .rectangle2_y(rectangle2_ys[674]), .rectangle2_width(rectangle2_widths[674]), .rectangle2_height(rectangle2_heights[674]), .rectangle2_weight(rectangle2_weights[674]), .rectangle3_x(rectangle3_xs[674]), .rectangle3_y(rectangle3_ys[674]), .rectangle3_width(rectangle3_widths[674]), .rectangle3_height(rectangle3_heights[674]), .rectangle3_weight(rectangle3_weights[674]), .feature_threshold(feature_thresholds[674]), .feature_above(feature_aboves[674]), .feature_below(feature_belows[674]), .scan_win_std_dev(scan_win_std_dev[674]), .feature_accum(feature_accums[674]));
  accum_calculator ac675(.scan_win(scan_win675), .rectangle1_x(rectangle1_xs[675]), .rectangle1_y(rectangle1_ys[675]), .rectangle1_width(rectangle1_widths[675]), .rectangle1_height(rectangle1_heights[675]), .rectangle1_weight(rectangle1_weights[675]), .rectangle2_x(rectangle2_xs[675]), .rectangle2_y(rectangle2_ys[675]), .rectangle2_width(rectangle2_widths[675]), .rectangle2_height(rectangle2_heights[675]), .rectangle2_weight(rectangle2_weights[675]), .rectangle3_x(rectangle3_xs[675]), .rectangle3_y(rectangle3_ys[675]), .rectangle3_width(rectangle3_widths[675]), .rectangle3_height(rectangle3_heights[675]), .rectangle3_weight(rectangle3_weights[675]), .feature_threshold(feature_thresholds[675]), .feature_above(feature_aboves[675]), .feature_below(feature_belows[675]), .scan_win_std_dev(scan_win_std_dev[675]), .feature_accum(feature_accums[675]));
  accum_calculator ac676(.scan_win(scan_win676), .rectangle1_x(rectangle1_xs[676]), .rectangle1_y(rectangle1_ys[676]), .rectangle1_width(rectangle1_widths[676]), .rectangle1_height(rectangle1_heights[676]), .rectangle1_weight(rectangle1_weights[676]), .rectangle2_x(rectangle2_xs[676]), .rectangle2_y(rectangle2_ys[676]), .rectangle2_width(rectangle2_widths[676]), .rectangle2_height(rectangle2_heights[676]), .rectangle2_weight(rectangle2_weights[676]), .rectangle3_x(rectangle3_xs[676]), .rectangle3_y(rectangle3_ys[676]), .rectangle3_width(rectangle3_widths[676]), .rectangle3_height(rectangle3_heights[676]), .rectangle3_weight(rectangle3_weights[676]), .feature_threshold(feature_thresholds[676]), .feature_above(feature_aboves[676]), .feature_below(feature_belows[676]), .scan_win_std_dev(scan_win_std_dev[676]), .feature_accum(feature_accums[676]));
  accum_calculator ac677(.scan_win(scan_win677), .rectangle1_x(rectangle1_xs[677]), .rectangle1_y(rectangle1_ys[677]), .rectangle1_width(rectangle1_widths[677]), .rectangle1_height(rectangle1_heights[677]), .rectangle1_weight(rectangle1_weights[677]), .rectangle2_x(rectangle2_xs[677]), .rectangle2_y(rectangle2_ys[677]), .rectangle2_width(rectangle2_widths[677]), .rectangle2_height(rectangle2_heights[677]), .rectangle2_weight(rectangle2_weights[677]), .rectangle3_x(rectangle3_xs[677]), .rectangle3_y(rectangle3_ys[677]), .rectangle3_width(rectangle3_widths[677]), .rectangle3_height(rectangle3_heights[677]), .rectangle3_weight(rectangle3_weights[677]), .feature_threshold(feature_thresholds[677]), .feature_above(feature_aboves[677]), .feature_below(feature_belows[677]), .scan_win_std_dev(scan_win_std_dev[677]), .feature_accum(feature_accums[677]));
  accum_calculator ac678(.scan_win(scan_win678), .rectangle1_x(rectangle1_xs[678]), .rectangle1_y(rectangle1_ys[678]), .rectangle1_width(rectangle1_widths[678]), .rectangle1_height(rectangle1_heights[678]), .rectangle1_weight(rectangle1_weights[678]), .rectangle2_x(rectangle2_xs[678]), .rectangle2_y(rectangle2_ys[678]), .rectangle2_width(rectangle2_widths[678]), .rectangle2_height(rectangle2_heights[678]), .rectangle2_weight(rectangle2_weights[678]), .rectangle3_x(rectangle3_xs[678]), .rectangle3_y(rectangle3_ys[678]), .rectangle3_width(rectangle3_widths[678]), .rectangle3_height(rectangle3_heights[678]), .rectangle3_weight(rectangle3_weights[678]), .feature_threshold(feature_thresholds[678]), .feature_above(feature_aboves[678]), .feature_below(feature_belows[678]), .scan_win_std_dev(scan_win_std_dev[678]), .feature_accum(feature_accums[678]));
  accum_calculator ac679(.scan_win(scan_win679), .rectangle1_x(rectangle1_xs[679]), .rectangle1_y(rectangle1_ys[679]), .rectangle1_width(rectangle1_widths[679]), .rectangle1_height(rectangle1_heights[679]), .rectangle1_weight(rectangle1_weights[679]), .rectangle2_x(rectangle2_xs[679]), .rectangle2_y(rectangle2_ys[679]), .rectangle2_width(rectangle2_widths[679]), .rectangle2_height(rectangle2_heights[679]), .rectangle2_weight(rectangle2_weights[679]), .rectangle3_x(rectangle3_xs[679]), .rectangle3_y(rectangle3_ys[679]), .rectangle3_width(rectangle3_widths[679]), .rectangle3_height(rectangle3_heights[679]), .rectangle3_weight(rectangle3_weights[679]), .feature_threshold(feature_thresholds[679]), .feature_above(feature_aboves[679]), .feature_below(feature_belows[679]), .scan_win_std_dev(scan_win_std_dev[679]), .feature_accum(feature_accums[679]));
  accum_calculator ac680(.scan_win(scan_win680), .rectangle1_x(rectangle1_xs[680]), .rectangle1_y(rectangle1_ys[680]), .rectangle1_width(rectangle1_widths[680]), .rectangle1_height(rectangle1_heights[680]), .rectangle1_weight(rectangle1_weights[680]), .rectangle2_x(rectangle2_xs[680]), .rectangle2_y(rectangle2_ys[680]), .rectangle2_width(rectangle2_widths[680]), .rectangle2_height(rectangle2_heights[680]), .rectangle2_weight(rectangle2_weights[680]), .rectangle3_x(rectangle3_xs[680]), .rectangle3_y(rectangle3_ys[680]), .rectangle3_width(rectangle3_widths[680]), .rectangle3_height(rectangle3_heights[680]), .rectangle3_weight(rectangle3_weights[680]), .feature_threshold(feature_thresholds[680]), .feature_above(feature_aboves[680]), .feature_below(feature_belows[680]), .scan_win_std_dev(scan_win_std_dev[680]), .feature_accum(feature_accums[680]));
  accum_calculator ac681(.scan_win(scan_win681), .rectangle1_x(rectangle1_xs[681]), .rectangle1_y(rectangle1_ys[681]), .rectangle1_width(rectangle1_widths[681]), .rectangle1_height(rectangle1_heights[681]), .rectangle1_weight(rectangle1_weights[681]), .rectangle2_x(rectangle2_xs[681]), .rectangle2_y(rectangle2_ys[681]), .rectangle2_width(rectangle2_widths[681]), .rectangle2_height(rectangle2_heights[681]), .rectangle2_weight(rectangle2_weights[681]), .rectangle3_x(rectangle3_xs[681]), .rectangle3_y(rectangle3_ys[681]), .rectangle3_width(rectangle3_widths[681]), .rectangle3_height(rectangle3_heights[681]), .rectangle3_weight(rectangle3_weights[681]), .feature_threshold(feature_thresholds[681]), .feature_above(feature_aboves[681]), .feature_below(feature_belows[681]), .scan_win_std_dev(scan_win_std_dev[681]), .feature_accum(feature_accums[681]));
  accum_calculator ac682(.scan_win(scan_win682), .rectangle1_x(rectangle1_xs[682]), .rectangle1_y(rectangle1_ys[682]), .rectangle1_width(rectangle1_widths[682]), .rectangle1_height(rectangle1_heights[682]), .rectangle1_weight(rectangle1_weights[682]), .rectangle2_x(rectangle2_xs[682]), .rectangle2_y(rectangle2_ys[682]), .rectangle2_width(rectangle2_widths[682]), .rectangle2_height(rectangle2_heights[682]), .rectangle2_weight(rectangle2_weights[682]), .rectangle3_x(rectangle3_xs[682]), .rectangle3_y(rectangle3_ys[682]), .rectangle3_width(rectangle3_widths[682]), .rectangle3_height(rectangle3_heights[682]), .rectangle3_weight(rectangle3_weights[682]), .feature_threshold(feature_thresholds[682]), .feature_above(feature_aboves[682]), .feature_below(feature_belows[682]), .scan_win_std_dev(scan_win_std_dev[682]), .feature_accum(feature_accums[682]));
  accum_calculator ac683(.scan_win(scan_win683), .rectangle1_x(rectangle1_xs[683]), .rectangle1_y(rectangle1_ys[683]), .rectangle1_width(rectangle1_widths[683]), .rectangle1_height(rectangle1_heights[683]), .rectangle1_weight(rectangle1_weights[683]), .rectangle2_x(rectangle2_xs[683]), .rectangle2_y(rectangle2_ys[683]), .rectangle2_width(rectangle2_widths[683]), .rectangle2_height(rectangle2_heights[683]), .rectangle2_weight(rectangle2_weights[683]), .rectangle3_x(rectangle3_xs[683]), .rectangle3_y(rectangle3_ys[683]), .rectangle3_width(rectangle3_widths[683]), .rectangle3_height(rectangle3_heights[683]), .rectangle3_weight(rectangle3_weights[683]), .feature_threshold(feature_thresholds[683]), .feature_above(feature_aboves[683]), .feature_below(feature_belows[683]), .scan_win_std_dev(scan_win_std_dev[683]), .feature_accum(feature_accums[683]));
  accum_calculator ac684(.scan_win(scan_win684), .rectangle1_x(rectangle1_xs[684]), .rectangle1_y(rectangle1_ys[684]), .rectangle1_width(rectangle1_widths[684]), .rectangle1_height(rectangle1_heights[684]), .rectangle1_weight(rectangle1_weights[684]), .rectangle2_x(rectangle2_xs[684]), .rectangle2_y(rectangle2_ys[684]), .rectangle2_width(rectangle2_widths[684]), .rectangle2_height(rectangle2_heights[684]), .rectangle2_weight(rectangle2_weights[684]), .rectangle3_x(rectangle3_xs[684]), .rectangle3_y(rectangle3_ys[684]), .rectangle3_width(rectangle3_widths[684]), .rectangle3_height(rectangle3_heights[684]), .rectangle3_weight(rectangle3_weights[684]), .feature_threshold(feature_thresholds[684]), .feature_above(feature_aboves[684]), .feature_below(feature_belows[684]), .scan_win_std_dev(scan_win_std_dev[684]), .feature_accum(feature_accums[684]));
  accum_calculator ac685(.scan_win(scan_win685), .rectangle1_x(rectangle1_xs[685]), .rectangle1_y(rectangle1_ys[685]), .rectangle1_width(rectangle1_widths[685]), .rectangle1_height(rectangle1_heights[685]), .rectangle1_weight(rectangle1_weights[685]), .rectangle2_x(rectangle2_xs[685]), .rectangle2_y(rectangle2_ys[685]), .rectangle2_width(rectangle2_widths[685]), .rectangle2_height(rectangle2_heights[685]), .rectangle2_weight(rectangle2_weights[685]), .rectangle3_x(rectangle3_xs[685]), .rectangle3_y(rectangle3_ys[685]), .rectangle3_width(rectangle3_widths[685]), .rectangle3_height(rectangle3_heights[685]), .rectangle3_weight(rectangle3_weights[685]), .feature_threshold(feature_thresholds[685]), .feature_above(feature_aboves[685]), .feature_below(feature_belows[685]), .scan_win_std_dev(scan_win_std_dev[685]), .feature_accum(feature_accums[685]));
  accum_calculator ac686(.scan_win(scan_win686), .rectangle1_x(rectangle1_xs[686]), .rectangle1_y(rectangle1_ys[686]), .rectangle1_width(rectangle1_widths[686]), .rectangle1_height(rectangle1_heights[686]), .rectangle1_weight(rectangle1_weights[686]), .rectangle2_x(rectangle2_xs[686]), .rectangle2_y(rectangle2_ys[686]), .rectangle2_width(rectangle2_widths[686]), .rectangle2_height(rectangle2_heights[686]), .rectangle2_weight(rectangle2_weights[686]), .rectangle3_x(rectangle3_xs[686]), .rectangle3_y(rectangle3_ys[686]), .rectangle3_width(rectangle3_widths[686]), .rectangle3_height(rectangle3_heights[686]), .rectangle3_weight(rectangle3_weights[686]), .feature_threshold(feature_thresholds[686]), .feature_above(feature_aboves[686]), .feature_below(feature_belows[686]), .scan_win_std_dev(scan_win_std_dev[686]), .feature_accum(feature_accums[686]));
  accum_calculator ac687(.scan_win(scan_win687), .rectangle1_x(rectangle1_xs[687]), .rectangle1_y(rectangle1_ys[687]), .rectangle1_width(rectangle1_widths[687]), .rectangle1_height(rectangle1_heights[687]), .rectangle1_weight(rectangle1_weights[687]), .rectangle2_x(rectangle2_xs[687]), .rectangle2_y(rectangle2_ys[687]), .rectangle2_width(rectangle2_widths[687]), .rectangle2_height(rectangle2_heights[687]), .rectangle2_weight(rectangle2_weights[687]), .rectangle3_x(rectangle3_xs[687]), .rectangle3_y(rectangle3_ys[687]), .rectangle3_width(rectangle3_widths[687]), .rectangle3_height(rectangle3_heights[687]), .rectangle3_weight(rectangle3_weights[687]), .feature_threshold(feature_thresholds[687]), .feature_above(feature_aboves[687]), .feature_below(feature_belows[687]), .scan_win_std_dev(scan_win_std_dev[687]), .feature_accum(feature_accums[687]));
  accum_calculator ac688(.scan_win(scan_win688), .rectangle1_x(rectangle1_xs[688]), .rectangle1_y(rectangle1_ys[688]), .rectangle1_width(rectangle1_widths[688]), .rectangle1_height(rectangle1_heights[688]), .rectangle1_weight(rectangle1_weights[688]), .rectangle2_x(rectangle2_xs[688]), .rectangle2_y(rectangle2_ys[688]), .rectangle2_width(rectangle2_widths[688]), .rectangle2_height(rectangle2_heights[688]), .rectangle2_weight(rectangle2_weights[688]), .rectangle3_x(rectangle3_xs[688]), .rectangle3_y(rectangle3_ys[688]), .rectangle3_width(rectangle3_widths[688]), .rectangle3_height(rectangle3_heights[688]), .rectangle3_weight(rectangle3_weights[688]), .feature_threshold(feature_thresholds[688]), .feature_above(feature_aboves[688]), .feature_below(feature_belows[688]), .scan_win_std_dev(scan_win_std_dev[688]), .feature_accum(feature_accums[688]));
  accum_calculator ac689(.scan_win(scan_win689), .rectangle1_x(rectangle1_xs[689]), .rectangle1_y(rectangle1_ys[689]), .rectangle1_width(rectangle1_widths[689]), .rectangle1_height(rectangle1_heights[689]), .rectangle1_weight(rectangle1_weights[689]), .rectangle2_x(rectangle2_xs[689]), .rectangle2_y(rectangle2_ys[689]), .rectangle2_width(rectangle2_widths[689]), .rectangle2_height(rectangle2_heights[689]), .rectangle2_weight(rectangle2_weights[689]), .rectangle3_x(rectangle3_xs[689]), .rectangle3_y(rectangle3_ys[689]), .rectangle3_width(rectangle3_widths[689]), .rectangle3_height(rectangle3_heights[689]), .rectangle3_weight(rectangle3_weights[689]), .feature_threshold(feature_thresholds[689]), .feature_above(feature_aboves[689]), .feature_below(feature_belows[689]), .scan_win_std_dev(scan_win_std_dev[689]), .feature_accum(feature_accums[689]));
  accum_calculator ac690(.scan_win(scan_win690), .rectangle1_x(rectangle1_xs[690]), .rectangle1_y(rectangle1_ys[690]), .rectangle1_width(rectangle1_widths[690]), .rectangle1_height(rectangle1_heights[690]), .rectangle1_weight(rectangle1_weights[690]), .rectangle2_x(rectangle2_xs[690]), .rectangle2_y(rectangle2_ys[690]), .rectangle2_width(rectangle2_widths[690]), .rectangle2_height(rectangle2_heights[690]), .rectangle2_weight(rectangle2_weights[690]), .rectangle3_x(rectangle3_xs[690]), .rectangle3_y(rectangle3_ys[690]), .rectangle3_width(rectangle3_widths[690]), .rectangle3_height(rectangle3_heights[690]), .rectangle3_weight(rectangle3_weights[690]), .feature_threshold(feature_thresholds[690]), .feature_above(feature_aboves[690]), .feature_below(feature_belows[690]), .scan_win_std_dev(scan_win_std_dev[690]), .feature_accum(feature_accums[690]));
  accum_calculator ac691(.scan_win(scan_win691), .rectangle1_x(rectangle1_xs[691]), .rectangle1_y(rectangle1_ys[691]), .rectangle1_width(rectangle1_widths[691]), .rectangle1_height(rectangle1_heights[691]), .rectangle1_weight(rectangle1_weights[691]), .rectangle2_x(rectangle2_xs[691]), .rectangle2_y(rectangle2_ys[691]), .rectangle2_width(rectangle2_widths[691]), .rectangle2_height(rectangle2_heights[691]), .rectangle2_weight(rectangle2_weights[691]), .rectangle3_x(rectangle3_xs[691]), .rectangle3_y(rectangle3_ys[691]), .rectangle3_width(rectangle3_widths[691]), .rectangle3_height(rectangle3_heights[691]), .rectangle3_weight(rectangle3_weights[691]), .feature_threshold(feature_thresholds[691]), .feature_above(feature_aboves[691]), .feature_below(feature_belows[691]), .scan_win_std_dev(scan_win_std_dev[691]), .feature_accum(feature_accums[691]));
  accum_calculator ac692(.scan_win(scan_win692), .rectangle1_x(rectangle1_xs[692]), .rectangle1_y(rectangle1_ys[692]), .rectangle1_width(rectangle1_widths[692]), .rectangle1_height(rectangle1_heights[692]), .rectangle1_weight(rectangle1_weights[692]), .rectangle2_x(rectangle2_xs[692]), .rectangle2_y(rectangle2_ys[692]), .rectangle2_width(rectangle2_widths[692]), .rectangle2_height(rectangle2_heights[692]), .rectangle2_weight(rectangle2_weights[692]), .rectangle3_x(rectangle3_xs[692]), .rectangle3_y(rectangle3_ys[692]), .rectangle3_width(rectangle3_widths[692]), .rectangle3_height(rectangle3_heights[692]), .rectangle3_weight(rectangle3_weights[692]), .feature_threshold(feature_thresholds[692]), .feature_above(feature_aboves[692]), .feature_below(feature_belows[692]), .scan_win_std_dev(scan_win_std_dev[692]), .feature_accum(feature_accums[692]));
  accum_calculator ac693(.scan_win(scan_win693), .rectangle1_x(rectangle1_xs[693]), .rectangle1_y(rectangle1_ys[693]), .rectangle1_width(rectangle1_widths[693]), .rectangle1_height(rectangle1_heights[693]), .rectangle1_weight(rectangle1_weights[693]), .rectangle2_x(rectangle2_xs[693]), .rectangle2_y(rectangle2_ys[693]), .rectangle2_width(rectangle2_widths[693]), .rectangle2_height(rectangle2_heights[693]), .rectangle2_weight(rectangle2_weights[693]), .rectangle3_x(rectangle3_xs[693]), .rectangle3_y(rectangle3_ys[693]), .rectangle3_width(rectangle3_widths[693]), .rectangle3_height(rectangle3_heights[693]), .rectangle3_weight(rectangle3_weights[693]), .feature_threshold(feature_thresholds[693]), .feature_above(feature_aboves[693]), .feature_below(feature_belows[693]), .scan_win_std_dev(scan_win_std_dev[693]), .feature_accum(feature_accums[693]));
  accum_calculator ac694(.scan_win(scan_win694), .rectangle1_x(rectangle1_xs[694]), .rectangle1_y(rectangle1_ys[694]), .rectangle1_width(rectangle1_widths[694]), .rectangle1_height(rectangle1_heights[694]), .rectangle1_weight(rectangle1_weights[694]), .rectangle2_x(rectangle2_xs[694]), .rectangle2_y(rectangle2_ys[694]), .rectangle2_width(rectangle2_widths[694]), .rectangle2_height(rectangle2_heights[694]), .rectangle2_weight(rectangle2_weights[694]), .rectangle3_x(rectangle3_xs[694]), .rectangle3_y(rectangle3_ys[694]), .rectangle3_width(rectangle3_widths[694]), .rectangle3_height(rectangle3_heights[694]), .rectangle3_weight(rectangle3_weights[694]), .feature_threshold(feature_thresholds[694]), .feature_above(feature_aboves[694]), .feature_below(feature_belows[694]), .scan_win_std_dev(scan_win_std_dev[694]), .feature_accum(feature_accums[694]));
  accum_calculator ac695(.scan_win(scan_win695), .rectangle1_x(rectangle1_xs[695]), .rectangle1_y(rectangle1_ys[695]), .rectangle1_width(rectangle1_widths[695]), .rectangle1_height(rectangle1_heights[695]), .rectangle1_weight(rectangle1_weights[695]), .rectangle2_x(rectangle2_xs[695]), .rectangle2_y(rectangle2_ys[695]), .rectangle2_width(rectangle2_widths[695]), .rectangle2_height(rectangle2_heights[695]), .rectangle2_weight(rectangle2_weights[695]), .rectangle3_x(rectangle3_xs[695]), .rectangle3_y(rectangle3_ys[695]), .rectangle3_width(rectangle3_widths[695]), .rectangle3_height(rectangle3_heights[695]), .rectangle3_weight(rectangle3_weights[695]), .feature_threshold(feature_thresholds[695]), .feature_above(feature_aboves[695]), .feature_below(feature_belows[695]), .scan_win_std_dev(scan_win_std_dev[695]), .feature_accum(feature_accums[695]));
  accum_calculator ac696(.scan_win(scan_win696), .rectangle1_x(rectangle1_xs[696]), .rectangle1_y(rectangle1_ys[696]), .rectangle1_width(rectangle1_widths[696]), .rectangle1_height(rectangle1_heights[696]), .rectangle1_weight(rectangle1_weights[696]), .rectangle2_x(rectangle2_xs[696]), .rectangle2_y(rectangle2_ys[696]), .rectangle2_width(rectangle2_widths[696]), .rectangle2_height(rectangle2_heights[696]), .rectangle2_weight(rectangle2_weights[696]), .rectangle3_x(rectangle3_xs[696]), .rectangle3_y(rectangle3_ys[696]), .rectangle3_width(rectangle3_widths[696]), .rectangle3_height(rectangle3_heights[696]), .rectangle3_weight(rectangle3_weights[696]), .feature_threshold(feature_thresholds[696]), .feature_above(feature_aboves[696]), .feature_below(feature_belows[696]), .scan_win_std_dev(scan_win_std_dev[696]), .feature_accum(feature_accums[696]));
  accum_calculator ac697(.scan_win(scan_win697), .rectangle1_x(rectangle1_xs[697]), .rectangle1_y(rectangle1_ys[697]), .rectangle1_width(rectangle1_widths[697]), .rectangle1_height(rectangle1_heights[697]), .rectangle1_weight(rectangle1_weights[697]), .rectangle2_x(rectangle2_xs[697]), .rectangle2_y(rectangle2_ys[697]), .rectangle2_width(rectangle2_widths[697]), .rectangle2_height(rectangle2_heights[697]), .rectangle2_weight(rectangle2_weights[697]), .rectangle3_x(rectangle3_xs[697]), .rectangle3_y(rectangle3_ys[697]), .rectangle3_width(rectangle3_widths[697]), .rectangle3_height(rectangle3_heights[697]), .rectangle3_weight(rectangle3_weights[697]), .feature_threshold(feature_thresholds[697]), .feature_above(feature_aboves[697]), .feature_below(feature_belows[697]), .scan_win_std_dev(scan_win_std_dev[697]), .feature_accum(feature_accums[697]));
  accum_calculator ac698(.scan_win(scan_win698), .rectangle1_x(rectangle1_xs[698]), .rectangle1_y(rectangle1_ys[698]), .rectangle1_width(rectangle1_widths[698]), .rectangle1_height(rectangle1_heights[698]), .rectangle1_weight(rectangle1_weights[698]), .rectangle2_x(rectangle2_xs[698]), .rectangle2_y(rectangle2_ys[698]), .rectangle2_width(rectangle2_widths[698]), .rectangle2_height(rectangle2_heights[698]), .rectangle2_weight(rectangle2_weights[698]), .rectangle3_x(rectangle3_xs[698]), .rectangle3_y(rectangle3_ys[698]), .rectangle3_width(rectangle3_widths[698]), .rectangle3_height(rectangle3_heights[698]), .rectangle3_weight(rectangle3_weights[698]), .feature_threshold(feature_thresholds[698]), .feature_above(feature_aboves[698]), .feature_below(feature_belows[698]), .scan_win_std_dev(scan_win_std_dev[698]), .feature_accum(feature_accums[698]));
  accum_calculator ac699(.scan_win(scan_win699), .rectangle1_x(rectangle1_xs[699]), .rectangle1_y(rectangle1_ys[699]), .rectangle1_width(rectangle1_widths[699]), .rectangle1_height(rectangle1_heights[699]), .rectangle1_weight(rectangle1_weights[699]), .rectangle2_x(rectangle2_xs[699]), .rectangle2_y(rectangle2_ys[699]), .rectangle2_width(rectangle2_widths[699]), .rectangle2_height(rectangle2_heights[699]), .rectangle2_weight(rectangle2_weights[699]), .rectangle3_x(rectangle3_xs[699]), .rectangle3_y(rectangle3_ys[699]), .rectangle3_width(rectangle3_widths[699]), .rectangle3_height(rectangle3_heights[699]), .rectangle3_weight(rectangle3_weights[699]), .feature_threshold(feature_thresholds[699]), .feature_above(feature_aboves[699]), .feature_below(feature_belows[699]), .scan_win_std_dev(scan_win_std_dev[699]), .feature_accum(feature_accums[699]));
  accum_calculator ac700(.scan_win(scan_win700), .rectangle1_x(rectangle1_xs[700]), .rectangle1_y(rectangle1_ys[700]), .rectangle1_width(rectangle1_widths[700]), .rectangle1_height(rectangle1_heights[700]), .rectangle1_weight(rectangle1_weights[700]), .rectangle2_x(rectangle2_xs[700]), .rectangle2_y(rectangle2_ys[700]), .rectangle2_width(rectangle2_widths[700]), .rectangle2_height(rectangle2_heights[700]), .rectangle2_weight(rectangle2_weights[700]), .rectangle3_x(rectangle3_xs[700]), .rectangle3_y(rectangle3_ys[700]), .rectangle3_width(rectangle3_widths[700]), .rectangle3_height(rectangle3_heights[700]), .rectangle3_weight(rectangle3_weights[700]), .feature_threshold(feature_thresholds[700]), .feature_above(feature_aboves[700]), .feature_below(feature_belows[700]), .scan_win_std_dev(scan_win_std_dev[700]), .feature_accum(feature_accums[700]));
  accum_calculator ac701(.scan_win(scan_win701), .rectangle1_x(rectangle1_xs[701]), .rectangle1_y(rectangle1_ys[701]), .rectangle1_width(rectangle1_widths[701]), .rectangle1_height(rectangle1_heights[701]), .rectangle1_weight(rectangle1_weights[701]), .rectangle2_x(rectangle2_xs[701]), .rectangle2_y(rectangle2_ys[701]), .rectangle2_width(rectangle2_widths[701]), .rectangle2_height(rectangle2_heights[701]), .rectangle2_weight(rectangle2_weights[701]), .rectangle3_x(rectangle3_xs[701]), .rectangle3_y(rectangle3_ys[701]), .rectangle3_width(rectangle3_widths[701]), .rectangle3_height(rectangle3_heights[701]), .rectangle3_weight(rectangle3_weights[701]), .feature_threshold(feature_thresholds[701]), .feature_above(feature_aboves[701]), .feature_below(feature_belows[701]), .scan_win_std_dev(scan_win_std_dev[701]), .feature_accum(feature_accums[701]));
  accum_calculator ac702(.scan_win(scan_win702), .rectangle1_x(rectangle1_xs[702]), .rectangle1_y(rectangle1_ys[702]), .rectangle1_width(rectangle1_widths[702]), .rectangle1_height(rectangle1_heights[702]), .rectangle1_weight(rectangle1_weights[702]), .rectangle2_x(rectangle2_xs[702]), .rectangle2_y(rectangle2_ys[702]), .rectangle2_width(rectangle2_widths[702]), .rectangle2_height(rectangle2_heights[702]), .rectangle2_weight(rectangle2_weights[702]), .rectangle3_x(rectangle3_xs[702]), .rectangle3_y(rectangle3_ys[702]), .rectangle3_width(rectangle3_widths[702]), .rectangle3_height(rectangle3_heights[702]), .rectangle3_weight(rectangle3_weights[702]), .feature_threshold(feature_thresholds[702]), .feature_above(feature_aboves[702]), .feature_below(feature_belows[702]), .scan_win_std_dev(scan_win_std_dev[702]), .feature_accum(feature_accums[702]));
  accum_calculator ac703(.scan_win(scan_win703), .rectangle1_x(rectangle1_xs[703]), .rectangle1_y(rectangle1_ys[703]), .rectangle1_width(rectangle1_widths[703]), .rectangle1_height(rectangle1_heights[703]), .rectangle1_weight(rectangle1_weights[703]), .rectangle2_x(rectangle2_xs[703]), .rectangle2_y(rectangle2_ys[703]), .rectangle2_width(rectangle2_widths[703]), .rectangle2_height(rectangle2_heights[703]), .rectangle2_weight(rectangle2_weights[703]), .rectangle3_x(rectangle3_xs[703]), .rectangle3_y(rectangle3_ys[703]), .rectangle3_width(rectangle3_widths[703]), .rectangle3_height(rectangle3_heights[703]), .rectangle3_weight(rectangle3_weights[703]), .feature_threshold(feature_thresholds[703]), .feature_above(feature_aboves[703]), .feature_below(feature_belows[703]), .scan_win_std_dev(scan_win_std_dev[703]), .feature_accum(feature_accums[703]));
  accum_calculator ac704(.scan_win(scan_win704), .rectangle1_x(rectangle1_xs[704]), .rectangle1_y(rectangle1_ys[704]), .rectangle1_width(rectangle1_widths[704]), .rectangle1_height(rectangle1_heights[704]), .rectangle1_weight(rectangle1_weights[704]), .rectangle2_x(rectangle2_xs[704]), .rectangle2_y(rectangle2_ys[704]), .rectangle2_width(rectangle2_widths[704]), .rectangle2_height(rectangle2_heights[704]), .rectangle2_weight(rectangle2_weights[704]), .rectangle3_x(rectangle3_xs[704]), .rectangle3_y(rectangle3_ys[704]), .rectangle3_width(rectangle3_widths[704]), .rectangle3_height(rectangle3_heights[704]), .rectangle3_weight(rectangle3_weights[704]), .feature_threshold(feature_thresholds[704]), .feature_above(feature_aboves[704]), .feature_below(feature_belows[704]), .scan_win_std_dev(scan_win_std_dev[704]), .feature_accum(feature_accums[704]));
  accum_calculator ac705(.scan_win(scan_win705), .rectangle1_x(rectangle1_xs[705]), .rectangle1_y(rectangle1_ys[705]), .rectangle1_width(rectangle1_widths[705]), .rectangle1_height(rectangle1_heights[705]), .rectangle1_weight(rectangle1_weights[705]), .rectangle2_x(rectangle2_xs[705]), .rectangle2_y(rectangle2_ys[705]), .rectangle2_width(rectangle2_widths[705]), .rectangle2_height(rectangle2_heights[705]), .rectangle2_weight(rectangle2_weights[705]), .rectangle3_x(rectangle3_xs[705]), .rectangle3_y(rectangle3_ys[705]), .rectangle3_width(rectangle3_widths[705]), .rectangle3_height(rectangle3_heights[705]), .rectangle3_weight(rectangle3_weights[705]), .feature_threshold(feature_thresholds[705]), .feature_above(feature_aboves[705]), .feature_below(feature_belows[705]), .scan_win_std_dev(scan_win_std_dev[705]), .feature_accum(feature_accums[705]));
  accum_calculator ac706(.scan_win(scan_win706), .rectangle1_x(rectangle1_xs[706]), .rectangle1_y(rectangle1_ys[706]), .rectangle1_width(rectangle1_widths[706]), .rectangle1_height(rectangle1_heights[706]), .rectangle1_weight(rectangle1_weights[706]), .rectangle2_x(rectangle2_xs[706]), .rectangle2_y(rectangle2_ys[706]), .rectangle2_width(rectangle2_widths[706]), .rectangle2_height(rectangle2_heights[706]), .rectangle2_weight(rectangle2_weights[706]), .rectangle3_x(rectangle3_xs[706]), .rectangle3_y(rectangle3_ys[706]), .rectangle3_width(rectangle3_widths[706]), .rectangle3_height(rectangle3_heights[706]), .rectangle3_weight(rectangle3_weights[706]), .feature_threshold(feature_thresholds[706]), .feature_above(feature_aboves[706]), .feature_below(feature_belows[706]), .scan_win_std_dev(scan_win_std_dev[706]), .feature_accum(feature_accums[706]));
  accum_calculator ac707(.scan_win(scan_win707), .rectangle1_x(rectangle1_xs[707]), .rectangle1_y(rectangle1_ys[707]), .rectangle1_width(rectangle1_widths[707]), .rectangle1_height(rectangle1_heights[707]), .rectangle1_weight(rectangle1_weights[707]), .rectangle2_x(rectangle2_xs[707]), .rectangle2_y(rectangle2_ys[707]), .rectangle2_width(rectangle2_widths[707]), .rectangle2_height(rectangle2_heights[707]), .rectangle2_weight(rectangle2_weights[707]), .rectangle3_x(rectangle3_xs[707]), .rectangle3_y(rectangle3_ys[707]), .rectangle3_width(rectangle3_widths[707]), .rectangle3_height(rectangle3_heights[707]), .rectangle3_weight(rectangle3_weights[707]), .feature_threshold(feature_thresholds[707]), .feature_above(feature_aboves[707]), .feature_below(feature_belows[707]), .scan_win_std_dev(scan_win_std_dev[707]), .feature_accum(feature_accums[707]));
  accum_calculator ac708(.scan_win(scan_win708), .rectangle1_x(rectangle1_xs[708]), .rectangle1_y(rectangle1_ys[708]), .rectangle1_width(rectangle1_widths[708]), .rectangle1_height(rectangle1_heights[708]), .rectangle1_weight(rectangle1_weights[708]), .rectangle2_x(rectangle2_xs[708]), .rectangle2_y(rectangle2_ys[708]), .rectangle2_width(rectangle2_widths[708]), .rectangle2_height(rectangle2_heights[708]), .rectangle2_weight(rectangle2_weights[708]), .rectangle3_x(rectangle3_xs[708]), .rectangle3_y(rectangle3_ys[708]), .rectangle3_width(rectangle3_widths[708]), .rectangle3_height(rectangle3_heights[708]), .rectangle3_weight(rectangle3_weights[708]), .feature_threshold(feature_thresholds[708]), .feature_above(feature_aboves[708]), .feature_below(feature_belows[708]), .scan_win_std_dev(scan_win_std_dev[708]), .feature_accum(feature_accums[708]));
  accum_calculator ac709(.scan_win(scan_win709), .rectangle1_x(rectangle1_xs[709]), .rectangle1_y(rectangle1_ys[709]), .rectangle1_width(rectangle1_widths[709]), .rectangle1_height(rectangle1_heights[709]), .rectangle1_weight(rectangle1_weights[709]), .rectangle2_x(rectangle2_xs[709]), .rectangle2_y(rectangle2_ys[709]), .rectangle2_width(rectangle2_widths[709]), .rectangle2_height(rectangle2_heights[709]), .rectangle2_weight(rectangle2_weights[709]), .rectangle3_x(rectangle3_xs[709]), .rectangle3_y(rectangle3_ys[709]), .rectangle3_width(rectangle3_widths[709]), .rectangle3_height(rectangle3_heights[709]), .rectangle3_weight(rectangle3_weights[709]), .feature_threshold(feature_thresholds[709]), .feature_above(feature_aboves[709]), .feature_below(feature_belows[709]), .scan_win_std_dev(scan_win_std_dev[709]), .feature_accum(feature_accums[709]));
  accum_calculator ac710(.scan_win(scan_win710), .rectangle1_x(rectangle1_xs[710]), .rectangle1_y(rectangle1_ys[710]), .rectangle1_width(rectangle1_widths[710]), .rectangle1_height(rectangle1_heights[710]), .rectangle1_weight(rectangle1_weights[710]), .rectangle2_x(rectangle2_xs[710]), .rectangle2_y(rectangle2_ys[710]), .rectangle2_width(rectangle2_widths[710]), .rectangle2_height(rectangle2_heights[710]), .rectangle2_weight(rectangle2_weights[710]), .rectangle3_x(rectangle3_xs[710]), .rectangle3_y(rectangle3_ys[710]), .rectangle3_width(rectangle3_widths[710]), .rectangle3_height(rectangle3_heights[710]), .rectangle3_weight(rectangle3_weights[710]), .feature_threshold(feature_thresholds[710]), .feature_above(feature_aboves[710]), .feature_below(feature_belows[710]), .scan_win_std_dev(scan_win_std_dev[710]), .feature_accum(feature_accums[710]));
  accum_calculator ac711(.scan_win(scan_win711), .rectangle1_x(rectangle1_xs[711]), .rectangle1_y(rectangle1_ys[711]), .rectangle1_width(rectangle1_widths[711]), .rectangle1_height(rectangle1_heights[711]), .rectangle1_weight(rectangle1_weights[711]), .rectangle2_x(rectangle2_xs[711]), .rectangle2_y(rectangle2_ys[711]), .rectangle2_width(rectangle2_widths[711]), .rectangle2_height(rectangle2_heights[711]), .rectangle2_weight(rectangle2_weights[711]), .rectangle3_x(rectangle3_xs[711]), .rectangle3_y(rectangle3_ys[711]), .rectangle3_width(rectangle3_widths[711]), .rectangle3_height(rectangle3_heights[711]), .rectangle3_weight(rectangle3_weights[711]), .feature_threshold(feature_thresholds[711]), .feature_above(feature_aboves[711]), .feature_below(feature_belows[711]), .scan_win_std_dev(scan_win_std_dev[711]), .feature_accum(feature_accums[711]));
  accum_calculator ac712(.scan_win(scan_win712), .rectangle1_x(rectangle1_xs[712]), .rectangle1_y(rectangle1_ys[712]), .rectangle1_width(rectangle1_widths[712]), .rectangle1_height(rectangle1_heights[712]), .rectangle1_weight(rectangle1_weights[712]), .rectangle2_x(rectangle2_xs[712]), .rectangle2_y(rectangle2_ys[712]), .rectangle2_width(rectangle2_widths[712]), .rectangle2_height(rectangle2_heights[712]), .rectangle2_weight(rectangle2_weights[712]), .rectangle3_x(rectangle3_xs[712]), .rectangle3_y(rectangle3_ys[712]), .rectangle3_width(rectangle3_widths[712]), .rectangle3_height(rectangle3_heights[712]), .rectangle3_weight(rectangle3_weights[712]), .feature_threshold(feature_thresholds[712]), .feature_above(feature_aboves[712]), .feature_below(feature_belows[712]), .scan_win_std_dev(scan_win_std_dev[712]), .feature_accum(feature_accums[712]));
  accum_calculator ac713(.scan_win(scan_win713), .rectangle1_x(rectangle1_xs[713]), .rectangle1_y(rectangle1_ys[713]), .rectangle1_width(rectangle1_widths[713]), .rectangle1_height(rectangle1_heights[713]), .rectangle1_weight(rectangle1_weights[713]), .rectangle2_x(rectangle2_xs[713]), .rectangle2_y(rectangle2_ys[713]), .rectangle2_width(rectangle2_widths[713]), .rectangle2_height(rectangle2_heights[713]), .rectangle2_weight(rectangle2_weights[713]), .rectangle3_x(rectangle3_xs[713]), .rectangle3_y(rectangle3_ys[713]), .rectangle3_width(rectangle3_widths[713]), .rectangle3_height(rectangle3_heights[713]), .rectangle3_weight(rectangle3_weights[713]), .feature_threshold(feature_thresholds[713]), .feature_above(feature_aboves[713]), .feature_below(feature_belows[713]), .scan_win_std_dev(scan_win_std_dev[713]), .feature_accum(feature_accums[713]));
  accum_calculator ac714(.scan_win(scan_win714), .rectangle1_x(rectangle1_xs[714]), .rectangle1_y(rectangle1_ys[714]), .rectangle1_width(rectangle1_widths[714]), .rectangle1_height(rectangle1_heights[714]), .rectangle1_weight(rectangle1_weights[714]), .rectangle2_x(rectangle2_xs[714]), .rectangle2_y(rectangle2_ys[714]), .rectangle2_width(rectangle2_widths[714]), .rectangle2_height(rectangle2_heights[714]), .rectangle2_weight(rectangle2_weights[714]), .rectangle3_x(rectangle3_xs[714]), .rectangle3_y(rectangle3_ys[714]), .rectangle3_width(rectangle3_widths[714]), .rectangle3_height(rectangle3_heights[714]), .rectangle3_weight(rectangle3_weights[714]), .feature_threshold(feature_thresholds[714]), .feature_above(feature_aboves[714]), .feature_below(feature_belows[714]), .scan_win_std_dev(scan_win_std_dev[714]), .feature_accum(feature_accums[714]));
  accum_calculator ac715(.scan_win(scan_win715), .rectangle1_x(rectangle1_xs[715]), .rectangle1_y(rectangle1_ys[715]), .rectangle1_width(rectangle1_widths[715]), .rectangle1_height(rectangle1_heights[715]), .rectangle1_weight(rectangle1_weights[715]), .rectangle2_x(rectangle2_xs[715]), .rectangle2_y(rectangle2_ys[715]), .rectangle2_width(rectangle2_widths[715]), .rectangle2_height(rectangle2_heights[715]), .rectangle2_weight(rectangle2_weights[715]), .rectangle3_x(rectangle3_xs[715]), .rectangle3_y(rectangle3_ys[715]), .rectangle3_width(rectangle3_widths[715]), .rectangle3_height(rectangle3_heights[715]), .rectangle3_weight(rectangle3_weights[715]), .feature_threshold(feature_thresholds[715]), .feature_above(feature_aboves[715]), .feature_below(feature_belows[715]), .scan_win_std_dev(scan_win_std_dev[715]), .feature_accum(feature_accums[715]));
  accum_calculator ac716(.scan_win(scan_win716), .rectangle1_x(rectangle1_xs[716]), .rectangle1_y(rectangle1_ys[716]), .rectangle1_width(rectangle1_widths[716]), .rectangle1_height(rectangle1_heights[716]), .rectangle1_weight(rectangle1_weights[716]), .rectangle2_x(rectangle2_xs[716]), .rectangle2_y(rectangle2_ys[716]), .rectangle2_width(rectangle2_widths[716]), .rectangle2_height(rectangle2_heights[716]), .rectangle2_weight(rectangle2_weights[716]), .rectangle3_x(rectangle3_xs[716]), .rectangle3_y(rectangle3_ys[716]), .rectangle3_width(rectangle3_widths[716]), .rectangle3_height(rectangle3_heights[716]), .rectangle3_weight(rectangle3_weights[716]), .feature_threshold(feature_thresholds[716]), .feature_above(feature_aboves[716]), .feature_below(feature_belows[716]), .scan_win_std_dev(scan_win_std_dev[716]), .feature_accum(feature_accums[716]));
  accum_calculator ac717(.scan_win(scan_win717), .rectangle1_x(rectangle1_xs[717]), .rectangle1_y(rectangle1_ys[717]), .rectangle1_width(rectangle1_widths[717]), .rectangle1_height(rectangle1_heights[717]), .rectangle1_weight(rectangle1_weights[717]), .rectangle2_x(rectangle2_xs[717]), .rectangle2_y(rectangle2_ys[717]), .rectangle2_width(rectangle2_widths[717]), .rectangle2_height(rectangle2_heights[717]), .rectangle2_weight(rectangle2_weights[717]), .rectangle3_x(rectangle3_xs[717]), .rectangle3_y(rectangle3_ys[717]), .rectangle3_width(rectangle3_widths[717]), .rectangle3_height(rectangle3_heights[717]), .rectangle3_weight(rectangle3_weights[717]), .feature_threshold(feature_thresholds[717]), .feature_above(feature_aboves[717]), .feature_below(feature_belows[717]), .scan_win_std_dev(scan_win_std_dev[717]), .feature_accum(feature_accums[717]));
  accum_calculator ac718(.scan_win(scan_win718), .rectangle1_x(rectangle1_xs[718]), .rectangle1_y(rectangle1_ys[718]), .rectangle1_width(rectangle1_widths[718]), .rectangle1_height(rectangle1_heights[718]), .rectangle1_weight(rectangle1_weights[718]), .rectangle2_x(rectangle2_xs[718]), .rectangle2_y(rectangle2_ys[718]), .rectangle2_width(rectangle2_widths[718]), .rectangle2_height(rectangle2_heights[718]), .rectangle2_weight(rectangle2_weights[718]), .rectangle3_x(rectangle3_xs[718]), .rectangle3_y(rectangle3_ys[718]), .rectangle3_width(rectangle3_widths[718]), .rectangle3_height(rectangle3_heights[718]), .rectangle3_weight(rectangle3_weights[718]), .feature_threshold(feature_thresholds[718]), .feature_above(feature_aboves[718]), .feature_below(feature_belows[718]), .scan_win_std_dev(scan_win_std_dev[718]), .feature_accum(feature_accums[718]));
  accum_calculator ac719(.scan_win(scan_win719), .rectangle1_x(rectangle1_xs[719]), .rectangle1_y(rectangle1_ys[719]), .rectangle1_width(rectangle1_widths[719]), .rectangle1_height(rectangle1_heights[719]), .rectangle1_weight(rectangle1_weights[719]), .rectangle2_x(rectangle2_xs[719]), .rectangle2_y(rectangle2_ys[719]), .rectangle2_width(rectangle2_widths[719]), .rectangle2_height(rectangle2_heights[719]), .rectangle2_weight(rectangle2_weights[719]), .rectangle3_x(rectangle3_xs[719]), .rectangle3_y(rectangle3_ys[719]), .rectangle3_width(rectangle3_widths[719]), .rectangle3_height(rectangle3_heights[719]), .rectangle3_weight(rectangle3_weights[719]), .feature_threshold(feature_thresholds[719]), .feature_above(feature_aboves[719]), .feature_below(feature_belows[719]), .scan_win_std_dev(scan_win_std_dev[719]), .feature_accum(feature_accums[719]));
  accum_calculator ac720(.scan_win(scan_win720), .rectangle1_x(rectangle1_xs[720]), .rectangle1_y(rectangle1_ys[720]), .rectangle1_width(rectangle1_widths[720]), .rectangle1_height(rectangle1_heights[720]), .rectangle1_weight(rectangle1_weights[720]), .rectangle2_x(rectangle2_xs[720]), .rectangle2_y(rectangle2_ys[720]), .rectangle2_width(rectangle2_widths[720]), .rectangle2_height(rectangle2_heights[720]), .rectangle2_weight(rectangle2_weights[720]), .rectangle3_x(rectangle3_xs[720]), .rectangle3_y(rectangle3_ys[720]), .rectangle3_width(rectangle3_widths[720]), .rectangle3_height(rectangle3_heights[720]), .rectangle3_weight(rectangle3_weights[720]), .feature_threshold(feature_thresholds[720]), .feature_above(feature_aboves[720]), .feature_below(feature_belows[720]), .scan_win_std_dev(scan_win_std_dev[720]), .feature_accum(feature_accums[720]));
  accum_calculator ac721(.scan_win(scan_win721), .rectangle1_x(rectangle1_xs[721]), .rectangle1_y(rectangle1_ys[721]), .rectangle1_width(rectangle1_widths[721]), .rectangle1_height(rectangle1_heights[721]), .rectangle1_weight(rectangle1_weights[721]), .rectangle2_x(rectangle2_xs[721]), .rectangle2_y(rectangle2_ys[721]), .rectangle2_width(rectangle2_widths[721]), .rectangle2_height(rectangle2_heights[721]), .rectangle2_weight(rectangle2_weights[721]), .rectangle3_x(rectangle3_xs[721]), .rectangle3_y(rectangle3_ys[721]), .rectangle3_width(rectangle3_widths[721]), .rectangle3_height(rectangle3_heights[721]), .rectangle3_weight(rectangle3_weights[721]), .feature_threshold(feature_thresholds[721]), .feature_above(feature_aboves[721]), .feature_below(feature_belows[721]), .scan_win_std_dev(scan_win_std_dev[721]), .feature_accum(feature_accums[721]));
  accum_calculator ac722(.scan_win(scan_win722), .rectangle1_x(rectangle1_xs[722]), .rectangle1_y(rectangle1_ys[722]), .rectangle1_width(rectangle1_widths[722]), .rectangle1_height(rectangle1_heights[722]), .rectangle1_weight(rectangle1_weights[722]), .rectangle2_x(rectangle2_xs[722]), .rectangle2_y(rectangle2_ys[722]), .rectangle2_width(rectangle2_widths[722]), .rectangle2_height(rectangle2_heights[722]), .rectangle2_weight(rectangle2_weights[722]), .rectangle3_x(rectangle3_xs[722]), .rectangle3_y(rectangle3_ys[722]), .rectangle3_width(rectangle3_widths[722]), .rectangle3_height(rectangle3_heights[722]), .rectangle3_weight(rectangle3_weights[722]), .feature_threshold(feature_thresholds[722]), .feature_above(feature_aboves[722]), .feature_below(feature_belows[722]), .scan_win_std_dev(scan_win_std_dev[722]), .feature_accum(feature_accums[722]));
  accum_calculator ac723(.scan_win(scan_win723), .rectangle1_x(rectangle1_xs[723]), .rectangle1_y(rectangle1_ys[723]), .rectangle1_width(rectangle1_widths[723]), .rectangle1_height(rectangle1_heights[723]), .rectangle1_weight(rectangle1_weights[723]), .rectangle2_x(rectangle2_xs[723]), .rectangle2_y(rectangle2_ys[723]), .rectangle2_width(rectangle2_widths[723]), .rectangle2_height(rectangle2_heights[723]), .rectangle2_weight(rectangle2_weights[723]), .rectangle3_x(rectangle3_xs[723]), .rectangle3_y(rectangle3_ys[723]), .rectangle3_width(rectangle3_widths[723]), .rectangle3_height(rectangle3_heights[723]), .rectangle3_weight(rectangle3_weights[723]), .feature_threshold(feature_thresholds[723]), .feature_above(feature_aboves[723]), .feature_below(feature_belows[723]), .scan_win_std_dev(scan_win_std_dev[723]), .feature_accum(feature_accums[723]));
  accum_calculator ac724(.scan_win(scan_win724), .rectangle1_x(rectangle1_xs[724]), .rectangle1_y(rectangle1_ys[724]), .rectangle1_width(rectangle1_widths[724]), .rectangle1_height(rectangle1_heights[724]), .rectangle1_weight(rectangle1_weights[724]), .rectangle2_x(rectangle2_xs[724]), .rectangle2_y(rectangle2_ys[724]), .rectangle2_width(rectangle2_widths[724]), .rectangle2_height(rectangle2_heights[724]), .rectangle2_weight(rectangle2_weights[724]), .rectangle3_x(rectangle3_xs[724]), .rectangle3_y(rectangle3_ys[724]), .rectangle3_width(rectangle3_widths[724]), .rectangle3_height(rectangle3_heights[724]), .rectangle3_weight(rectangle3_weights[724]), .feature_threshold(feature_thresholds[724]), .feature_above(feature_aboves[724]), .feature_below(feature_belows[724]), .scan_win_std_dev(scan_win_std_dev[724]), .feature_accum(feature_accums[724]));
  accum_calculator ac725(.scan_win(scan_win725), .rectangle1_x(rectangle1_xs[725]), .rectangle1_y(rectangle1_ys[725]), .rectangle1_width(rectangle1_widths[725]), .rectangle1_height(rectangle1_heights[725]), .rectangle1_weight(rectangle1_weights[725]), .rectangle2_x(rectangle2_xs[725]), .rectangle2_y(rectangle2_ys[725]), .rectangle2_width(rectangle2_widths[725]), .rectangle2_height(rectangle2_heights[725]), .rectangle2_weight(rectangle2_weights[725]), .rectangle3_x(rectangle3_xs[725]), .rectangle3_y(rectangle3_ys[725]), .rectangle3_width(rectangle3_widths[725]), .rectangle3_height(rectangle3_heights[725]), .rectangle3_weight(rectangle3_weights[725]), .feature_threshold(feature_thresholds[725]), .feature_above(feature_aboves[725]), .feature_below(feature_belows[725]), .scan_win_std_dev(scan_win_std_dev[725]), .feature_accum(feature_accums[725]));
  accum_calculator ac726(.scan_win(scan_win726), .rectangle1_x(rectangle1_xs[726]), .rectangle1_y(rectangle1_ys[726]), .rectangle1_width(rectangle1_widths[726]), .rectangle1_height(rectangle1_heights[726]), .rectangle1_weight(rectangle1_weights[726]), .rectangle2_x(rectangle2_xs[726]), .rectangle2_y(rectangle2_ys[726]), .rectangle2_width(rectangle2_widths[726]), .rectangle2_height(rectangle2_heights[726]), .rectangle2_weight(rectangle2_weights[726]), .rectangle3_x(rectangle3_xs[726]), .rectangle3_y(rectangle3_ys[726]), .rectangle3_width(rectangle3_widths[726]), .rectangle3_height(rectangle3_heights[726]), .rectangle3_weight(rectangle3_weights[726]), .feature_threshold(feature_thresholds[726]), .feature_above(feature_aboves[726]), .feature_below(feature_belows[726]), .scan_win_std_dev(scan_win_std_dev[726]), .feature_accum(feature_accums[726]));
  accum_calculator ac727(.scan_win(scan_win727), .rectangle1_x(rectangle1_xs[727]), .rectangle1_y(rectangle1_ys[727]), .rectangle1_width(rectangle1_widths[727]), .rectangle1_height(rectangle1_heights[727]), .rectangle1_weight(rectangle1_weights[727]), .rectangle2_x(rectangle2_xs[727]), .rectangle2_y(rectangle2_ys[727]), .rectangle2_width(rectangle2_widths[727]), .rectangle2_height(rectangle2_heights[727]), .rectangle2_weight(rectangle2_weights[727]), .rectangle3_x(rectangle3_xs[727]), .rectangle3_y(rectangle3_ys[727]), .rectangle3_width(rectangle3_widths[727]), .rectangle3_height(rectangle3_heights[727]), .rectangle3_weight(rectangle3_weights[727]), .feature_threshold(feature_thresholds[727]), .feature_above(feature_aboves[727]), .feature_below(feature_belows[727]), .scan_win_std_dev(scan_win_std_dev[727]), .feature_accum(feature_accums[727]));
  accum_calculator ac728(.scan_win(scan_win728), .rectangle1_x(rectangle1_xs[728]), .rectangle1_y(rectangle1_ys[728]), .rectangle1_width(rectangle1_widths[728]), .rectangle1_height(rectangle1_heights[728]), .rectangle1_weight(rectangle1_weights[728]), .rectangle2_x(rectangle2_xs[728]), .rectangle2_y(rectangle2_ys[728]), .rectangle2_width(rectangle2_widths[728]), .rectangle2_height(rectangle2_heights[728]), .rectangle2_weight(rectangle2_weights[728]), .rectangle3_x(rectangle3_xs[728]), .rectangle3_y(rectangle3_ys[728]), .rectangle3_width(rectangle3_widths[728]), .rectangle3_height(rectangle3_heights[728]), .rectangle3_weight(rectangle3_weights[728]), .feature_threshold(feature_thresholds[728]), .feature_above(feature_aboves[728]), .feature_below(feature_belows[728]), .scan_win_std_dev(scan_win_std_dev[728]), .feature_accum(feature_accums[728]));
  accum_calculator ac729(.scan_win(scan_win729), .rectangle1_x(rectangle1_xs[729]), .rectangle1_y(rectangle1_ys[729]), .rectangle1_width(rectangle1_widths[729]), .rectangle1_height(rectangle1_heights[729]), .rectangle1_weight(rectangle1_weights[729]), .rectangle2_x(rectangle2_xs[729]), .rectangle2_y(rectangle2_ys[729]), .rectangle2_width(rectangle2_widths[729]), .rectangle2_height(rectangle2_heights[729]), .rectangle2_weight(rectangle2_weights[729]), .rectangle3_x(rectangle3_xs[729]), .rectangle3_y(rectangle3_ys[729]), .rectangle3_width(rectangle3_widths[729]), .rectangle3_height(rectangle3_heights[729]), .rectangle3_weight(rectangle3_weights[729]), .feature_threshold(feature_thresholds[729]), .feature_above(feature_aboves[729]), .feature_below(feature_belows[729]), .scan_win_std_dev(scan_win_std_dev[729]), .feature_accum(feature_accums[729]));
  accum_calculator ac730(.scan_win(scan_win730), .rectangle1_x(rectangle1_xs[730]), .rectangle1_y(rectangle1_ys[730]), .rectangle1_width(rectangle1_widths[730]), .rectangle1_height(rectangle1_heights[730]), .rectangle1_weight(rectangle1_weights[730]), .rectangle2_x(rectangle2_xs[730]), .rectangle2_y(rectangle2_ys[730]), .rectangle2_width(rectangle2_widths[730]), .rectangle2_height(rectangle2_heights[730]), .rectangle2_weight(rectangle2_weights[730]), .rectangle3_x(rectangle3_xs[730]), .rectangle3_y(rectangle3_ys[730]), .rectangle3_width(rectangle3_widths[730]), .rectangle3_height(rectangle3_heights[730]), .rectangle3_weight(rectangle3_weights[730]), .feature_threshold(feature_thresholds[730]), .feature_above(feature_aboves[730]), .feature_below(feature_belows[730]), .scan_win_std_dev(scan_win_std_dev[730]), .feature_accum(feature_accums[730]));
  accum_calculator ac731(.scan_win(scan_win731), .rectangle1_x(rectangle1_xs[731]), .rectangle1_y(rectangle1_ys[731]), .rectangle1_width(rectangle1_widths[731]), .rectangle1_height(rectangle1_heights[731]), .rectangle1_weight(rectangle1_weights[731]), .rectangle2_x(rectangle2_xs[731]), .rectangle2_y(rectangle2_ys[731]), .rectangle2_width(rectangle2_widths[731]), .rectangle2_height(rectangle2_heights[731]), .rectangle2_weight(rectangle2_weights[731]), .rectangle3_x(rectangle3_xs[731]), .rectangle3_y(rectangle3_ys[731]), .rectangle3_width(rectangle3_widths[731]), .rectangle3_height(rectangle3_heights[731]), .rectangle3_weight(rectangle3_weights[731]), .feature_threshold(feature_thresholds[731]), .feature_above(feature_aboves[731]), .feature_below(feature_belows[731]), .scan_win_std_dev(scan_win_std_dev[731]), .feature_accum(feature_accums[731]));
  accum_calculator ac732(.scan_win(scan_win732), .rectangle1_x(rectangle1_xs[732]), .rectangle1_y(rectangle1_ys[732]), .rectangle1_width(rectangle1_widths[732]), .rectangle1_height(rectangle1_heights[732]), .rectangle1_weight(rectangle1_weights[732]), .rectangle2_x(rectangle2_xs[732]), .rectangle2_y(rectangle2_ys[732]), .rectangle2_width(rectangle2_widths[732]), .rectangle2_height(rectangle2_heights[732]), .rectangle2_weight(rectangle2_weights[732]), .rectangle3_x(rectangle3_xs[732]), .rectangle3_y(rectangle3_ys[732]), .rectangle3_width(rectangle3_widths[732]), .rectangle3_height(rectangle3_heights[732]), .rectangle3_weight(rectangle3_weights[732]), .feature_threshold(feature_thresholds[732]), .feature_above(feature_aboves[732]), .feature_below(feature_belows[732]), .scan_win_std_dev(scan_win_std_dev[732]), .feature_accum(feature_accums[732]));
  accum_calculator ac733(.scan_win(scan_win733), .rectangle1_x(rectangle1_xs[733]), .rectangle1_y(rectangle1_ys[733]), .rectangle1_width(rectangle1_widths[733]), .rectangle1_height(rectangle1_heights[733]), .rectangle1_weight(rectangle1_weights[733]), .rectangle2_x(rectangle2_xs[733]), .rectangle2_y(rectangle2_ys[733]), .rectangle2_width(rectangle2_widths[733]), .rectangle2_height(rectangle2_heights[733]), .rectangle2_weight(rectangle2_weights[733]), .rectangle3_x(rectangle3_xs[733]), .rectangle3_y(rectangle3_ys[733]), .rectangle3_width(rectangle3_widths[733]), .rectangle3_height(rectangle3_heights[733]), .rectangle3_weight(rectangle3_weights[733]), .feature_threshold(feature_thresholds[733]), .feature_above(feature_aboves[733]), .feature_below(feature_belows[733]), .scan_win_std_dev(scan_win_std_dev[733]), .feature_accum(feature_accums[733]));
  accum_calculator ac734(.scan_win(scan_win734), .rectangle1_x(rectangle1_xs[734]), .rectangle1_y(rectangle1_ys[734]), .rectangle1_width(rectangle1_widths[734]), .rectangle1_height(rectangle1_heights[734]), .rectangle1_weight(rectangle1_weights[734]), .rectangle2_x(rectangle2_xs[734]), .rectangle2_y(rectangle2_ys[734]), .rectangle2_width(rectangle2_widths[734]), .rectangle2_height(rectangle2_heights[734]), .rectangle2_weight(rectangle2_weights[734]), .rectangle3_x(rectangle3_xs[734]), .rectangle3_y(rectangle3_ys[734]), .rectangle3_width(rectangle3_widths[734]), .rectangle3_height(rectangle3_heights[734]), .rectangle3_weight(rectangle3_weights[734]), .feature_threshold(feature_thresholds[734]), .feature_above(feature_aboves[734]), .feature_below(feature_belows[734]), .scan_win_std_dev(scan_win_std_dev[734]), .feature_accum(feature_accums[734]));
  accum_calculator ac735(.scan_win(scan_win735), .rectangle1_x(rectangle1_xs[735]), .rectangle1_y(rectangle1_ys[735]), .rectangle1_width(rectangle1_widths[735]), .rectangle1_height(rectangle1_heights[735]), .rectangle1_weight(rectangle1_weights[735]), .rectangle2_x(rectangle2_xs[735]), .rectangle2_y(rectangle2_ys[735]), .rectangle2_width(rectangle2_widths[735]), .rectangle2_height(rectangle2_heights[735]), .rectangle2_weight(rectangle2_weights[735]), .rectangle3_x(rectangle3_xs[735]), .rectangle3_y(rectangle3_ys[735]), .rectangle3_width(rectangle3_widths[735]), .rectangle3_height(rectangle3_heights[735]), .rectangle3_weight(rectangle3_weights[735]), .feature_threshold(feature_thresholds[735]), .feature_above(feature_aboves[735]), .feature_below(feature_belows[735]), .scan_win_std_dev(scan_win_std_dev[735]), .feature_accum(feature_accums[735]));
  accum_calculator ac736(.scan_win(scan_win736), .rectangle1_x(rectangle1_xs[736]), .rectangle1_y(rectangle1_ys[736]), .rectangle1_width(rectangle1_widths[736]), .rectangle1_height(rectangle1_heights[736]), .rectangle1_weight(rectangle1_weights[736]), .rectangle2_x(rectangle2_xs[736]), .rectangle2_y(rectangle2_ys[736]), .rectangle2_width(rectangle2_widths[736]), .rectangle2_height(rectangle2_heights[736]), .rectangle2_weight(rectangle2_weights[736]), .rectangle3_x(rectangle3_xs[736]), .rectangle3_y(rectangle3_ys[736]), .rectangle3_width(rectangle3_widths[736]), .rectangle3_height(rectangle3_heights[736]), .rectangle3_weight(rectangle3_weights[736]), .feature_threshold(feature_thresholds[736]), .feature_above(feature_aboves[736]), .feature_below(feature_belows[736]), .scan_win_std_dev(scan_win_std_dev[736]), .feature_accum(feature_accums[736]));
  accum_calculator ac737(.scan_win(scan_win737), .rectangle1_x(rectangle1_xs[737]), .rectangle1_y(rectangle1_ys[737]), .rectangle1_width(rectangle1_widths[737]), .rectangle1_height(rectangle1_heights[737]), .rectangle1_weight(rectangle1_weights[737]), .rectangle2_x(rectangle2_xs[737]), .rectangle2_y(rectangle2_ys[737]), .rectangle2_width(rectangle2_widths[737]), .rectangle2_height(rectangle2_heights[737]), .rectangle2_weight(rectangle2_weights[737]), .rectangle3_x(rectangle3_xs[737]), .rectangle3_y(rectangle3_ys[737]), .rectangle3_width(rectangle3_widths[737]), .rectangle3_height(rectangle3_heights[737]), .rectangle3_weight(rectangle3_weights[737]), .feature_threshold(feature_thresholds[737]), .feature_above(feature_aboves[737]), .feature_below(feature_belows[737]), .scan_win_std_dev(scan_win_std_dev[737]), .feature_accum(feature_accums[737]));
  accum_calculator ac738(.scan_win(scan_win738), .rectangle1_x(rectangle1_xs[738]), .rectangle1_y(rectangle1_ys[738]), .rectangle1_width(rectangle1_widths[738]), .rectangle1_height(rectangle1_heights[738]), .rectangle1_weight(rectangle1_weights[738]), .rectangle2_x(rectangle2_xs[738]), .rectangle2_y(rectangle2_ys[738]), .rectangle2_width(rectangle2_widths[738]), .rectangle2_height(rectangle2_heights[738]), .rectangle2_weight(rectangle2_weights[738]), .rectangle3_x(rectangle3_xs[738]), .rectangle3_y(rectangle3_ys[738]), .rectangle3_width(rectangle3_widths[738]), .rectangle3_height(rectangle3_heights[738]), .rectangle3_weight(rectangle3_weights[738]), .feature_threshold(feature_thresholds[738]), .feature_above(feature_aboves[738]), .feature_below(feature_belows[738]), .scan_win_std_dev(scan_win_std_dev[738]), .feature_accum(feature_accums[738]));
  accum_calculator ac739(.scan_win(scan_win739), .rectangle1_x(rectangle1_xs[739]), .rectangle1_y(rectangle1_ys[739]), .rectangle1_width(rectangle1_widths[739]), .rectangle1_height(rectangle1_heights[739]), .rectangle1_weight(rectangle1_weights[739]), .rectangle2_x(rectangle2_xs[739]), .rectangle2_y(rectangle2_ys[739]), .rectangle2_width(rectangle2_widths[739]), .rectangle2_height(rectangle2_heights[739]), .rectangle2_weight(rectangle2_weights[739]), .rectangle3_x(rectangle3_xs[739]), .rectangle3_y(rectangle3_ys[739]), .rectangle3_width(rectangle3_widths[739]), .rectangle3_height(rectangle3_heights[739]), .rectangle3_weight(rectangle3_weights[739]), .feature_threshold(feature_thresholds[739]), .feature_above(feature_aboves[739]), .feature_below(feature_belows[739]), .scan_win_std_dev(scan_win_std_dev[739]), .feature_accum(feature_accums[739]));
  accum_calculator ac740(.scan_win(scan_win740), .rectangle1_x(rectangle1_xs[740]), .rectangle1_y(rectangle1_ys[740]), .rectangle1_width(rectangle1_widths[740]), .rectangle1_height(rectangle1_heights[740]), .rectangle1_weight(rectangle1_weights[740]), .rectangle2_x(rectangle2_xs[740]), .rectangle2_y(rectangle2_ys[740]), .rectangle2_width(rectangle2_widths[740]), .rectangle2_height(rectangle2_heights[740]), .rectangle2_weight(rectangle2_weights[740]), .rectangle3_x(rectangle3_xs[740]), .rectangle3_y(rectangle3_ys[740]), .rectangle3_width(rectangle3_widths[740]), .rectangle3_height(rectangle3_heights[740]), .rectangle3_weight(rectangle3_weights[740]), .feature_threshold(feature_thresholds[740]), .feature_above(feature_aboves[740]), .feature_below(feature_belows[740]), .scan_win_std_dev(scan_win_std_dev[740]), .feature_accum(feature_accums[740]));
  accum_calculator ac741(.scan_win(scan_win741), .rectangle1_x(rectangle1_xs[741]), .rectangle1_y(rectangle1_ys[741]), .rectangle1_width(rectangle1_widths[741]), .rectangle1_height(rectangle1_heights[741]), .rectangle1_weight(rectangle1_weights[741]), .rectangle2_x(rectangle2_xs[741]), .rectangle2_y(rectangle2_ys[741]), .rectangle2_width(rectangle2_widths[741]), .rectangle2_height(rectangle2_heights[741]), .rectangle2_weight(rectangle2_weights[741]), .rectangle3_x(rectangle3_xs[741]), .rectangle3_y(rectangle3_ys[741]), .rectangle3_width(rectangle3_widths[741]), .rectangle3_height(rectangle3_heights[741]), .rectangle3_weight(rectangle3_weights[741]), .feature_threshold(feature_thresholds[741]), .feature_above(feature_aboves[741]), .feature_below(feature_belows[741]), .scan_win_std_dev(scan_win_std_dev[741]), .feature_accum(feature_accums[741]));
  accum_calculator ac742(.scan_win(scan_win742), .rectangle1_x(rectangle1_xs[742]), .rectangle1_y(rectangle1_ys[742]), .rectangle1_width(rectangle1_widths[742]), .rectangle1_height(rectangle1_heights[742]), .rectangle1_weight(rectangle1_weights[742]), .rectangle2_x(rectangle2_xs[742]), .rectangle2_y(rectangle2_ys[742]), .rectangle2_width(rectangle2_widths[742]), .rectangle2_height(rectangle2_heights[742]), .rectangle2_weight(rectangle2_weights[742]), .rectangle3_x(rectangle3_xs[742]), .rectangle3_y(rectangle3_ys[742]), .rectangle3_width(rectangle3_widths[742]), .rectangle3_height(rectangle3_heights[742]), .rectangle3_weight(rectangle3_weights[742]), .feature_threshold(feature_thresholds[742]), .feature_above(feature_aboves[742]), .feature_below(feature_belows[742]), .scan_win_std_dev(scan_win_std_dev[742]), .feature_accum(feature_accums[742]));
  accum_calculator ac743(.scan_win(scan_win743), .rectangle1_x(rectangle1_xs[743]), .rectangle1_y(rectangle1_ys[743]), .rectangle1_width(rectangle1_widths[743]), .rectangle1_height(rectangle1_heights[743]), .rectangle1_weight(rectangle1_weights[743]), .rectangle2_x(rectangle2_xs[743]), .rectangle2_y(rectangle2_ys[743]), .rectangle2_width(rectangle2_widths[743]), .rectangle2_height(rectangle2_heights[743]), .rectangle2_weight(rectangle2_weights[743]), .rectangle3_x(rectangle3_xs[743]), .rectangle3_y(rectangle3_ys[743]), .rectangle3_width(rectangle3_widths[743]), .rectangle3_height(rectangle3_heights[743]), .rectangle3_weight(rectangle3_weights[743]), .feature_threshold(feature_thresholds[743]), .feature_above(feature_aboves[743]), .feature_below(feature_belows[743]), .scan_win_std_dev(scan_win_std_dev[743]), .feature_accum(feature_accums[743]));
  accum_calculator ac744(.scan_win(scan_win744), .rectangle1_x(rectangle1_xs[744]), .rectangle1_y(rectangle1_ys[744]), .rectangle1_width(rectangle1_widths[744]), .rectangle1_height(rectangle1_heights[744]), .rectangle1_weight(rectangle1_weights[744]), .rectangle2_x(rectangle2_xs[744]), .rectangle2_y(rectangle2_ys[744]), .rectangle2_width(rectangle2_widths[744]), .rectangle2_height(rectangle2_heights[744]), .rectangle2_weight(rectangle2_weights[744]), .rectangle3_x(rectangle3_xs[744]), .rectangle3_y(rectangle3_ys[744]), .rectangle3_width(rectangle3_widths[744]), .rectangle3_height(rectangle3_heights[744]), .rectangle3_weight(rectangle3_weights[744]), .feature_threshold(feature_thresholds[744]), .feature_above(feature_aboves[744]), .feature_below(feature_belows[744]), .scan_win_std_dev(scan_win_std_dev[744]), .feature_accum(feature_accums[744]));
  accum_calculator ac745(.scan_win(scan_win745), .rectangle1_x(rectangle1_xs[745]), .rectangle1_y(rectangle1_ys[745]), .rectangle1_width(rectangle1_widths[745]), .rectangle1_height(rectangle1_heights[745]), .rectangle1_weight(rectangle1_weights[745]), .rectangle2_x(rectangle2_xs[745]), .rectangle2_y(rectangle2_ys[745]), .rectangle2_width(rectangle2_widths[745]), .rectangle2_height(rectangle2_heights[745]), .rectangle2_weight(rectangle2_weights[745]), .rectangle3_x(rectangle3_xs[745]), .rectangle3_y(rectangle3_ys[745]), .rectangle3_width(rectangle3_widths[745]), .rectangle3_height(rectangle3_heights[745]), .rectangle3_weight(rectangle3_weights[745]), .feature_threshold(feature_thresholds[745]), .feature_above(feature_aboves[745]), .feature_below(feature_belows[745]), .scan_win_std_dev(scan_win_std_dev[745]), .feature_accum(feature_accums[745]));
  accum_calculator ac746(.scan_win(scan_win746), .rectangle1_x(rectangle1_xs[746]), .rectangle1_y(rectangle1_ys[746]), .rectangle1_width(rectangle1_widths[746]), .rectangle1_height(rectangle1_heights[746]), .rectangle1_weight(rectangle1_weights[746]), .rectangle2_x(rectangle2_xs[746]), .rectangle2_y(rectangle2_ys[746]), .rectangle2_width(rectangle2_widths[746]), .rectangle2_height(rectangle2_heights[746]), .rectangle2_weight(rectangle2_weights[746]), .rectangle3_x(rectangle3_xs[746]), .rectangle3_y(rectangle3_ys[746]), .rectangle3_width(rectangle3_widths[746]), .rectangle3_height(rectangle3_heights[746]), .rectangle3_weight(rectangle3_weights[746]), .feature_threshold(feature_thresholds[746]), .feature_above(feature_aboves[746]), .feature_below(feature_belows[746]), .scan_win_std_dev(scan_win_std_dev[746]), .feature_accum(feature_accums[746]));
  accum_calculator ac747(.scan_win(scan_win747), .rectangle1_x(rectangle1_xs[747]), .rectangle1_y(rectangle1_ys[747]), .rectangle1_width(rectangle1_widths[747]), .rectangle1_height(rectangle1_heights[747]), .rectangle1_weight(rectangle1_weights[747]), .rectangle2_x(rectangle2_xs[747]), .rectangle2_y(rectangle2_ys[747]), .rectangle2_width(rectangle2_widths[747]), .rectangle2_height(rectangle2_heights[747]), .rectangle2_weight(rectangle2_weights[747]), .rectangle3_x(rectangle3_xs[747]), .rectangle3_y(rectangle3_ys[747]), .rectangle3_width(rectangle3_widths[747]), .rectangle3_height(rectangle3_heights[747]), .rectangle3_weight(rectangle3_weights[747]), .feature_threshold(feature_thresholds[747]), .feature_above(feature_aboves[747]), .feature_below(feature_belows[747]), .scan_win_std_dev(scan_win_std_dev[747]), .feature_accum(feature_accums[747]));
  accum_calculator ac748(.scan_win(scan_win748), .rectangle1_x(rectangle1_xs[748]), .rectangle1_y(rectangle1_ys[748]), .rectangle1_width(rectangle1_widths[748]), .rectangle1_height(rectangle1_heights[748]), .rectangle1_weight(rectangle1_weights[748]), .rectangle2_x(rectangle2_xs[748]), .rectangle2_y(rectangle2_ys[748]), .rectangle2_width(rectangle2_widths[748]), .rectangle2_height(rectangle2_heights[748]), .rectangle2_weight(rectangle2_weights[748]), .rectangle3_x(rectangle3_xs[748]), .rectangle3_y(rectangle3_ys[748]), .rectangle3_width(rectangle3_widths[748]), .rectangle3_height(rectangle3_heights[748]), .rectangle3_weight(rectangle3_weights[748]), .feature_threshold(feature_thresholds[748]), .feature_above(feature_aboves[748]), .feature_below(feature_belows[748]), .scan_win_std_dev(scan_win_std_dev[748]), .feature_accum(feature_accums[748]));
  accum_calculator ac749(.scan_win(scan_win749), .rectangle1_x(rectangle1_xs[749]), .rectangle1_y(rectangle1_ys[749]), .rectangle1_width(rectangle1_widths[749]), .rectangle1_height(rectangle1_heights[749]), .rectangle1_weight(rectangle1_weights[749]), .rectangle2_x(rectangle2_xs[749]), .rectangle2_y(rectangle2_ys[749]), .rectangle2_width(rectangle2_widths[749]), .rectangle2_height(rectangle2_heights[749]), .rectangle2_weight(rectangle2_weights[749]), .rectangle3_x(rectangle3_xs[749]), .rectangle3_y(rectangle3_ys[749]), .rectangle3_width(rectangle3_widths[749]), .rectangle3_height(rectangle3_heights[749]), .rectangle3_weight(rectangle3_weights[749]), .feature_threshold(feature_thresholds[749]), .feature_above(feature_aboves[749]), .feature_below(feature_belows[749]), .scan_win_std_dev(scan_win_std_dev[749]), .feature_accum(feature_accums[749]));
  accum_calculator ac750(.scan_win(scan_win750), .rectangle1_x(rectangle1_xs[750]), .rectangle1_y(rectangle1_ys[750]), .rectangle1_width(rectangle1_widths[750]), .rectangle1_height(rectangle1_heights[750]), .rectangle1_weight(rectangle1_weights[750]), .rectangle2_x(rectangle2_xs[750]), .rectangle2_y(rectangle2_ys[750]), .rectangle2_width(rectangle2_widths[750]), .rectangle2_height(rectangle2_heights[750]), .rectangle2_weight(rectangle2_weights[750]), .rectangle3_x(rectangle3_xs[750]), .rectangle3_y(rectangle3_ys[750]), .rectangle3_width(rectangle3_widths[750]), .rectangle3_height(rectangle3_heights[750]), .rectangle3_weight(rectangle3_weights[750]), .feature_threshold(feature_thresholds[750]), .feature_above(feature_aboves[750]), .feature_below(feature_belows[750]), .scan_win_std_dev(scan_win_std_dev[750]), .feature_accum(feature_accums[750]));
  accum_calculator ac751(.scan_win(scan_win751), .rectangle1_x(rectangle1_xs[751]), .rectangle1_y(rectangle1_ys[751]), .rectangle1_width(rectangle1_widths[751]), .rectangle1_height(rectangle1_heights[751]), .rectangle1_weight(rectangle1_weights[751]), .rectangle2_x(rectangle2_xs[751]), .rectangle2_y(rectangle2_ys[751]), .rectangle2_width(rectangle2_widths[751]), .rectangle2_height(rectangle2_heights[751]), .rectangle2_weight(rectangle2_weights[751]), .rectangle3_x(rectangle3_xs[751]), .rectangle3_y(rectangle3_ys[751]), .rectangle3_width(rectangle3_widths[751]), .rectangle3_height(rectangle3_heights[751]), .rectangle3_weight(rectangle3_weights[751]), .feature_threshold(feature_thresholds[751]), .feature_above(feature_aboves[751]), .feature_below(feature_belows[751]), .scan_win_std_dev(scan_win_std_dev[751]), .feature_accum(feature_accums[751]));
  accum_calculator ac752(.scan_win(scan_win752), .rectangle1_x(rectangle1_xs[752]), .rectangle1_y(rectangle1_ys[752]), .rectangle1_width(rectangle1_widths[752]), .rectangle1_height(rectangle1_heights[752]), .rectangle1_weight(rectangle1_weights[752]), .rectangle2_x(rectangle2_xs[752]), .rectangle2_y(rectangle2_ys[752]), .rectangle2_width(rectangle2_widths[752]), .rectangle2_height(rectangle2_heights[752]), .rectangle2_weight(rectangle2_weights[752]), .rectangle3_x(rectangle3_xs[752]), .rectangle3_y(rectangle3_ys[752]), .rectangle3_width(rectangle3_widths[752]), .rectangle3_height(rectangle3_heights[752]), .rectangle3_weight(rectangle3_weights[752]), .feature_threshold(feature_thresholds[752]), .feature_above(feature_aboves[752]), .feature_below(feature_belows[752]), .scan_win_std_dev(scan_win_std_dev[752]), .feature_accum(feature_accums[752]));
  accum_calculator ac753(.scan_win(scan_win753), .rectangle1_x(rectangle1_xs[753]), .rectangle1_y(rectangle1_ys[753]), .rectangle1_width(rectangle1_widths[753]), .rectangle1_height(rectangle1_heights[753]), .rectangle1_weight(rectangle1_weights[753]), .rectangle2_x(rectangle2_xs[753]), .rectangle2_y(rectangle2_ys[753]), .rectangle2_width(rectangle2_widths[753]), .rectangle2_height(rectangle2_heights[753]), .rectangle2_weight(rectangle2_weights[753]), .rectangle3_x(rectangle3_xs[753]), .rectangle3_y(rectangle3_ys[753]), .rectangle3_width(rectangle3_widths[753]), .rectangle3_height(rectangle3_heights[753]), .rectangle3_weight(rectangle3_weights[753]), .feature_threshold(feature_thresholds[753]), .feature_above(feature_aboves[753]), .feature_below(feature_belows[753]), .scan_win_std_dev(scan_win_std_dev[753]), .feature_accum(feature_accums[753]));
  accum_calculator ac754(.scan_win(scan_win754), .rectangle1_x(rectangle1_xs[754]), .rectangle1_y(rectangle1_ys[754]), .rectangle1_width(rectangle1_widths[754]), .rectangle1_height(rectangle1_heights[754]), .rectangle1_weight(rectangle1_weights[754]), .rectangle2_x(rectangle2_xs[754]), .rectangle2_y(rectangle2_ys[754]), .rectangle2_width(rectangle2_widths[754]), .rectangle2_height(rectangle2_heights[754]), .rectangle2_weight(rectangle2_weights[754]), .rectangle3_x(rectangle3_xs[754]), .rectangle3_y(rectangle3_ys[754]), .rectangle3_width(rectangle3_widths[754]), .rectangle3_height(rectangle3_heights[754]), .rectangle3_weight(rectangle3_weights[754]), .feature_threshold(feature_thresholds[754]), .feature_above(feature_aboves[754]), .feature_below(feature_belows[754]), .scan_win_std_dev(scan_win_std_dev[754]), .feature_accum(feature_accums[754]));
  accum_calculator ac755(.scan_win(scan_win755), .rectangle1_x(rectangle1_xs[755]), .rectangle1_y(rectangle1_ys[755]), .rectangle1_width(rectangle1_widths[755]), .rectangle1_height(rectangle1_heights[755]), .rectangle1_weight(rectangle1_weights[755]), .rectangle2_x(rectangle2_xs[755]), .rectangle2_y(rectangle2_ys[755]), .rectangle2_width(rectangle2_widths[755]), .rectangle2_height(rectangle2_heights[755]), .rectangle2_weight(rectangle2_weights[755]), .rectangle3_x(rectangle3_xs[755]), .rectangle3_y(rectangle3_ys[755]), .rectangle3_width(rectangle3_widths[755]), .rectangle3_height(rectangle3_heights[755]), .rectangle3_weight(rectangle3_weights[755]), .feature_threshold(feature_thresholds[755]), .feature_above(feature_aboves[755]), .feature_below(feature_belows[755]), .scan_win_std_dev(scan_win_std_dev[755]), .feature_accum(feature_accums[755]));
  accum_calculator ac756(.scan_win(scan_win756), .rectangle1_x(rectangle1_xs[756]), .rectangle1_y(rectangle1_ys[756]), .rectangle1_width(rectangle1_widths[756]), .rectangle1_height(rectangle1_heights[756]), .rectangle1_weight(rectangle1_weights[756]), .rectangle2_x(rectangle2_xs[756]), .rectangle2_y(rectangle2_ys[756]), .rectangle2_width(rectangle2_widths[756]), .rectangle2_height(rectangle2_heights[756]), .rectangle2_weight(rectangle2_weights[756]), .rectangle3_x(rectangle3_xs[756]), .rectangle3_y(rectangle3_ys[756]), .rectangle3_width(rectangle3_widths[756]), .rectangle3_height(rectangle3_heights[756]), .rectangle3_weight(rectangle3_weights[756]), .feature_threshold(feature_thresholds[756]), .feature_above(feature_aboves[756]), .feature_below(feature_belows[756]), .scan_win_std_dev(scan_win_std_dev[756]), .feature_accum(feature_accums[756]));
  accum_calculator ac757(.scan_win(scan_win757), .rectangle1_x(rectangle1_xs[757]), .rectangle1_y(rectangle1_ys[757]), .rectangle1_width(rectangle1_widths[757]), .rectangle1_height(rectangle1_heights[757]), .rectangle1_weight(rectangle1_weights[757]), .rectangle2_x(rectangle2_xs[757]), .rectangle2_y(rectangle2_ys[757]), .rectangle2_width(rectangle2_widths[757]), .rectangle2_height(rectangle2_heights[757]), .rectangle2_weight(rectangle2_weights[757]), .rectangle3_x(rectangle3_xs[757]), .rectangle3_y(rectangle3_ys[757]), .rectangle3_width(rectangle3_widths[757]), .rectangle3_height(rectangle3_heights[757]), .rectangle3_weight(rectangle3_weights[757]), .feature_threshold(feature_thresholds[757]), .feature_above(feature_aboves[757]), .feature_below(feature_belows[757]), .scan_win_std_dev(scan_win_std_dev[757]), .feature_accum(feature_accums[757]));
  accum_calculator ac758(.scan_win(scan_win758), .rectangle1_x(rectangle1_xs[758]), .rectangle1_y(rectangle1_ys[758]), .rectangle1_width(rectangle1_widths[758]), .rectangle1_height(rectangle1_heights[758]), .rectangle1_weight(rectangle1_weights[758]), .rectangle2_x(rectangle2_xs[758]), .rectangle2_y(rectangle2_ys[758]), .rectangle2_width(rectangle2_widths[758]), .rectangle2_height(rectangle2_heights[758]), .rectangle2_weight(rectangle2_weights[758]), .rectangle3_x(rectangle3_xs[758]), .rectangle3_y(rectangle3_ys[758]), .rectangle3_width(rectangle3_widths[758]), .rectangle3_height(rectangle3_heights[758]), .rectangle3_weight(rectangle3_weights[758]), .feature_threshold(feature_thresholds[758]), .feature_above(feature_aboves[758]), .feature_below(feature_belows[758]), .scan_win_std_dev(scan_win_std_dev[758]), .feature_accum(feature_accums[758]));
  accum_calculator ac759(.scan_win(scan_win759), .rectangle1_x(rectangle1_xs[759]), .rectangle1_y(rectangle1_ys[759]), .rectangle1_width(rectangle1_widths[759]), .rectangle1_height(rectangle1_heights[759]), .rectangle1_weight(rectangle1_weights[759]), .rectangle2_x(rectangle2_xs[759]), .rectangle2_y(rectangle2_ys[759]), .rectangle2_width(rectangle2_widths[759]), .rectangle2_height(rectangle2_heights[759]), .rectangle2_weight(rectangle2_weights[759]), .rectangle3_x(rectangle3_xs[759]), .rectangle3_y(rectangle3_ys[759]), .rectangle3_width(rectangle3_widths[759]), .rectangle3_height(rectangle3_heights[759]), .rectangle3_weight(rectangle3_weights[759]), .feature_threshold(feature_thresholds[759]), .feature_above(feature_aboves[759]), .feature_below(feature_belows[759]), .scan_win_std_dev(scan_win_std_dev[759]), .feature_accum(feature_accums[759]));
  accum_calculator ac760(.scan_win(scan_win760), .rectangle1_x(rectangle1_xs[760]), .rectangle1_y(rectangle1_ys[760]), .rectangle1_width(rectangle1_widths[760]), .rectangle1_height(rectangle1_heights[760]), .rectangle1_weight(rectangle1_weights[760]), .rectangle2_x(rectangle2_xs[760]), .rectangle2_y(rectangle2_ys[760]), .rectangle2_width(rectangle2_widths[760]), .rectangle2_height(rectangle2_heights[760]), .rectangle2_weight(rectangle2_weights[760]), .rectangle3_x(rectangle3_xs[760]), .rectangle3_y(rectangle3_ys[760]), .rectangle3_width(rectangle3_widths[760]), .rectangle3_height(rectangle3_heights[760]), .rectangle3_weight(rectangle3_weights[760]), .feature_threshold(feature_thresholds[760]), .feature_above(feature_aboves[760]), .feature_below(feature_belows[760]), .scan_win_std_dev(scan_win_std_dev[760]), .feature_accum(feature_accums[760]));
  accum_calculator ac761(.scan_win(scan_win761), .rectangle1_x(rectangle1_xs[761]), .rectangle1_y(rectangle1_ys[761]), .rectangle1_width(rectangle1_widths[761]), .rectangle1_height(rectangle1_heights[761]), .rectangle1_weight(rectangle1_weights[761]), .rectangle2_x(rectangle2_xs[761]), .rectangle2_y(rectangle2_ys[761]), .rectangle2_width(rectangle2_widths[761]), .rectangle2_height(rectangle2_heights[761]), .rectangle2_weight(rectangle2_weights[761]), .rectangle3_x(rectangle3_xs[761]), .rectangle3_y(rectangle3_ys[761]), .rectangle3_width(rectangle3_widths[761]), .rectangle3_height(rectangle3_heights[761]), .rectangle3_weight(rectangle3_weights[761]), .feature_threshold(feature_thresholds[761]), .feature_above(feature_aboves[761]), .feature_below(feature_belows[761]), .scan_win_std_dev(scan_win_std_dev[761]), .feature_accum(feature_accums[761]));
  accum_calculator ac762(.scan_win(scan_win762), .rectangle1_x(rectangle1_xs[762]), .rectangle1_y(rectangle1_ys[762]), .rectangle1_width(rectangle1_widths[762]), .rectangle1_height(rectangle1_heights[762]), .rectangle1_weight(rectangle1_weights[762]), .rectangle2_x(rectangle2_xs[762]), .rectangle2_y(rectangle2_ys[762]), .rectangle2_width(rectangle2_widths[762]), .rectangle2_height(rectangle2_heights[762]), .rectangle2_weight(rectangle2_weights[762]), .rectangle3_x(rectangle3_xs[762]), .rectangle3_y(rectangle3_ys[762]), .rectangle3_width(rectangle3_widths[762]), .rectangle3_height(rectangle3_heights[762]), .rectangle3_weight(rectangle3_weights[762]), .feature_threshold(feature_thresholds[762]), .feature_above(feature_aboves[762]), .feature_below(feature_belows[762]), .scan_win_std_dev(scan_win_std_dev[762]), .feature_accum(feature_accums[762]));
  accum_calculator ac763(.scan_win(scan_win763), .rectangle1_x(rectangle1_xs[763]), .rectangle1_y(rectangle1_ys[763]), .rectangle1_width(rectangle1_widths[763]), .rectangle1_height(rectangle1_heights[763]), .rectangle1_weight(rectangle1_weights[763]), .rectangle2_x(rectangle2_xs[763]), .rectangle2_y(rectangle2_ys[763]), .rectangle2_width(rectangle2_widths[763]), .rectangle2_height(rectangle2_heights[763]), .rectangle2_weight(rectangle2_weights[763]), .rectangle3_x(rectangle3_xs[763]), .rectangle3_y(rectangle3_ys[763]), .rectangle3_width(rectangle3_widths[763]), .rectangle3_height(rectangle3_heights[763]), .rectangle3_weight(rectangle3_weights[763]), .feature_threshold(feature_thresholds[763]), .feature_above(feature_aboves[763]), .feature_below(feature_belows[763]), .scan_win_std_dev(scan_win_std_dev[763]), .feature_accum(feature_accums[763]));
  accum_calculator ac764(.scan_win(scan_win764), .rectangle1_x(rectangle1_xs[764]), .rectangle1_y(rectangle1_ys[764]), .rectangle1_width(rectangle1_widths[764]), .rectangle1_height(rectangle1_heights[764]), .rectangle1_weight(rectangle1_weights[764]), .rectangle2_x(rectangle2_xs[764]), .rectangle2_y(rectangle2_ys[764]), .rectangle2_width(rectangle2_widths[764]), .rectangle2_height(rectangle2_heights[764]), .rectangle2_weight(rectangle2_weights[764]), .rectangle3_x(rectangle3_xs[764]), .rectangle3_y(rectangle3_ys[764]), .rectangle3_width(rectangle3_widths[764]), .rectangle3_height(rectangle3_heights[764]), .rectangle3_weight(rectangle3_weights[764]), .feature_threshold(feature_thresholds[764]), .feature_above(feature_aboves[764]), .feature_below(feature_belows[764]), .scan_win_std_dev(scan_win_std_dev[764]), .feature_accum(feature_accums[764]));
  accum_calculator ac765(.scan_win(scan_win765), .rectangle1_x(rectangle1_xs[765]), .rectangle1_y(rectangle1_ys[765]), .rectangle1_width(rectangle1_widths[765]), .rectangle1_height(rectangle1_heights[765]), .rectangle1_weight(rectangle1_weights[765]), .rectangle2_x(rectangle2_xs[765]), .rectangle2_y(rectangle2_ys[765]), .rectangle2_width(rectangle2_widths[765]), .rectangle2_height(rectangle2_heights[765]), .rectangle2_weight(rectangle2_weights[765]), .rectangle3_x(rectangle3_xs[765]), .rectangle3_y(rectangle3_ys[765]), .rectangle3_width(rectangle3_widths[765]), .rectangle3_height(rectangle3_heights[765]), .rectangle3_weight(rectangle3_weights[765]), .feature_threshold(feature_thresholds[765]), .feature_above(feature_aboves[765]), .feature_below(feature_belows[765]), .scan_win_std_dev(scan_win_std_dev[765]), .feature_accum(feature_accums[765]));
  accum_calculator ac766(.scan_win(scan_win766), .rectangle1_x(rectangle1_xs[766]), .rectangle1_y(rectangle1_ys[766]), .rectangle1_width(rectangle1_widths[766]), .rectangle1_height(rectangle1_heights[766]), .rectangle1_weight(rectangle1_weights[766]), .rectangle2_x(rectangle2_xs[766]), .rectangle2_y(rectangle2_ys[766]), .rectangle2_width(rectangle2_widths[766]), .rectangle2_height(rectangle2_heights[766]), .rectangle2_weight(rectangle2_weights[766]), .rectangle3_x(rectangle3_xs[766]), .rectangle3_y(rectangle3_ys[766]), .rectangle3_width(rectangle3_widths[766]), .rectangle3_height(rectangle3_heights[766]), .rectangle3_weight(rectangle3_weights[766]), .feature_threshold(feature_thresholds[766]), .feature_above(feature_aboves[766]), .feature_below(feature_belows[766]), .scan_win_std_dev(scan_win_std_dev[766]), .feature_accum(feature_accums[766]));
  accum_calculator ac767(.scan_win(scan_win767), .rectangle1_x(rectangle1_xs[767]), .rectangle1_y(rectangle1_ys[767]), .rectangle1_width(rectangle1_widths[767]), .rectangle1_height(rectangle1_heights[767]), .rectangle1_weight(rectangle1_weights[767]), .rectangle2_x(rectangle2_xs[767]), .rectangle2_y(rectangle2_ys[767]), .rectangle2_width(rectangle2_widths[767]), .rectangle2_height(rectangle2_heights[767]), .rectangle2_weight(rectangle2_weights[767]), .rectangle3_x(rectangle3_xs[767]), .rectangle3_y(rectangle3_ys[767]), .rectangle3_width(rectangle3_widths[767]), .rectangle3_height(rectangle3_heights[767]), .rectangle3_weight(rectangle3_weights[767]), .feature_threshold(feature_thresholds[767]), .feature_above(feature_aboves[767]), .feature_below(feature_belows[767]), .scan_win_std_dev(scan_win_std_dev[767]), .feature_accum(feature_accums[767]));
  accum_calculator ac768(.scan_win(scan_win768), .rectangle1_x(rectangle1_xs[768]), .rectangle1_y(rectangle1_ys[768]), .rectangle1_width(rectangle1_widths[768]), .rectangle1_height(rectangle1_heights[768]), .rectangle1_weight(rectangle1_weights[768]), .rectangle2_x(rectangle2_xs[768]), .rectangle2_y(rectangle2_ys[768]), .rectangle2_width(rectangle2_widths[768]), .rectangle2_height(rectangle2_heights[768]), .rectangle2_weight(rectangle2_weights[768]), .rectangle3_x(rectangle3_xs[768]), .rectangle3_y(rectangle3_ys[768]), .rectangle3_width(rectangle3_widths[768]), .rectangle3_height(rectangle3_heights[768]), .rectangle3_weight(rectangle3_weights[768]), .feature_threshold(feature_thresholds[768]), .feature_above(feature_aboves[768]), .feature_below(feature_belows[768]), .scan_win_std_dev(scan_win_std_dev[768]), .feature_accum(feature_accums[768]));
  accum_calculator ac769(.scan_win(scan_win769), .rectangle1_x(rectangle1_xs[769]), .rectangle1_y(rectangle1_ys[769]), .rectangle1_width(rectangle1_widths[769]), .rectangle1_height(rectangle1_heights[769]), .rectangle1_weight(rectangle1_weights[769]), .rectangle2_x(rectangle2_xs[769]), .rectangle2_y(rectangle2_ys[769]), .rectangle2_width(rectangle2_widths[769]), .rectangle2_height(rectangle2_heights[769]), .rectangle2_weight(rectangle2_weights[769]), .rectangle3_x(rectangle3_xs[769]), .rectangle3_y(rectangle3_ys[769]), .rectangle3_width(rectangle3_widths[769]), .rectangle3_height(rectangle3_heights[769]), .rectangle3_weight(rectangle3_weights[769]), .feature_threshold(feature_thresholds[769]), .feature_above(feature_aboves[769]), .feature_below(feature_belows[769]), .scan_win_std_dev(scan_win_std_dev[769]), .feature_accum(feature_accums[769]));
  accum_calculator ac770(.scan_win(scan_win770), .rectangle1_x(rectangle1_xs[770]), .rectangle1_y(rectangle1_ys[770]), .rectangle1_width(rectangle1_widths[770]), .rectangle1_height(rectangle1_heights[770]), .rectangle1_weight(rectangle1_weights[770]), .rectangle2_x(rectangle2_xs[770]), .rectangle2_y(rectangle2_ys[770]), .rectangle2_width(rectangle2_widths[770]), .rectangle2_height(rectangle2_heights[770]), .rectangle2_weight(rectangle2_weights[770]), .rectangle3_x(rectangle3_xs[770]), .rectangle3_y(rectangle3_ys[770]), .rectangle3_width(rectangle3_widths[770]), .rectangle3_height(rectangle3_heights[770]), .rectangle3_weight(rectangle3_weights[770]), .feature_threshold(feature_thresholds[770]), .feature_above(feature_aboves[770]), .feature_below(feature_belows[770]), .scan_win_std_dev(scan_win_std_dev[770]), .feature_accum(feature_accums[770]));
  accum_calculator ac771(.scan_win(scan_win771), .rectangle1_x(rectangle1_xs[771]), .rectangle1_y(rectangle1_ys[771]), .rectangle1_width(rectangle1_widths[771]), .rectangle1_height(rectangle1_heights[771]), .rectangle1_weight(rectangle1_weights[771]), .rectangle2_x(rectangle2_xs[771]), .rectangle2_y(rectangle2_ys[771]), .rectangle2_width(rectangle2_widths[771]), .rectangle2_height(rectangle2_heights[771]), .rectangle2_weight(rectangle2_weights[771]), .rectangle3_x(rectangle3_xs[771]), .rectangle3_y(rectangle3_ys[771]), .rectangle3_width(rectangle3_widths[771]), .rectangle3_height(rectangle3_heights[771]), .rectangle3_weight(rectangle3_weights[771]), .feature_threshold(feature_thresholds[771]), .feature_above(feature_aboves[771]), .feature_below(feature_belows[771]), .scan_win_std_dev(scan_win_std_dev[771]), .feature_accum(feature_accums[771]));
  accum_calculator ac772(.scan_win(scan_win772), .rectangle1_x(rectangle1_xs[772]), .rectangle1_y(rectangle1_ys[772]), .rectangle1_width(rectangle1_widths[772]), .rectangle1_height(rectangle1_heights[772]), .rectangle1_weight(rectangle1_weights[772]), .rectangle2_x(rectangle2_xs[772]), .rectangle2_y(rectangle2_ys[772]), .rectangle2_width(rectangle2_widths[772]), .rectangle2_height(rectangle2_heights[772]), .rectangle2_weight(rectangle2_weights[772]), .rectangle3_x(rectangle3_xs[772]), .rectangle3_y(rectangle3_ys[772]), .rectangle3_width(rectangle3_widths[772]), .rectangle3_height(rectangle3_heights[772]), .rectangle3_weight(rectangle3_weights[772]), .feature_threshold(feature_thresholds[772]), .feature_above(feature_aboves[772]), .feature_below(feature_belows[772]), .scan_win_std_dev(scan_win_std_dev[772]), .feature_accum(feature_accums[772]));
  accum_calculator ac773(.scan_win(scan_win773), .rectangle1_x(rectangle1_xs[773]), .rectangle1_y(rectangle1_ys[773]), .rectangle1_width(rectangle1_widths[773]), .rectangle1_height(rectangle1_heights[773]), .rectangle1_weight(rectangle1_weights[773]), .rectangle2_x(rectangle2_xs[773]), .rectangle2_y(rectangle2_ys[773]), .rectangle2_width(rectangle2_widths[773]), .rectangle2_height(rectangle2_heights[773]), .rectangle2_weight(rectangle2_weights[773]), .rectangle3_x(rectangle3_xs[773]), .rectangle3_y(rectangle3_ys[773]), .rectangle3_width(rectangle3_widths[773]), .rectangle3_height(rectangle3_heights[773]), .rectangle3_weight(rectangle3_weights[773]), .feature_threshold(feature_thresholds[773]), .feature_above(feature_aboves[773]), .feature_below(feature_belows[773]), .scan_win_std_dev(scan_win_std_dev[773]), .feature_accum(feature_accums[773]));
  accum_calculator ac774(.scan_win(scan_win774), .rectangle1_x(rectangle1_xs[774]), .rectangle1_y(rectangle1_ys[774]), .rectangle1_width(rectangle1_widths[774]), .rectangle1_height(rectangle1_heights[774]), .rectangle1_weight(rectangle1_weights[774]), .rectangle2_x(rectangle2_xs[774]), .rectangle2_y(rectangle2_ys[774]), .rectangle2_width(rectangle2_widths[774]), .rectangle2_height(rectangle2_heights[774]), .rectangle2_weight(rectangle2_weights[774]), .rectangle3_x(rectangle3_xs[774]), .rectangle3_y(rectangle3_ys[774]), .rectangle3_width(rectangle3_widths[774]), .rectangle3_height(rectangle3_heights[774]), .rectangle3_weight(rectangle3_weights[774]), .feature_threshold(feature_thresholds[774]), .feature_above(feature_aboves[774]), .feature_below(feature_belows[774]), .scan_win_std_dev(scan_win_std_dev[774]), .feature_accum(feature_accums[774]));
  accum_calculator ac775(.scan_win(scan_win775), .rectangle1_x(rectangle1_xs[775]), .rectangle1_y(rectangle1_ys[775]), .rectangle1_width(rectangle1_widths[775]), .rectangle1_height(rectangle1_heights[775]), .rectangle1_weight(rectangle1_weights[775]), .rectangle2_x(rectangle2_xs[775]), .rectangle2_y(rectangle2_ys[775]), .rectangle2_width(rectangle2_widths[775]), .rectangle2_height(rectangle2_heights[775]), .rectangle2_weight(rectangle2_weights[775]), .rectangle3_x(rectangle3_xs[775]), .rectangle3_y(rectangle3_ys[775]), .rectangle3_width(rectangle3_widths[775]), .rectangle3_height(rectangle3_heights[775]), .rectangle3_weight(rectangle3_weights[775]), .feature_threshold(feature_thresholds[775]), .feature_above(feature_aboves[775]), .feature_below(feature_belows[775]), .scan_win_std_dev(scan_win_std_dev[775]), .feature_accum(feature_accums[775]));
  accum_calculator ac776(.scan_win(scan_win776), .rectangle1_x(rectangle1_xs[776]), .rectangle1_y(rectangle1_ys[776]), .rectangle1_width(rectangle1_widths[776]), .rectangle1_height(rectangle1_heights[776]), .rectangle1_weight(rectangle1_weights[776]), .rectangle2_x(rectangle2_xs[776]), .rectangle2_y(rectangle2_ys[776]), .rectangle2_width(rectangle2_widths[776]), .rectangle2_height(rectangle2_heights[776]), .rectangle2_weight(rectangle2_weights[776]), .rectangle3_x(rectangle3_xs[776]), .rectangle3_y(rectangle3_ys[776]), .rectangle3_width(rectangle3_widths[776]), .rectangle3_height(rectangle3_heights[776]), .rectangle3_weight(rectangle3_weights[776]), .feature_threshold(feature_thresholds[776]), .feature_above(feature_aboves[776]), .feature_below(feature_belows[776]), .scan_win_std_dev(scan_win_std_dev[776]), .feature_accum(feature_accums[776]));
  accum_calculator ac777(.scan_win(scan_win777), .rectangle1_x(rectangle1_xs[777]), .rectangle1_y(rectangle1_ys[777]), .rectangle1_width(rectangle1_widths[777]), .rectangle1_height(rectangle1_heights[777]), .rectangle1_weight(rectangle1_weights[777]), .rectangle2_x(rectangle2_xs[777]), .rectangle2_y(rectangle2_ys[777]), .rectangle2_width(rectangle2_widths[777]), .rectangle2_height(rectangle2_heights[777]), .rectangle2_weight(rectangle2_weights[777]), .rectangle3_x(rectangle3_xs[777]), .rectangle3_y(rectangle3_ys[777]), .rectangle3_width(rectangle3_widths[777]), .rectangle3_height(rectangle3_heights[777]), .rectangle3_weight(rectangle3_weights[777]), .feature_threshold(feature_thresholds[777]), .feature_above(feature_aboves[777]), .feature_below(feature_belows[777]), .scan_win_std_dev(scan_win_std_dev[777]), .feature_accum(feature_accums[777]));
  accum_calculator ac778(.scan_win(scan_win778), .rectangle1_x(rectangle1_xs[778]), .rectangle1_y(rectangle1_ys[778]), .rectangle1_width(rectangle1_widths[778]), .rectangle1_height(rectangle1_heights[778]), .rectangle1_weight(rectangle1_weights[778]), .rectangle2_x(rectangle2_xs[778]), .rectangle2_y(rectangle2_ys[778]), .rectangle2_width(rectangle2_widths[778]), .rectangle2_height(rectangle2_heights[778]), .rectangle2_weight(rectangle2_weights[778]), .rectangle3_x(rectangle3_xs[778]), .rectangle3_y(rectangle3_ys[778]), .rectangle3_width(rectangle3_widths[778]), .rectangle3_height(rectangle3_heights[778]), .rectangle3_weight(rectangle3_weights[778]), .feature_threshold(feature_thresholds[778]), .feature_above(feature_aboves[778]), .feature_below(feature_belows[778]), .scan_win_std_dev(scan_win_std_dev[778]), .feature_accum(feature_accums[778]));
  accum_calculator ac779(.scan_win(scan_win779), .rectangle1_x(rectangle1_xs[779]), .rectangle1_y(rectangle1_ys[779]), .rectangle1_width(rectangle1_widths[779]), .rectangle1_height(rectangle1_heights[779]), .rectangle1_weight(rectangle1_weights[779]), .rectangle2_x(rectangle2_xs[779]), .rectangle2_y(rectangle2_ys[779]), .rectangle2_width(rectangle2_widths[779]), .rectangle2_height(rectangle2_heights[779]), .rectangle2_weight(rectangle2_weights[779]), .rectangle3_x(rectangle3_xs[779]), .rectangle3_y(rectangle3_ys[779]), .rectangle3_width(rectangle3_widths[779]), .rectangle3_height(rectangle3_heights[779]), .rectangle3_weight(rectangle3_weights[779]), .feature_threshold(feature_thresholds[779]), .feature_above(feature_aboves[779]), .feature_below(feature_belows[779]), .scan_win_std_dev(scan_win_std_dev[779]), .feature_accum(feature_accums[779]));
  accum_calculator ac780(.scan_win(scan_win780), .rectangle1_x(rectangle1_xs[780]), .rectangle1_y(rectangle1_ys[780]), .rectangle1_width(rectangle1_widths[780]), .rectangle1_height(rectangle1_heights[780]), .rectangle1_weight(rectangle1_weights[780]), .rectangle2_x(rectangle2_xs[780]), .rectangle2_y(rectangle2_ys[780]), .rectangle2_width(rectangle2_widths[780]), .rectangle2_height(rectangle2_heights[780]), .rectangle2_weight(rectangle2_weights[780]), .rectangle3_x(rectangle3_xs[780]), .rectangle3_y(rectangle3_ys[780]), .rectangle3_width(rectangle3_widths[780]), .rectangle3_height(rectangle3_heights[780]), .rectangle3_weight(rectangle3_weights[780]), .feature_threshold(feature_thresholds[780]), .feature_above(feature_aboves[780]), .feature_below(feature_belows[780]), .scan_win_std_dev(scan_win_std_dev[780]), .feature_accum(feature_accums[780]));
  accum_calculator ac781(.scan_win(scan_win781), .rectangle1_x(rectangle1_xs[781]), .rectangle1_y(rectangle1_ys[781]), .rectangle1_width(rectangle1_widths[781]), .rectangle1_height(rectangle1_heights[781]), .rectangle1_weight(rectangle1_weights[781]), .rectangle2_x(rectangle2_xs[781]), .rectangle2_y(rectangle2_ys[781]), .rectangle2_width(rectangle2_widths[781]), .rectangle2_height(rectangle2_heights[781]), .rectangle2_weight(rectangle2_weights[781]), .rectangle3_x(rectangle3_xs[781]), .rectangle3_y(rectangle3_ys[781]), .rectangle3_width(rectangle3_widths[781]), .rectangle3_height(rectangle3_heights[781]), .rectangle3_weight(rectangle3_weights[781]), .feature_threshold(feature_thresholds[781]), .feature_above(feature_aboves[781]), .feature_below(feature_belows[781]), .scan_win_std_dev(scan_win_std_dev[781]), .feature_accum(feature_accums[781]));
  accum_calculator ac782(.scan_win(scan_win782), .rectangle1_x(rectangle1_xs[782]), .rectangle1_y(rectangle1_ys[782]), .rectangle1_width(rectangle1_widths[782]), .rectangle1_height(rectangle1_heights[782]), .rectangle1_weight(rectangle1_weights[782]), .rectangle2_x(rectangle2_xs[782]), .rectangle2_y(rectangle2_ys[782]), .rectangle2_width(rectangle2_widths[782]), .rectangle2_height(rectangle2_heights[782]), .rectangle2_weight(rectangle2_weights[782]), .rectangle3_x(rectangle3_xs[782]), .rectangle3_y(rectangle3_ys[782]), .rectangle3_width(rectangle3_widths[782]), .rectangle3_height(rectangle3_heights[782]), .rectangle3_weight(rectangle3_weights[782]), .feature_threshold(feature_thresholds[782]), .feature_above(feature_aboves[782]), .feature_below(feature_belows[782]), .scan_win_std_dev(scan_win_std_dev[782]), .feature_accum(feature_accums[782]));
  accum_calculator ac783(.scan_win(scan_win783), .rectangle1_x(rectangle1_xs[783]), .rectangle1_y(rectangle1_ys[783]), .rectangle1_width(rectangle1_widths[783]), .rectangle1_height(rectangle1_heights[783]), .rectangle1_weight(rectangle1_weights[783]), .rectangle2_x(rectangle2_xs[783]), .rectangle2_y(rectangle2_ys[783]), .rectangle2_width(rectangle2_widths[783]), .rectangle2_height(rectangle2_heights[783]), .rectangle2_weight(rectangle2_weights[783]), .rectangle3_x(rectangle3_xs[783]), .rectangle3_y(rectangle3_ys[783]), .rectangle3_width(rectangle3_widths[783]), .rectangle3_height(rectangle3_heights[783]), .rectangle3_weight(rectangle3_weights[783]), .feature_threshold(feature_thresholds[783]), .feature_above(feature_aboves[783]), .feature_below(feature_belows[783]), .scan_win_std_dev(scan_win_std_dev[783]), .feature_accum(feature_accums[783]));
  accum_calculator ac784(.scan_win(scan_win784), .rectangle1_x(rectangle1_xs[784]), .rectangle1_y(rectangle1_ys[784]), .rectangle1_width(rectangle1_widths[784]), .rectangle1_height(rectangle1_heights[784]), .rectangle1_weight(rectangle1_weights[784]), .rectangle2_x(rectangle2_xs[784]), .rectangle2_y(rectangle2_ys[784]), .rectangle2_width(rectangle2_widths[784]), .rectangle2_height(rectangle2_heights[784]), .rectangle2_weight(rectangle2_weights[784]), .rectangle3_x(rectangle3_xs[784]), .rectangle3_y(rectangle3_ys[784]), .rectangle3_width(rectangle3_widths[784]), .rectangle3_height(rectangle3_heights[784]), .rectangle3_weight(rectangle3_weights[784]), .feature_threshold(feature_thresholds[784]), .feature_above(feature_aboves[784]), .feature_below(feature_belows[784]), .scan_win_std_dev(scan_win_std_dev[784]), .feature_accum(feature_accums[784]));
  accum_calculator ac785(.scan_win(scan_win785), .rectangle1_x(rectangle1_xs[785]), .rectangle1_y(rectangle1_ys[785]), .rectangle1_width(rectangle1_widths[785]), .rectangle1_height(rectangle1_heights[785]), .rectangle1_weight(rectangle1_weights[785]), .rectangle2_x(rectangle2_xs[785]), .rectangle2_y(rectangle2_ys[785]), .rectangle2_width(rectangle2_widths[785]), .rectangle2_height(rectangle2_heights[785]), .rectangle2_weight(rectangle2_weights[785]), .rectangle3_x(rectangle3_xs[785]), .rectangle3_y(rectangle3_ys[785]), .rectangle3_width(rectangle3_widths[785]), .rectangle3_height(rectangle3_heights[785]), .rectangle3_weight(rectangle3_weights[785]), .feature_threshold(feature_thresholds[785]), .feature_above(feature_aboves[785]), .feature_below(feature_belows[785]), .scan_win_std_dev(scan_win_std_dev[785]), .feature_accum(feature_accums[785]));
  accum_calculator ac786(.scan_win(scan_win786), .rectangle1_x(rectangle1_xs[786]), .rectangle1_y(rectangle1_ys[786]), .rectangle1_width(rectangle1_widths[786]), .rectangle1_height(rectangle1_heights[786]), .rectangle1_weight(rectangle1_weights[786]), .rectangle2_x(rectangle2_xs[786]), .rectangle2_y(rectangle2_ys[786]), .rectangle2_width(rectangle2_widths[786]), .rectangle2_height(rectangle2_heights[786]), .rectangle2_weight(rectangle2_weights[786]), .rectangle3_x(rectangle3_xs[786]), .rectangle3_y(rectangle3_ys[786]), .rectangle3_width(rectangle3_widths[786]), .rectangle3_height(rectangle3_heights[786]), .rectangle3_weight(rectangle3_weights[786]), .feature_threshold(feature_thresholds[786]), .feature_above(feature_aboves[786]), .feature_below(feature_belows[786]), .scan_win_std_dev(scan_win_std_dev[786]), .feature_accum(feature_accums[786]));
  accum_calculator ac787(.scan_win(scan_win787), .rectangle1_x(rectangle1_xs[787]), .rectangle1_y(rectangle1_ys[787]), .rectangle1_width(rectangle1_widths[787]), .rectangle1_height(rectangle1_heights[787]), .rectangle1_weight(rectangle1_weights[787]), .rectangle2_x(rectangle2_xs[787]), .rectangle2_y(rectangle2_ys[787]), .rectangle2_width(rectangle2_widths[787]), .rectangle2_height(rectangle2_heights[787]), .rectangle2_weight(rectangle2_weights[787]), .rectangle3_x(rectangle3_xs[787]), .rectangle3_y(rectangle3_ys[787]), .rectangle3_width(rectangle3_widths[787]), .rectangle3_height(rectangle3_heights[787]), .rectangle3_weight(rectangle3_weights[787]), .feature_threshold(feature_thresholds[787]), .feature_above(feature_aboves[787]), .feature_below(feature_belows[787]), .scan_win_std_dev(scan_win_std_dev[787]), .feature_accum(feature_accums[787]));
  accum_calculator ac788(.scan_win(scan_win788), .rectangle1_x(rectangle1_xs[788]), .rectangle1_y(rectangle1_ys[788]), .rectangle1_width(rectangle1_widths[788]), .rectangle1_height(rectangle1_heights[788]), .rectangle1_weight(rectangle1_weights[788]), .rectangle2_x(rectangle2_xs[788]), .rectangle2_y(rectangle2_ys[788]), .rectangle2_width(rectangle2_widths[788]), .rectangle2_height(rectangle2_heights[788]), .rectangle2_weight(rectangle2_weights[788]), .rectangle3_x(rectangle3_xs[788]), .rectangle3_y(rectangle3_ys[788]), .rectangle3_width(rectangle3_widths[788]), .rectangle3_height(rectangle3_heights[788]), .rectangle3_weight(rectangle3_weights[788]), .feature_threshold(feature_thresholds[788]), .feature_above(feature_aboves[788]), .feature_below(feature_belows[788]), .scan_win_std_dev(scan_win_std_dev[788]), .feature_accum(feature_accums[788]));
  accum_calculator ac789(.scan_win(scan_win789), .rectangle1_x(rectangle1_xs[789]), .rectangle1_y(rectangle1_ys[789]), .rectangle1_width(rectangle1_widths[789]), .rectangle1_height(rectangle1_heights[789]), .rectangle1_weight(rectangle1_weights[789]), .rectangle2_x(rectangle2_xs[789]), .rectangle2_y(rectangle2_ys[789]), .rectangle2_width(rectangle2_widths[789]), .rectangle2_height(rectangle2_heights[789]), .rectangle2_weight(rectangle2_weights[789]), .rectangle3_x(rectangle3_xs[789]), .rectangle3_y(rectangle3_ys[789]), .rectangle3_width(rectangle3_widths[789]), .rectangle3_height(rectangle3_heights[789]), .rectangle3_weight(rectangle3_weights[789]), .feature_threshold(feature_thresholds[789]), .feature_above(feature_aboves[789]), .feature_below(feature_belows[789]), .scan_win_std_dev(scan_win_std_dev[789]), .feature_accum(feature_accums[789]));
  accum_calculator ac790(.scan_win(scan_win790), .rectangle1_x(rectangle1_xs[790]), .rectangle1_y(rectangle1_ys[790]), .rectangle1_width(rectangle1_widths[790]), .rectangle1_height(rectangle1_heights[790]), .rectangle1_weight(rectangle1_weights[790]), .rectangle2_x(rectangle2_xs[790]), .rectangle2_y(rectangle2_ys[790]), .rectangle2_width(rectangle2_widths[790]), .rectangle2_height(rectangle2_heights[790]), .rectangle2_weight(rectangle2_weights[790]), .rectangle3_x(rectangle3_xs[790]), .rectangle3_y(rectangle3_ys[790]), .rectangle3_width(rectangle3_widths[790]), .rectangle3_height(rectangle3_heights[790]), .rectangle3_weight(rectangle3_weights[790]), .feature_threshold(feature_thresholds[790]), .feature_above(feature_aboves[790]), .feature_below(feature_belows[790]), .scan_win_std_dev(scan_win_std_dev[790]), .feature_accum(feature_accums[790]));
  accum_calculator ac791(.scan_win(scan_win791), .rectangle1_x(rectangle1_xs[791]), .rectangle1_y(rectangle1_ys[791]), .rectangle1_width(rectangle1_widths[791]), .rectangle1_height(rectangle1_heights[791]), .rectangle1_weight(rectangle1_weights[791]), .rectangle2_x(rectangle2_xs[791]), .rectangle2_y(rectangle2_ys[791]), .rectangle2_width(rectangle2_widths[791]), .rectangle2_height(rectangle2_heights[791]), .rectangle2_weight(rectangle2_weights[791]), .rectangle3_x(rectangle3_xs[791]), .rectangle3_y(rectangle3_ys[791]), .rectangle3_width(rectangle3_widths[791]), .rectangle3_height(rectangle3_heights[791]), .rectangle3_weight(rectangle3_weights[791]), .feature_threshold(feature_thresholds[791]), .feature_above(feature_aboves[791]), .feature_below(feature_belows[791]), .scan_win_std_dev(scan_win_std_dev[791]), .feature_accum(feature_accums[791]));
  accum_calculator ac792(.scan_win(scan_win792), .rectangle1_x(rectangle1_xs[792]), .rectangle1_y(rectangle1_ys[792]), .rectangle1_width(rectangle1_widths[792]), .rectangle1_height(rectangle1_heights[792]), .rectangle1_weight(rectangle1_weights[792]), .rectangle2_x(rectangle2_xs[792]), .rectangle2_y(rectangle2_ys[792]), .rectangle2_width(rectangle2_widths[792]), .rectangle2_height(rectangle2_heights[792]), .rectangle2_weight(rectangle2_weights[792]), .rectangle3_x(rectangle3_xs[792]), .rectangle3_y(rectangle3_ys[792]), .rectangle3_width(rectangle3_widths[792]), .rectangle3_height(rectangle3_heights[792]), .rectangle3_weight(rectangle3_weights[792]), .feature_threshold(feature_thresholds[792]), .feature_above(feature_aboves[792]), .feature_below(feature_belows[792]), .scan_win_std_dev(scan_win_std_dev[792]), .feature_accum(feature_accums[792]));
  accum_calculator ac793(.scan_win(scan_win793), .rectangle1_x(rectangle1_xs[793]), .rectangle1_y(rectangle1_ys[793]), .rectangle1_width(rectangle1_widths[793]), .rectangle1_height(rectangle1_heights[793]), .rectangle1_weight(rectangle1_weights[793]), .rectangle2_x(rectangle2_xs[793]), .rectangle2_y(rectangle2_ys[793]), .rectangle2_width(rectangle2_widths[793]), .rectangle2_height(rectangle2_heights[793]), .rectangle2_weight(rectangle2_weights[793]), .rectangle3_x(rectangle3_xs[793]), .rectangle3_y(rectangle3_ys[793]), .rectangle3_width(rectangle3_widths[793]), .rectangle3_height(rectangle3_heights[793]), .rectangle3_weight(rectangle3_weights[793]), .feature_threshold(feature_thresholds[793]), .feature_above(feature_aboves[793]), .feature_below(feature_belows[793]), .scan_win_std_dev(scan_win_std_dev[793]), .feature_accum(feature_accums[793]));
  accum_calculator ac794(.scan_win(scan_win794), .rectangle1_x(rectangle1_xs[794]), .rectangle1_y(rectangle1_ys[794]), .rectangle1_width(rectangle1_widths[794]), .rectangle1_height(rectangle1_heights[794]), .rectangle1_weight(rectangle1_weights[794]), .rectangle2_x(rectangle2_xs[794]), .rectangle2_y(rectangle2_ys[794]), .rectangle2_width(rectangle2_widths[794]), .rectangle2_height(rectangle2_heights[794]), .rectangle2_weight(rectangle2_weights[794]), .rectangle3_x(rectangle3_xs[794]), .rectangle3_y(rectangle3_ys[794]), .rectangle3_width(rectangle3_widths[794]), .rectangle3_height(rectangle3_heights[794]), .rectangle3_weight(rectangle3_weights[794]), .feature_threshold(feature_thresholds[794]), .feature_above(feature_aboves[794]), .feature_below(feature_belows[794]), .scan_win_std_dev(scan_win_std_dev[794]), .feature_accum(feature_accums[794]));
  accum_calculator ac795(.scan_win(scan_win795), .rectangle1_x(rectangle1_xs[795]), .rectangle1_y(rectangle1_ys[795]), .rectangle1_width(rectangle1_widths[795]), .rectangle1_height(rectangle1_heights[795]), .rectangle1_weight(rectangle1_weights[795]), .rectangle2_x(rectangle2_xs[795]), .rectangle2_y(rectangle2_ys[795]), .rectangle2_width(rectangle2_widths[795]), .rectangle2_height(rectangle2_heights[795]), .rectangle2_weight(rectangle2_weights[795]), .rectangle3_x(rectangle3_xs[795]), .rectangle3_y(rectangle3_ys[795]), .rectangle3_width(rectangle3_widths[795]), .rectangle3_height(rectangle3_heights[795]), .rectangle3_weight(rectangle3_weights[795]), .feature_threshold(feature_thresholds[795]), .feature_above(feature_aboves[795]), .feature_below(feature_belows[795]), .scan_win_std_dev(scan_win_std_dev[795]), .feature_accum(feature_accums[795]));
  accum_calculator ac796(.scan_win(scan_win796), .rectangle1_x(rectangle1_xs[796]), .rectangle1_y(rectangle1_ys[796]), .rectangle1_width(rectangle1_widths[796]), .rectangle1_height(rectangle1_heights[796]), .rectangle1_weight(rectangle1_weights[796]), .rectangle2_x(rectangle2_xs[796]), .rectangle2_y(rectangle2_ys[796]), .rectangle2_width(rectangle2_widths[796]), .rectangle2_height(rectangle2_heights[796]), .rectangle2_weight(rectangle2_weights[796]), .rectangle3_x(rectangle3_xs[796]), .rectangle3_y(rectangle3_ys[796]), .rectangle3_width(rectangle3_widths[796]), .rectangle3_height(rectangle3_heights[796]), .rectangle3_weight(rectangle3_weights[796]), .feature_threshold(feature_thresholds[796]), .feature_above(feature_aboves[796]), .feature_below(feature_belows[796]), .scan_win_std_dev(scan_win_std_dev[796]), .feature_accum(feature_accums[796]));
  accum_calculator ac797(.scan_win(scan_win797), .rectangle1_x(rectangle1_xs[797]), .rectangle1_y(rectangle1_ys[797]), .rectangle1_width(rectangle1_widths[797]), .rectangle1_height(rectangle1_heights[797]), .rectangle1_weight(rectangle1_weights[797]), .rectangle2_x(rectangle2_xs[797]), .rectangle2_y(rectangle2_ys[797]), .rectangle2_width(rectangle2_widths[797]), .rectangle2_height(rectangle2_heights[797]), .rectangle2_weight(rectangle2_weights[797]), .rectangle3_x(rectangle3_xs[797]), .rectangle3_y(rectangle3_ys[797]), .rectangle3_width(rectangle3_widths[797]), .rectangle3_height(rectangle3_heights[797]), .rectangle3_weight(rectangle3_weights[797]), .feature_threshold(feature_thresholds[797]), .feature_above(feature_aboves[797]), .feature_below(feature_belows[797]), .scan_win_std_dev(scan_win_std_dev[797]), .feature_accum(feature_accums[797]));
  accum_calculator ac798(.scan_win(scan_win798), .rectangle1_x(rectangle1_xs[798]), .rectangle1_y(rectangle1_ys[798]), .rectangle1_width(rectangle1_widths[798]), .rectangle1_height(rectangle1_heights[798]), .rectangle1_weight(rectangle1_weights[798]), .rectangle2_x(rectangle2_xs[798]), .rectangle2_y(rectangle2_ys[798]), .rectangle2_width(rectangle2_widths[798]), .rectangle2_height(rectangle2_heights[798]), .rectangle2_weight(rectangle2_weights[798]), .rectangle3_x(rectangle3_xs[798]), .rectangle3_y(rectangle3_ys[798]), .rectangle3_width(rectangle3_widths[798]), .rectangle3_height(rectangle3_heights[798]), .rectangle3_weight(rectangle3_weights[798]), .feature_threshold(feature_thresholds[798]), .feature_above(feature_aboves[798]), .feature_below(feature_belows[798]), .scan_win_std_dev(scan_win_std_dev[798]), .feature_accum(feature_accums[798]));
  accum_calculator ac799(.scan_win(scan_win799), .rectangle1_x(rectangle1_xs[799]), .rectangle1_y(rectangle1_ys[799]), .rectangle1_width(rectangle1_widths[799]), .rectangle1_height(rectangle1_heights[799]), .rectangle1_weight(rectangle1_weights[799]), .rectangle2_x(rectangle2_xs[799]), .rectangle2_y(rectangle2_ys[799]), .rectangle2_width(rectangle2_widths[799]), .rectangle2_height(rectangle2_heights[799]), .rectangle2_weight(rectangle2_weights[799]), .rectangle3_x(rectangle3_xs[799]), .rectangle3_y(rectangle3_ys[799]), .rectangle3_width(rectangle3_widths[799]), .rectangle3_height(rectangle3_heights[799]), .rectangle3_weight(rectangle3_weights[799]), .feature_threshold(feature_thresholds[799]), .feature_above(feature_aboves[799]), .feature_below(feature_belows[799]), .scan_win_std_dev(scan_win_std_dev[799]), .feature_accum(feature_accums[799]));
  accum_calculator ac800(.scan_win(scan_win800), .rectangle1_x(rectangle1_xs[800]), .rectangle1_y(rectangle1_ys[800]), .rectangle1_width(rectangle1_widths[800]), .rectangle1_height(rectangle1_heights[800]), .rectangle1_weight(rectangle1_weights[800]), .rectangle2_x(rectangle2_xs[800]), .rectangle2_y(rectangle2_ys[800]), .rectangle2_width(rectangle2_widths[800]), .rectangle2_height(rectangle2_heights[800]), .rectangle2_weight(rectangle2_weights[800]), .rectangle3_x(rectangle3_xs[800]), .rectangle3_y(rectangle3_ys[800]), .rectangle3_width(rectangle3_widths[800]), .rectangle3_height(rectangle3_heights[800]), .rectangle3_weight(rectangle3_weights[800]), .feature_threshold(feature_thresholds[800]), .feature_above(feature_aboves[800]), .feature_below(feature_belows[800]), .scan_win_std_dev(scan_win_std_dev[800]), .feature_accum(feature_accums[800]));
  accum_calculator ac801(.scan_win(scan_win801), .rectangle1_x(rectangle1_xs[801]), .rectangle1_y(rectangle1_ys[801]), .rectangle1_width(rectangle1_widths[801]), .rectangle1_height(rectangle1_heights[801]), .rectangle1_weight(rectangle1_weights[801]), .rectangle2_x(rectangle2_xs[801]), .rectangle2_y(rectangle2_ys[801]), .rectangle2_width(rectangle2_widths[801]), .rectangle2_height(rectangle2_heights[801]), .rectangle2_weight(rectangle2_weights[801]), .rectangle3_x(rectangle3_xs[801]), .rectangle3_y(rectangle3_ys[801]), .rectangle3_width(rectangle3_widths[801]), .rectangle3_height(rectangle3_heights[801]), .rectangle3_weight(rectangle3_weights[801]), .feature_threshold(feature_thresholds[801]), .feature_above(feature_aboves[801]), .feature_below(feature_belows[801]), .scan_win_std_dev(scan_win_std_dev[801]), .feature_accum(feature_accums[801]));
  accum_calculator ac802(.scan_win(scan_win802), .rectangle1_x(rectangle1_xs[802]), .rectangle1_y(rectangle1_ys[802]), .rectangle1_width(rectangle1_widths[802]), .rectangle1_height(rectangle1_heights[802]), .rectangle1_weight(rectangle1_weights[802]), .rectangle2_x(rectangle2_xs[802]), .rectangle2_y(rectangle2_ys[802]), .rectangle2_width(rectangle2_widths[802]), .rectangle2_height(rectangle2_heights[802]), .rectangle2_weight(rectangle2_weights[802]), .rectangle3_x(rectangle3_xs[802]), .rectangle3_y(rectangle3_ys[802]), .rectangle3_width(rectangle3_widths[802]), .rectangle3_height(rectangle3_heights[802]), .rectangle3_weight(rectangle3_weights[802]), .feature_threshold(feature_thresholds[802]), .feature_above(feature_aboves[802]), .feature_below(feature_belows[802]), .scan_win_std_dev(scan_win_std_dev[802]), .feature_accum(feature_accums[802]));
  accum_calculator ac803(.scan_win(scan_win803), .rectangle1_x(rectangle1_xs[803]), .rectangle1_y(rectangle1_ys[803]), .rectangle1_width(rectangle1_widths[803]), .rectangle1_height(rectangle1_heights[803]), .rectangle1_weight(rectangle1_weights[803]), .rectangle2_x(rectangle2_xs[803]), .rectangle2_y(rectangle2_ys[803]), .rectangle2_width(rectangle2_widths[803]), .rectangle2_height(rectangle2_heights[803]), .rectangle2_weight(rectangle2_weights[803]), .rectangle3_x(rectangle3_xs[803]), .rectangle3_y(rectangle3_ys[803]), .rectangle3_width(rectangle3_widths[803]), .rectangle3_height(rectangle3_heights[803]), .rectangle3_weight(rectangle3_weights[803]), .feature_threshold(feature_thresholds[803]), .feature_above(feature_aboves[803]), .feature_below(feature_belows[803]), .scan_win_std_dev(scan_win_std_dev[803]), .feature_accum(feature_accums[803]));
  accum_calculator ac804(.scan_win(scan_win804), .rectangle1_x(rectangle1_xs[804]), .rectangle1_y(rectangle1_ys[804]), .rectangle1_width(rectangle1_widths[804]), .rectangle1_height(rectangle1_heights[804]), .rectangle1_weight(rectangle1_weights[804]), .rectangle2_x(rectangle2_xs[804]), .rectangle2_y(rectangle2_ys[804]), .rectangle2_width(rectangle2_widths[804]), .rectangle2_height(rectangle2_heights[804]), .rectangle2_weight(rectangle2_weights[804]), .rectangle3_x(rectangle3_xs[804]), .rectangle3_y(rectangle3_ys[804]), .rectangle3_width(rectangle3_widths[804]), .rectangle3_height(rectangle3_heights[804]), .rectangle3_weight(rectangle3_weights[804]), .feature_threshold(feature_thresholds[804]), .feature_above(feature_aboves[804]), .feature_below(feature_belows[804]), .scan_win_std_dev(scan_win_std_dev[804]), .feature_accum(feature_accums[804]));
  accum_calculator ac805(.scan_win(scan_win805), .rectangle1_x(rectangle1_xs[805]), .rectangle1_y(rectangle1_ys[805]), .rectangle1_width(rectangle1_widths[805]), .rectangle1_height(rectangle1_heights[805]), .rectangle1_weight(rectangle1_weights[805]), .rectangle2_x(rectangle2_xs[805]), .rectangle2_y(rectangle2_ys[805]), .rectangle2_width(rectangle2_widths[805]), .rectangle2_height(rectangle2_heights[805]), .rectangle2_weight(rectangle2_weights[805]), .rectangle3_x(rectangle3_xs[805]), .rectangle3_y(rectangle3_ys[805]), .rectangle3_width(rectangle3_widths[805]), .rectangle3_height(rectangle3_heights[805]), .rectangle3_weight(rectangle3_weights[805]), .feature_threshold(feature_thresholds[805]), .feature_above(feature_aboves[805]), .feature_below(feature_belows[805]), .scan_win_std_dev(scan_win_std_dev[805]), .feature_accum(feature_accums[805]));
  accum_calculator ac806(.scan_win(scan_win806), .rectangle1_x(rectangle1_xs[806]), .rectangle1_y(rectangle1_ys[806]), .rectangle1_width(rectangle1_widths[806]), .rectangle1_height(rectangle1_heights[806]), .rectangle1_weight(rectangle1_weights[806]), .rectangle2_x(rectangle2_xs[806]), .rectangle2_y(rectangle2_ys[806]), .rectangle2_width(rectangle2_widths[806]), .rectangle2_height(rectangle2_heights[806]), .rectangle2_weight(rectangle2_weights[806]), .rectangle3_x(rectangle3_xs[806]), .rectangle3_y(rectangle3_ys[806]), .rectangle3_width(rectangle3_widths[806]), .rectangle3_height(rectangle3_heights[806]), .rectangle3_weight(rectangle3_weights[806]), .feature_threshold(feature_thresholds[806]), .feature_above(feature_aboves[806]), .feature_below(feature_belows[806]), .scan_win_std_dev(scan_win_std_dev[806]), .feature_accum(feature_accums[806]));
  accum_calculator ac807(.scan_win(scan_win807), .rectangle1_x(rectangle1_xs[807]), .rectangle1_y(rectangle1_ys[807]), .rectangle1_width(rectangle1_widths[807]), .rectangle1_height(rectangle1_heights[807]), .rectangle1_weight(rectangle1_weights[807]), .rectangle2_x(rectangle2_xs[807]), .rectangle2_y(rectangle2_ys[807]), .rectangle2_width(rectangle2_widths[807]), .rectangle2_height(rectangle2_heights[807]), .rectangle2_weight(rectangle2_weights[807]), .rectangle3_x(rectangle3_xs[807]), .rectangle3_y(rectangle3_ys[807]), .rectangle3_width(rectangle3_widths[807]), .rectangle3_height(rectangle3_heights[807]), .rectangle3_weight(rectangle3_weights[807]), .feature_threshold(feature_thresholds[807]), .feature_above(feature_aboves[807]), .feature_below(feature_belows[807]), .scan_win_std_dev(scan_win_std_dev[807]), .feature_accum(feature_accums[807]));
  accum_calculator ac808(.scan_win(scan_win808), .rectangle1_x(rectangle1_xs[808]), .rectangle1_y(rectangle1_ys[808]), .rectangle1_width(rectangle1_widths[808]), .rectangle1_height(rectangle1_heights[808]), .rectangle1_weight(rectangle1_weights[808]), .rectangle2_x(rectangle2_xs[808]), .rectangle2_y(rectangle2_ys[808]), .rectangle2_width(rectangle2_widths[808]), .rectangle2_height(rectangle2_heights[808]), .rectangle2_weight(rectangle2_weights[808]), .rectangle3_x(rectangle3_xs[808]), .rectangle3_y(rectangle3_ys[808]), .rectangle3_width(rectangle3_widths[808]), .rectangle3_height(rectangle3_heights[808]), .rectangle3_weight(rectangle3_weights[808]), .feature_threshold(feature_thresholds[808]), .feature_above(feature_aboves[808]), .feature_below(feature_belows[808]), .scan_win_std_dev(scan_win_std_dev[808]), .feature_accum(feature_accums[808]));
  accum_calculator ac809(.scan_win(scan_win809), .rectangle1_x(rectangle1_xs[809]), .rectangle1_y(rectangle1_ys[809]), .rectangle1_width(rectangle1_widths[809]), .rectangle1_height(rectangle1_heights[809]), .rectangle1_weight(rectangle1_weights[809]), .rectangle2_x(rectangle2_xs[809]), .rectangle2_y(rectangle2_ys[809]), .rectangle2_width(rectangle2_widths[809]), .rectangle2_height(rectangle2_heights[809]), .rectangle2_weight(rectangle2_weights[809]), .rectangle3_x(rectangle3_xs[809]), .rectangle3_y(rectangle3_ys[809]), .rectangle3_width(rectangle3_widths[809]), .rectangle3_height(rectangle3_heights[809]), .rectangle3_weight(rectangle3_weights[809]), .feature_threshold(feature_thresholds[809]), .feature_above(feature_aboves[809]), .feature_below(feature_belows[809]), .scan_win_std_dev(scan_win_std_dev[809]), .feature_accum(feature_accums[809]));
  accum_calculator ac810(.scan_win(scan_win810), .rectangle1_x(rectangle1_xs[810]), .rectangle1_y(rectangle1_ys[810]), .rectangle1_width(rectangle1_widths[810]), .rectangle1_height(rectangle1_heights[810]), .rectangle1_weight(rectangle1_weights[810]), .rectangle2_x(rectangle2_xs[810]), .rectangle2_y(rectangle2_ys[810]), .rectangle2_width(rectangle2_widths[810]), .rectangle2_height(rectangle2_heights[810]), .rectangle2_weight(rectangle2_weights[810]), .rectangle3_x(rectangle3_xs[810]), .rectangle3_y(rectangle3_ys[810]), .rectangle3_width(rectangle3_widths[810]), .rectangle3_height(rectangle3_heights[810]), .rectangle3_weight(rectangle3_weights[810]), .feature_threshold(feature_thresholds[810]), .feature_above(feature_aboves[810]), .feature_below(feature_belows[810]), .scan_win_std_dev(scan_win_std_dev[810]), .feature_accum(feature_accums[810]));
  accum_calculator ac811(.scan_win(scan_win811), .rectangle1_x(rectangle1_xs[811]), .rectangle1_y(rectangle1_ys[811]), .rectangle1_width(rectangle1_widths[811]), .rectangle1_height(rectangle1_heights[811]), .rectangle1_weight(rectangle1_weights[811]), .rectangle2_x(rectangle2_xs[811]), .rectangle2_y(rectangle2_ys[811]), .rectangle2_width(rectangle2_widths[811]), .rectangle2_height(rectangle2_heights[811]), .rectangle2_weight(rectangle2_weights[811]), .rectangle3_x(rectangle3_xs[811]), .rectangle3_y(rectangle3_ys[811]), .rectangle3_width(rectangle3_widths[811]), .rectangle3_height(rectangle3_heights[811]), .rectangle3_weight(rectangle3_weights[811]), .feature_threshold(feature_thresholds[811]), .feature_above(feature_aboves[811]), .feature_below(feature_belows[811]), .scan_win_std_dev(scan_win_std_dev[811]), .feature_accum(feature_accums[811]));
  accum_calculator ac812(.scan_win(scan_win812), .rectangle1_x(rectangle1_xs[812]), .rectangle1_y(rectangle1_ys[812]), .rectangle1_width(rectangle1_widths[812]), .rectangle1_height(rectangle1_heights[812]), .rectangle1_weight(rectangle1_weights[812]), .rectangle2_x(rectangle2_xs[812]), .rectangle2_y(rectangle2_ys[812]), .rectangle2_width(rectangle2_widths[812]), .rectangle2_height(rectangle2_heights[812]), .rectangle2_weight(rectangle2_weights[812]), .rectangle3_x(rectangle3_xs[812]), .rectangle3_y(rectangle3_ys[812]), .rectangle3_width(rectangle3_widths[812]), .rectangle3_height(rectangle3_heights[812]), .rectangle3_weight(rectangle3_weights[812]), .feature_threshold(feature_thresholds[812]), .feature_above(feature_aboves[812]), .feature_below(feature_belows[812]), .scan_win_std_dev(scan_win_std_dev[812]), .feature_accum(feature_accums[812]));
  accum_calculator ac813(.scan_win(scan_win813), .rectangle1_x(rectangle1_xs[813]), .rectangle1_y(rectangle1_ys[813]), .rectangle1_width(rectangle1_widths[813]), .rectangle1_height(rectangle1_heights[813]), .rectangle1_weight(rectangle1_weights[813]), .rectangle2_x(rectangle2_xs[813]), .rectangle2_y(rectangle2_ys[813]), .rectangle2_width(rectangle2_widths[813]), .rectangle2_height(rectangle2_heights[813]), .rectangle2_weight(rectangle2_weights[813]), .rectangle3_x(rectangle3_xs[813]), .rectangle3_y(rectangle3_ys[813]), .rectangle3_width(rectangle3_widths[813]), .rectangle3_height(rectangle3_heights[813]), .rectangle3_weight(rectangle3_weights[813]), .feature_threshold(feature_thresholds[813]), .feature_above(feature_aboves[813]), .feature_below(feature_belows[813]), .scan_win_std_dev(scan_win_std_dev[813]), .feature_accum(feature_accums[813]));
  accum_calculator ac814(.scan_win(scan_win814), .rectangle1_x(rectangle1_xs[814]), .rectangle1_y(rectangle1_ys[814]), .rectangle1_width(rectangle1_widths[814]), .rectangle1_height(rectangle1_heights[814]), .rectangle1_weight(rectangle1_weights[814]), .rectangle2_x(rectangle2_xs[814]), .rectangle2_y(rectangle2_ys[814]), .rectangle2_width(rectangle2_widths[814]), .rectangle2_height(rectangle2_heights[814]), .rectangle2_weight(rectangle2_weights[814]), .rectangle3_x(rectangle3_xs[814]), .rectangle3_y(rectangle3_ys[814]), .rectangle3_width(rectangle3_widths[814]), .rectangle3_height(rectangle3_heights[814]), .rectangle3_weight(rectangle3_weights[814]), .feature_threshold(feature_thresholds[814]), .feature_above(feature_aboves[814]), .feature_below(feature_belows[814]), .scan_win_std_dev(scan_win_std_dev[814]), .feature_accum(feature_accums[814]));
  accum_calculator ac815(.scan_win(scan_win815), .rectangle1_x(rectangle1_xs[815]), .rectangle1_y(rectangle1_ys[815]), .rectangle1_width(rectangle1_widths[815]), .rectangle1_height(rectangle1_heights[815]), .rectangle1_weight(rectangle1_weights[815]), .rectangle2_x(rectangle2_xs[815]), .rectangle2_y(rectangle2_ys[815]), .rectangle2_width(rectangle2_widths[815]), .rectangle2_height(rectangle2_heights[815]), .rectangle2_weight(rectangle2_weights[815]), .rectangle3_x(rectangle3_xs[815]), .rectangle3_y(rectangle3_ys[815]), .rectangle3_width(rectangle3_widths[815]), .rectangle3_height(rectangle3_heights[815]), .rectangle3_weight(rectangle3_weights[815]), .feature_threshold(feature_thresholds[815]), .feature_above(feature_aboves[815]), .feature_below(feature_belows[815]), .scan_win_std_dev(scan_win_std_dev[815]), .feature_accum(feature_accums[815]));
  accum_calculator ac816(.scan_win(scan_win816), .rectangle1_x(rectangle1_xs[816]), .rectangle1_y(rectangle1_ys[816]), .rectangle1_width(rectangle1_widths[816]), .rectangle1_height(rectangle1_heights[816]), .rectangle1_weight(rectangle1_weights[816]), .rectangle2_x(rectangle2_xs[816]), .rectangle2_y(rectangle2_ys[816]), .rectangle2_width(rectangle2_widths[816]), .rectangle2_height(rectangle2_heights[816]), .rectangle2_weight(rectangle2_weights[816]), .rectangle3_x(rectangle3_xs[816]), .rectangle3_y(rectangle3_ys[816]), .rectangle3_width(rectangle3_widths[816]), .rectangle3_height(rectangle3_heights[816]), .rectangle3_weight(rectangle3_weights[816]), .feature_threshold(feature_thresholds[816]), .feature_above(feature_aboves[816]), .feature_below(feature_belows[816]), .scan_win_std_dev(scan_win_std_dev[816]), .feature_accum(feature_accums[816]));
  accum_calculator ac817(.scan_win(scan_win817), .rectangle1_x(rectangle1_xs[817]), .rectangle1_y(rectangle1_ys[817]), .rectangle1_width(rectangle1_widths[817]), .rectangle1_height(rectangle1_heights[817]), .rectangle1_weight(rectangle1_weights[817]), .rectangle2_x(rectangle2_xs[817]), .rectangle2_y(rectangle2_ys[817]), .rectangle2_width(rectangle2_widths[817]), .rectangle2_height(rectangle2_heights[817]), .rectangle2_weight(rectangle2_weights[817]), .rectangle3_x(rectangle3_xs[817]), .rectangle3_y(rectangle3_ys[817]), .rectangle3_width(rectangle3_widths[817]), .rectangle3_height(rectangle3_heights[817]), .rectangle3_weight(rectangle3_weights[817]), .feature_threshold(feature_thresholds[817]), .feature_above(feature_aboves[817]), .feature_below(feature_belows[817]), .scan_win_std_dev(scan_win_std_dev[817]), .feature_accum(feature_accums[817]));
  accum_calculator ac818(.scan_win(scan_win818), .rectangle1_x(rectangle1_xs[818]), .rectangle1_y(rectangle1_ys[818]), .rectangle1_width(rectangle1_widths[818]), .rectangle1_height(rectangle1_heights[818]), .rectangle1_weight(rectangle1_weights[818]), .rectangle2_x(rectangle2_xs[818]), .rectangle2_y(rectangle2_ys[818]), .rectangle2_width(rectangle2_widths[818]), .rectangle2_height(rectangle2_heights[818]), .rectangle2_weight(rectangle2_weights[818]), .rectangle3_x(rectangle3_xs[818]), .rectangle3_y(rectangle3_ys[818]), .rectangle3_width(rectangle3_widths[818]), .rectangle3_height(rectangle3_heights[818]), .rectangle3_weight(rectangle3_weights[818]), .feature_threshold(feature_thresholds[818]), .feature_above(feature_aboves[818]), .feature_below(feature_belows[818]), .scan_win_std_dev(scan_win_std_dev[818]), .feature_accum(feature_accums[818]));
  accum_calculator ac819(.scan_win(scan_win819), .rectangle1_x(rectangle1_xs[819]), .rectangle1_y(rectangle1_ys[819]), .rectangle1_width(rectangle1_widths[819]), .rectangle1_height(rectangle1_heights[819]), .rectangle1_weight(rectangle1_weights[819]), .rectangle2_x(rectangle2_xs[819]), .rectangle2_y(rectangle2_ys[819]), .rectangle2_width(rectangle2_widths[819]), .rectangle2_height(rectangle2_heights[819]), .rectangle2_weight(rectangle2_weights[819]), .rectangle3_x(rectangle3_xs[819]), .rectangle3_y(rectangle3_ys[819]), .rectangle3_width(rectangle3_widths[819]), .rectangle3_height(rectangle3_heights[819]), .rectangle3_weight(rectangle3_weights[819]), .feature_threshold(feature_thresholds[819]), .feature_above(feature_aboves[819]), .feature_below(feature_belows[819]), .scan_win_std_dev(scan_win_std_dev[819]), .feature_accum(feature_accums[819]));
  accum_calculator ac820(.scan_win(scan_win820), .rectangle1_x(rectangle1_xs[820]), .rectangle1_y(rectangle1_ys[820]), .rectangle1_width(rectangle1_widths[820]), .rectangle1_height(rectangle1_heights[820]), .rectangle1_weight(rectangle1_weights[820]), .rectangle2_x(rectangle2_xs[820]), .rectangle2_y(rectangle2_ys[820]), .rectangle2_width(rectangle2_widths[820]), .rectangle2_height(rectangle2_heights[820]), .rectangle2_weight(rectangle2_weights[820]), .rectangle3_x(rectangle3_xs[820]), .rectangle3_y(rectangle3_ys[820]), .rectangle3_width(rectangle3_widths[820]), .rectangle3_height(rectangle3_heights[820]), .rectangle3_weight(rectangle3_weights[820]), .feature_threshold(feature_thresholds[820]), .feature_above(feature_aboves[820]), .feature_below(feature_belows[820]), .scan_win_std_dev(scan_win_std_dev[820]), .feature_accum(feature_accums[820]));
  accum_calculator ac821(.scan_win(scan_win821), .rectangle1_x(rectangle1_xs[821]), .rectangle1_y(rectangle1_ys[821]), .rectangle1_width(rectangle1_widths[821]), .rectangle1_height(rectangle1_heights[821]), .rectangle1_weight(rectangle1_weights[821]), .rectangle2_x(rectangle2_xs[821]), .rectangle2_y(rectangle2_ys[821]), .rectangle2_width(rectangle2_widths[821]), .rectangle2_height(rectangle2_heights[821]), .rectangle2_weight(rectangle2_weights[821]), .rectangle3_x(rectangle3_xs[821]), .rectangle3_y(rectangle3_ys[821]), .rectangle3_width(rectangle3_widths[821]), .rectangle3_height(rectangle3_heights[821]), .rectangle3_weight(rectangle3_weights[821]), .feature_threshold(feature_thresholds[821]), .feature_above(feature_aboves[821]), .feature_below(feature_belows[821]), .scan_win_std_dev(scan_win_std_dev[821]), .feature_accum(feature_accums[821]));
  accum_calculator ac822(.scan_win(scan_win822), .rectangle1_x(rectangle1_xs[822]), .rectangle1_y(rectangle1_ys[822]), .rectangle1_width(rectangle1_widths[822]), .rectangle1_height(rectangle1_heights[822]), .rectangle1_weight(rectangle1_weights[822]), .rectangle2_x(rectangle2_xs[822]), .rectangle2_y(rectangle2_ys[822]), .rectangle2_width(rectangle2_widths[822]), .rectangle2_height(rectangle2_heights[822]), .rectangle2_weight(rectangle2_weights[822]), .rectangle3_x(rectangle3_xs[822]), .rectangle3_y(rectangle3_ys[822]), .rectangle3_width(rectangle3_widths[822]), .rectangle3_height(rectangle3_heights[822]), .rectangle3_weight(rectangle3_weights[822]), .feature_threshold(feature_thresholds[822]), .feature_above(feature_aboves[822]), .feature_below(feature_belows[822]), .scan_win_std_dev(scan_win_std_dev[822]), .feature_accum(feature_accums[822]));
  accum_calculator ac823(.scan_win(scan_win823), .rectangle1_x(rectangle1_xs[823]), .rectangle1_y(rectangle1_ys[823]), .rectangle1_width(rectangle1_widths[823]), .rectangle1_height(rectangle1_heights[823]), .rectangle1_weight(rectangle1_weights[823]), .rectangle2_x(rectangle2_xs[823]), .rectangle2_y(rectangle2_ys[823]), .rectangle2_width(rectangle2_widths[823]), .rectangle2_height(rectangle2_heights[823]), .rectangle2_weight(rectangle2_weights[823]), .rectangle3_x(rectangle3_xs[823]), .rectangle3_y(rectangle3_ys[823]), .rectangle3_width(rectangle3_widths[823]), .rectangle3_height(rectangle3_heights[823]), .rectangle3_weight(rectangle3_weights[823]), .feature_threshold(feature_thresholds[823]), .feature_above(feature_aboves[823]), .feature_below(feature_belows[823]), .scan_win_std_dev(scan_win_std_dev[823]), .feature_accum(feature_accums[823]));
  accum_calculator ac824(.scan_win(scan_win824), .rectangle1_x(rectangle1_xs[824]), .rectangle1_y(rectangle1_ys[824]), .rectangle1_width(rectangle1_widths[824]), .rectangle1_height(rectangle1_heights[824]), .rectangle1_weight(rectangle1_weights[824]), .rectangle2_x(rectangle2_xs[824]), .rectangle2_y(rectangle2_ys[824]), .rectangle2_width(rectangle2_widths[824]), .rectangle2_height(rectangle2_heights[824]), .rectangle2_weight(rectangle2_weights[824]), .rectangle3_x(rectangle3_xs[824]), .rectangle3_y(rectangle3_ys[824]), .rectangle3_width(rectangle3_widths[824]), .rectangle3_height(rectangle3_heights[824]), .rectangle3_weight(rectangle3_weights[824]), .feature_threshold(feature_thresholds[824]), .feature_above(feature_aboves[824]), .feature_below(feature_belows[824]), .scan_win_std_dev(scan_win_std_dev[824]), .feature_accum(feature_accums[824]));
  accum_calculator ac825(.scan_win(scan_win825), .rectangle1_x(rectangle1_xs[825]), .rectangle1_y(rectangle1_ys[825]), .rectangle1_width(rectangle1_widths[825]), .rectangle1_height(rectangle1_heights[825]), .rectangle1_weight(rectangle1_weights[825]), .rectangle2_x(rectangle2_xs[825]), .rectangle2_y(rectangle2_ys[825]), .rectangle2_width(rectangle2_widths[825]), .rectangle2_height(rectangle2_heights[825]), .rectangle2_weight(rectangle2_weights[825]), .rectangle3_x(rectangle3_xs[825]), .rectangle3_y(rectangle3_ys[825]), .rectangle3_width(rectangle3_widths[825]), .rectangle3_height(rectangle3_heights[825]), .rectangle3_weight(rectangle3_weights[825]), .feature_threshold(feature_thresholds[825]), .feature_above(feature_aboves[825]), .feature_below(feature_belows[825]), .scan_win_std_dev(scan_win_std_dev[825]), .feature_accum(feature_accums[825]));
  accum_calculator ac826(.scan_win(scan_win826), .rectangle1_x(rectangle1_xs[826]), .rectangle1_y(rectangle1_ys[826]), .rectangle1_width(rectangle1_widths[826]), .rectangle1_height(rectangle1_heights[826]), .rectangle1_weight(rectangle1_weights[826]), .rectangle2_x(rectangle2_xs[826]), .rectangle2_y(rectangle2_ys[826]), .rectangle2_width(rectangle2_widths[826]), .rectangle2_height(rectangle2_heights[826]), .rectangle2_weight(rectangle2_weights[826]), .rectangle3_x(rectangle3_xs[826]), .rectangle3_y(rectangle3_ys[826]), .rectangle3_width(rectangle3_widths[826]), .rectangle3_height(rectangle3_heights[826]), .rectangle3_weight(rectangle3_weights[826]), .feature_threshold(feature_thresholds[826]), .feature_above(feature_aboves[826]), .feature_below(feature_belows[826]), .scan_win_std_dev(scan_win_std_dev[826]), .feature_accum(feature_accums[826]));
  accum_calculator ac827(.scan_win(scan_win827), .rectangle1_x(rectangle1_xs[827]), .rectangle1_y(rectangle1_ys[827]), .rectangle1_width(rectangle1_widths[827]), .rectangle1_height(rectangle1_heights[827]), .rectangle1_weight(rectangle1_weights[827]), .rectangle2_x(rectangle2_xs[827]), .rectangle2_y(rectangle2_ys[827]), .rectangle2_width(rectangle2_widths[827]), .rectangle2_height(rectangle2_heights[827]), .rectangle2_weight(rectangle2_weights[827]), .rectangle3_x(rectangle3_xs[827]), .rectangle3_y(rectangle3_ys[827]), .rectangle3_width(rectangle3_widths[827]), .rectangle3_height(rectangle3_heights[827]), .rectangle3_weight(rectangle3_weights[827]), .feature_threshold(feature_thresholds[827]), .feature_above(feature_aboves[827]), .feature_below(feature_belows[827]), .scan_win_std_dev(scan_win_std_dev[827]), .feature_accum(feature_accums[827]));
  accum_calculator ac828(.scan_win(scan_win828), .rectangle1_x(rectangle1_xs[828]), .rectangle1_y(rectangle1_ys[828]), .rectangle1_width(rectangle1_widths[828]), .rectangle1_height(rectangle1_heights[828]), .rectangle1_weight(rectangle1_weights[828]), .rectangle2_x(rectangle2_xs[828]), .rectangle2_y(rectangle2_ys[828]), .rectangle2_width(rectangle2_widths[828]), .rectangle2_height(rectangle2_heights[828]), .rectangle2_weight(rectangle2_weights[828]), .rectangle3_x(rectangle3_xs[828]), .rectangle3_y(rectangle3_ys[828]), .rectangle3_width(rectangle3_widths[828]), .rectangle3_height(rectangle3_heights[828]), .rectangle3_weight(rectangle3_weights[828]), .feature_threshold(feature_thresholds[828]), .feature_above(feature_aboves[828]), .feature_below(feature_belows[828]), .scan_win_std_dev(scan_win_std_dev[828]), .feature_accum(feature_accums[828]));
  accum_calculator ac829(.scan_win(scan_win829), .rectangle1_x(rectangle1_xs[829]), .rectangle1_y(rectangle1_ys[829]), .rectangle1_width(rectangle1_widths[829]), .rectangle1_height(rectangle1_heights[829]), .rectangle1_weight(rectangle1_weights[829]), .rectangle2_x(rectangle2_xs[829]), .rectangle2_y(rectangle2_ys[829]), .rectangle2_width(rectangle2_widths[829]), .rectangle2_height(rectangle2_heights[829]), .rectangle2_weight(rectangle2_weights[829]), .rectangle3_x(rectangle3_xs[829]), .rectangle3_y(rectangle3_ys[829]), .rectangle3_width(rectangle3_widths[829]), .rectangle3_height(rectangle3_heights[829]), .rectangle3_weight(rectangle3_weights[829]), .feature_threshold(feature_thresholds[829]), .feature_above(feature_aboves[829]), .feature_below(feature_belows[829]), .scan_win_std_dev(scan_win_std_dev[829]), .feature_accum(feature_accums[829]));
  accum_calculator ac830(.scan_win(scan_win830), .rectangle1_x(rectangle1_xs[830]), .rectangle1_y(rectangle1_ys[830]), .rectangle1_width(rectangle1_widths[830]), .rectangle1_height(rectangle1_heights[830]), .rectangle1_weight(rectangle1_weights[830]), .rectangle2_x(rectangle2_xs[830]), .rectangle2_y(rectangle2_ys[830]), .rectangle2_width(rectangle2_widths[830]), .rectangle2_height(rectangle2_heights[830]), .rectangle2_weight(rectangle2_weights[830]), .rectangle3_x(rectangle3_xs[830]), .rectangle3_y(rectangle3_ys[830]), .rectangle3_width(rectangle3_widths[830]), .rectangle3_height(rectangle3_heights[830]), .rectangle3_weight(rectangle3_weights[830]), .feature_threshold(feature_thresholds[830]), .feature_above(feature_aboves[830]), .feature_below(feature_belows[830]), .scan_win_std_dev(scan_win_std_dev[830]), .feature_accum(feature_accums[830]));
  accum_calculator ac831(.scan_win(scan_win831), .rectangle1_x(rectangle1_xs[831]), .rectangle1_y(rectangle1_ys[831]), .rectangle1_width(rectangle1_widths[831]), .rectangle1_height(rectangle1_heights[831]), .rectangle1_weight(rectangle1_weights[831]), .rectangle2_x(rectangle2_xs[831]), .rectangle2_y(rectangle2_ys[831]), .rectangle2_width(rectangle2_widths[831]), .rectangle2_height(rectangle2_heights[831]), .rectangle2_weight(rectangle2_weights[831]), .rectangle3_x(rectangle3_xs[831]), .rectangle3_y(rectangle3_ys[831]), .rectangle3_width(rectangle3_widths[831]), .rectangle3_height(rectangle3_heights[831]), .rectangle3_weight(rectangle3_weights[831]), .feature_threshold(feature_thresholds[831]), .feature_above(feature_aboves[831]), .feature_below(feature_belows[831]), .scan_win_std_dev(scan_win_std_dev[831]), .feature_accum(feature_accums[831]));
  accum_calculator ac832(.scan_win(scan_win832), .rectangle1_x(rectangle1_xs[832]), .rectangle1_y(rectangle1_ys[832]), .rectangle1_width(rectangle1_widths[832]), .rectangle1_height(rectangle1_heights[832]), .rectangle1_weight(rectangle1_weights[832]), .rectangle2_x(rectangle2_xs[832]), .rectangle2_y(rectangle2_ys[832]), .rectangle2_width(rectangle2_widths[832]), .rectangle2_height(rectangle2_heights[832]), .rectangle2_weight(rectangle2_weights[832]), .rectangle3_x(rectangle3_xs[832]), .rectangle3_y(rectangle3_ys[832]), .rectangle3_width(rectangle3_widths[832]), .rectangle3_height(rectangle3_heights[832]), .rectangle3_weight(rectangle3_weights[832]), .feature_threshold(feature_thresholds[832]), .feature_above(feature_aboves[832]), .feature_below(feature_belows[832]), .scan_win_std_dev(scan_win_std_dev[832]), .feature_accum(feature_accums[832]));
  accum_calculator ac833(.scan_win(scan_win833), .rectangle1_x(rectangle1_xs[833]), .rectangle1_y(rectangle1_ys[833]), .rectangle1_width(rectangle1_widths[833]), .rectangle1_height(rectangle1_heights[833]), .rectangle1_weight(rectangle1_weights[833]), .rectangle2_x(rectangle2_xs[833]), .rectangle2_y(rectangle2_ys[833]), .rectangle2_width(rectangle2_widths[833]), .rectangle2_height(rectangle2_heights[833]), .rectangle2_weight(rectangle2_weights[833]), .rectangle3_x(rectangle3_xs[833]), .rectangle3_y(rectangle3_ys[833]), .rectangle3_width(rectangle3_widths[833]), .rectangle3_height(rectangle3_heights[833]), .rectangle3_weight(rectangle3_weights[833]), .feature_threshold(feature_thresholds[833]), .feature_above(feature_aboves[833]), .feature_below(feature_belows[833]), .scan_win_std_dev(scan_win_std_dev[833]), .feature_accum(feature_accums[833]));
  accum_calculator ac834(.scan_win(scan_win834), .rectangle1_x(rectangle1_xs[834]), .rectangle1_y(rectangle1_ys[834]), .rectangle1_width(rectangle1_widths[834]), .rectangle1_height(rectangle1_heights[834]), .rectangle1_weight(rectangle1_weights[834]), .rectangle2_x(rectangle2_xs[834]), .rectangle2_y(rectangle2_ys[834]), .rectangle2_width(rectangle2_widths[834]), .rectangle2_height(rectangle2_heights[834]), .rectangle2_weight(rectangle2_weights[834]), .rectangle3_x(rectangle3_xs[834]), .rectangle3_y(rectangle3_ys[834]), .rectangle3_width(rectangle3_widths[834]), .rectangle3_height(rectangle3_heights[834]), .rectangle3_weight(rectangle3_weights[834]), .feature_threshold(feature_thresholds[834]), .feature_above(feature_aboves[834]), .feature_below(feature_belows[834]), .scan_win_std_dev(scan_win_std_dev[834]), .feature_accum(feature_accums[834]));
  accum_calculator ac835(.scan_win(scan_win835), .rectangle1_x(rectangle1_xs[835]), .rectangle1_y(rectangle1_ys[835]), .rectangle1_width(rectangle1_widths[835]), .rectangle1_height(rectangle1_heights[835]), .rectangle1_weight(rectangle1_weights[835]), .rectangle2_x(rectangle2_xs[835]), .rectangle2_y(rectangle2_ys[835]), .rectangle2_width(rectangle2_widths[835]), .rectangle2_height(rectangle2_heights[835]), .rectangle2_weight(rectangle2_weights[835]), .rectangle3_x(rectangle3_xs[835]), .rectangle3_y(rectangle3_ys[835]), .rectangle3_width(rectangle3_widths[835]), .rectangle3_height(rectangle3_heights[835]), .rectangle3_weight(rectangle3_weights[835]), .feature_threshold(feature_thresholds[835]), .feature_above(feature_aboves[835]), .feature_below(feature_belows[835]), .scan_win_std_dev(scan_win_std_dev[835]), .feature_accum(feature_accums[835]));
  accum_calculator ac836(.scan_win(scan_win836), .rectangle1_x(rectangle1_xs[836]), .rectangle1_y(rectangle1_ys[836]), .rectangle1_width(rectangle1_widths[836]), .rectangle1_height(rectangle1_heights[836]), .rectangle1_weight(rectangle1_weights[836]), .rectangle2_x(rectangle2_xs[836]), .rectangle2_y(rectangle2_ys[836]), .rectangle2_width(rectangle2_widths[836]), .rectangle2_height(rectangle2_heights[836]), .rectangle2_weight(rectangle2_weights[836]), .rectangle3_x(rectangle3_xs[836]), .rectangle3_y(rectangle3_ys[836]), .rectangle3_width(rectangle3_widths[836]), .rectangle3_height(rectangle3_heights[836]), .rectangle3_weight(rectangle3_weights[836]), .feature_threshold(feature_thresholds[836]), .feature_above(feature_aboves[836]), .feature_below(feature_belows[836]), .scan_win_std_dev(scan_win_std_dev[836]), .feature_accum(feature_accums[836]));
  accum_calculator ac837(.scan_win(scan_win837), .rectangle1_x(rectangle1_xs[837]), .rectangle1_y(rectangle1_ys[837]), .rectangle1_width(rectangle1_widths[837]), .rectangle1_height(rectangle1_heights[837]), .rectangle1_weight(rectangle1_weights[837]), .rectangle2_x(rectangle2_xs[837]), .rectangle2_y(rectangle2_ys[837]), .rectangle2_width(rectangle2_widths[837]), .rectangle2_height(rectangle2_heights[837]), .rectangle2_weight(rectangle2_weights[837]), .rectangle3_x(rectangle3_xs[837]), .rectangle3_y(rectangle3_ys[837]), .rectangle3_width(rectangle3_widths[837]), .rectangle3_height(rectangle3_heights[837]), .rectangle3_weight(rectangle3_weights[837]), .feature_threshold(feature_thresholds[837]), .feature_above(feature_aboves[837]), .feature_below(feature_belows[837]), .scan_win_std_dev(scan_win_std_dev[837]), .feature_accum(feature_accums[837]));
  accum_calculator ac838(.scan_win(scan_win838), .rectangle1_x(rectangle1_xs[838]), .rectangle1_y(rectangle1_ys[838]), .rectangle1_width(rectangle1_widths[838]), .rectangle1_height(rectangle1_heights[838]), .rectangle1_weight(rectangle1_weights[838]), .rectangle2_x(rectangle2_xs[838]), .rectangle2_y(rectangle2_ys[838]), .rectangle2_width(rectangle2_widths[838]), .rectangle2_height(rectangle2_heights[838]), .rectangle2_weight(rectangle2_weights[838]), .rectangle3_x(rectangle3_xs[838]), .rectangle3_y(rectangle3_ys[838]), .rectangle3_width(rectangle3_widths[838]), .rectangle3_height(rectangle3_heights[838]), .rectangle3_weight(rectangle3_weights[838]), .feature_threshold(feature_thresholds[838]), .feature_above(feature_aboves[838]), .feature_below(feature_belows[838]), .scan_win_std_dev(scan_win_std_dev[838]), .feature_accum(feature_accums[838]));
  accum_calculator ac839(.scan_win(scan_win839), .rectangle1_x(rectangle1_xs[839]), .rectangle1_y(rectangle1_ys[839]), .rectangle1_width(rectangle1_widths[839]), .rectangle1_height(rectangle1_heights[839]), .rectangle1_weight(rectangle1_weights[839]), .rectangle2_x(rectangle2_xs[839]), .rectangle2_y(rectangle2_ys[839]), .rectangle2_width(rectangle2_widths[839]), .rectangle2_height(rectangle2_heights[839]), .rectangle2_weight(rectangle2_weights[839]), .rectangle3_x(rectangle3_xs[839]), .rectangle3_y(rectangle3_ys[839]), .rectangle3_width(rectangle3_widths[839]), .rectangle3_height(rectangle3_heights[839]), .rectangle3_weight(rectangle3_weights[839]), .feature_threshold(feature_thresholds[839]), .feature_above(feature_aboves[839]), .feature_below(feature_belows[839]), .scan_win_std_dev(scan_win_std_dev[839]), .feature_accum(feature_accums[839]));
  accum_calculator ac840(.scan_win(scan_win840), .rectangle1_x(rectangle1_xs[840]), .rectangle1_y(rectangle1_ys[840]), .rectangle1_width(rectangle1_widths[840]), .rectangle1_height(rectangle1_heights[840]), .rectangle1_weight(rectangle1_weights[840]), .rectangle2_x(rectangle2_xs[840]), .rectangle2_y(rectangle2_ys[840]), .rectangle2_width(rectangle2_widths[840]), .rectangle2_height(rectangle2_heights[840]), .rectangle2_weight(rectangle2_weights[840]), .rectangle3_x(rectangle3_xs[840]), .rectangle3_y(rectangle3_ys[840]), .rectangle3_width(rectangle3_widths[840]), .rectangle3_height(rectangle3_heights[840]), .rectangle3_weight(rectangle3_weights[840]), .feature_threshold(feature_thresholds[840]), .feature_above(feature_aboves[840]), .feature_below(feature_belows[840]), .scan_win_std_dev(scan_win_std_dev[840]), .feature_accum(feature_accums[840]));
  accum_calculator ac841(.scan_win(scan_win841), .rectangle1_x(rectangle1_xs[841]), .rectangle1_y(rectangle1_ys[841]), .rectangle1_width(rectangle1_widths[841]), .rectangle1_height(rectangle1_heights[841]), .rectangle1_weight(rectangle1_weights[841]), .rectangle2_x(rectangle2_xs[841]), .rectangle2_y(rectangle2_ys[841]), .rectangle2_width(rectangle2_widths[841]), .rectangle2_height(rectangle2_heights[841]), .rectangle2_weight(rectangle2_weights[841]), .rectangle3_x(rectangle3_xs[841]), .rectangle3_y(rectangle3_ys[841]), .rectangle3_width(rectangle3_widths[841]), .rectangle3_height(rectangle3_heights[841]), .rectangle3_weight(rectangle3_weights[841]), .feature_threshold(feature_thresholds[841]), .feature_above(feature_aboves[841]), .feature_below(feature_belows[841]), .scan_win_std_dev(scan_win_std_dev[841]), .feature_accum(feature_accums[841]));
  accum_calculator ac842(.scan_win(scan_win842), .rectangle1_x(rectangle1_xs[842]), .rectangle1_y(rectangle1_ys[842]), .rectangle1_width(rectangle1_widths[842]), .rectangle1_height(rectangle1_heights[842]), .rectangle1_weight(rectangle1_weights[842]), .rectangle2_x(rectangle2_xs[842]), .rectangle2_y(rectangle2_ys[842]), .rectangle2_width(rectangle2_widths[842]), .rectangle2_height(rectangle2_heights[842]), .rectangle2_weight(rectangle2_weights[842]), .rectangle3_x(rectangle3_xs[842]), .rectangle3_y(rectangle3_ys[842]), .rectangle3_width(rectangle3_widths[842]), .rectangle3_height(rectangle3_heights[842]), .rectangle3_weight(rectangle3_weights[842]), .feature_threshold(feature_thresholds[842]), .feature_above(feature_aboves[842]), .feature_below(feature_belows[842]), .scan_win_std_dev(scan_win_std_dev[842]), .feature_accum(feature_accums[842]));
  accum_calculator ac843(.scan_win(scan_win843), .rectangle1_x(rectangle1_xs[843]), .rectangle1_y(rectangle1_ys[843]), .rectangle1_width(rectangle1_widths[843]), .rectangle1_height(rectangle1_heights[843]), .rectangle1_weight(rectangle1_weights[843]), .rectangle2_x(rectangle2_xs[843]), .rectangle2_y(rectangle2_ys[843]), .rectangle2_width(rectangle2_widths[843]), .rectangle2_height(rectangle2_heights[843]), .rectangle2_weight(rectangle2_weights[843]), .rectangle3_x(rectangle3_xs[843]), .rectangle3_y(rectangle3_ys[843]), .rectangle3_width(rectangle3_widths[843]), .rectangle3_height(rectangle3_heights[843]), .rectangle3_weight(rectangle3_weights[843]), .feature_threshold(feature_thresholds[843]), .feature_above(feature_aboves[843]), .feature_below(feature_belows[843]), .scan_win_std_dev(scan_win_std_dev[843]), .feature_accum(feature_accums[843]));
  accum_calculator ac844(.scan_win(scan_win844), .rectangle1_x(rectangle1_xs[844]), .rectangle1_y(rectangle1_ys[844]), .rectangle1_width(rectangle1_widths[844]), .rectangle1_height(rectangle1_heights[844]), .rectangle1_weight(rectangle1_weights[844]), .rectangle2_x(rectangle2_xs[844]), .rectangle2_y(rectangle2_ys[844]), .rectangle2_width(rectangle2_widths[844]), .rectangle2_height(rectangle2_heights[844]), .rectangle2_weight(rectangle2_weights[844]), .rectangle3_x(rectangle3_xs[844]), .rectangle3_y(rectangle3_ys[844]), .rectangle3_width(rectangle3_widths[844]), .rectangle3_height(rectangle3_heights[844]), .rectangle3_weight(rectangle3_weights[844]), .feature_threshold(feature_thresholds[844]), .feature_above(feature_aboves[844]), .feature_below(feature_belows[844]), .scan_win_std_dev(scan_win_std_dev[844]), .feature_accum(feature_accums[844]));
  accum_calculator ac845(.scan_win(scan_win845), .rectangle1_x(rectangle1_xs[845]), .rectangle1_y(rectangle1_ys[845]), .rectangle1_width(rectangle1_widths[845]), .rectangle1_height(rectangle1_heights[845]), .rectangle1_weight(rectangle1_weights[845]), .rectangle2_x(rectangle2_xs[845]), .rectangle2_y(rectangle2_ys[845]), .rectangle2_width(rectangle2_widths[845]), .rectangle2_height(rectangle2_heights[845]), .rectangle2_weight(rectangle2_weights[845]), .rectangle3_x(rectangle3_xs[845]), .rectangle3_y(rectangle3_ys[845]), .rectangle3_width(rectangle3_widths[845]), .rectangle3_height(rectangle3_heights[845]), .rectangle3_weight(rectangle3_weights[845]), .feature_threshold(feature_thresholds[845]), .feature_above(feature_aboves[845]), .feature_below(feature_belows[845]), .scan_win_std_dev(scan_win_std_dev[845]), .feature_accum(feature_accums[845]));
  accum_calculator ac846(.scan_win(scan_win846), .rectangle1_x(rectangle1_xs[846]), .rectangle1_y(rectangle1_ys[846]), .rectangle1_width(rectangle1_widths[846]), .rectangle1_height(rectangle1_heights[846]), .rectangle1_weight(rectangle1_weights[846]), .rectangle2_x(rectangle2_xs[846]), .rectangle2_y(rectangle2_ys[846]), .rectangle2_width(rectangle2_widths[846]), .rectangle2_height(rectangle2_heights[846]), .rectangle2_weight(rectangle2_weights[846]), .rectangle3_x(rectangle3_xs[846]), .rectangle3_y(rectangle3_ys[846]), .rectangle3_width(rectangle3_widths[846]), .rectangle3_height(rectangle3_heights[846]), .rectangle3_weight(rectangle3_weights[846]), .feature_threshold(feature_thresholds[846]), .feature_above(feature_aboves[846]), .feature_below(feature_belows[846]), .scan_win_std_dev(scan_win_std_dev[846]), .feature_accum(feature_accums[846]));
  accum_calculator ac847(.scan_win(scan_win847), .rectangle1_x(rectangle1_xs[847]), .rectangle1_y(rectangle1_ys[847]), .rectangle1_width(rectangle1_widths[847]), .rectangle1_height(rectangle1_heights[847]), .rectangle1_weight(rectangle1_weights[847]), .rectangle2_x(rectangle2_xs[847]), .rectangle2_y(rectangle2_ys[847]), .rectangle2_width(rectangle2_widths[847]), .rectangle2_height(rectangle2_heights[847]), .rectangle2_weight(rectangle2_weights[847]), .rectangle3_x(rectangle3_xs[847]), .rectangle3_y(rectangle3_ys[847]), .rectangle3_width(rectangle3_widths[847]), .rectangle3_height(rectangle3_heights[847]), .rectangle3_weight(rectangle3_weights[847]), .feature_threshold(feature_thresholds[847]), .feature_above(feature_aboves[847]), .feature_below(feature_belows[847]), .scan_win_std_dev(scan_win_std_dev[847]), .feature_accum(feature_accums[847]));
  accum_calculator ac848(.scan_win(scan_win848), .rectangle1_x(rectangle1_xs[848]), .rectangle1_y(rectangle1_ys[848]), .rectangle1_width(rectangle1_widths[848]), .rectangle1_height(rectangle1_heights[848]), .rectangle1_weight(rectangle1_weights[848]), .rectangle2_x(rectangle2_xs[848]), .rectangle2_y(rectangle2_ys[848]), .rectangle2_width(rectangle2_widths[848]), .rectangle2_height(rectangle2_heights[848]), .rectangle2_weight(rectangle2_weights[848]), .rectangle3_x(rectangle3_xs[848]), .rectangle3_y(rectangle3_ys[848]), .rectangle3_width(rectangle3_widths[848]), .rectangle3_height(rectangle3_heights[848]), .rectangle3_weight(rectangle3_weights[848]), .feature_threshold(feature_thresholds[848]), .feature_above(feature_aboves[848]), .feature_below(feature_belows[848]), .scan_win_std_dev(scan_win_std_dev[848]), .feature_accum(feature_accums[848]));
  accum_calculator ac849(.scan_win(scan_win849), .rectangle1_x(rectangle1_xs[849]), .rectangle1_y(rectangle1_ys[849]), .rectangle1_width(rectangle1_widths[849]), .rectangle1_height(rectangle1_heights[849]), .rectangle1_weight(rectangle1_weights[849]), .rectangle2_x(rectangle2_xs[849]), .rectangle2_y(rectangle2_ys[849]), .rectangle2_width(rectangle2_widths[849]), .rectangle2_height(rectangle2_heights[849]), .rectangle2_weight(rectangle2_weights[849]), .rectangle3_x(rectangle3_xs[849]), .rectangle3_y(rectangle3_ys[849]), .rectangle3_width(rectangle3_widths[849]), .rectangle3_height(rectangle3_heights[849]), .rectangle3_weight(rectangle3_weights[849]), .feature_threshold(feature_thresholds[849]), .feature_above(feature_aboves[849]), .feature_below(feature_belows[849]), .scan_win_std_dev(scan_win_std_dev[849]), .feature_accum(feature_accums[849]));
  accum_calculator ac850(.scan_win(scan_win850), .rectangle1_x(rectangle1_xs[850]), .rectangle1_y(rectangle1_ys[850]), .rectangle1_width(rectangle1_widths[850]), .rectangle1_height(rectangle1_heights[850]), .rectangle1_weight(rectangle1_weights[850]), .rectangle2_x(rectangle2_xs[850]), .rectangle2_y(rectangle2_ys[850]), .rectangle2_width(rectangle2_widths[850]), .rectangle2_height(rectangle2_heights[850]), .rectangle2_weight(rectangle2_weights[850]), .rectangle3_x(rectangle3_xs[850]), .rectangle3_y(rectangle3_ys[850]), .rectangle3_width(rectangle3_widths[850]), .rectangle3_height(rectangle3_heights[850]), .rectangle3_weight(rectangle3_weights[850]), .feature_threshold(feature_thresholds[850]), .feature_above(feature_aboves[850]), .feature_below(feature_belows[850]), .scan_win_std_dev(scan_win_std_dev[850]), .feature_accum(feature_accums[850]));
  accum_calculator ac851(.scan_win(scan_win851), .rectangle1_x(rectangle1_xs[851]), .rectangle1_y(rectangle1_ys[851]), .rectangle1_width(rectangle1_widths[851]), .rectangle1_height(rectangle1_heights[851]), .rectangle1_weight(rectangle1_weights[851]), .rectangle2_x(rectangle2_xs[851]), .rectangle2_y(rectangle2_ys[851]), .rectangle2_width(rectangle2_widths[851]), .rectangle2_height(rectangle2_heights[851]), .rectangle2_weight(rectangle2_weights[851]), .rectangle3_x(rectangle3_xs[851]), .rectangle3_y(rectangle3_ys[851]), .rectangle3_width(rectangle3_widths[851]), .rectangle3_height(rectangle3_heights[851]), .rectangle3_weight(rectangle3_weights[851]), .feature_threshold(feature_thresholds[851]), .feature_above(feature_aboves[851]), .feature_below(feature_belows[851]), .scan_win_std_dev(scan_win_std_dev[851]), .feature_accum(feature_accums[851]));
  accum_calculator ac852(.scan_win(scan_win852), .rectangle1_x(rectangle1_xs[852]), .rectangle1_y(rectangle1_ys[852]), .rectangle1_width(rectangle1_widths[852]), .rectangle1_height(rectangle1_heights[852]), .rectangle1_weight(rectangle1_weights[852]), .rectangle2_x(rectangle2_xs[852]), .rectangle2_y(rectangle2_ys[852]), .rectangle2_width(rectangle2_widths[852]), .rectangle2_height(rectangle2_heights[852]), .rectangle2_weight(rectangle2_weights[852]), .rectangle3_x(rectangle3_xs[852]), .rectangle3_y(rectangle3_ys[852]), .rectangle3_width(rectangle3_widths[852]), .rectangle3_height(rectangle3_heights[852]), .rectangle3_weight(rectangle3_weights[852]), .feature_threshold(feature_thresholds[852]), .feature_above(feature_aboves[852]), .feature_below(feature_belows[852]), .scan_win_std_dev(scan_win_std_dev[852]), .feature_accum(feature_accums[852]));
  accum_calculator ac853(.scan_win(scan_win853), .rectangle1_x(rectangle1_xs[853]), .rectangle1_y(rectangle1_ys[853]), .rectangle1_width(rectangle1_widths[853]), .rectangle1_height(rectangle1_heights[853]), .rectangle1_weight(rectangle1_weights[853]), .rectangle2_x(rectangle2_xs[853]), .rectangle2_y(rectangle2_ys[853]), .rectangle2_width(rectangle2_widths[853]), .rectangle2_height(rectangle2_heights[853]), .rectangle2_weight(rectangle2_weights[853]), .rectangle3_x(rectangle3_xs[853]), .rectangle3_y(rectangle3_ys[853]), .rectangle3_width(rectangle3_widths[853]), .rectangle3_height(rectangle3_heights[853]), .rectangle3_weight(rectangle3_weights[853]), .feature_threshold(feature_thresholds[853]), .feature_above(feature_aboves[853]), .feature_below(feature_belows[853]), .scan_win_std_dev(scan_win_std_dev[853]), .feature_accum(feature_accums[853]));
  accum_calculator ac854(.scan_win(scan_win854), .rectangle1_x(rectangle1_xs[854]), .rectangle1_y(rectangle1_ys[854]), .rectangle1_width(rectangle1_widths[854]), .rectangle1_height(rectangle1_heights[854]), .rectangle1_weight(rectangle1_weights[854]), .rectangle2_x(rectangle2_xs[854]), .rectangle2_y(rectangle2_ys[854]), .rectangle2_width(rectangle2_widths[854]), .rectangle2_height(rectangle2_heights[854]), .rectangle2_weight(rectangle2_weights[854]), .rectangle3_x(rectangle3_xs[854]), .rectangle3_y(rectangle3_ys[854]), .rectangle3_width(rectangle3_widths[854]), .rectangle3_height(rectangle3_heights[854]), .rectangle3_weight(rectangle3_weights[854]), .feature_threshold(feature_thresholds[854]), .feature_above(feature_aboves[854]), .feature_below(feature_belows[854]), .scan_win_std_dev(scan_win_std_dev[854]), .feature_accum(feature_accums[854]));
  accum_calculator ac855(.scan_win(scan_win855), .rectangle1_x(rectangle1_xs[855]), .rectangle1_y(rectangle1_ys[855]), .rectangle1_width(rectangle1_widths[855]), .rectangle1_height(rectangle1_heights[855]), .rectangle1_weight(rectangle1_weights[855]), .rectangle2_x(rectangle2_xs[855]), .rectangle2_y(rectangle2_ys[855]), .rectangle2_width(rectangle2_widths[855]), .rectangle2_height(rectangle2_heights[855]), .rectangle2_weight(rectangle2_weights[855]), .rectangle3_x(rectangle3_xs[855]), .rectangle3_y(rectangle3_ys[855]), .rectangle3_width(rectangle3_widths[855]), .rectangle3_height(rectangle3_heights[855]), .rectangle3_weight(rectangle3_weights[855]), .feature_threshold(feature_thresholds[855]), .feature_above(feature_aboves[855]), .feature_below(feature_belows[855]), .scan_win_std_dev(scan_win_std_dev[855]), .feature_accum(feature_accums[855]));
  accum_calculator ac856(.scan_win(scan_win856), .rectangle1_x(rectangle1_xs[856]), .rectangle1_y(rectangle1_ys[856]), .rectangle1_width(rectangle1_widths[856]), .rectangle1_height(rectangle1_heights[856]), .rectangle1_weight(rectangle1_weights[856]), .rectangle2_x(rectangle2_xs[856]), .rectangle2_y(rectangle2_ys[856]), .rectangle2_width(rectangle2_widths[856]), .rectangle2_height(rectangle2_heights[856]), .rectangle2_weight(rectangle2_weights[856]), .rectangle3_x(rectangle3_xs[856]), .rectangle3_y(rectangle3_ys[856]), .rectangle3_width(rectangle3_widths[856]), .rectangle3_height(rectangle3_heights[856]), .rectangle3_weight(rectangle3_weights[856]), .feature_threshold(feature_thresholds[856]), .feature_above(feature_aboves[856]), .feature_below(feature_belows[856]), .scan_win_std_dev(scan_win_std_dev[856]), .feature_accum(feature_accums[856]));
  accum_calculator ac857(.scan_win(scan_win857), .rectangle1_x(rectangle1_xs[857]), .rectangle1_y(rectangle1_ys[857]), .rectangle1_width(rectangle1_widths[857]), .rectangle1_height(rectangle1_heights[857]), .rectangle1_weight(rectangle1_weights[857]), .rectangle2_x(rectangle2_xs[857]), .rectangle2_y(rectangle2_ys[857]), .rectangle2_width(rectangle2_widths[857]), .rectangle2_height(rectangle2_heights[857]), .rectangle2_weight(rectangle2_weights[857]), .rectangle3_x(rectangle3_xs[857]), .rectangle3_y(rectangle3_ys[857]), .rectangle3_width(rectangle3_widths[857]), .rectangle3_height(rectangle3_heights[857]), .rectangle3_weight(rectangle3_weights[857]), .feature_threshold(feature_thresholds[857]), .feature_above(feature_aboves[857]), .feature_below(feature_belows[857]), .scan_win_std_dev(scan_win_std_dev[857]), .feature_accum(feature_accums[857]));
  accum_calculator ac858(.scan_win(scan_win858), .rectangle1_x(rectangle1_xs[858]), .rectangle1_y(rectangle1_ys[858]), .rectangle1_width(rectangle1_widths[858]), .rectangle1_height(rectangle1_heights[858]), .rectangle1_weight(rectangle1_weights[858]), .rectangle2_x(rectangle2_xs[858]), .rectangle2_y(rectangle2_ys[858]), .rectangle2_width(rectangle2_widths[858]), .rectangle2_height(rectangle2_heights[858]), .rectangle2_weight(rectangle2_weights[858]), .rectangle3_x(rectangle3_xs[858]), .rectangle3_y(rectangle3_ys[858]), .rectangle3_width(rectangle3_widths[858]), .rectangle3_height(rectangle3_heights[858]), .rectangle3_weight(rectangle3_weights[858]), .feature_threshold(feature_thresholds[858]), .feature_above(feature_aboves[858]), .feature_below(feature_belows[858]), .scan_win_std_dev(scan_win_std_dev[858]), .feature_accum(feature_accums[858]));
  accum_calculator ac859(.scan_win(scan_win859), .rectangle1_x(rectangle1_xs[859]), .rectangle1_y(rectangle1_ys[859]), .rectangle1_width(rectangle1_widths[859]), .rectangle1_height(rectangle1_heights[859]), .rectangle1_weight(rectangle1_weights[859]), .rectangle2_x(rectangle2_xs[859]), .rectangle2_y(rectangle2_ys[859]), .rectangle2_width(rectangle2_widths[859]), .rectangle2_height(rectangle2_heights[859]), .rectangle2_weight(rectangle2_weights[859]), .rectangle3_x(rectangle3_xs[859]), .rectangle3_y(rectangle3_ys[859]), .rectangle3_width(rectangle3_widths[859]), .rectangle3_height(rectangle3_heights[859]), .rectangle3_weight(rectangle3_weights[859]), .feature_threshold(feature_thresholds[859]), .feature_above(feature_aboves[859]), .feature_below(feature_belows[859]), .scan_win_std_dev(scan_win_std_dev[859]), .feature_accum(feature_accums[859]));
  accum_calculator ac860(.scan_win(scan_win860), .rectangle1_x(rectangle1_xs[860]), .rectangle1_y(rectangle1_ys[860]), .rectangle1_width(rectangle1_widths[860]), .rectangle1_height(rectangle1_heights[860]), .rectangle1_weight(rectangle1_weights[860]), .rectangle2_x(rectangle2_xs[860]), .rectangle2_y(rectangle2_ys[860]), .rectangle2_width(rectangle2_widths[860]), .rectangle2_height(rectangle2_heights[860]), .rectangle2_weight(rectangle2_weights[860]), .rectangle3_x(rectangle3_xs[860]), .rectangle3_y(rectangle3_ys[860]), .rectangle3_width(rectangle3_widths[860]), .rectangle3_height(rectangle3_heights[860]), .rectangle3_weight(rectangle3_weights[860]), .feature_threshold(feature_thresholds[860]), .feature_above(feature_aboves[860]), .feature_below(feature_belows[860]), .scan_win_std_dev(scan_win_std_dev[860]), .feature_accum(feature_accums[860]));
  accum_calculator ac861(.scan_win(scan_win861), .rectangle1_x(rectangle1_xs[861]), .rectangle1_y(rectangle1_ys[861]), .rectangle1_width(rectangle1_widths[861]), .rectangle1_height(rectangle1_heights[861]), .rectangle1_weight(rectangle1_weights[861]), .rectangle2_x(rectangle2_xs[861]), .rectangle2_y(rectangle2_ys[861]), .rectangle2_width(rectangle2_widths[861]), .rectangle2_height(rectangle2_heights[861]), .rectangle2_weight(rectangle2_weights[861]), .rectangle3_x(rectangle3_xs[861]), .rectangle3_y(rectangle3_ys[861]), .rectangle3_width(rectangle3_widths[861]), .rectangle3_height(rectangle3_heights[861]), .rectangle3_weight(rectangle3_weights[861]), .feature_threshold(feature_thresholds[861]), .feature_above(feature_aboves[861]), .feature_below(feature_belows[861]), .scan_win_std_dev(scan_win_std_dev[861]), .feature_accum(feature_accums[861]));
  accum_calculator ac862(.scan_win(scan_win862), .rectangle1_x(rectangle1_xs[862]), .rectangle1_y(rectangle1_ys[862]), .rectangle1_width(rectangle1_widths[862]), .rectangle1_height(rectangle1_heights[862]), .rectangle1_weight(rectangle1_weights[862]), .rectangle2_x(rectangle2_xs[862]), .rectangle2_y(rectangle2_ys[862]), .rectangle2_width(rectangle2_widths[862]), .rectangle2_height(rectangle2_heights[862]), .rectangle2_weight(rectangle2_weights[862]), .rectangle3_x(rectangle3_xs[862]), .rectangle3_y(rectangle3_ys[862]), .rectangle3_width(rectangle3_widths[862]), .rectangle3_height(rectangle3_heights[862]), .rectangle3_weight(rectangle3_weights[862]), .feature_threshold(feature_thresholds[862]), .feature_above(feature_aboves[862]), .feature_below(feature_belows[862]), .scan_win_std_dev(scan_win_std_dev[862]), .feature_accum(feature_accums[862]));
  accum_calculator ac863(.scan_win(scan_win863), .rectangle1_x(rectangle1_xs[863]), .rectangle1_y(rectangle1_ys[863]), .rectangle1_width(rectangle1_widths[863]), .rectangle1_height(rectangle1_heights[863]), .rectangle1_weight(rectangle1_weights[863]), .rectangle2_x(rectangle2_xs[863]), .rectangle2_y(rectangle2_ys[863]), .rectangle2_width(rectangle2_widths[863]), .rectangle2_height(rectangle2_heights[863]), .rectangle2_weight(rectangle2_weights[863]), .rectangle3_x(rectangle3_xs[863]), .rectangle3_y(rectangle3_ys[863]), .rectangle3_width(rectangle3_widths[863]), .rectangle3_height(rectangle3_heights[863]), .rectangle3_weight(rectangle3_weights[863]), .feature_threshold(feature_thresholds[863]), .feature_above(feature_aboves[863]), .feature_below(feature_belows[863]), .scan_win_std_dev(scan_win_std_dev[863]), .feature_accum(feature_accums[863]));
  accum_calculator ac864(.scan_win(scan_win864), .rectangle1_x(rectangle1_xs[864]), .rectangle1_y(rectangle1_ys[864]), .rectangle1_width(rectangle1_widths[864]), .rectangle1_height(rectangle1_heights[864]), .rectangle1_weight(rectangle1_weights[864]), .rectangle2_x(rectangle2_xs[864]), .rectangle2_y(rectangle2_ys[864]), .rectangle2_width(rectangle2_widths[864]), .rectangle2_height(rectangle2_heights[864]), .rectangle2_weight(rectangle2_weights[864]), .rectangle3_x(rectangle3_xs[864]), .rectangle3_y(rectangle3_ys[864]), .rectangle3_width(rectangle3_widths[864]), .rectangle3_height(rectangle3_heights[864]), .rectangle3_weight(rectangle3_weights[864]), .feature_threshold(feature_thresholds[864]), .feature_above(feature_aboves[864]), .feature_below(feature_belows[864]), .scan_win_std_dev(scan_win_std_dev[864]), .feature_accum(feature_accums[864]));
  accum_calculator ac865(.scan_win(scan_win865), .rectangle1_x(rectangle1_xs[865]), .rectangle1_y(rectangle1_ys[865]), .rectangle1_width(rectangle1_widths[865]), .rectangle1_height(rectangle1_heights[865]), .rectangle1_weight(rectangle1_weights[865]), .rectangle2_x(rectangle2_xs[865]), .rectangle2_y(rectangle2_ys[865]), .rectangle2_width(rectangle2_widths[865]), .rectangle2_height(rectangle2_heights[865]), .rectangle2_weight(rectangle2_weights[865]), .rectangle3_x(rectangle3_xs[865]), .rectangle3_y(rectangle3_ys[865]), .rectangle3_width(rectangle3_widths[865]), .rectangle3_height(rectangle3_heights[865]), .rectangle3_weight(rectangle3_weights[865]), .feature_threshold(feature_thresholds[865]), .feature_above(feature_aboves[865]), .feature_below(feature_belows[865]), .scan_win_std_dev(scan_win_std_dev[865]), .feature_accum(feature_accums[865]));
  accum_calculator ac866(.scan_win(scan_win866), .rectangle1_x(rectangle1_xs[866]), .rectangle1_y(rectangle1_ys[866]), .rectangle1_width(rectangle1_widths[866]), .rectangle1_height(rectangle1_heights[866]), .rectangle1_weight(rectangle1_weights[866]), .rectangle2_x(rectangle2_xs[866]), .rectangle2_y(rectangle2_ys[866]), .rectangle2_width(rectangle2_widths[866]), .rectangle2_height(rectangle2_heights[866]), .rectangle2_weight(rectangle2_weights[866]), .rectangle3_x(rectangle3_xs[866]), .rectangle3_y(rectangle3_ys[866]), .rectangle3_width(rectangle3_widths[866]), .rectangle3_height(rectangle3_heights[866]), .rectangle3_weight(rectangle3_weights[866]), .feature_threshold(feature_thresholds[866]), .feature_above(feature_aboves[866]), .feature_below(feature_belows[866]), .scan_win_std_dev(scan_win_std_dev[866]), .feature_accum(feature_accums[866]));
  accum_calculator ac867(.scan_win(scan_win867), .rectangle1_x(rectangle1_xs[867]), .rectangle1_y(rectangle1_ys[867]), .rectangle1_width(rectangle1_widths[867]), .rectangle1_height(rectangle1_heights[867]), .rectangle1_weight(rectangle1_weights[867]), .rectangle2_x(rectangle2_xs[867]), .rectangle2_y(rectangle2_ys[867]), .rectangle2_width(rectangle2_widths[867]), .rectangle2_height(rectangle2_heights[867]), .rectangle2_weight(rectangle2_weights[867]), .rectangle3_x(rectangle3_xs[867]), .rectangle3_y(rectangle3_ys[867]), .rectangle3_width(rectangle3_widths[867]), .rectangle3_height(rectangle3_heights[867]), .rectangle3_weight(rectangle3_weights[867]), .feature_threshold(feature_thresholds[867]), .feature_above(feature_aboves[867]), .feature_below(feature_belows[867]), .scan_win_std_dev(scan_win_std_dev[867]), .feature_accum(feature_accums[867]));
  accum_calculator ac868(.scan_win(scan_win868), .rectangle1_x(rectangle1_xs[868]), .rectangle1_y(rectangle1_ys[868]), .rectangle1_width(rectangle1_widths[868]), .rectangle1_height(rectangle1_heights[868]), .rectangle1_weight(rectangle1_weights[868]), .rectangle2_x(rectangle2_xs[868]), .rectangle2_y(rectangle2_ys[868]), .rectangle2_width(rectangle2_widths[868]), .rectangle2_height(rectangle2_heights[868]), .rectangle2_weight(rectangle2_weights[868]), .rectangle3_x(rectangle3_xs[868]), .rectangle3_y(rectangle3_ys[868]), .rectangle3_width(rectangle3_widths[868]), .rectangle3_height(rectangle3_heights[868]), .rectangle3_weight(rectangle3_weights[868]), .feature_threshold(feature_thresholds[868]), .feature_above(feature_aboves[868]), .feature_below(feature_belows[868]), .scan_win_std_dev(scan_win_std_dev[868]), .feature_accum(feature_accums[868]));
  accum_calculator ac869(.scan_win(scan_win869), .rectangle1_x(rectangle1_xs[869]), .rectangle1_y(rectangle1_ys[869]), .rectangle1_width(rectangle1_widths[869]), .rectangle1_height(rectangle1_heights[869]), .rectangle1_weight(rectangle1_weights[869]), .rectangle2_x(rectangle2_xs[869]), .rectangle2_y(rectangle2_ys[869]), .rectangle2_width(rectangle2_widths[869]), .rectangle2_height(rectangle2_heights[869]), .rectangle2_weight(rectangle2_weights[869]), .rectangle3_x(rectangle3_xs[869]), .rectangle3_y(rectangle3_ys[869]), .rectangle3_width(rectangle3_widths[869]), .rectangle3_height(rectangle3_heights[869]), .rectangle3_weight(rectangle3_weights[869]), .feature_threshold(feature_thresholds[869]), .feature_above(feature_aboves[869]), .feature_below(feature_belows[869]), .scan_win_std_dev(scan_win_std_dev[869]), .feature_accum(feature_accums[869]));
  accum_calculator ac870(.scan_win(scan_win870), .rectangle1_x(rectangle1_xs[870]), .rectangle1_y(rectangle1_ys[870]), .rectangle1_width(rectangle1_widths[870]), .rectangle1_height(rectangle1_heights[870]), .rectangle1_weight(rectangle1_weights[870]), .rectangle2_x(rectangle2_xs[870]), .rectangle2_y(rectangle2_ys[870]), .rectangle2_width(rectangle2_widths[870]), .rectangle2_height(rectangle2_heights[870]), .rectangle2_weight(rectangle2_weights[870]), .rectangle3_x(rectangle3_xs[870]), .rectangle3_y(rectangle3_ys[870]), .rectangle3_width(rectangle3_widths[870]), .rectangle3_height(rectangle3_heights[870]), .rectangle3_weight(rectangle3_weights[870]), .feature_threshold(feature_thresholds[870]), .feature_above(feature_aboves[870]), .feature_below(feature_belows[870]), .scan_win_std_dev(scan_win_std_dev[870]), .feature_accum(feature_accums[870]));
  accum_calculator ac871(.scan_win(scan_win871), .rectangle1_x(rectangle1_xs[871]), .rectangle1_y(rectangle1_ys[871]), .rectangle1_width(rectangle1_widths[871]), .rectangle1_height(rectangle1_heights[871]), .rectangle1_weight(rectangle1_weights[871]), .rectangle2_x(rectangle2_xs[871]), .rectangle2_y(rectangle2_ys[871]), .rectangle2_width(rectangle2_widths[871]), .rectangle2_height(rectangle2_heights[871]), .rectangle2_weight(rectangle2_weights[871]), .rectangle3_x(rectangle3_xs[871]), .rectangle3_y(rectangle3_ys[871]), .rectangle3_width(rectangle3_widths[871]), .rectangle3_height(rectangle3_heights[871]), .rectangle3_weight(rectangle3_weights[871]), .feature_threshold(feature_thresholds[871]), .feature_above(feature_aboves[871]), .feature_below(feature_belows[871]), .scan_win_std_dev(scan_win_std_dev[871]), .feature_accum(feature_accums[871]));
  accum_calculator ac872(.scan_win(scan_win872), .rectangle1_x(rectangle1_xs[872]), .rectangle1_y(rectangle1_ys[872]), .rectangle1_width(rectangle1_widths[872]), .rectangle1_height(rectangle1_heights[872]), .rectangle1_weight(rectangle1_weights[872]), .rectangle2_x(rectangle2_xs[872]), .rectangle2_y(rectangle2_ys[872]), .rectangle2_width(rectangle2_widths[872]), .rectangle2_height(rectangle2_heights[872]), .rectangle2_weight(rectangle2_weights[872]), .rectangle3_x(rectangle3_xs[872]), .rectangle3_y(rectangle3_ys[872]), .rectangle3_width(rectangle3_widths[872]), .rectangle3_height(rectangle3_heights[872]), .rectangle3_weight(rectangle3_weights[872]), .feature_threshold(feature_thresholds[872]), .feature_above(feature_aboves[872]), .feature_below(feature_belows[872]), .scan_win_std_dev(scan_win_std_dev[872]), .feature_accum(feature_accums[872]));
  accum_calculator ac873(.scan_win(scan_win873), .rectangle1_x(rectangle1_xs[873]), .rectangle1_y(rectangle1_ys[873]), .rectangle1_width(rectangle1_widths[873]), .rectangle1_height(rectangle1_heights[873]), .rectangle1_weight(rectangle1_weights[873]), .rectangle2_x(rectangle2_xs[873]), .rectangle2_y(rectangle2_ys[873]), .rectangle2_width(rectangle2_widths[873]), .rectangle2_height(rectangle2_heights[873]), .rectangle2_weight(rectangle2_weights[873]), .rectangle3_x(rectangle3_xs[873]), .rectangle3_y(rectangle3_ys[873]), .rectangle3_width(rectangle3_widths[873]), .rectangle3_height(rectangle3_heights[873]), .rectangle3_weight(rectangle3_weights[873]), .feature_threshold(feature_thresholds[873]), .feature_above(feature_aboves[873]), .feature_below(feature_belows[873]), .scan_win_std_dev(scan_win_std_dev[873]), .feature_accum(feature_accums[873]));
  accum_calculator ac874(.scan_win(scan_win874), .rectangle1_x(rectangle1_xs[874]), .rectangle1_y(rectangle1_ys[874]), .rectangle1_width(rectangle1_widths[874]), .rectangle1_height(rectangle1_heights[874]), .rectangle1_weight(rectangle1_weights[874]), .rectangle2_x(rectangle2_xs[874]), .rectangle2_y(rectangle2_ys[874]), .rectangle2_width(rectangle2_widths[874]), .rectangle2_height(rectangle2_heights[874]), .rectangle2_weight(rectangle2_weights[874]), .rectangle3_x(rectangle3_xs[874]), .rectangle3_y(rectangle3_ys[874]), .rectangle3_width(rectangle3_widths[874]), .rectangle3_height(rectangle3_heights[874]), .rectangle3_weight(rectangle3_weights[874]), .feature_threshold(feature_thresholds[874]), .feature_above(feature_aboves[874]), .feature_below(feature_belows[874]), .scan_win_std_dev(scan_win_std_dev[874]), .feature_accum(feature_accums[874]));
  accum_calculator ac875(.scan_win(scan_win875), .rectangle1_x(rectangle1_xs[875]), .rectangle1_y(rectangle1_ys[875]), .rectangle1_width(rectangle1_widths[875]), .rectangle1_height(rectangle1_heights[875]), .rectangle1_weight(rectangle1_weights[875]), .rectangle2_x(rectangle2_xs[875]), .rectangle2_y(rectangle2_ys[875]), .rectangle2_width(rectangle2_widths[875]), .rectangle2_height(rectangle2_heights[875]), .rectangle2_weight(rectangle2_weights[875]), .rectangle3_x(rectangle3_xs[875]), .rectangle3_y(rectangle3_ys[875]), .rectangle3_width(rectangle3_widths[875]), .rectangle3_height(rectangle3_heights[875]), .rectangle3_weight(rectangle3_weights[875]), .feature_threshold(feature_thresholds[875]), .feature_above(feature_aboves[875]), .feature_below(feature_belows[875]), .scan_win_std_dev(scan_win_std_dev[875]), .feature_accum(feature_accums[875]));
  accum_calculator ac876(.scan_win(scan_win876), .rectangle1_x(rectangle1_xs[876]), .rectangle1_y(rectangle1_ys[876]), .rectangle1_width(rectangle1_widths[876]), .rectangle1_height(rectangle1_heights[876]), .rectangle1_weight(rectangle1_weights[876]), .rectangle2_x(rectangle2_xs[876]), .rectangle2_y(rectangle2_ys[876]), .rectangle2_width(rectangle2_widths[876]), .rectangle2_height(rectangle2_heights[876]), .rectangle2_weight(rectangle2_weights[876]), .rectangle3_x(rectangle3_xs[876]), .rectangle3_y(rectangle3_ys[876]), .rectangle3_width(rectangle3_widths[876]), .rectangle3_height(rectangle3_heights[876]), .rectangle3_weight(rectangle3_weights[876]), .feature_threshold(feature_thresholds[876]), .feature_above(feature_aboves[876]), .feature_below(feature_belows[876]), .scan_win_std_dev(scan_win_std_dev[876]), .feature_accum(feature_accums[876]));
  accum_calculator ac877(.scan_win(scan_win877), .rectangle1_x(rectangle1_xs[877]), .rectangle1_y(rectangle1_ys[877]), .rectangle1_width(rectangle1_widths[877]), .rectangle1_height(rectangle1_heights[877]), .rectangle1_weight(rectangle1_weights[877]), .rectangle2_x(rectangle2_xs[877]), .rectangle2_y(rectangle2_ys[877]), .rectangle2_width(rectangle2_widths[877]), .rectangle2_height(rectangle2_heights[877]), .rectangle2_weight(rectangle2_weights[877]), .rectangle3_x(rectangle3_xs[877]), .rectangle3_y(rectangle3_ys[877]), .rectangle3_width(rectangle3_widths[877]), .rectangle3_height(rectangle3_heights[877]), .rectangle3_weight(rectangle3_weights[877]), .feature_threshold(feature_thresholds[877]), .feature_above(feature_aboves[877]), .feature_below(feature_belows[877]), .scan_win_std_dev(scan_win_std_dev[877]), .feature_accum(feature_accums[877]));
  accum_calculator ac878(.scan_win(scan_win878), .rectangle1_x(rectangle1_xs[878]), .rectangle1_y(rectangle1_ys[878]), .rectangle1_width(rectangle1_widths[878]), .rectangle1_height(rectangle1_heights[878]), .rectangle1_weight(rectangle1_weights[878]), .rectangle2_x(rectangle2_xs[878]), .rectangle2_y(rectangle2_ys[878]), .rectangle2_width(rectangle2_widths[878]), .rectangle2_height(rectangle2_heights[878]), .rectangle2_weight(rectangle2_weights[878]), .rectangle3_x(rectangle3_xs[878]), .rectangle3_y(rectangle3_ys[878]), .rectangle3_width(rectangle3_widths[878]), .rectangle3_height(rectangle3_heights[878]), .rectangle3_weight(rectangle3_weights[878]), .feature_threshold(feature_thresholds[878]), .feature_above(feature_aboves[878]), .feature_below(feature_belows[878]), .scan_win_std_dev(scan_win_std_dev[878]), .feature_accum(feature_accums[878]));
  accum_calculator ac879(.scan_win(scan_win879), .rectangle1_x(rectangle1_xs[879]), .rectangle1_y(rectangle1_ys[879]), .rectangle1_width(rectangle1_widths[879]), .rectangle1_height(rectangle1_heights[879]), .rectangle1_weight(rectangle1_weights[879]), .rectangle2_x(rectangle2_xs[879]), .rectangle2_y(rectangle2_ys[879]), .rectangle2_width(rectangle2_widths[879]), .rectangle2_height(rectangle2_heights[879]), .rectangle2_weight(rectangle2_weights[879]), .rectangle3_x(rectangle3_xs[879]), .rectangle3_y(rectangle3_ys[879]), .rectangle3_width(rectangle3_widths[879]), .rectangle3_height(rectangle3_heights[879]), .rectangle3_weight(rectangle3_weights[879]), .feature_threshold(feature_thresholds[879]), .feature_above(feature_aboves[879]), .feature_below(feature_belows[879]), .scan_win_std_dev(scan_win_std_dev[879]), .feature_accum(feature_accums[879]));
  accum_calculator ac880(.scan_win(scan_win880), .rectangle1_x(rectangle1_xs[880]), .rectangle1_y(rectangle1_ys[880]), .rectangle1_width(rectangle1_widths[880]), .rectangle1_height(rectangle1_heights[880]), .rectangle1_weight(rectangle1_weights[880]), .rectangle2_x(rectangle2_xs[880]), .rectangle2_y(rectangle2_ys[880]), .rectangle2_width(rectangle2_widths[880]), .rectangle2_height(rectangle2_heights[880]), .rectangle2_weight(rectangle2_weights[880]), .rectangle3_x(rectangle3_xs[880]), .rectangle3_y(rectangle3_ys[880]), .rectangle3_width(rectangle3_widths[880]), .rectangle3_height(rectangle3_heights[880]), .rectangle3_weight(rectangle3_weights[880]), .feature_threshold(feature_thresholds[880]), .feature_above(feature_aboves[880]), .feature_below(feature_belows[880]), .scan_win_std_dev(scan_win_std_dev[880]), .feature_accum(feature_accums[880]));
  accum_calculator ac881(.scan_win(scan_win881), .rectangle1_x(rectangle1_xs[881]), .rectangle1_y(rectangle1_ys[881]), .rectangle1_width(rectangle1_widths[881]), .rectangle1_height(rectangle1_heights[881]), .rectangle1_weight(rectangle1_weights[881]), .rectangle2_x(rectangle2_xs[881]), .rectangle2_y(rectangle2_ys[881]), .rectangle2_width(rectangle2_widths[881]), .rectangle2_height(rectangle2_heights[881]), .rectangle2_weight(rectangle2_weights[881]), .rectangle3_x(rectangle3_xs[881]), .rectangle3_y(rectangle3_ys[881]), .rectangle3_width(rectangle3_widths[881]), .rectangle3_height(rectangle3_heights[881]), .rectangle3_weight(rectangle3_weights[881]), .feature_threshold(feature_thresholds[881]), .feature_above(feature_aboves[881]), .feature_below(feature_belows[881]), .scan_win_std_dev(scan_win_std_dev[881]), .feature_accum(feature_accums[881]));
  accum_calculator ac882(.scan_win(scan_win882), .rectangle1_x(rectangle1_xs[882]), .rectangle1_y(rectangle1_ys[882]), .rectangle1_width(rectangle1_widths[882]), .rectangle1_height(rectangle1_heights[882]), .rectangle1_weight(rectangle1_weights[882]), .rectangle2_x(rectangle2_xs[882]), .rectangle2_y(rectangle2_ys[882]), .rectangle2_width(rectangle2_widths[882]), .rectangle2_height(rectangle2_heights[882]), .rectangle2_weight(rectangle2_weights[882]), .rectangle3_x(rectangle3_xs[882]), .rectangle3_y(rectangle3_ys[882]), .rectangle3_width(rectangle3_widths[882]), .rectangle3_height(rectangle3_heights[882]), .rectangle3_weight(rectangle3_weights[882]), .feature_threshold(feature_thresholds[882]), .feature_above(feature_aboves[882]), .feature_below(feature_belows[882]), .scan_win_std_dev(scan_win_std_dev[882]), .feature_accum(feature_accums[882]));
  accum_calculator ac883(.scan_win(scan_win883), .rectangle1_x(rectangle1_xs[883]), .rectangle1_y(rectangle1_ys[883]), .rectangle1_width(rectangle1_widths[883]), .rectangle1_height(rectangle1_heights[883]), .rectangle1_weight(rectangle1_weights[883]), .rectangle2_x(rectangle2_xs[883]), .rectangle2_y(rectangle2_ys[883]), .rectangle2_width(rectangle2_widths[883]), .rectangle2_height(rectangle2_heights[883]), .rectangle2_weight(rectangle2_weights[883]), .rectangle3_x(rectangle3_xs[883]), .rectangle3_y(rectangle3_ys[883]), .rectangle3_width(rectangle3_widths[883]), .rectangle3_height(rectangle3_heights[883]), .rectangle3_weight(rectangle3_weights[883]), .feature_threshold(feature_thresholds[883]), .feature_above(feature_aboves[883]), .feature_below(feature_belows[883]), .scan_win_std_dev(scan_win_std_dev[883]), .feature_accum(feature_accums[883]));
  accum_calculator ac884(.scan_win(scan_win884), .rectangle1_x(rectangle1_xs[884]), .rectangle1_y(rectangle1_ys[884]), .rectangle1_width(rectangle1_widths[884]), .rectangle1_height(rectangle1_heights[884]), .rectangle1_weight(rectangle1_weights[884]), .rectangle2_x(rectangle2_xs[884]), .rectangle2_y(rectangle2_ys[884]), .rectangle2_width(rectangle2_widths[884]), .rectangle2_height(rectangle2_heights[884]), .rectangle2_weight(rectangle2_weights[884]), .rectangle3_x(rectangle3_xs[884]), .rectangle3_y(rectangle3_ys[884]), .rectangle3_width(rectangle3_widths[884]), .rectangle3_height(rectangle3_heights[884]), .rectangle3_weight(rectangle3_weights[884]), .feature_threshold(feature_thresholds[884]), .feature_above(feature_aboves[884]), .feature_below(feature_belows[884]), .scan_win_std_dev(scan_win_std_dev[884]), .feature_accum(feature_accums[884]));
  accum_calculator ac885(.scan_win(scan_win885), .rectangle1_x(rectangle1_xs[885]), .rectangle1_y(rectangle1_ys[885]), .rectangle1_width(rectangle1_widths[885]), .rectangle1_height(rectangle1_heights[885]), .rectangle1_weight(rectangle1_weights[885]), .rectangle2_x(rectangle2_xs[885]), .rectangle2_y(rectangle2_ys[885]), .rectangle2_width(rectangle2_widths[885]), .rectangle2_height(rectangle2_heights[885]), .rectangle2_weight(rectangle2_weights[885]), .rectangle3_x(rectangle3_xs[885]), .rectangle3_y(rectangle3_ys[885]), .rectangle3_width(rectangle3_widths[885]), .rectangle3_height(rectangle3_heights[885]), .rectangle3_weight(rectangle3_weights[885]), .feature_threshold(feature_thresholds[885]), .feature_above(feature_aboves[885]), .feature_below(feature_belows[885]), .scan_win_std_dev(scan_win_std_dev[885]), .feature_accum(feature_accums[885]));
  accum_calculator ac886(.scan_win(scan_win886), .rectangle1_x(rectangle1_xs[886]), .rectangle1_y(rectangle1_ys[886]), .rectangle1_width(rectangle1_widths[886]), .rectangle1_height(rectangle1_heights[886]), .rectangle1_weight(rectangle1_weights[886]), .rectangle2_x(rectangle2_xs[886]), .rectangle2_y(rectangle2_ys[886]), .rectangle2_width(rectangle2_widths[886]), .rectangle2_height(rectangle2_heights[886]), .rectangle2_weight(rectangle2_weights[886]), .rectangle3_x(rectangle3_xs[886]), .rectangle3_y(rectangle3_ys[886]), .rectangle3_width(rectangle3_widths[886]), .rectangle3_height(rectangle3_heights[886]), .rectangle3_weight(rectangle3_weights[886]), .feature_threshold(feature_thresholds[886]), .feature_above(feature_aboves[886]), .feature_below(feature_belows[886]), .scan_win_std_dev(scan_win_std_dev[886]), .feature_accum(feature_accums[886]));
  accum_calculator ac887(.scan_win(scan_win887), .rectangle1_x(rectangle1_xs[887]), .rectangle1_y(rectangle1_ys[887]), .rectangle1_width(rectangle1_widths[887]), .rectangle1_height(rectangle1_heights[887]), .rectangle1_weight(rectangle1_weights[887]), .rectangle2_x(rectangle2_xs[887]), .rectangle2_y(rectangle2_ys[887]), .rectangle2_width(rectangle2_widths[887]), .rectangle2_height(rectangle2_heights[887]), .rectangle2_weight(rectangle2_weights[887]), .rectangle3_x(rectangle3_xs[887]), .rectangle3_y(rectangle3_ys[887]), .rectangle3_width(rectangle3_widths[887]), .rectangle3_height(rectangle3_heights[887]), .rectangle3_weight(rectangle3_weights[887]), .feature_threshold(feature_thresholds[887]), .feature_above(feature_aboves[887]), .feature_below(feature_belows[887]), .scan_win_std_dev(scan_win_std_dev[887]), .feature_accum(feature_accums[887]));
  accum_calculator ac888(.scan_win(scan_win888), .rectangle1_x(rectangle1_xs[888]), .rectangle1_y(rectangle1_ys[888]), .rectangle1_width(rectangle1_widths[888]), .rectangle1_height(rectangle1_heights[888]), .rectangle1_weight(rectangle1_weights[888]), .rectangle2_x(rectangle2_xs[888]), .rectangle2_y(rectangle2_ys[888]), .rectangle2_width(rectangle2_widths[888]), .rectangle2_height(rectangle2_heights[888]), .rectangle2_weight(rectangle2_weights[888]), .rectangle3_x(rectangle3_xs[888]), .rectangle3_y(rectangle3_ys[888]), .rectangle3_width(rectangle3_widths[888]), .rectangle3_height(rectangle3_heights[888]), .rectangle3_weight(rectangle3_weights[888]), .feature_threshold(feature_thresholds[888]), .feature_above(feature_aboves[888]), .feature_below(feature_belows[888]), .scan_win_std_dev(scan_win_std_dev[888]), .feature_accum(feature_accums[888]));
  accum_calculator ac889(.scan_win(scan_win889), .rectangle1_x(rectangle1_xs[889]), .rectangle1_y(rectangle1_ys[889]), .rectangle1_width(rectangle1_widths[889]), .rectangle1_height(rectangle1_heights[889]), .rectangle1_weight(rectangle1_weights[889]), .rectangle2_x(rectangle2_xs[889]), .rectangle2_y(rectangle2_ys[889]), .rectangle2_width(rectangle2_widths[889]), .rectangle2_height(rectangle2_heights[889]), .rectangle2_weight(rectangle2_weights[889]), .rectangle3_x(rectangle3_xs[889]), .rectangle3_y(rectangle3_ys[889]), .rectangle3_width(rectangle3_widths[889]), .rectangle3_height(rectangle3_heights[889]), .rectangle3_weight(rectangle3_weights[889]), .feature_threshold(feature_thresholds[889]), .feature_above(feature_aboves[889]), .feature_below(feature_belows[889]), .scan_win_std_dev(scan_win_std_dev[889]), .feature_accum(feature_accums[889]));
  accum_calculator ac890(.scan_win(scan_win890), .rectangle1_x(rectangle1_xs[890]), .rectangle1_y(rectangle1_ys[890]), .rectangle1_width(rectangle1_widths[890]), .rectangle1_height(rectangle1_heights[890]), .rectangle1_weight(rectangle1_weights[890]), .rectangle2_x(rectangle2_xs[890]), .rectangle2_y(rectangle2_ys[890]), .rectangle2_width(rectangle2_widths[890]), .rectangle2_height(rectangle2_heights[890]), .rectangle2_weight(rectangle2_weights[890]), .rectangle3_x(rectangle3_xs[890]), .rectangle3_y(rectangle3_ys[890]), .rectangle3_width(rectangle3_widths[890]), .rectangle3_height(rectangle3_heights[890]), .rectangle3_weight(rectangle3_weights[890]), .feature_threshold(feature_thresholds[890]), .feature_above(feature_aboves[890]), .feature_below(feature_belows[890]), .scan_win_std_dev(scan_win_std_dev[890]), .feature_accum(feature_accums[890]));
  accum_calculator ac891(.scan_win(scan_win891), .rectangle1_x(rectangle1_xs[891]), .rectangle1_y(rectangle1_ys[891]), .rectangle1_width(rectangle1_widths[891]), .rectangle1_height(rectangle1_heights[891]), .rectangle1_weight(rectangle1_weights[891]), .rectangle2_x(rectangle2_xs[891]), .rectangle2_y(rectangle2_ys[891]), .rectangle2_width(rectangle2_widths[891]), .rectangle2_height(rectangle2_heights[891]), .rectangle2_weight(rectangle2_weights[891]), .rectangle3_x(rectangle3_xs[891]), .rectangle3_y(rectangle3_ys[891]), .rectangle3_width(rectangle3_widths[891]), .rectangle3_height(rectangle3_heights[891]), .rectangle3_weight(rectangle3_weights[891]), .feature_threshold(feature_thresholds[891]), .feature_above(feature_aboves[891]), .feature_below(feature_belows[891]), .scan_win_std_dev(scan_win_std_dev[891]), .feature_accum(feature_accums[891]));
  accum_calculator ac892(.scan_win(scan_win892), .rectangle1_x(rectangle1_xs[892]), .rectangle1_y(rectangle1_ys[892]), .rectangle1_width(rectangle1_widths[892]), .rectangle1_height(rectangle1_heights[892]), .rectangle1_weight(rectangle1_weights[892]), .rectangle2_x(rectangle2_xs[892]), .rectangle2_y(rectangle2_ys[892]), .rectangle2_width(rectangle2_widths[892]), .rectangle2_height(rectangle2_heights[892]), .rectangle2_weight(rectangle2_weights[892]), .rectangle3_x(rectangle3_xs[892]), .rectangle3_y(rectangle3_ys[892]), .rectangle3_width(rectangle3_widths[892]), .rectangle3_height(rectangle3_heights[892]), .rectangle3_weight(rectangle3_weights[892]), .feature_threshold(feature_thresholds[892]), .feature_above(feature_aboves[892]), .feature_below(feature_belows[892]), .scan_win_std_dev(scan_win_std_dev[892]), .feature_accum(feature_accums[892]));
  accum_calculator ac893(.scan_win(scan_win893), .rectangle1_x(rectangle1_xs[893]), .rectangle1_y(rectangle1_ys[893]), .rectangle1_width(rectangle1_widths[893]), .rectangle1_height(rectangle1_heights[893]), .rectangle1_weight(rectangle1_weights[893]), .rectangle2_x(rectangle2_xs[893]), .rectangle2_y(rectangle2_ys[893]), .rectangle2_width(rectangle2_widths[893]), .rectangle2_height(rectangle2_heights[893]), .rectangle2_weight(rectangle2_weights[893]), .rectangle3_x(rectangle3_xs[893]), .rectangle3_y(rectangle3_ys[893]), .rectangle3_width(rectangle3_widths[893]), .rectangle3_height(rectangle3_heights[893]), .rectangle3_weight(rectangle3_weights[893]), .feature_threshold(feature_thresholds[893]), .feature_above(feature_aboves[893]), .feature_below(feature_belows[893]), .scan_win_std_dev(scan_win_std_dev[893]), .feature_accum(feature_accums[893]));
  accum_calculator ac894(.scan_win(scan_win894), .rectangle1_x(rectangle1_xs[894]), .rectangle1_y(rectangle1_ys[894]), .rectangle1_width(rectangle1_widths[894]), .rectangle1_height(rectangle1_heights[894]), .rectangle1_weight(rectangle1_weights[894]), .rectangle2_x(rectangle2_xs[894]), .rectangle2_y(rectangle2_ys[894]), .rectangle2_width(rectangle2_widths[894]), .rectangle2_height(rectangle2_heights[894]), .rectangle2_weight(rectangle2_weights[894]), .rectangle3_x(rectangle3_xs[894]), .rectangle3_y(rectangle3_ys[894]), .rectangle3_width(rectangle3_widths[894]), .rectangle3_height(rectangle3_heights[894]), .rectangle3_weight(rectangle3_weights[894]), .feature_threshold(feature_thresholds[894]), .feature_above(feature_aboves[894]), .feature_below(feature_belows[894]), .scan_win_std_dev(scan_win_std_dev[894]), .feature_accum(feature_accums[894]));
  accum_calculator ac895(.scan_win(scan_win895), .rectangle1_x(rectangle1_xs[895]), .rectangle1_y(rectangle1_ys[895]), .rectangle1_width(rectangle1_widths[895]), .rectangle1_height(rectangle1_heights[895]), .rectangle1_weight(rectangle1_weights[895]), .rectangle2_x(rectangle2_xs[895]), .rectangle2_y(rectangle2_ys[895]), .rectangle2_width(rectangle2_widths[895]), .rectangle2_height(rectangle2_heights[895]), .rectangle2_weight(rectangle2_weights[895]), .rectangle3_x(rectangle3_xs[895]), .rectangle3_y(rectangle3_ys[895]), .rectangle3_width(rectangle3_widths[895]), .rectangle3_height(rectangle3_heights[895]), .rectangle3_weight(rectangle3_weights[895]), .feature_threshold(feature_thresholds[895]), .feature_above(feature_aboves[895]), .feature_below(feature_belows[895]), .scan_win_std_dev(scan_win_std_dev[895]), .feature_accum(feature_accums[895]));
  accum_calculator ac896(.scan_win(scan_win896), .rectangle1_x(rectangle1_xs[896]), .rectangle1_y(rectangle1_ys[896]), .rectangle1_width(rectangle1_widths[896]), .rectangle1_height(rectangle1_heights[896]), .rectangle1_weight(rectangle1_weights[896]), .rectangle2_x(rectangle2_xs[896]), .rectangle2_y(rectangle2_ys[896]), .rectangle2_width(rectangle2_widths[896]), .rectangle2_height(rectangle2_heights[896]), .rectangle2_weight(rectangle2_weights[896]), .rectangle3_x(rectangle3_xs[896]), .rectangle3_y(rectangle3_ys[896]), .rectangle3_width(rectangle3_widths[896]), .rectangle3_height(rectangle3_heights[896]), .rectangle3_weight(rectangle3_weights[896]), .feature_threshold(feature_thresholds[896]), .feature_above(feature_aboves[896]), .feature_below(feature_belows[896]), .scan_win_std_dev(scan_win_std_dev[896]), .feature_accum(feature_accums[896]));
  accum_calculator ac897(.scan_win(scan_win897), .rectangle1_x(rectangle1_xs[897]), .rectangle1_y(rectangle1_ys[897]), .rectangle1_width(rectangle1_widths[897]), .rectangle1_height(rectangle1_heights[897]), .rectangle1_weight(rectangle1_weights[897]), .rectangle2_x(rectangle2_xs[897]), .rectangle2_y(rectangle2_ys[897]), .rectangle2_width(rectangle2_widths[897]), .rectangle2_height(rectangle2_heights[897]), .rectangle2_weight(rectangle2_weights[897]), .rectangle3_x(rectangle3_xs[897]), .rectangle3_y(rectangle3_ys[897]), .rectangle3_width(rectangle3_widths[897]), .rectangle3_height(rectangle3_heights[897]), .rectangle3_weight(rectangle3_weights[897]), .feature_threshold(feature_thresholds[897]), .feature_above(feature_aboves[897]), .feature_below(feature_belows[897]), .scan_win_std_dev(scan_win_std_dev[897]), .feature_accum(feature_accums[897]));
  accum_calculator ac898(.scan_win(scan_win898), .rectangle1_x(rectangle1_xs[898]), .rectangle1_y(rectangle1_ys[898]), .rectangle1_width(rectangle1_widths[898]), .rectangle1_height(rectangle1_heights[898]), .rectangle1_weight(rectangle1_weights[898]), .rectangle2_x(rectangle2_xs[898]), .rectangle2_y(rectangle2_ys[898]), .rectangle2_width(rectangle2_widths[898]), .rectangle2_height(rectangle2_heights[898]), .rectangle2_weight(rectangle2_weights[898]), .rectangle3_x(rectangle3_xs[898]), .rectangle3_y(rectangle3_ys[898]), .rectangle3_width(rectangle3_widths[898]), .rectangle3_height(rectangle3_heights[898]), .rectangle3_weight(rectangle3_weights[898]), .feature_threshold(feature_thresholds[898]), .feature_above(feature_aboves[898]), .feature_below(feature_belows[898]), .scan_win_std_dev(scan_win_std_dev[898]), .feature_accum(feature_accums[898]));
  accum_calculator ac899(.scan_win(scan_win899), .rectangle1_x(rectangle1_xs[899]), .rectangle1_y(rectangle1_ys[899]), .rectangle1_width(rectangle1_widths[899]), .rectangle1_height(rectangle1_heights[899]), .rectangle1_weight(rectangle1_weights[899]), .rectangle2_x(rectangle2_xs[899]), .rectangle2_y(rectangle2_ys[899]), .rectangle2_width(rectangle2_widths[899]), .rectangle2_height(rectangle2_heights[899]), .rectangle2_weight(rectangle2_weights[899]), .rectangle3_x(rectangle3_xs[899]), .rectangle3_y(rectangle3_ys[899]), .rectangle3_width(rectangle3_widths[899]), .rectangle3_height(rectangle3_heights[899]), .rectangle3_weight(rectangle3_weights[899]), .feature_threshold(feature_thresholds[899]), .feature_above(feature_aboves[899]), .feature_below(feature_belows[899]), .scan_win_std_dev(scan_win_std_dev[899]), .feature_accum(feature_accums[899]));
  accum_calculator ac900(.scan_win(scan_win900), .rectangle1_x(rectangle1_xs[900]), .rectangle1_y(rectangle1_ys[900]), .rectangle1_width(rectangle1_widths[900]), .rectangle1_height(rectangle1_heights[900]), .rectangle1_weight(rectangle1_weights[900]), .rectangle2_x(rectangle2_xs[900]), .rectangle2_y(rectangle2_ys[900]), .rectangle2_width(rectangle2_widths[900]), .rectangle2_height(rectangle2_heights[900]), .rectangle2_weight(rectangle2_weights[900]), .rectangle3_x(rectangle3_xs[900]), .rectangle3_y(rectangle3_ys[900]), .rectangle3_width(rectangle3_widths[900]), .rectangle3_height(rectangle3_heights[900]), .rectangle3_weight(rectangle3_weights[900]), .feature_threshold(feature_thresholds[900]), .feature_above(feature_aboves[900]), .feature_below(feature_belows[900]), .scan_win_std_dev(scan_win_std_dev[900]), .feature_accum(feature_accums[900]));
  accum_calculator ac901(.scan_win(scan_win901), .rectangle1_x(rectangle1_xs[901]), .rectangle1_y(rectangle1_ys[901]), .rectangle1_width(rectangle1_widths[901]), .rectangle1_height(rectangle1_heights[901]), .rectangle1_weight(rectangle1_weights[901]), .rectangle2_x(rectangle2_xs[901]), .rectangle2_y(rectangle2_ys[901]), .rectangle2_width(rectangle2_widths[901]), .rectangle2_height(rectangle2_heights[901]), .rectangle2_weight(rectangle2_weights[901]), .rectangle3_x(rectangle3_xs[901]), .rectangle3_y(rectangle3_ys[901]), .rectangle3_width(rectangle3_widths[901]), .rectangle3_height(rectangle3_heights[901]), .rectangle3_weight(rectangle3_weights[901]), .feature_threshold(feature_thresholds[901]), .feature_above(feature_aboves[901]), .feature_below(feature_belows[901]), .scan_win_std_dev(scan_win_std_dev[901]), .feature_accum(feature_accums[901]));
  accum_calculator ac902(.scan_win(scan_win902), .rectangle1_x(rectangle1_xs[902]), .rectangle1_y(rectangle1_ys[902]), .rectangle1_width(rectangle1_widths[902]), .rectangle1_height(rectangle1_heights[902]), .rectangle1_weight(rectangle1_weights[902]), .rectangle2_x(rectangle2_xs[902]), .rectangle2_y(rectangle2_ys[902]), .rectangle2_width(rectangle2_widths[902]), .rectangle2_height(rectangle2_heights[902]), .rectangle2_weight(rectangle2_weights[902]), .rectangle3_x(rectangle3_xs[902]), .rectangle3_y(rectangle3_ys[902]), .rectangle3_width(rectangle3_widths[902]), .rectangle3_height(rectangle3_heights[902]), .rectangle3_weight(rectangle3_weights[902]), .feature_threshold(feature_thresholds[902]), .feature_above(feature_aboves[902]), .feature_below(feature_belows[902]), .scan_win_std_dev(scan_win_std_dev[902]), .feature_accum(feature_accums[902]));
  accum_calculator ac903(.scan_win(scan_win903), .rectangle1_x(rectangle1_xs[903]), .rectangle1_y(rectangle1_ys[903]), .rectangle1_width(rectangle1_widths[903]), .rectangle1_height(rectangle1_heights[903]), .rectangle1_weight(rectangle1_weights[903]), .rectangle2_x(rectangle2_xs[903]), .rectangle2_y(rectangle2_ys[903]), .rectangle2_width(rectangle2_widths[903]), .rectangle2_height(rectangle2_heights[903]), .rectangle2_weight(rectangle2_weights[903]), .rectangle3_x(rectangle3_xs[903]), .rectangle3_y(rectangle3_ys[903]), .rectangle3_width(rectangle3_widths[903]), .rectangle3_height(rectangle3_heights[903]), .rectangle3_weight(rectangle3_weights[903]), .feature_threshold(feature_thresholds[903]), .feature_above(feature_aboves[903]), .feature_below(feature_belows[903]), .scan_win_std_dev(scan_win_std_dev[903]), .feature_accum(feature_accums[903]));
  accum_calculator ac904(.scan_win(scan_win904), .rectangle1_x(rectangle1_xs[904]), .rectangle1_y(rectangle1_ys[904]), .rectangle1_width(rectangle1_widths[904]), .rectangle1_height(rectangle1_heights[904]), .rectangle1_weight(rectangle1_weights[904]), .rectangle2_x(rectangle2_xs[904]), .rectangle2_y(rectangle2_ys[904]), .rectangle2_width(rectangle2_widths[904]), .rectangle2_height(rectangle2_heights[904]), .rectangle2_weight(rectangle2_weights[904]), .rectangle3_x(rectangle3_xs[904]), .rectangle3_y(rectangle3_ys[904]), .rectangle3_width(rectangle3_widths[904]), .rectangle3_height(rectangle3_heights[904]), .rectangle3_weight(rectangle3_weights[904]), .feature_threshold(feature_thresholds[904]), .feature_above(feature_aboves[904]), .feature_below(feature_belows[904]), .scan_win_std_dev(scan_win_std_dev[904]), .feature_accum(feature_accums[904]));
  accum_calculator ac905(.scan_win(scan_win905), .rectangle1_x(rectangle1_xs[905]), .rectangle1_y(rectangle1_ys[905]), .rectangle1_width(rectangle1_widths[905]), .rectangle1_height(rectangle1_heights[905]), .rectangle1_weight(rectangle1_weights[905]), .rectangle2_x(rectangle2_xs[905]), .rectangle2_y(rectangle2_ys[905]), .rectangle2_width(rectangle2_widths[905]), .rectangle2_height(rectangle2_heights[905]), .rectangle2_weight(rectangle2_weights[905]), .rectangle3_x(rectangle3_xs[905]), .rectangle3_y(rectangle3_ys[905]), .rectangle3_width(rectangle3_widths[905]), .rectangle3_height(rectangle3_heights[905]), .rectangle3_weight(rectangle3_weights[905]), .feature_threshold(feature_thresholds[905]), .feature_above(feature_aboves[905]), .feature_below(feature_belows[905]), .scan_win_std_dev(scan_win_std_dev[905]), .feature_accum(feature_accums[905]));
  accum_calculator ac906(.scan_win(scan_win906), .rectangle1_x(rectangle1_xs[906]), .rectangle1_y(rectangle1_ys[906]), .rectangle1_width(rectangle1_widths[906]), .rectangle1_height(rectangle1_heights[906]), .rectangle1_weight(rectangle1_weights[906]), .rectangle2_x(rectangle2_xs[906]), .rectangle2_y(rectangle2_ys[906]), .rectangle2_width(rectangle2_widths[906]), .rectangle2_height(rectangle2_heights[906]), .rectangle2_weight(rectangle2_weights[906]), .rectangle3_x(rectangle3_xs[906]), .rectangle3_y(rectangle3_ys[906]), .rectangle3_width(rectangle3_widths[906]), .rectangle3_height(rectangle3_heights[906]), .rectangle3_weight(rectangle3_weights[906]), .feature_threshold(feature_thresholds[906]), .feature_above(feature_aboves[906]), .feature_below(feature_belows[906]), .scan_win_std_dev(scan_win_std_dev[906]), .feature_accum(feature_accums[906]));
  accum_calculator ac907(.scan_win(scan_win907), .rectangle1_x(rectangle1_xs[907]), .rectangle1_y(rectangle1_ys[907]), .rectangle1_width(rectangle1_widths[907]), .rectangle1_height(rectangle1_heights[907]), .rectangle1_weight(rectangle1_weights[907]), .rectangle2_x(rectangle2_xs[907]), .rectangle2_y(rectangle2_ys[907]), .rectangle2_width(rectangle2_widths[907]), .rectangle2_height(rectangle2_heights[907]), .rectangle2_weight(rectangle2_weights[907]), .rectangle3_x(rectangle3_xs[907]), .rectangle3_y(rectangle3_ys[907]), .rectangle3_width(rectangle3_widths[907]), .rectangle3_height(rectangle3_heights[907]), .rectangle3_weight(rectangle3_weights[907]), .feature_threshold(feature_thresholds[907]), .feature_above(feature_aboves[907]), .feature_below(feature_belows[907]), .scan_win_std_dev(scan_win_std_dev[907]), .feature_accum(feature_accums[907]));
  accum_calculator ac908(.scan_win(scan_win908), .rectangle1_x(rectangle1_xs[908]), .rectangle1_y(rectangle1_ys[908]), .rectangle1_width(rectangle1_widths[908]), .rectangle1_height(rectangle1_heights[908]), .rectangle1_weight(rectangle1_weights[908]), .rectangle2_x(rectangle2_xs[908]), .rectangle2_y(rectangle2_ys[908]), .rectangle2_width(rectangle2_widths[908]), .rectangle2_height(rectangle2_heights[908]), .rectangle2_weight(rectangle2_weights[908]), .rectangle3_x(rectangle3_xs[908]), .rectangle3_y(rectangle3_ys[908]), .rectangle3_width(rectangle3_widths[908]), .rectangle3_height(rectangle3_heights[908]), .rectangle3_weight(rectangle3_weights[908]), .feature_threshold(feature_thresholds[908]), .feature_above(feature_aboves[908]), .feature_below(feature_belows[908]), .scan_win_std_dev(scan_win_std_dev[908]), .feature_accum(feature_accums[908]));
  accum_calculator ac909(.scan_win(scan_win909), .rectangle1_x(rectangle1_xs[909]), .rectangle1_y(rectangle1_ys[909]), .rectangle1_width(rectangle1_widths[909]), .rectangle1_height(rectangle1_heights[909]), .rectangle1_weight(rectangle1_weights[909]), .rectangle2_x(rectangle2_xs[909]), .rectangle2_y(rectangle2_ys[909]), .rectangle2_width(rectangle2_widths[909]), .rectangle2_height(rectangle2_heights[909]), .rectangle2_weight(rectangle2_weights[909]), .rectangle3_x(rectangle3_xs[909]), .rectangle3_y(rectangle3_ys[909]), .rectangle3_width(rectangle3_widths[909]), .rectangle3_height(rectangle3_heights[909]), .rectangle3_weight(rectangle3_weights[909]), .feature_threshold(feature_thresholds[909]), .feature_above(feature_aboves[909]), .feature_below(feature_belows[909]), .scan_win_std_dev(scan_win_std_dev[909]), .feature_accum(feature_accums[909]));
  accum_calculator ac910(.scan_win(scan_win910), .rectangle1_x(rectangle1_xs[910]), .rectangle1_y(rectangle1_ys[910]), .rectangle1_width(rectangle1_widths[910]), .rectangle1_height(rectangle1_heights[910]), .rectangle1_weight(rectangle1_weights[910]), .rectangle2_x(rectangle2_xs[910]), .rectangle2_y(rectangle2_ys[910]), .rectangle2_width(rectangle2_widths[910]), .rectangle2_height(rectangle2_heights[910]), .rectangle2_weight(rectangle2_weights[910]), .rectangle3_x(rectangle3_xs[910]), .rectangle3_y(rectangle3_ys[910]), .rectangle3_width(rectangle3_widths[910]), .rectangle3_height(rectangle3_heights[910]), .rectangle3_weight(rectangle3_weights[910]), .feature_threshold(feature_thresholds[910]), .feature_above(feature_aboves[910]), .feature_below(feature_belows[910]), .scan_win_std_dev(scan_win_std_dev[910]), .feature_accum(feature_accums[910]));
  accum_calculator ac911(.scan_win(scan_win911), .rectangle1_x(rectangle1_xs[911]), .rectangle1_y(rectangle1_ys[911]), .rectangle1_width(rectangle1_widths[911]), .rectangle1_height(rectangle1_heights[911]), .rectangle1_weight(rectangle1_weights[911]), .rectangle2_x(rectangle2_xs[911]), .rectangle2_y(rectangle2_ys[911]), .rectangle2_width(rectangle2_widths[911]), .rectangle2_height(rectangle2_heights[911]), .rectangle2_weight(rectangle2_weights[911]), .rectangle3_x(rectangle3_xs[911]), .rectangle3_y(rectangle3_ys[911]), .rectangle3_width(rectangle3_widths[911]), .rectangle3_height(rectangle3_heights[911]), .rectangle3_weight(rectangle3_weights[911]), .feature_threshold(feature_thresholds[911]), .feature_above(feature_aboves[911]), .feature_below(feature_belows[911]), .scan_win_std_dev(scan_win_std_dev[911]), .feature_accum(feature_accums[911]));
  accum_calculator ac912(.scan_win(scan_win912), .rectangle1_x(rectangle1_xs[912]), .rectangle1_y(rectangle1_ys[912]), .rectangle1_width(rectangle1_widths[912]), .rectangle1_height(rectangle1_heights[912]), .rectangle1_weight(rectangle1_weights[912]), .rectangle2_x(rectangle2_xs[912]), .rectangle2_y(rectangle2_ys[912]), .rectangle2_width(rectangle2_widths[912]), .rectangle2_height(rectangle2_heights[912]), .rectangle2_weight(rectangle2_weights[912]), .rectangle3_x(rectangle3_xs[912]), .rectangle3_y(rectangle3_ys[912]), .rectangle3_width(rectangle3_widths[912]), .rectangle3_height(rectangle3_heights[912]), .rectangle3_weight(rectangle3_weights[912]), .feature_threshold(feature_thresholds[912]), .feature_above(feature_aboves[912]), .feature_below(feature_belows[912]), .scan_win_std_dev(scan_win_std_dev[912]), .feature_accum(feature_accums[912]));
  accum_calculator ac913(.scan_win(scan_win913), .rectangle1_x(rectangle1_xs[913]), .rectangle1_y(rectangle1_ys[913]), .rectangle1_width(rectangle1_widths[913]), .rectangle1_height(rectangle1_heights[913]), .rectangle1_weight(rectangle1_weights[913]), .rectangle2_x(rectangle2_xs[913]), .rectangle2_y(rectangle2_ys[913]), .rectangle2_width(rectangle2_widths[913]), .rectangle2_height(rectangle2_heights[913]), .rectangle2_weight(rectangle2_weights[913]), .rectangle3_x(rectangle3_xs[913]), .rectangle3_y(rectangle3_ys[913]), .rectangle3_width(rectangle3_widths[913]), .rectangle3_height(rectangle3_heights[913]), .rectangle3_weight(rectangle3_weights[913]), .feature_threshold(feature_thresholds[913]), .feature_above(feature_aboves[913]), .feature_below(feature_belows[913]), .scan_win_std_dev(scan_win_std_dev[913]), .feature_accum(feature_accums[913]));
  accum_calculator ac914(.scan_win(scan_win914), .rectangle1_x(rectangle1_xs[914]), .rectangle1_y(rectangle1_ys[914]), .rectangle1_width(rectangle1_widths[914]), .rectangle1_height(rectangle1_heights[914]), .rectangle1_weight(rectangle1_weights[914]), .rectangle2_x(rectangle2_xs[914]), .rectangle2_y(rectangle2_ys[914]), .rectangle2_width(rectangle2_widths[914]), .rectangle2_height(rectangle2_heights[914]), .rectangle2_weight(rectangle2_weights[914]), .rectangle3_x(rectangle3_xs[914]), .rectangle3_y(rectangle3_ys[914]), .rectangle3_width(rectangle3_widths[914]), .rectangle3_height(rectangle3_heights[914]), .rectangle3_weight(rectangle3_weights[914]), .feature_threshold(feature_thresholds[914]), .feature_above(feature_aboves[914]), .feature_below(feature_belows[914]), .scan_win_std_dev(scan_win_std_dev[914]), .feature_accum(feature_accums[914]));
  accum_calculator ac915(.scan_win(scan_win915), .rectangle1_x(rectangle1_xs[915]), .rectangle1_y(rectangle1_ys[915]), .rectangle1_width(rectangle1_widths[915]), .rectangle1_height(rectangle1_heights[915]), .rectangle1_weight(rectangle1_weights[915]), .rectangle2_x(rectangle2_xs[915]), .rectangle2_y(rectangle2_ys[915]), .rectangle2_width(rectangle2_widths[915]), .rectangle2_height(rectangle2_heights[915]), .rectangle2_weight(rectangle2_weights[915]), .rectangle3_x(rectangle3_xs[915]), .rectangle3_y(rectangle3_ys[915]), .rectangle3_width(rectangle3_widths[915]), .rectangle3_height(rectangle3_heights[915]), .rectangle3_weight(rectangle3_weights[915]), .feature_threshold(feature_thresholds[915]), .feature_above(feature_aboves[915]), .feature_below(feature_belows[915]), .scan_win_std_dev(scan_win_std_dev[915]), .feature_accum(feature_accums[915]));
  accum_calculator ac916(.scan_win(scan_win916), .rectangle1_x(rectangle1_xs[916]), .rectangle1_y(rectangle1_ys[916]), .rectangle1_width(rectangle1_widths[916]), .rectangle1_height(rectangle1_heights[916]), .rectangle1_weight(rectangle1_weights[916]), .rectangle2_x(rectangle2_xs[916]), .rectangle2_y(rectangle2_ys[916]), .rectangle2_width(rectangle2_widths[916]), .rectangle2_height(rectangle2_heights[916]), .rectangle2_weight(rectangle2_weights[916]), .rectangle3_x(rectangle3_xs[916]), .rectangle3_y(rectangle3_ys[916]), .rectangle3_width(rectangle3_widths[916]), .rectangle3_height(rectangle3_heights[916]), .rectangle3_weight(rectangle3_weights[916]), .feature_threshold(feature_thresholds[916]), .feature_above(feature_aboves[916]), .feature_below(feature_belows[916]), .scan_win_std_dev(scan_win_std_dev[916]), .feature_accum(feature_accums[916]));
  accum_calculator ac917(.scan_win(scan_win917), .rectangle1_x(rectangle1_xs[917]), .rectangle1_y(rectangle1_ys[917]), .rectangle1_width(rectangle1_widths[917]), .rectangle1_height(rectangle1_heights[917]), .rectangle1_weight(rectangle1_weights[917]), .rectangle2_x(rectangle2_xs[917]), .rectangle2_y(rectangle2_ys[917]), .rectangle2_width(rectangle2_widths[917]), .rectangle2_height(rectangle2_heights[917]), .rectangle2_weight(rectangle2_weights[917]), .rectangle3_x(rectangle3_xs[917]), .rectangle3_y(rectangle3_ys[917]), .rectangle3_width(rectangle3_widths[917]), .rectangle3_height(rectangle3_heights[917]), .rectangle3_weight(rectangle3_weights[917]), .feature_threshold(feature_thresholds[917]), .feature_above(feature_aboves[917]), .feature_below(feature_belows[917]), .scan_win_std_dev(scan_win_std_dev[917]), .feature_accum(feature_accums[917]));
  accum_calculator ac918(.scan_win(scan_win918), .rectangle1_x(rectangle1_xs[918]), .rectangle1_y(rectangle1_ys[918]), .rectangle1_width(rectangle1_widths[918]), .rectangle1_height(rectangle1_heights[918]), .rectangle1_weight(rectangle1_weights[918]), .rectangle2_x(rectangle2_xs[918]), .rectangle2_y(rectangle2_ys[918]), .rectangle2_width(rectangle2_widths[918]), .rectangle2_height(rectangle2_heights[918]), .rectangle2_weight(rectangle2_weights[918]), .rectangle3_x(rectangle3_xs[918]), .rectangle3_y(rectangle3_ys[918]), .rectangle3_width(rectangle3_widths[918]), .rectangle3_height(rectangle3_heights[918]), .rectangle3_weight(rectangle3_weights[918]), .feature_threshold(feature_thresholds[918]), .feature_above(feature_aboves[918]), .feature_below(feature_belows[918]), .scan_win_std_dev(scan_win_std_dev[918]), .feature_accum(feature_accums[918]));
  accum_calculator ac919(.scan_win(scan_win919), .rectangle1_x(rectangle1_xs[919]), .rectangle1_y(rectangle1_ys[919]), .rectangle1_width(rectangle1_widths[919]), .rectangle1_height(rectangle1_heights[919]), .rectangle1_weight(rectangle1_weights[919]), .rectangle2_x(rectangle2_xs[919]), .rectangle2_y(rectangle2_ys[919]), .rectangle2_width(rectangle2_widths[919]), .rectangle2_height(rectangle2_heights[919]), .rectangle2_weight(rectangle2_weights[919]), .rectangle3_x(rectangle3_xs[919]), .rectangle3_y(rectangle3_ys[919]), .rectangle3_width(rectangle3_widths[919]), .rectangle3_height(rectangle3_heights[919]), .rectangle3_weight(rectangle3_weights[919]), .feature_threshold(feature_thresholds[919]), .feature_above(feature_aboves[919]), .feature_below(feature_belows[919]), .scan_win_std_dev(scan_win_std_dev[919]), .feature_accum(feature_accums[919]));
  accum_calculator ac920(.scan_win(scan_win920), .rectangle1_x(rectangle1_xs[920]), .rectangle1_y(rectangle1_ys[920]), .rectangle1_width(rectangle1_widths[920]), .rectangle1_height(rectangle1_heights[920]), .rectangle1_weight(rectangle1_weights[920]), .rectangle2_x(rectangle2_xs[920]), .rectangle2_y(rectangle2_ys[920]), .rectangle2_width(rectangle2_widths[920]), .rectangle2_height(rectangle2_heights[920]), .rectangle2_weight(rectangle2_weights[920]), .rectangle3_x(rectangle3_xs[920]), .rectangle3_y(rectangle3_ys[920]), .rectangle3_width(rectangle3_widths[920]), .rectangle3_height(rectangle3_heights[920]), .rectangle3_weight(rectangle3_weights[920]), .feature_threshold(feature_thresholds[920]), .feature_above(feature_aboves[920]), .feature_below(feature_belows[920]), .scan_win_std_dev(scan_win_std_dev[920]), .feature_accum(feature_accums[920]));
  accum_calculator ac921(.scan_win(scan_win921), .rectangle1_x(rectangle1_xs[921]), .rectangle1_y(rectangle1_ys[921]), .rectangle1_width(rectangle1_widths[921]), .rectangle1_height(rectangle1_heights[921]), .rectangle1_weight(rectangle1_weights[921]), .rectangle2_x(rectangle2_xs[921]), .rectangle2_y(rectangle2_ys[921]), .rectangle2_width(rectangle2_widths[921]), .rectangle2_height(rectangle2_heights[921]), .rectangle2_weight(rectangle2_weights[921]), .rectangle3_x(rectangle3_xs[921]), .rectangle3_y(rectangle3_ys[921]), .rectangle3_width(rectangle3_widths[921]), .rectangle3_height(rectangle3_heights[921]), .rectangle3_weight(rectangle3_weights[921]), .feature_threshold(feature_thresholds[921]), .feature_above(feature_aboves[921]), .feature_below(feature_belows[921]), .scan_win_std_dev(scan_win_std_dev[921]), .feature_accum(feature_accums[921]));
  accum_calculator ac922(.scan_win(scan_win922), .rectangle1_x(rectangle1_xs[922]), .rectangle1_y(rectangle1_ys[922]), .rectangle1_width(rectangle1_widths[922]), .rectangle1_height(rectangle1_heights[922]), .rectangle1_weight(rectangle1_weights[922]), .rectangle2_x(rectangle2_xs[922]), .rectangle2_y(rectangle2_ys[922]), .rectangle2_width(rectangle2_widths[922]), .rectangle2_height(rectangle2_heights[922]), .rectangle2_weight(rectangle2_weights[922]), .rectangle3_x(rectangle3_xs[922]), .rectangle3_y(rectangle3_ys[922]), .rectangle3_width(rectangle3_widths[922]), .rectangle3_height(rectangle3_heights[922]), .rectangle3_weight(rectangle3_weights[922]), .feature_threshold(feature_thresholds[922]), .feature_above(feature_aboves[922]), .feature_below(feature_belows[922]), .scan_win_std_dev(scan_win_std_dev[922]), .feature_accum(feature_accums[922]));
  accum_calculator ac923(.scan_win(scan_win923), .rectangle1_x(rectangle1_xs[923]), .rectangle1_y(rectangle1_ys[923]), .rectangle1_width(rectangle1_widths[923]), .rectangle1_height(rectangle1_heights[923]), .rectangle1_weight(rectangle1_weights[923]), .rectangle2_x(rectangle2_xs[923]), .rectangle2_y(rectangle2_ys[923]), .rectangle2_width(rectangle2_widths[923]), .rectangle2_height(rectangle2_heights[923]), .rectangle2_weight(rectangle2_weights[923]), .rectangle3_x(rectangle3_xs[923]), .rectangle3_y(rectangle3_ys[923]), .rectangle3_width(rectangle3_widths[923]), .rectangle3_height(rectangle3_heights[923]), .rectangle3_weight(rectangle3_weights[923]), .feature_threshold(feature_thresholds[923]), .feature_above(feature_aboves[923]), .feature_below(feature_belows[923]), .scan_win_std_dev(scan_win_std_dev[923]), .feature_accum(feature_accums[923]));
  accum_calculator ac924(.scan_win(scan_win924), .rectangle1_x(rectangle1_xs[924]), .rectangle1_y(rectangle1_ys[924]), .rectangle1_width(rectangle1_widths[924]), .rectangle1_height(rectangle1_heights[924]), .rectangle1_weight(rectangle1_weights[924]), .rectangle2_x(rectangle2_xs[924]), .rectangle2_y(rectangle2_ys[924]), .rectangle2_width(rectangle2_widths[924]), .rectangle2_height(rectangle2_heights[924]), .rectangle2_weight(rectangle2_weights[924]), .rectangle3_x(rectangle3_xs[924]), .rectangle3_y(rectangle3_ys[924]), .rectangle3_width(rectangle3_widths[924]), .rectangle3_height(rectangle3_heights[924]), .rectangle3_weight(rectangle3_weights[924]), .feature_threshold(feature_thresholds[924]), .feature_above(feature_aboves[924]), .feature_below(feature_belows[924]), .scan_win_std_dev(scan_win_std_dev[924]), .feature_accum(feature_accums[924]));
  accum_calculator ac925(.scan_win(scan_win925), .rectangle1_x(rectangle1_xs[925]), .rectangle1_y(rectangle1_ys[925]), .rectangle1_width(rectangle1_widths[925]), .rectangle1_height(rectangle1_heights[925]), .rectangle1_weight(rectangle1_weights[925]), .rectangle2_x(rectangle2_xs[925]), .rectangle2_y(rectangle2_ys[925]), .rectangle2_width(rectangle2_widths[925]), .rectangle2_height(rectangle2_heights[925]), .rectangle2_weight(rectangle2_weights[925]), .rectangle3_x(rectangle3_xs[925]), .rectangle3_y(rectangle3_ys[925]), .rectangle3_width(rectangle3_widths[925]), .rectangle3_height(rectangle3_heights[925]), .rectangle3_weight(rectangle3_weights[925]), .feature_threshold(feature_thresholds[925]), .feature_above(feature_aboves[925]), .feature_below(feature_belows[925]), .scan_win_std_dev(scan_win_std_dev[925]), .feature_accum(feature_accums[925]));
  accum_calculator ac926(.scan_win(scan_win926), .rectangle1_x(rectangle1_xs[926]), .rectangle1_y(rectangle1_ys[926]), .rectangle1_width(rectangle1_widths[926]), .rectangle1_height(rectangle1_heights[926]), .rectangle1_weight(rectangle1_weights[926]), .rectangle2_x(rectangle2_xs[926]), .rectangle2_y(rectangle2_ys[926]), .rectangle2_width(rectangle2_widths[926]), .rectangle2_height(rectangle2_heights[926]), .rectangle2_weight(rectangle2_weights[926]), .rectangle3_x(rectangle3_xs[926]), .rectangle3_y(rectangle3_ys[926]), .rectangle3_width(rectangle3_widths[926]), .rectangle3_height(rectangle3_heights[926]), .rectangle3_weight(rectangle3_weights[926]), .feature_threshold(feature_thresholds[926]), .feature_above(feature_aboves[926]), .feature_below(feature_belows[926]), .scan_win_std_dev(scan_win_std_dev[926]), .feature_accum(feature_accums[926]));
  accum_calculator ac927(.scan_win(scan_win927), .rectangle1_x(rectangle1_xs[927]), .rectangle1_y(rectangle1_ys[927]), .rectangle1_width(rectangle1_widths[927]), .rectangle1_height(rectangle1_heights[927]), .rectangle1_weight(rectangle1_weights[927]), .rectangle2_x(rectangle2_xs[927]), .rectangle2_y(rectangle2_ys[927]), .rectangle2_width(rectangle2_widths[927]), .rectangle2_height(rectangle2_heights[927]), .rectangle2_weight(rectangle2_weights[927]), .rectangle3_x(rectangle3_xs[927]), .rectangle3_y(rectangle3_ys[927]), .rectangle3_width(rectangle3_widths[927]), .rectangle3_height(rectangle3_heights[927]), .rectangle3_weight(rectangle3_weights[927]), .feature_threshold(feature_thresholds[927]), .feature_above(feature_aboves[927]), .feature_below(feature_belows[927]), .scan_win_std_dev(scan_win_std_dev[927]), .feature_accum(feature_accums[927]));
  accum_calculator ac928(.scan_win(scan_win928), .rectangle1_x(rectangle1_xs[928]), .rectangle1_y(rectangle1_ys[928]), .rectangle1_width(rectangle1_widths[928]), .rectangle1_height(rectangle1_heights[928]), .rectangle1_weight(rectangle1_weights[928]), .rectangle2_x(rectangle2_xs[928]), .rectangle2_y(rectangle2_ys[928]), .rectangle2_width(rectangle2_widths[928]), .rectangle2_height(rectangle2_heights[928]), .rectangle2_weight(rectangle2_weights[928]), .rectangle3_x(rectangle3_xs[928]), .rectangle3_y(rectangle3_ys[928]), .rectangle3_width(rectangle3_widths[928]), .rectangle3_height(rectangle3_heights[928]), .rectangle3_weight(rectangle3_weights[928]), .feature_threshold(feature_thresholds[928]), .feature_above(feature_aboves[928]), .feature_below(feature_belows[928]), .scan_win_std_dev(scan_win_std_dev[928]), .feature_accum(feature_accums[928]));
  accum_calculator ac929(.scan_win(scan_win929), .rectangle1_x(rectangle1_xs[929]), .rectangle1_y(rectangle1_ys[929]), .rectangle1_width(rectangle1_widths[929]), .rectangle1_height(rectangle1_heights[929]), .rectangle1_weight(rectangle1_weights[929]), .rectangle2_x(rectangle2_xs[929]), .rectangle2_y(rectangle2_ys[929]), .rectangle2_width(rectangle2_widths[929]), .rectangle2_height(rectangle2_heights[929]), .rectangle2_weight(rectangle2_weights[929]), .rectangle3_x(rectangle3_xs[929]), .rectangle3_y(rectangle3_ys[929]), .rectangle3_width(rectangle3_widths[929]), .rectangle3_height(rectangle3_heights[929]), .rectangle3_weight(rectangle3_weights[929]), .feature_threshold(feature_thresholds[929]), .feature_above(feature_aboves[929]), .feature_below(feature_belows[929]), .scan_win_std_dev(scan_win_std_dev[929]), .feature_accum(feature_accums[929]));
  accum_calculator ac930(.scan_win(scan_win930), .rectangle1_x(rectangle1_xs[930]), .rectangle1_y(rectangle1_ys[930]), .rectangle1_width(rectangle1_widths[930]), .rectangle1_height(rectangle1_heights[930]), .rectangle1_weight(rectangle1_weights[930]), .rectangle2_x(rectangle2_xs[930]), .rectangle2_y(rectangle2_ys[930]), .rectangle2_width(rectangle2_widths[930]), .rectangle2_height(rectangle2_heights[930]), .rectangle2_weight(rectangle2_weights[930]), .rectangle3_x(rectangle3_xs[930]), .rectangle3_y(rectangle3_ys[930]), .rectangle3_width(rectangle3_widths[930]), .rectangle3_height(rectangle3_heights[930]), .rectangle3_weight(rectangle3_weights[930]), .feature_threshold(feature_thresholds[930]), .feature_above(feature_aboves[930]), .feature_below(feature_belows[930]), .scan_win_std_dev(scan_win_std_dev[930]), .feature_accum(feature_accums[930]));
  accum_calculator ac931(.scan_win(scan_win931), .rectangle1_x(rectangle1_xs[931]), .rectangle1_y(rectangle1_ys[931]), .rectangle1_width(rectangle1_widths[931]), .rectangle1_height(rectangle1_heights[931]), .rectangle1_weight(rectangle1_weights[931]), .rectangle2_x(rectangle2_xs[931]), .rectangle2_y(rectangle2_ys[931]), .rectangle2_width(rectangle2_widths[931]), .rectangle2_height(rectangle2_heights[931]), .rectangle2_weight(rectangle2_weights[931]), .rectangle3_x(rectangle3_xs[931]), .rectangle3_y(rectangle3_ys[931]), .rectangle3_width(rectangle3_widths[931]), .rectangle3_height(rectangle3_heights[931]), .rectangle3_weight(rectangle3_weights[931]), .feature_threshold(feature_thresholds[931]), .feature_above(feature_aboves[931]), .feature_below(feature_belows[931]), .scan_win_std_dev(scan_win_std_dev[931]), .feature_accum(feature_accums[931]));
  accum_calculator ac932(.scan_win(scan_win932), .rectangle1_x(rectangle1_xs[932]), .rectangle1_y(rectangle1_ys[932]), .rectangle1_width(rectangle1_widths[932]), .rectangle1_height(rectangle1_heights[932]), .rectangle1_weight(rectangle1_weights[932]), .rectangle2_x(rectangle2_xs[932]), .rectangle2_y(rectangle2_ys[932]), .rectangle2_width(rectangle2_widths[932]), .rectangle2_height(rectangle2_heights[932]), .rectangle2_weight(rectangle2_weights[932]), .rectangle3_x(rectangle3_xs[932]), .rectangle3_y(rectangle3_ys[932]), .rectangle3_width(rectangle3_widths[932]), .rectangle3_height(rectangle3_heights[932]), .rectangle3_weight(rectangle3_weights[932]), .feature_threshold(feature_thresholds[932]), .feature_above(feature_aboves[932]), .feature_below(feature_belows[932]), .scan_win_std_dev(scan_win_std_dev[932]), .feature_accum(feature_accums[932]));
  accum_calculator ac933(.scan_win(scan_win933), .rectangle1_x(rectangle1_xs[933]), .rectangle1_y(rectangle1_ys[933]), .rectangle1_width(rectangle1_widths[933]), .rectangle1_height(rectangle1_heights[933]), .rectangle1_weight(rectangle1_weights[933]), .rectangle2_x(rectangle2_xs[933]), .rectangle2_y(rectangle2_ys[933]), .rectangle2_width(rectangle2_widths[933]), .rectangle2_height(rectangle2_heights[933]), .rectangle2_weight(rectangle2_weights[933]), .rectangle3_x(rectangle3_xs[933]), .rectangle3_y(rectangle3_ys[933]), .rectangle3_width(rectangle3_widths[933]), .rectangle3_height(rectangle3_heights[933]), .rectangle3_weight(rectangle3_weights[933]), .feature_threshold(feature_thresholds[933]), .feature_above(feature_aboves[933]), .feature_below(feature_belows[933]), .scan_win_std_dev(scan_win_std_dev[933]), .feature_accum(feature_accums[933]));
  accum_calculator ac934(.scan_win(scan_win934), .rectangle1_x(rectangle1_xs[934]), .rectangle1_y(rectangle1_ys[934]), .rectangle1_width(rectangle1_widths[934]), .rectangle1_height(rectangle1_heights[934]), .rectangle1_weight(rectangle1_weights[934]), .rectangle2_x(rectangle2_xs[934]), .rectangle2_y(rectangle2_ys[934]), .rectangle2_width(rectangle2_widths[934]), .rectangle2_height(rectangle2_heights[934]), .rectangle2_weight(rectangle2_weights[934]), .rectangle3_x(rectangle3_xs[934]), .rectangle3_y(rectangle3_ys[934]), .rectangle3_width(rectangle3_widths[934]), .rectangle3_height(rectangle3_heights[934]), .rectangle3_weight(rectangle3_weights[934]), .feature_threshold(feature_thresholds[934]), .feature_above(feature_aboves[934]), .feature_below(feature_belows[934]), .scan_win_std_dev(scan_win_std_dev[934]), .feature_accum(feature_accums[934]));
  accum_calculator ac935(.scan_win(scan_win935), .rectangle1_x(rectangle1_xs[935]), .rectangle1_y(rectangle1_ys[935]), .rectangle1_width(rectangle1_widths[935]), .rectangle1_height(rectangle1_heights[935]), .rectangle1_weight(rectangle1_weights[935]), .rectangle2_x(rectangle2_xs[935]), .rectangle2_y(rectangle2_ys[935]), .rectangle2_width(rectangle2_widths[935]), .rectangle2_height(rectangle2_heights[935]), .rectangle2_weight(rectangle2_weights[935]), .rectangle3_x(rectangle3_xs[935]), .rectangle3_y(rectangle3_ys[935]), .rectangle3_width(rectangle3_widths[935]), .rectangle3_height(rectangle3_heights[935]), .rectangle3_weight(rectangle3_weights[935]), .feature_threshold(feature_thresholds[935]), .feature_above(feature_aboves[935]), .feature_below(feature_belows[935]), .scan_win_std_dev(scan_win_std_dev[935]), .feature_accum(feature_accums[935]));
  accum_calculator ac936(.scan_win(scan_win936), .rectangle1_x(rectangle1_xs[936]), .rectangle1_y(rectangle1_ys[936]), .rectangle1_width(rectangle1_widths[936]), .rectangle1_height(rectangle1_heights[936]), .rectangle1_weight(rectangle1_weights[936]), .rectangle2_x(rectangle2_xs[936]), .rectangle2_y(rectangle2_ys[936]), .rectangle2_width(rectangle2_widths[936]), .rectangle2_height(rectangle2_heights[936]), .rectangle2_weight(rectangle2_weights[936]), .rectangle3_x(rectangle3_xs[936]), .rectangle3_y(rectangle3_ys[936]), .rectangle3_width(rectangle3_widths[936]), .rectangle3_height(rectangle3_heights[936]), .rectangle3_weight(rectangle3_weights[936]), .feature_threshold(feature_thresholds[936]), .feature_above(feature_aboves[936]), .feature_below(feature_belows[936]), .scan_win_std_dev(scan_win_std_dev[936]), .feature_accum(feature_accums[936]));
  accum_calculator ac937(.scan_win(scan_win937), .rectangle1_x(rectangle1_xs[937]), .rectangle1_y(rectangle1_ys[937]), .rectangle1_width(rectangle1_widths[937]), .rectangle1_height(rectangle1_heights[937]), .rectangle1_weight(rectangle1_weights[937]), .rectangle2_x(rectangle2_xs[937]), .rectangle2_y(rectangle2_ys[937]), .rectangle2_width(rectangle2_widths[937]), .rectangle2_height(rectangle2_heights[937]), .rectangle2_weight(rectangle2_weights[937]), .rectangle3_x(rectangle3_xs[937]), .rectangle3_y(rectangle3_ys[937]), .rectangle3_width(rectangle3_widths[937]), .rectangle3_height(rectangle3_heights[937]), .rectangle3_weight(rectangle3_weights[937]), .feature_threshold(feature_thresholds[937]), .feature_above(feature_aboves[937]), .feature_below(feature_belows[937]), .scan_win_std_dev(scan_win_std_dev[937]), .feature_accum(feature_accums[937]));
  accum_calculator ac938(.scan_win(scan_win938), .rectangle1_x(rectangle1_xs[938]), .rectangle1_y(rectangle1_ys[938]), .rectangle1_width(rectangle1_widths[938]), .rectangle1_height(rectangle1_heights[938]), .rectangle1_weight(rectangle1_weights[938]), .rectangle2_x(rectangle2_xs[938]), .rectangle2_y(rectangle2_ys[938]), .rectangle2_width(rectangle2_widths[938]), .rectangle2_height(rectangle2_heights[938]), .rectangle2_weight(rectangle2_weights[938]), .rectangle3_x(rectangle3_xs[938]), .rectangle3_y(rectangle3_ys[938]), .rectangle3_width(rectangle3_widths[938]), .rectangle3_height(rectangle3_heights[938]), .rectangle3_weight(rectangle3_weights[938]), .feature_threshold(feature_thresholds[938]), .feature_above(feature_aboves[938]), .feature_below(feature_belows[938]), .scan_win_std_dev(scan_win_std_dev[938]), .feature_accum(feature_accums[938]));
  accum_calculator ac939(.scan_win(scan_win939), .rectangle1_x(rectangle1_xs[939]), .rectangle1_y(rectangle1_ys[939]), .rectangle1_width(rectangle1_widths[939]), .rectangle1_height(rectangle1_heights[939]), .rectangle1_weight(rectangle1_weights[939]), .rectangle2_x(rectangle2_xs[939]), .rectangle2_y(rectangle2_ys[939]), .rectangle2_width(rectangle2_widths[939]), .rectangle2_height(rectangle2_heights[939]), .rectangle2_weight(rectangle2_weights[939]), .rectangle3_x(rectangle3_xs[939]), .rectangle3_y(rectangle3_ys[939]), .rectangle3_width(rectangle3_widths[939]), .rectangle3_height(rectangle3_heights[939]), .rectangle3_weight(rectangle3_weights[939]), .feature_threshold(feature_thresholds[939]), .feature_above(feature_aboves[939]), .feature_below(feature_belows[939]), .scan_win_std_dev(scan_win_std_dev[939]), .feature_accum(feature_accums[939]));
  accum_calculator ac940(.scan_win(scan_win940), .rectangle1_x(rectangle1_xs[940]), .rectangle1_y(rectangle1_ys[940]), .rectangle1_width(rectangle1_widths[940]), .rectangle1_height(rectangle1_heights[940]), .rectangle1_weight(rectangle1_weights[940]), .rectangle2_x(rectangle2_xs[940]), .rectangle2_y(rectangle2_ys[940]), .rectangle2_width(rectangle2_widths[940]), .rectangle2_height(rectangle2_heights[940]), .rectangle2_weight(rectangle2_weights[940]), .rectangle3_x(rectangle3_xs[940]), .rectangle3_y(rectangle3_ys[940]), .rectangle3_width(rectangle3_widths[940]), .rectangle3_height(rectangle3_heights[940]), .rectangle3_weight(rectangle3_weights[940]), .feature_threshold(feature_thresholds[940]), .feature_above(feature_aboves[940]), .feature_below(feature_belows[940]), .scan_win_std_dev(scan_win_std_dev[940]), .feature_accum(feature_accums[940]));
  accum_calculator ac941(.scan_win(scan_win941), .rectangle1_x(rectangle1_xs[941]), .rectangle1_y(rectangle1_ys[941]), .rectangle1_width(rectangle1_widths[941]), .rectangle1_height(rectangle1_heights[941]), .rectangle1_weight(rectangle1_weights[941]), .rectangle2_x(rectangle2_xs[941]), .rectangle2_y(rectangle2_ys[941]), .rectangle2_width(rectangle2_widths[941]), .rectangle2_height(rectangle2_heights[941]), .rectangle2_weight(rectangle2_weights[941]), .rectangle3_x(rectangle3_xs[941]), .rectangle3_y(rectangle3_ys[941]), .rectangle3_width(rectangle3_widths[941]), .rectangle3_height(rectangle3_heights[941]), .rectangle3_weight(rectangle3_weights[941]), .feature_threshold(feature_thresholds[941]), .feature_above(feature_aboves[941]), .feature_below(feature_belows[941]), .scan_win_std_dev(scan_win_std_dev[941]), .feature_accum(feature_accums[941]));
  accum_calculator ac942(.scan_win(scan_win942), .rectangle1_x(rectangle1_xs[942]), .rectangle1_y(rectangle1_ys[942]), .rectangle1_width(rectangle1_widths[942]), .rectangle1_height(rectangle1_heights[942]), .rectangle1_weight(rectangle1_weights[942]), .rectangle2_x(rectangle2_xs[942]), .rectangle2_y(rectangle2_ys[942]), .rectangle2_width(rectangle2_widths[942]), .rectangle2_height(rectangle2_heights[942]), .rectangle2_weight(rectangle2_weights[942]), .rectangle3_x(rectangle3_xs[942]), .rectangle3_y(rectangle3_ys[942]), .rectangle3_width(rectangle3_widths[942]), .rectangle3_height(rectangle3_heights[942]), .rectangle3_weight(rectangle3_weights[942]), .feature_threshold(feature_thresholds[942]), .feature_above(feature_aboves[942]), .feature_below(feature_belows[942]), .scan_win_std_dev(scan_win_std_dev[942]), .feature_accum(feature_accums[942]));
  accum_calculator ac943(.scan_win(scan_win943), .rectangle1_x(rectangle1_xs[943]), .rectangle1_y(rectangle1_ys[943]), .rectangle1_width(rectangle1_widths[943]), .rectangle1_height(rectangle1_heights[943]), .rectangle1_weight(rectangle1_weights[943]), .rectangle2_x(rectangle2_xs[943]), .rectangle2_y(rectangle2_ys[943]), .rectangle2_width(rectangle2_widths[943]), .rectangle2_height(rectangle2_heights[943]), .rectangle2_weight(rectangle2_weights[943]), .rectangle3_x(rectangle3_xs[943]), .rectangle3_y(rectangle3_ys[943]), .rectangle3_width(rectangle3_widths[943]), .rectangle3_height(rectangle3_heights[943]), .rectangle3_weight(rectangle3_weights[943]), .feature_threshold(feature_thresholds[943]), .feature_above(feature_aboves[943]), .feature_below(feature_belows[943]), .scan_win_std_dev(scan_win_std_dev[943]), .feature_accum(feature_accums[943]));
  accum_calculator ac944(.scan_win(scan_win944), .rectangle1_x(rectangle1_xs[944]), .rectangle1_y(rectangle1_ys[944]), .rectangle1_width(rectangle1_widths[944]), .rectangle1_height(rectangle1_heights[944]), .rectangle1_weight(rectangle1_weights[944]), .rectangle2_x(rectangle2_xs[944]), .rectangle2_y(rectangle2_ys[944]), .rectangle2_width(rectangle2_widths[944]), .rectangle2_height(rectangle2_heights[944]), .rectangle2_weight(rectangle2_weights[944]), .rectangle3_x(rectangle3_xs[944]), .rectangle3_y(rectangle3_ys[944]), .rectangle3_width(rectangle3_widths[944]), .rectangle3_height(rectangle3_heights[944]), .rectangle3_weight(rectangle3_weights[944]), .feature_threshold(feature_thresholds[944]), .feature_above(feature_aboves[944]), .feature_below(feature_belows[944]), .scan_win_std_dev(scan_win_std_dev[944]), .feature_accum(feature_accums[944]));
  accum_calculator ac945(.scan_win(scan_win945), .rectangle1_x(rectangle1_xs[945]), .rectangle1_y(rectangle1_ys[945]), .rectangle1_width(rectangle1_widths[945]), .rectangle1_height(rectangle1_heights[945]), .rectangle1_weight(rectangle1_weights[945]), .rectangle2_x(rectangle2_xs[945]), .rectangle2_y(rectangle2_ys[945]), .rectangle2_width(rectangle2_widths[945]), .rectangle2_height(rectangle2_heights[945]), .rectangle2_weight(rectangle2_weights[945]), .rectangle3_x(rectangle3_xs[945]), .rectangle3_y(rectangle3_ys[945]), .rectangle3_width(rectangle3_widths[945]), .rectangle3_height(rectangle3_heights[945]), .rectangle3_weight(rectangle3_weights[945]), .feature_threshold(feature_thresholds[945]), .feature_above(feature_aboves[945]), .feature_below(feature_belows[945]), .scan_win_std_dev(scan_win_std_dev[945]), .feature_accum(feature_accums[945]));
  accum_calculator ac946(.scan_win(scan_win946), .rectangle1_x(rectangle1_xs[946]), .rectangle1_y(rectangle1_ys[946]), .rectangle1_width(rectangle1_widths[946]), .rectangle1_height(rectangle1_heights[946]), .rectangle1_weight(rectangle1_weights[946]), .rectangle2_x(rectangle2_xs[946]), .rectangle2_y(rectangle2_ys[946]), .rectangle2_width(rectangle2_widths[946]), .rectangle2_height(rectangle2_heights[946]), .rectangle2_weight(rectangle2_weights[946]), .rectangle3_x(rectangle3_xs[946]), .rectangle3_y(rectangle3_ys[946]), .rectangle3_width(rectangle3_widths[946]), .rectangle3_height(rectangle3_heights[946]), .rectangle3_weight(rectangle3_weights[946]), .feature_threshold(feature_thresholds[946]), .feature_above(feature_aboves[946]), .feature_below(feature_belows[946]), .scan_win_std_dev(scan_win_std_dev[946]), .feature_accum(feature_accums[946]));
  accum_calculator ac947(.scan_win(scan_win947), .rectangle1_x(rectangle1_xs[947]), .rectangle1_y(rectangle1_ys[947]), .rectangle1_width(rectangle1_widths[947]), .rectangle1_height(rectangle1_heights[947]), .rectangle1_weight(rectangle1_weights[947]), .rectangle2_x(rectangle2_xs[947]), .rectangle2_y(rectangle2_ys[947]), .rectangle2_width(rectangle2_widths[947]), .rectangle2_height(rectangle2_heights[947]), .rectangle2_weight(rectangle2_weights[947]), .rectangle3_x(rectangle3_xs[947]), .rectangle3_y(rectangle3_ys[947]), .rectangle3_width(rectangle3_widths[947]), .rectangle3_height(rectangle3_heights[947]), .rectangle3_weight(rectangle3_weights[947]), .feature_threshold(feature_thresholds[947]), .feature_above(feature_aboves[947]), .feature_below(feature_belows[947]), .scan_win_std_dev(scan_win_std_dev[947]), .feature_accum(feature_accums[947]));
  accum_calculator ac948(.scan_win(scan_win948), .rectangle1_x(rectangle1_xs[948]), .rectangle1_y(rectangle1_ys[948]), .rectangle1_width(rectangle1_widths[948]), .rectangle1_height(rectangle1_heights[948]), .rectangle1_weight(rectangle1_weights[948]), .rectangle2_x(rectangle2_xs[948]), .rectangle2_y(rectangle2_ys[948]), .rectangle2_width(rectangle2_widths[948]), .rectangle2_height(rectangle2_heights[948]), .rectangle2_weight(rectangle2_weights[948]), .rectangle3_x(rectangle3_xs[948]), .rectangle3_y(rectangle3_ys[948]), .rectangle3_width(rectangle3_widths[948]), .rectangle3_height(rectangle3_heights[948]), .rectangle3_weight(rectangle3_weights[948]), .feature_threshold(feature_thresholds[948]), .feature_above(feature_aboves[948]), .feature_below(feature_belows[948]), .scan_win_std_dev(scan_win_std_dev[948]), .feature_accum(feature_accums[948]));
  accum_calculator ac949(.scan_win(scan_win949), .rectangle1_x(rectangle1_xs[949]), .rectangle1_y(rectangle1_ys[949]), .rectangle1_width(rectangle1_widths[949]), .rectangle1_height(rectangle1_heights[949]), .rectangle1_weight(rectangle1_weights[949]), .rectangle2_x(rectangle2_xs[949]), .rectangle2_y(rectangle2_ys[949]), .rectangle2_width(rectangle2_widths[949]), .rectangle2_height(rectangle2_heights[949]), .rectangle2_weight(rectangle2_weights[949]), .rectangle3_x(rectangle3_xs[949]), .rectangle3_y(rectangle3_ys[949]), .rectangle3_width(rectangle3_widths[949]), .rectangle3_height(rectangle3_heights[949]), .rectangle3_weight(rectangle3_weights[949]), .feature_threshold(feature_thresholds[949]), .feature_above(feature_aboves[949]), .feature_below(feature_belows[949]), .scan_win_std_dev(scan_win_std_dev[949]), .feature_accum(feature_accums[949]));
  accum_calculator ac950(.scan_win(scan_win950), .rectangle1_x(rectangle1_xs[950]), .rectangle1_y(rectangle1_ys[950]), .rectangle1_width(rectangle1_widths[950]), .rectangle1_height(rectangle1_heights[950]), .rectangle1_weight(rectangle1_weights[950]), .rectangle2_x(rectangle2_xs[950]), .rectangle2_y(rectangle2_ys[950]), .rectangle2_width(rectangle2_widths[950]), .rectangle2_height(rectangle2_heights[950]), .rectangle2_weight(rectangle2_weights[950]), .rectangle3_x(rectangle3_xs[950]), .rectangle3_y(rectangle3_ys[950]), .rectangle3_width(rectangle3_widths[950]), .rectangle3_height(rectangle3_heights[950]), .rectangle3_weight(rectangle3_weights[950]), .feature_threshold(feature_thresholds[950]), .feature_above(feature_aboves[950]), .feature_below(feature_belows[950]), .scan_win_std_dev(scan_win_std_dev[950]), .feature_accum(feature_accums[950]));
  accum_calculator ac951(.scan_win(scan_win951), .rectangle1_x(rectangle1_xs[951]), .rectangle1_y(rectangle1_ys[951]), .rectangle1_width(rectangle1_widths[951]), .rectangle1_height(rectangle1_heights[951]), .rectangle1_weight(rectangle1_weights[951]), .rectangle2_x(rectangle2_xs[951]), .rectangle2_y(rectangle2_ys[951]), .rectangle2_width(rectangle2_widths[951]), .rectangle2_height(rectangle2_heights[951]), .rectangle2_weight(rectangle2_weights[951]), .rectangle3_x(rectangle3_xs[951]), .rectangle3_y(rectangle3_ys[951]), .rectangle3_width(rectangle3_widths[951]), .rectangle3_height(rectangle3_heights[951]), .rectangle3_weight(rectangle3_weights[951]), .feature_threshold(feature_thresholds[951]), .feature_above(feature_aboves[951]), .feature_below(feature_belows[951]), .scan_win_std_dev(scan_win_std_dev[951]), .feature_accum(feature_accums[951]));
  accum_calculator ac952(.scan_win(scan_win952), .rectangle1_x(rectangle1_xs[952]), .rectangle1_y(rectangle1_ys[952]), .rectangle1_width(rectangle1_widths[952]), .rectangle1_height(rectangle1_heights[952]), .rectangle1_weight(rectangle1_weights[952]), .rectangle2_x(rectangle2_xs[952]), .rectangle2_y(rectangle2_ys[952]), .rectangle2_width(rectangle2_widths[952]), .rectangle2_height(rectangle2_heights[952]), .rectangle2_weight(rectangle2_weights[952]), .rectangle3_x(rectangle3_xs[952]), .rectangle3_y(rectangle3_ys[952]), .rectangle3_width(rectangle3_widths[952]), .rectangle3_height(rectangle3_heights[952]), .rectangle3_weight(rectangle3_weights[952]), .feature_threshold(feature_thresholds[952]), .feature_above(feature_aboves[952]), .feature_below(feature_belows[952]), .scan_win_std_dev(scan_win_std_dev[952]), .feature_accum(feature_accums[952]));
  accum_calculator ac953(.scan_win(scan_win953), .rectangle1_x(rectangle1_xs[953]), .rectangle1_y(rectangle1_ys[953]), .rectangle1_width(rectangle1_widths[953]), .rectangle1_height(rectangle1_heights[953]), .rectangle1_weight(rectangle1_weights[953]), .rectangle2_x(rectangle2_xs[953]), .rectangle2_y(rectangle2_ys[953]), .rectangle2_width(rectangle2_widths[953]), .rectangle2_height(rectangle2_heights[953]), .rectangle2_weight(rectangle2_weights[953]), .rectangle3_x(rectangle3_xs[953]), .rectangle3_y(rectangle3_ys[953]), .rectangle3_width(rectangle3_widths[953]), .rectangle3_height(rectangle3_heights[953]), .rectangle3_weight(rectangle3_weights[953]), .feature_threshold(feature_thresholds[953]), .feature_above(feature_aboves[953]), .feature_below(feature_belows[953]), .scan_win_std_dev(scan_win_std_dev[953]), .feature_accum(feature_accums[953]));
  accum_calculator ac954(.scan_win(scan_win954), .rectangle1_x(rectangle1_xs[954]), .rectangle1_y(rectangle1_ys[954]), .rectangle1_width(rectangle1_widths[954]), .rectangle1_height(rectangle1_heights[954]), .rectangle1_weight(rectangle1_weights[954]), .rectangle2_x(rectangle2_xs[954]), .rectangle2_y(rectangle2_ys[954]), .rectangle2_width(rectangle2_widths[954]), .rectangle2_height(rectangle2_heights[954]), .rectangle2_weight(rectangle2_weights[954]), .rectangle3_x(rectangle3_xs[954]), .rectangle3_y(rectangle3_ys[954]), .rectangle3_width(rectangle3_widths[954]), .rectangle3_height(rectangle3_heights[954]), .rectangle3_weight(rectangle3_weights[954]), .feature_threshold(feature_thresholds[954]), .feature_above(feature_aboves[954]), .feature_below(feature_belows[954]), .scan_win_std_dev(scan_win_std_dev[954]), .feature_accum(feature_accums[954]));
  accum_calculator ac955(.scan_win(scan_win955), .rectangle1_x(rectangle1_xs[955]), .rectangle1_y(rectangle1_ys[955]), .rectangle1_width(rectangle1_widths[955]), .rectangle1_height(rectangle1_heights[955]), .rectangle1_weight(rectangle1_weights[955]), .rectangle2_x(rectangle2_xs[955]), .rectangle2_y(rectangle2_ys[955]), .rectangle2_width(rectangle2_widths[955]), .rectangle2_height(rectangle2_heights[955]), .rectangle2_weight(rectangle2_weights[955]), .rectangle3_x(rectangle3_xs[955]), .rectangle3_y(rectangle3_ys[955]), .rectangle3_width(rectangle3_widths[955]), .rectangle3_height(rectangle3_heights[955]), .rectangle3_weight(rectangle3_weights[955]), .feature_threshold(feature_thresholds[955]), .feature_above(feature_aboves[955]), .feature_below(feature_belows[955]), .scan_win_std_dev(scan_win_std_dev[955]), .feature_accum(feature_accums[955]));
  accum_calculator ac956(.scan_win(scan_win956), .rectangle1_x(rectangle1_xs[956]), .rectangle1_y(rectangle1_ys[956]), .rectangle1_width(rectangle1_widths[956]), .rectangle1_height(rectangle1_heights[956]), .rectangle1_weight(rectangle1_weights[956]), .rectangle2_x(rectangle2_xs[956]), .rectangle2_y(rectangle2_ys[956]), .rectangle2_width(rectangle2_widths[956]), .rectangle2_height(rectangle2_heights[956]), .rectangle2_weight(rectangle2_weights[956]), .rectangle3_x(rectangle3_xs[956]), .rectangle3_y(rectangle3_ys[956]), .rectangle3_width(rectangle3_widths[956]), .rectangle3_height(rectangle3_heights[956]), .rectangle3_weight(rectangle3_weights[956]), .feature_threshold(feature_thresholds[956]), .feature_above(feature_aboves[956]), .feature_below(feature_belows[956]), .scan_win_std_dev(scan_win_std_dev[956]), .feature_accum(feature_accums[956]));
  accum_calculator ac957(.scan_win(scan_win957), .rectangle1_x(rectangle1_xs[957]), .rectangle1_y(rectangle1_ys[957]), .rectangle1_width(rectangle1_widths[957]), .rectangle1_height(rectangle1_heights[957]), .rectangle1_weight(rectangle1_weights[957]), .rectangle2_x(rectangle2_xs[957]), .rectangle2_y(rectangle2_ys[957]), .rectangle2_width(rectangle2_widths[957]), .rectangle2_height(rectangle2_heights[957]), .rectangle2_weight(rectangle2_weights[957]), .rectangle3_x(rectangle3_xs[957]), .rectangle3_y(rectangle3_ys[957]), .rectangle3_width(rectangle3_widths[957]), .rectangle3_height(rectangle3_heights[957]), .rectangle3_weight(rectangle3_weights[957]), .feature_threshold(feature_thresholds[957]), .feature_above(feature_aboves[957]), .feature_below(feature_belows[957]), .scan_win_std_dev(scan_win_std_dev[957]), .feature_accum(feature_accums[957]));
  accum_calculator ac958(.scan_win(scan_win958), .rectangle1_x(rectangle1_xs[958]), .rectangle1_y(rectangle1_ys[958]), .rectangle1_width(rectangle1_widths[958]), .rectangle1_height(rectangle1_heights[958]), .rectangle1_weight(rectangle1_weights[958]), .rectangle2_x(rectangle2_xs[958]), .rectangle2_y(rectangle2_ys[958]), .rectangle2_width(rectangle2_widths[958]), .rectangle2_height(rectangle2_heights[958]), .rectangle2_weight(rectangle2_weights[958]), .rectangle3_x(rectangle3_xs[958]), .rectangle3_y(rectangle3_ys[958]), .rectangle3_width(rectangle3_widths[958]), .rectangle3_height(rectangle3_heights[958]), .rectangle3_weight(rectangle3_weights[958]), .feature_threshold(feature_thresholds[958]), .feature_above(feature_aboves[958]), .feature_below(feature_belows[958]), .scan_win_std_dev(scan_win_std_dev[958]), .feature_accum(feature_accums[958]));
  accum_calculator ac959(.scan_win(scan_win959), .rectangle1_x(rectangle1_xs[959]), .rectangle1_y(rectangle1_ys[959]), .rectangle1_width(rectangle1_widths[959]), .rectangle1_height(rectangle1_heights[959]), .rectangle1_weight(rectangle1_weights[959]), .rectangle2_x(rectangle2_xs[959]), .rectangle2_y(rectangle2_ys[959]), .rectangle2_width(rectangle2_widths[959]), .rectangle2_height(rectangle2_heights[959]), .rectangle2_weight(rectangle2_weights[959]), .rectangle3_x(rectangle3_xs[959]), .rectangle3_y(rectangle3_ys[959]), .rectangle3_width(rectangle3_widths[959]), .rectangle3_height(rectangle3_heights[959]), .rectangle3_weight(rectangle3_weights[959]), .feature_threshold(feature_thresholds[959]), .feature_above(feature_aboves[959]), .feature_below(feature_belows[959]), .scan_win_std_dev(scan_win_std_dev[959]), .feature_accum(feature_accums[959]));
  accum_calculator ac960(.scan_win(scan_win960), .rectangle1_x(rectangle1_xs[960]), .rectangle1_y(rectangle1_ys[960]), .rectangle1_width(rectangle1_widths[960]), .rectangle1_height(rectangle1_heights[960]), .rectangle1_weight(rectangle1_weights[960]), .rectangle2_x(rectangle2_xs[960]), .rectangle2_y(rectangle2_ys[960]), .rectangle2_width(rectangle2_widths[960]), .rectangle2_height(rectangle2_heights[960]), .rectangle2_weight(rectangle2_weights[960]), .rectangle3_x(rectangle3_xs[960]), .rectangle3_y(rectangle3_ys[960]), .rectangle3_width(rectangle3_widths[960]), .rectangle3_height(rectangle3_heights[960]), .rectangle3_weight(rectangle3_weights[960]), .feature_threshold(feature_thresholds[960]), .feature_above(feature_aboves[960]), .feature_below(feature_belows[960]), .scan_win_std_dev(scan_win_std_dev[960]), .feature_accum(feature_accums[960]));
  accum_calculator ac961(.scan_win(scan_win961), .rectangle1_x(rectangle1_xs[961]), .rectangle1_y(rectangle1_ys[961]), .rectangle1_width(rectangle1_widths[961]), .rectangle1_height(rectangle1_heights[961]), .rectangle1_weight(rectangle1_weights[961]), .rectangle2_x(rectangle2_xs[961]), .rectangle2_y(rectangle2_ys[961]), .rectangle2_width(rectangle2_widths[961]), .rectangle2_height(rectangle2_heights[961]), .rectangle2_weight(rectangle2_weights[961]), .rectangle3_x(rectangle3_xs[961]), .rectangle3_y(rectangle3_ys[961]), .rectangle3_width(rectangle3_widths[961]), .rectangle3_height(rectangle3_heights[961]), .rectangle3_weight(rectangle3_weights[961]), .feature_threshold(feature_thresholds[961]), .feature_above(feature_aboves[961]), .feature_below(feature_belows[961]), .scan_win_std_dev(scan_win_std_dev[961]), .feature_accum(feature_accums[961]));
  accum_calculator ac962(.scan_win(scan_win962), .rectangle1_x(rectangle1_xs[962]), .rectangle1_y(rectangle1_ys[962]), .rectangle1_width(rectangle1_widths[962]), .rectangle1_height(rectangle1_heights[962]), .rectangle1_weight(rectangle1_weights[962]), .rectangle2_x(rectangle2_xs[962]), .rectangle2_y(rectangle2_ys[962]), .rectangle2_width(rectangle2_widths[962]), .rectangle2_height(rectangle2_heights[962]), .rectangle2_weight(rectangle2_weights[962]), .rectangle3_x(rectangle3_xs[962]), .rectangle3_y(rectangle3_ys[962]), .rectangle3_width(rectangle3_widths[962]), .rectangle3_height(rectangle3_heights[962]), .rectangle3_weight(rectangle3_weights[962]), .feature_threshold(feature_thresholds[962]), .feature_above(feature_aboves[962]), .feature_below(feature_belows[962]), .scan_win_std_dev(scan_win_std_dev[962]), .feature_accum(feature_accums[962]));
  accum_calculator ac963(.scan_win(scan_win963), .rectangle1_x(rectangle1_xs[963]), .rectangle1_y(rectangle1_ys[963]), .rectangle1_width(rectangle1_widths[963]), .rectangle1_height(rectangle1_heights[963]), .rectangle1_weight(rectangle1_weights[963]), .rectangle2_x(rectangle2_xs[963]), .rectangle2_y(rectangle2_ys[963]), .rectangle2_width(rectangle2_widths[963]), .rectangle2_height(rectangle2_heights[963]), .rectangle2_weight(rectangle2_weights[963]), .rectangle3_x(rectangle3_xs[963]), .rectangle3_y(rectangle3_ys[963]), .rectangle3_width(rectangle3_widths[963]), .rectangle3_height(rectangle3_heights[963]), .rectangle3_weight(rectangle3_weights[963]), .feature_threshold(feature_thresholds[963]), .feature_above(feature_aboves[963]), .feature_below(feature_belows[963]), .scan_win_std_dev(scan_win_std_dev[963]), .feature_accum(feature_accums[963]));
  accum_calculator ac964(.scan_win(scan_win964), .rectangle1_x(rectangle1_xs[964]), .rectangle1_y(rectangle1_ys[964]), .rectangle1_width(rectangle1_widths[964]), .rectangle1_height(rectangle1_heights[964]), .rectangle1_weight(rectangle1_weights[964]), .rectangle2_x(rectangle2_xs[964]), .rectangle2_y(rectangle2_ys[964]), .rectangle2_width(rectangle2_widths[964]), .rectangle2_height(rectangle2_heights[964]), .rectangle2_weight(rectangle2_weights[964]), .rectangle3_x(rectangle3_xs[964]), .rectangle3_y(rectangle3_ys[964]), .rectangle3_width(rectangle3_widths[964]), .rectangle3_height(rectangle3_heights[964]), .rectangle3_weight(rectangle3_weights[964]), .feature_threshold(feature_thresholds[964]), .feature_above(feature_aboves[964]), .feature_below(feature_belows[964]), .scan_win_std_dev(scan_win_std_dev[964]), .feature_accum(feature_accums[964]));
  accum_calculator ac965(.scan_win(scan_win965), .rectangle1_x(rectangle1_xs[965]), .rectangle1_y(rectangle1_ys[965]), .rectangle1_width(rectangle1_widths[965]), .rectangle1_height(rectangle1_heights[965]), .rectangle1_weight(rectangle1_weights[965]), .rectangle2_x(rectangle2_xs[965]), .rectangle2_y(rectangle2_ys[965]), .rectangle2_width(rectangle2_widths[965]), .rectangle2_height(rectangle2_heights[965]), .rectangle2_weight(rectangle2_weights[965]), .rectangle3_x(rectangle3_xs[965]), .rectangle3_y(rectangle3_ys[965]), .rectangle3_width(rectangle3_widths[965]), .rectangle3_height(rectangle3_heights[965]), .rectangle3_weight(rectangle3_weights[965]), .feature_threshold(feature_thresholds[965]), .feature_above(feature_aboves[965]), .feature_below(feature_belows[965]), .scan_win_std_dev(scan_win_std_dev[965]), .feature_accum(feature_accums[965]));
  accum_calculator ac966(.scan_win(scan_win966), .rectangle1_x(rectangle1_xs[966]), .rectangle1_y(rectangle1_ys[966]), .rectangle1_width(rectangle1_widths[966]), .rectangle1_height(rectangle1_heights[966]), .rectangle1_weight(rectangle1_weights[966]), .rectangle2_x(rectangle2_xs[966]), .rectangle2_y(rectangle2_ys[966]), .rectangle2_width(rectangle2_widths[966]), .rectangle2_height(rectangle2_heights[966]), .rectangle2_weight(rectangle2_weights[966]), .rectangle3_x(rectangle3_xs[966]), .rectangle3_y(rectangle3_ys[966]), .rectangle3_width(rectangle3_widths[966]), .rectangle3_height(rectangle3_heights[966]), .rectangle3_weight(rectangle3_weights[966]), .feature_threshold(feature_thresholds[966]), .feature_above(feature_aboves[966]), .feature_below(feature_belows[966]), .scan_win_std_dev(scan_win_std_dev[966]), .feature_accum(feature_accums[966]));
  accum_calculator ac967(.scan_win(scan_win967), .rectangle1_x(rectangle1_xs[967]), .rectangle1_y(rectangle1_ys[967]), .rectangle1_width(rectangle1_widths[967]), .rectangle1_height(rectangle1_heights[967]), .rectangle1_weight(rectangle1_weights[967]), .rectangle2_x(rectangle2_xs[967]), .rectangle2_y(rectangle2_ys[967]), .rectangle2_width(rectangle2_widths[967]), .rectangle2_height(rectangle2_heights[967]), .rectangle2_weight(rectangle2_weights[967]), .rectangle3_x(rectangle3_xs[967]), .rectangle3_y(rectangle3_ys[967]), .rectangle3_width(rectangle3_widths[967]), .rectangle3_height(rectangle3_heights[967]), .rectangle3_weight(rectangle3_weights[967]), .feature_threshold(feature_thresholds[967]), .feature_above(feature_aboves[967]), .feature_below(feature_belows[967]), .scan_win_std_dev(scan_win_std_dev[967]), .feature_accum(feature_accums[967]));
  accum_calculator ac968(.scan_win(scan_win968), .rectangle1_x(rectangle1_xs[968]), .rectangle1_y(rectangle1_ys[968]), .rectangle1_width(rectangle1_widths[968]), .rectangle1_height(rectangle1_heights[968]), .rectangle1_weight(rectangle1_weights[968]), .rectangle2_x(rectangle2_xs[968]), .rectangle2_y(rectangle2_ys[968]), .rectangle2_width(rectangle2_widths[968]), .rectangle2_height(rectangle2_heights[968]), .rectangle2_weight(rectangle2_weights[968]), .rectangle3_x(rectangle3_xs[968]), .rectangle3_y(rectangle3_ys[968]), .rectangle3_width(rectangle3_widths[968]), .rectangle3_height(rectangle3_heights[968]), .rectangle3_weight(rectangle3_weights[968]), .feature_threshold(feature_thresholds[968]), .feature_above(feature_aboves[968]), .feature_below(feature_belows[968]), .scan_win_std_dev(scan_win_std_dev[968]), .feature_accum(feature_accums[968]));
  accum_calculator ac969(.scan_win(scan_win969), .rectangle1_x(rectangle1_xs[969]), .rectangle1_y(rectangle1_ys[969]), .rectangle1_width(rectangle1_widths[969]), .rectangle1_height(rectangle1_heights[969]), .rectangle1_weight(rectangle1_weights[969]), .rectangle2_x(rectangle2_xs[969]), .rectangle2_y(rectangle2_ys[969]), .rectangle2_width(rectangle2_widths[969]), .rectangle2_height(rectangle2_heights[969]), .rectangle2_weight(rectangle2_weights[969]), .rectangle3_x(rectangle3_xs[969]), .rectangle3_y(rectangle3_ys[969]), .rectangle3_width(rectangle3_widths[969]), .rectangle3_height(rectangle3_heights[969]), .rectangle3_weight(rectangle3_weights[969]), .feature_threshold(feature_thresholds[969]), .feature_above(feature_aboves[969]), .feature_below(feature_belows[969]), .scan_win_std_dev(scan_win_std_dev[969]), .feature_accum(feature_accums[969]));
  accum_calculator ac970(.scan_win(scan_win970), .rectangle1_x(rectangle1_xs[970]), .rectangle1_y(rectangle1_ys[970]), .rectangle1_width(rectangle1_widths[970]), .rectangle1_height(rectangle1_heights[970]), .rectangle1_weight(rectangle1_weights[970]), .rectangle2_x(rectangle2_xs[970]), .rectangle2_y(rectangle2_ys[970]), .rectangle2_width(rectangle2_widths[970]), .rectangle2_height(rectangle2_heights[970]), .rectangle2_weight(rectangle2_weights[970]), .rectangle3_x(rectangle3_xs[970]), .rectangle3_y(rectangle3_ys[970]), .rectangle3_width(rectangle3_widths[970]), .rectangle3_height(rectangle3_heights[970]), .rectangle3_weight(rectangle3_weights[970]), .feature_threshold(feature_thresholds[970]), .feature_above(feature_aboves[970]), .feature_below(feature_belows[970]), .scan_win_std_dev(scan_win_std_dev[970]), .feature_accum(feature_accums[970]));
  accum_calculator ac971(.scan_win(scan_win971), .rectangle1_x(rectangle1_xs[971]), .rectangle1_y(rectangle1_ys[971]), .rectangle1_width(rectangle1_widths[971]), .rectangle1_height(rectangle1_heights[971]), .rectangle1_weight(rectangle1_weights[971]), .rectangle2_x(rectangle2_xs[971]), .rectangle2_y(rectangle2_ys[971]), .rectangle2_width(rectangle2_widths[971]), .rectangle2_height(rectangle2_heights[971]), .rectangle2_weight(rectangle2_weights[971]), .rectangle3_x(rectangle3_xs[971]), .rectangle3_y(rectangle3_ys[971]), .rectangle3_width(rectangle3_widths[971]), .rectangle3_height(rectangle3_heights[971]), .rectangle3_weight(rectangle3_weights[971]), .feature_threshold(feature_thresholds[971]), .feature_above(feature_aboves[971]), .feature_below(feature_belows[971]), .scan_win_std_dev(scan_win_std_dev[971]), .feature_accum(feature_accums[971]));
  accum_calculator ac972(.scan_win(scan_win972), .rectangle1_x(rectangle1_xs[972]), .rectangle1_y(rectangle1_ys[972]), .rectangle1_width(rectangle1_widths[972]), .rectangle1_height(rectangle1_heights[972]), .rectangle1_weight(rectangle1_weights[972]), .rectangle2_x(rectangle2_xs[972]), .rectangle2_y(rectangle2_ys[972]), .rectangle2_width(rectangle2_widths[972]), .rectangle2_height(rectangle2_heights[972]), .rectangle2_weight(rectangle2_weights[972]), .rectangle3_x(rectangle3_xs[972]), .rectangle3_y(rectangle3_ys[972]), .rectangle3_width(rectangle3_widths[972]), .rectangle3_height(rectangle3_heights[972]), .rectangle3_weight(rectangle3_weights[972]), .feature_threshold(feature_thresholds[972]), .feature_above(feature_aboves[972]), .feature_below(feature_belows[972]), .scan_win_std_dev(scan_win_std_dev[972]), .feature_accum(feature_accums[972]));
  accum_calculator ac973(.scan_win(scan_win973), .rectangle1_x(rectangle1_xs[973]), .rectangle1_y(rectangle1_ys[973]), .rectangle1_width(rectangle1_widths[973]), .rectangle1_height(rectangle1_heights[973]), .rectangle1_weight(rectangle1_weights[973]), .rectangle2_x(rectangle2_xs[973]), .rectangle2_y(rectangle2_ys[973]), .rectangle2_width(rectangle2_widths[973]), .rectangle2_height(rectangle2_heights[973]), .rectangle2_weight(rectangle2_weights[973]), .rectangle3_x(rectangle3_xs[973]), .rectangle3_y(rectangle3_ys[973]), .rectangle3_width(rectangle3_widths[973]), .rectangle3_height(rectangle3_heights[973]), .rectangle3_weight(rectangle3_weights[973]), .feature_threshold(feature_thresholds[973]), .feature_above(feature_aboves[973]), .feature_below(feature_belows[973]), .scan_win_std_dev(scan_win_std_dev[973]), .feature_accum(feature_accums[973]));
  accum_calculator ac974(.scan_win(scan_win974), .rectangle1_x(rectangle1_xs[974]), .rectangle1_y(rectangle1_ys[974]), .rectangle1_width(rectangle1_widths[974]), .rectangle1_height(rectangle1_heights[974]), .rectangle1_weight(rectangle1_weights[974]), .rectangle2_x(rectangle2_xs[974]), .rectangle2_y(rectangle2_ys[974]), .rectangle2_width(rectangle2_widths[974]), .rectangle2_height(rectangle2_heights[974]), .rectangle2_weight(rectangle2_weights[974]), .rectangle3_x(rectangle3_xs[974]), .rectangle3_y(rectangle3_ys[974]), .rectangle3_width(rectangle3_widths[974]), .rectangle3_height(rectangle3_heights[974]), .rectangle3_weight(rectangle3_weights[974]), .feature_threshold(feature_thresholds[974]), .feature_above(feature_aboves[974]), .feature_below(feature_belows[974]), .scan_win_std_dev(scan_win_std_dev[974]), .feature_accum(feature_accums[974]));
  accum_calculator ac975(.scan_win(scan_win975), .rectangle1_x(rectangle1_xs[975]), .rectangle1_y(rectangle1_ys[975]), .rectangle1_width(rectangle1_widths[975]), .rectangle1_height(rectangle1_heights[975]), .rectangle1_weight(rectangle1_weights[975]), .rectangle2_x(rectangle2_xs[975]), .rectangle2_y(rectangle2_ys[975]), .rectangle2_width(rectangle2_widths[975]), .rectangle2_height(rectangle2_heights[975]), .rectangle2_weight(rectangle2_weights[975]), .rectangle3_x(rectangle3_xs[975]), .rectangle3_y(rectangle3_ys[975]), .rectangle3_width(rectangle3_widths[975]), .rectangle3_height(rectangle3_heights[975]), .rectangle3_weight(rectangle3_weights[975]), .feature_threshold(feature_thresholds[975]), .feature_above(feature_aboves[975]), .feature_below(feature_belows[975]), .scan_win_std_dev(scan_win_std_dev[975]), .feature_accum(feature_accums[975]));
  accum_calculator ac976(.scan_win(scan_win976), .rectangle1_x(rectangle1_xs[976]), .rectangle1_y(rectangle1_ys[976]), .rectangle1_width(rectangle1_widths[976]), .rectangle1_height(rectangle1_heights[976]), .rectangle1_weight(rectangle1_weights[976]), .rectangle2_x(rectangle2_xs[976]), .rectangle2_y(rectangle2_ys[976]), .rectangle2_width(rectangle2_widths[976]), .rectangle2_height(rectangle2_heights[976]), .rectangle2_weight(rectangle2_weights[976]), .rectangle3_x(rectangle3_xs[976]), .rectangle3_y(rectangle3_ys[976]), .rectangle3_width(rectangle3_widths[976]), .rectangle3_height(rectangle3_heights[976]), .rectangle3_weight(rectangle3_weights[976]), .feature_threshold(feature_thresholds[976]), .feature_above(feature_aboves[976]), .feature_below(feature_belows[976]), .scan_win_std_dev(scan_win_std_dev[976]), .feature_accum(feature_accums[976]));
  accum_calculator ac977(.scan_win(scan_win977), .rectangle1_x(rectangle1_xs[977]), .rectangle1_y(rectangle1_ys[977]), .rectangle1_width(rectangle1_widths[977]), .rectangle1_height(rectangle1_heights[977]), .rectangle1_weight(rectangle1_weights[977]), .rectangle2_x(rectangle2_xs[977]), .rectangle2_y(rectangle2_ys[977]), .rectangle2_width(rectangle2_widths[977]), .rectangle2_height(rectangle2_heights[977]), .rectangle2_weight(rectangle2_weights[977]), .rectangle3_x(rectangle3_xs[977]), .rectangle3_y(rectangle3_ys[977]), .rectangle3_width(rectangle3_widths[977]), .rectangle3_height(rectangle3_heights[977]), .rectangle3_weight(rectangle3_weights[977]), .feature_threshold(feature_thresholds[977]), .feature_above(feature_aboves[977]), .feature_below(feature_belows[977]), .scan_win_std_dev(scan_win_std_dev[977]), .feature_accum(feature_accums[977]));
  accum_calculator ac978(.scan_win(scan_win978), .rectangle1_x(rectangle1_xs[978]), .rectangle1_y(rectangle1_ys[978]), .rectangle1_width(rectangle1_widths[978]), .rectangle1_height(rectangle1_heights[978]), .rectangle1_weight(rectangle1_weights[978]), .rectangle2_x(rectangle2_xs[978]), .rectangle2_y(rectangle2_ys[978]), .rectangle2_width(rectangle2_widths[978]), .rectangle2_height(rectangle2_heights[978]), .rectangle2_weight(rectangle2_weights[978]), .rectangle3_x(rectangle3_xs[978]), .rectangle3_y(rectangle3_ys[978]), .rectangle3_width(rectangle3_widths[978]), .rectangle3_height(rectangle3_heights[978]), .rectangle3_weight(rectangle3_weights[978]), .feature_threshold(feature_thresholds[978]), .feature_above(feature_aboves[978]), .feature_below(feature_belows[978]), .scan_win_std_dev(scan_win_std_dev[978]), .feature_accum(feature_accums[978]));
  accum_calculator ac979(.scan_win(scan_win979), .rectangle1_x(rectangle1_xs[979]), .rectangle1_y(rectangle1_ys[979]), .rectangle1_width(rectangle1_widths[979]), .rectangle1_height(rectangle1_heights[979]), .rectangle1_weight(rectangle1_weights[979]), .rectangle2_x(rectangle2_xs[979]), .rectangle2_y(rectangle2_ys[979]), .rectangle2_width(rectangle2_widths[979]), .rectangle2_height(rectangle2_heights[979]), .rectangle2_weight(rectangle2_weights[979]), .rectangle3_x(rectangle3_xs[979]), .rectangle3_y(rectangle3_ys[979]), .rectangle3_width(rectangle3_widths[979]), .rectangle3_height(rectangle3_heights[979]), .rectangle3_weight(rectangle3_weights[979]), .feature_threshold(feature_thresholds[979]), .feature_above(feature_aboves[979]), .feature_below(feature_belows[979]), .scan_win_std_dev(scan_win_std_dev[979]), .feature_accum(feature_accums[979]));
  accum_calculator ac980(.scan_win(scan_win980), .rectangle1_x(rectangle1_xs[980]), .rectangle1_y(rectangle1_ys[980]), .rectangle1_width(rectangle1_widths[980]), .rectangle1_height(rectangle1_heights[980]), .rectangle1_weight(rectangle1_weights[980]), .rectangle2_x(rectangle2_xs[980]), .rectangle2_y(rectangle2_ys[980]), .rectangle2_width(rectangle2_widths[980]), .rectangle2_height(rectangle2_heights[980]), .rectangle2_weight(rectangle2_weights[980]), .rectangle3_x(rectangle3_xs[980]), .rectangle3_y(rectangle3_ys[980]), .rectangle3_width(rectangle3_widths[980]), .rectangle3_height(rectangle3_heights[980]), .rectangle3_weight(rectangle3_weights[980]), .feature_threshold(feature_thresholds[980]), .feature_above(feature_aboves[980]), .feature_below(feature_belows[980]), .scan_win_std_dev(scan_win_std_dev[980]), .feature_accum(feature_accums[980]));
  accum_calculator ac981(.scan_win(scan_win981), .rectangle1_x(rectangle1_xs[981]), .rectangle1_y(rectangle1_ys[981]), .rectangle1_width(rectangle1_widths[981]), .rectangle1_height(rectangle1_heights[981]), .rectangle1_weight(rectangle1_weights[981]), .rectangle2_x(rectangle2_xs[981]), .rectangle2_y(rectangle2_ys[981]), .rectangle2_width(rectangle2_widths[981]), .rectangle2_height(rectangle2_heights[981]), .rectangle2_weight(rectangle2_weights[981]), .rectangle3_x(rectangle3_xs[981]), .rectangle3_y(rectangle3_ys[981]), .rectangle3_width(rectangle3_widths[981]), .rectangle3_height(rectangle3_heights[981]), .rectangle3_weight(rectangle3_weights[981]), .feature_threshold(feature_thresholds[981]), .feature_above(feature_aboves[981]), .feature_below(feature_belows[981]), .scan_win_std_dev(scan_win_std_dev[981]), .feature_accum(feature_accums[981]));
  accum_calculator ac982(.scan_win(scan_win982), .rectangle1_x(rectangle1_xs[982]), .rectangle1_y(rectangle1_ys[982]), .rectangle1_width(rectangle1_widths[982]), .rectangle1_height(rectangle1_heights[982]), .rectangle1_weight(rectangle1_weights[982]), .rectangle2_x(rectangle2_xs[982]), .rectangle2_y(rectangle2_ys[982]), .rectangle2_width(rectangle2_widths[982]), .rectangle2_height(rectangle2_heights[982]), .rectangle2_weight(rectangle2_weights[982]), .rectangle3_x(rectangle3_xs[982]), .rectangle3_y(rectangle3_ys[982]), .rectangle3_width(rectangle3_widths[982]), .rectangle3_height(rectangle3_heights[982]), .rectangle3_weight(rectangle3_weights[982]), .feature_threshold(feature_thresholds[982]), .feature_above(feature_aboves[982]), .feature_below(feature_belows[982]), .scan_win_std_dev(scan_win_std_dev[982]), .feature_accum(feature_accums[982]));
  accum_calculator ac983(.scan_win(scan_win983), .rectangle1_x(rectangle1_xs[983]), .rectangle1_y(rectangle1_ys[983]), .rectangle1_width(rectangle1_widths[983]), .rectangle1_height(rectangle1_heights[983]), .rectangle1_weight(rectangle1_weights[983]), .rectangle2_x(rectangle2_xs[983]), .rectangle2_y(rectangle2_ys[983]), .rectangle2_width(rectangle2_widths[983]), .rectangle2_height(rectangle2_heights[983]), .rectangle2_weight(rectangle2_weights[983]), .rectangle3_x(rectangle3_xs[983]), .rectangle3_y(rectangle3_ys[983]), .rectangle3_width(rectangle3_widths[983]), .rectangle3_height(rectangle3_heights[983]), .rectangle3_weight(rectangle3_weights[983]), .feature_threshold(feature_thresholds[983]), .feature_above(feature_aboves[983]), .feature_below(feature_belows[983]), .scan_win_std_dev(scan_win_std_dev[983]), .feature_accum(feature_accums[983]));
  accum_calculator ac984(.scan_win(scan_win984), .rectangle1_x(rectangle1_xs[984]), .rectangle1_y(rectangle1_ys[984]), .rectangle1_width(rectangle1_widths[984]), .rectangle1_height(rectangle1_heights[984]), .rectangle1_weight(rectangle1_weights[984]), .rectangle2_x(rectangle2_xs[984]), .rectangle2_y(rectangle2_ys[984]), .rectangle2_width(rectangle2_widths[984]), .rectangle2_height(rectangle2_heights[984]), .rectangle2_weight(rectangle2_weights[984]), .rectangle3_x(rectangle3_xs[984]), .rectangle3_y(rectangle3_ys[984]), .rectangle3_width(rectangle3_widths[984]), .rectangle3_height(rectangle3_heights[984]), .rectangle3_weight(rectangle3_weights[984]), .feature_threshold(feature_thresholds[984]), .feature_above(feature_aboves[984]), .feature_below(feature_belows[984]), .scan_win_std_dev(scan_win_std_dev[984]), .feature_accum(feature_accums[984]));
  accum_calculator ac985(.scan_win(scan_win985), .rectangle1_x(rectangle1_xs[985]), .rectangle1_y(rectangle1_ys[985]), .rectangle1_width(rectangle1_widths[985]), .rectangle1_height(rectangle1_heights[985]), .rectangle1_weight(rectangle1_weights[985]), .rectangle2_x(rectangle2_xs[985]), .rectangle2_y(rectangle2_ys[985]), .rectangle2_width(rectangle2_widths[985]), .rectangle2_height(rectangle2_heights[985]), .rectangle2_weight(rectangle2_weights[985]), .rectangle3_x(rectangle3_xs[985]), .rectangle3_y(rectangle3_ys[985]), .rectangle3_width(rectangle3_widths[985]), .rectangle3_height(rectangle3_heights[985]), .rectangle3_weight(rectangle3_weights[985]), .feature_threshold(feature_thresholds[985]), .feature_above(feature_aboves[985]), .feature_below(feature_belows[985]), .scan_win_std_dev(scan_win_std_dev[985]), .feature_accum(feature_accums[985]));
  accum_calculator ac986(.scan_win(scan_win986), .rectangle1_x(rectangle1_xs[986]), .rectangle1_y(rectangle1_ys[986]), .rectangle1_width(rectangle1_widths[986]), .rectangle1_height(rectangle1_heights[986]), .rectangle1_weight(rectangle1_weights[986]), .rectangle2_x(rectangle2_xs[986]), .rectangle2_y(rectangle2_ys[986]), .rectangle2_width(rectangle2_widths[986]), .rectangle2_height(rectangle2_heights[986]), .rectangle2_weight(rectangle2_weights[986]), .rectangle3_x(rectangle3_xs[986]), .rectangle3_y(rectangle3_ys[986]), .rectangle3_width(rectangle3_widths[986]), .rectangle3_height(rectangle3_heights[986]), .rectangle3_weight(rectangle3_weights[986]), .feature_threshold(feature_thresholds[986]), .feature_above(feature_aboves[986]), .feature_below(feature_belows[986]), .scan_win_std_dev(scan_win_std_dev[986]), .feature_accum(feature_accums[986]));
  accum_calculator ac987(.scan_win(scan_win987), .rectangle1_x(rectangle1_xs[987]), .rectangle1_y(rectangle1_ys[987]), .rectangle1_width(rectangle1_widths[987]), .rectangle1_height(rectangle1_heights[987]), .rectangle1_weight(rectangle1_weights[987]), .rectangle2_x(rectangle2_xs[987]), .rectangle2_y(rectangle2_ys[987]), .rectangle2_width(rectangle2_widths[987]), .rectangle2_height(rectangle2_heights[987]), .rectangle2_weight(rectangle2_weights[987]), .rectangle3_x(rectangle3_xs[987]), .rectangle3_y(rectangle3_ys[987]), .rectangle3_width(rectangle3_widths[987]), .rectangle3_height(rectangle3_heights[987]), .rectangle3_weight(rectangle3_weights[987]), .feature_threshold(feature_thresholds[987]), .feature_above(feature_aboves[987]), .feature_below(feature_belows[987]), .scan_win_std_dev(scan_win_std_dev[987]), .feature_accum(feature_accums[987]));
  accum_calculator ac988(.scan_win(scan_win988), .rectangle1_x(rectangle1_xs[988]), .rectangle1_y(rectangle1_ys[988]), .rectangle1_width(rectangle1_widths[988]), .rectangle1_height(rectangle1_heights[988]), .rectangle1_weight(rectangle1_weights[988]), .rectangle2_x(rectangle2_xs[988]), .rectangle2_y(rectangle2_ys[988]), .rectangle2_width(rectangle2_widths[988]), .rectangle2_height(rectangle2_heights[988]), .rectangle2_weight(rectangle2_weights[988]), .rectangle3_x(rectangle3_xs[988]), .rectangle3_y(rectangle3_ys[988]), .rectangle3_width(rectangle3_widths[988]), .rectangle3_height(rectangle3_heights[988]), .rectangle3_weight(rectangle3_weights[988]), .feature_threshold(feature_thresholds[988]), .feature_above(feature_aboves[988]), .feature_below(feature_belows[988]), .scan_win_std_dev(scan_win_std_dev[988]), .feature_accum(feature_accums[988]));
  accum_calculator ac989(.scan_win(scan_win989), .rectangle1_x(rectangle1_xs[989]), .rectangle1_y(rectangle1_ys[989]), .rectangle1_width(rectangle1_widths[989]), .rectangle1_height(rectangle1_heights[989]), .rectangle1_weight(rectangle1_weights[989]), .rectangle2_x(rectangle2_xs[989]), .rectangle2_y(rectangle2_ys[989]), .rectangle2_width(rectangle2_widths[989]), .rectangle2_height(rectangle2_heights[989]), .rectangle2_weight(rectangle2_weights[989]), .rectangle3_x(rectangle3_xs[989]), .rectangle3_y(rectangle3_ys[989]), .rectangle3_width(rectangle3_widths[989]), .rectangle3_height(rectangle3_heights[989]), .rectangle3_weight(rectangle3_weights[989]), .feature_threshold(feature_thresholds[989]), .feature_above(feature_aboves[989]), .feature_below(feature_belows[989]), .scan_win_std_dev(scan_win_std_dev[989]), .feature_accum(feature_accums[989]));
  accum_calculator ac990(.scan_win(scan_win990), .rectangle1_x(rectangle1_xs[990]), .rectangle1_y(rectangle1_ys[990]), .rectangle1_width(rectangle1_widths[990]), .rectangle1_height(rectangle1_heights[990]), .rectangle1_weight(rectangle1_weights[990]), .rectangle2_x(rectangle2_xs[990]), .rectangle2_y(rectangle2_ys[990]), .rectangle2_width(rectangle2_widths[990]), .rectangle2_height(rectangle2_heights[990]), .rectangle2_weight(rectangle2_weights[990]), .rectangle3_x(rectangle3_xs[990]), .rectangle3_y(rectangle3_ys[990]), .rectangle3_width(rectangle3_widths[990]), .rectangle3_height(rectangle3_heights[990]), .rectangle3_weight(rectangle3_weights[990]), .feature_threshold(feature_thresholds[990]), .feature_above(feature_aboves[990]), .feature_below(feature_belows[990]), .scan_win_std_dev(scan_win_std_dev[990]), .feature_accum(feature_accums[990]));
  accum_calculator ac991(.scan_win(scan_win991), .rectangle1_x(rectangle1_xs[991]), .rectangle1_y(rectangle1_ys[991]), .rectangle1_width(rectangle1_widths[991]), .rectangle1_height(rectangle1_heights[991]), .rectangle1_weight(rectangle1_weights[991]), .rectangle2_x(rectangle2_xs[991]), .rectangle2_y(rectangle2_ys[991]), .rectangle2_width(rectangle2_widths[991]), .rectangle2_height(rectangle2_heights[991]), .rectangle2_weight(rectangle2_weights[991]), .rectangle3_x(rectangle3_xs[991]), .rectangle3_y(rectangle3_ys[991]), .rectangle3_width(rectangle3_widths[991]), .rectangle3_height(rectangle3_heights[991]), .rectangle3_weight(rectangle3_weights[991]), .feature_threshold(feature_thresholds[991]), .feature_above(feature_aboves[991]), .feature_below(feature_belows[991]), .scan_win_std_dev(scan_win_std_dev[991]), .feature_accum(feature_accums[991]));
  accum_calculator ac992(.scan_win(scan_win992), .rectangle1_x(rectangle1_xs[992]), .rectangle1_y(rectangle1_ys[992]), .rectangle1_width(rectangle1_widths[992]), .rectangle1_height(rectangle1_heights[992]), .rectangle1_weight(rectangle1_weights[992]), .rectangle2_x(rectangle2_xs[992]), .rectangle2_y(rectangle2_ys[992]), .rectangle2_width(rectangle2_widths[992]), .rectangle2_height(rectangle2_heights[992]), .rectangle2_weight(rectangle2_weights[992]), .rectangle3_x(rectangle3_xs[992]), .rectangle3_y(rectangle3_ys[992]), .rectangle3_width(rectangle3_widths[992]), .rectangle3_height(rectangle3_heights[992]), .rectangle3_weight(rectangle3_weights[992]), .feature_threshold(feature_thresholds[992]), .feature_above(feature_aboves[992]), .feature_below(feature_belows[992]), .scan_win_std_dev(scan_win_std_dev[992]), .feature_accum(feature_accums[992]));
  accum_calculator ac993(.scan_win(scan_win993), .rectangle1_x(rectangle1_xs[993]), .rectangle1_y(rectangle1_ys[993]), .rectangle1_width(rectangle1_widths[993]), .rectangle1_height(rectangle1_heights[993]), .rectangle1_weight(rectangle1_weights[993]), .rectangle2_x(rectangle2_xs[993]), .rectangle2_y(rectangle2_ys[993]), .rectangle2_width(rectangle2_widths[993]), .rectangle2_height(rectangle2_heights[993]), .rectangle2_weight(rectangle2_weights[993]), .rectangle3_x(rectangle3_xs[993]), .rectangle3_y(rectangle3_ys[993]), .rectangle3_width(rectangle3_widths[993]), .rectangle3_height(rectangle3_heights[993]), .rectangle3_weight(rectangle3_weights[993]), .feature_threshold(feature_thresholds[993]), .feature_above(feature_aboves[993]), .feature_below(feature_belows[993]), .scan_win_std_dev(scan_win_std_dev[993]), .feature_accum(feature_accums[993]));
  accum_calculator ac994(.scan_win(scan_win994), .rectangle1_x(rectangle1_xs[994]), .rectangle1_y(rectangle1_ys[994]), .rectangle1_width(rectangle1_widths[994]), .rectangle1_height(rectangle1_heights[994]), .rectangle1_weight(rectangle1_weights[994]), .rectangle2_x(rectangle2_xs[994]), .rectangle2_y(rectangle2_ys[994]), .rectangle2_width(rectangle2_widths[994]), .rectangle2_height(rectangle2_heights[994]), .rectangle2_weight(rectangle2_weights[994]), .rectangle3_x(rectangle3_xs[994]), .rectangle3_y(rectangle3_ys[994]), .rectangle3_width(rectangle3_widths[994]), .rectangle3_height(rectangle3_heights[994]), .rectangle3_weight(rectangle3_weights[994]), .feature_threshold(feature_thresholds[994]), .feature_above(feature_aboves[994]), .feature_below(feature_belows[994]), .scan_win_std_dev(scan_win_std_dev[994]), .feature_accum(feature_accums[994]));
  accum_calculator ac995(.scan_win(scan_win995), .rectangle1_x(rectangle1_xs[995]), .rectangle1_y(rectangle1_ys[995]), .rectangle1_width(rectangle1_widths[995]), .rectangle1_height(rectangle1_heights[995]), .rectangle1_weight(rectangle1_weights[995]), .rectangle2_x(rectangle2_xs[995]), .rectangle2_y(rectangle2_ys[995]), .rectangle2_width(rectangle2_widths[995]), .rectangle2_height(rectangle2_heights[995]), .rectangle2_weight(rectangle2_weights[995]), .rectangle3_x(rectangle3_xs[995]), .rectangle3_y(rectangle3_ys[995]), .rectangle3_width(rectangle3_widths[995]), .rectangle3_height(rectangle3_heights[995]), .rectangle3_weight(rectangle3_weights[995]), .feature_threshold(feature_thresholds[995]), .feature_above(feature_aboves[995]), .feature_below(feature_belows[995]), .scan_win_std_dev(scan_win_std_dev[995]), .feature_accum(feature_accums[995]));
  accum_calculator ac996(.scan_win(scan_win996), .rectangle1_x(rectangle1_xs[996]), .rectangle1_y(rectangle1_ys[996]), .rectangle1_width(rectangle1_widths[996]), .rectangle1_height(rectangle1_heights[996]), .rectangle1_weight(rectangle1_weights[996]), .rectangle2_x(rectangle2_xs[996]), .rectangle2_y(rectangle2_ys[996]), .rectangle2_width(rectangle2_widths[996]), .rectangle2_height(rectangle2_heights[996]), .rectangle2_weight(rectangle2_weights[996]), .rectangle3_x(rectangle3_xs[996]), .rectangle3_y(rectangle3_ys[996]), .rectangle3_width(rectangle3_widths[996]), .rectangle3_height(rectangle3_heights[996]), .rectangle3_weight(rectangle3_weights[996]), .feature_threshold(feature_thresholds[996]), .feature_above(feature_aboves[996]), .feature_below(feature_belows[996]), .scan_win_std_dev(scan_win_std_dev[996]), .feature_accum(feature_accums[996]));
  accum_calculator ac997(.scan_win(scan_win997), .rectangle1_x(rectangle1_xs[997]), .rectangle1_y(rectangle1_ys[997]), .rectangle1_width(rectangle1_widths[997]), .rectangle1_height(rectangle1_heights[997]), .rectangle1_weight(rectangle1_weights[997]), .rectangle2_x(rectangle2_xs[997]), .rectangle2_y(rectangle2_ys[997]), .rectangle2_width(rectangle2_widths[997]), .rectangle2_height(rectangle2_heights[997]), .rectangle2_weight(rectangle2_weights[997]), .rectangle3_x(rectangle3_xs[997]), .rectangle3_y(rectangle3_ys[997]), .rectangle3_width(rectangle3_widths[997]), .rectangle3_height(rectangle3_heights[997]), .rectangle3_weight(rectangle3_weights[997]), .feature_threshold(feature_thresholds[997]), .feature_above(feature_aboves[997]), .feature_below(feature_belows[997]), .scan_win_std_dev(scan_win_std_dev[997]), .feature_accum(feature_accums[997]));
  accum_calculator ac998(.scan_win(scan_win998), .rectangle1_x(rectangle1_xs[998]), .rectangle1_y(rectangle1_ys[998]), .rectangle1_width(rectangle1_widths[998]), .rectangle1_height(rectangle1_heights[998]), .rectangle1_weight(rectangle1_weights[998]), .rectangle2_x(rectangle2_xs[998]), .rectangle2_y(rectangle2_ys[998]), .rectangle2_width(rectangle2_widths[998]), .rectangle2_height(rectangle2_heights[998]), .rectangle2_weight(rectangle2_weights[998]), .rectangle3_x(rectangle3_xs[998]), .rectangle3_y(rectangle3_ys[998]), .rectangle3_width(rectangle3_widths[998]), .rectangle3_height(rectangle3_heights[998]), .rectangle3_weight(rectangle3_weights[998]), .feature_threshold(feature_thresholds[998]), .feature_above(feature_aboves[998]), .feature_below(feature_belows[998]), .scan_win_std_dev(scan_win_std_dev[998]), .feature_accum(feature_accums[998]));
  accum_calculator ac999(.scan_win(scan_win999), .rectangle1_x(rectangle1_xs[999]), .rectangle1_y(rectangle1_ys[999]), .rectangle1_width(rectangle1_widths[999]), .rectangle1_height(rectangle1_heights[999]), .rectangle1_weight(rectangle1_weights[999]), .rectangle2_x(rectangle2_xs[999]), .rectangle2_y(rectangle2_ys[999]), .rectangle2_width(rectangle2_widths[999]), .rectangle2_height(rectangle2_heights[999]), .rectangle2_weight(rectangle2_weights[999]), .rectangle3_x(rectangle3_xs[999]), .rectangle3_y(rectangle3_ys[999]), .rectangle3_width(rectangle3_widths[999]), .rectangle3_height(rectangle3_heights[999]), .rectangle3_weight(rectangle3_weights[999]), .feature_threshold(feature_thresholds[999]), .feature_above(feature_aboves[999]), .feature_below(feature_belows[999]), .scan_win_std_dev(scan_win_std_dev[999]), .feature_accum(feature_accums[999]));
  accum_calculator ac1000(.scan_win(scan_win1000), .rectangle1_x(rectangle1_xs[1000]), .rectangle1_y(rectangle1_ys[1000]), .rectangle1_width(rectangle1_widths[1000]), .rectangle1_height(rectangle1_heights[1000]), .rectangle1_weight(rectangle1_weights[1000]), .rectangle2_x(rectangle2_xs[1000]), .rectangle2_y(rectangle2_ys[1000]), .rectangle2_width(rectangle2_widths[1000]), .rectangle2_height(rectangle2_heights[1000]), .rectangle2_weight(rectangle2_weights[1000]), .rectangle3_x(rectangle3_xs[1000]), .rectangle3_y(rectangle3_ys[1000]), .rectangle3_width(rectangle3_widths[1000]), .rectangle3_height(rectangle3_heights[1000]), .rectangle3_weight(rectangle3_weights[1000]), .feature_threshold(feature_thresholds[1000]), .feature_above(feature_aboves[1000]), .feature_below(feature_belows[1000]), .scan_win_std_dev(scan_win_std_dev[1000]), .feature_accum(feature_accums[1000]));
  accum_calculator ac1001(.scan_win(scan_win1001), .rectangle1_x(rectangle1_xs[1001]), .rectangle1_y(rectangle1_ys[1001]), .rectangle1_width(rectangle1_widths[1001]), .rectangle1_height(rectangle1_heights[1001]), .rectangle1_weight(rectangle1_weights[1001]), .rectangle2_x(rectangle2_xs[1001]), .rectangle2_y(rectangle2_ys[1001]), .rectangle2_width(rectangle2_widths[1001]), .rectangle2_height(rectangle2_heights[1001]), .rectangle2_weight(rectangle2_weights[1001]), .rectangle3_x(rectangle3_xs[1001]), .rectangle3_y(rectangle3_ys[1001]), .rectangle3_width(rectangle3_widths[1001]), .rectangle3_height(rectangle3_heights[1001]), .rectangle3_weight(rectangle3_weights[1001]), .feature_threshold(feature_thresholds[1001]), .feature_above(feature_aboves[1001]), .feature_below(feature_belows[1001]), .scan_win_std_dev(scan_win_std_dev[1001]), .feature_accum(feature_accums[1001]));
  accum_calculator ac1002(.scan_win(scan_win1002), .rectangle1_x(rectangle1_xs[1002]), .rectangle1_y(rectangle1_ys[1002]), .rectangle1_width(rectangle1_widths[1002]), .rectangle1_height(rectangle1_heights[1002]), .rectangle1_weight(rectangle1_weights[1002]), .rectangle2_x(rectangle2_xs[1002]), .rectangle2_y(rectangle2_ys[1002]), .rectangle2_width(rectangle2_widths[1002]), .rectangle2_height(rectangle2_heights[1002]), .rectangle2_weight(rectangle2_weights[1002]), .rectangle3_x(rectangle3_xs[1002]), .rectangle3_y(rectangle3_ys[1002]), .rectangle3_width(rectangle3_widths[1002]), .rectangle3_height(rectangle3_heights[1002]), .rectangle3_weight(rectangle3_weights[1002]), .feature_threshold(feature_thresholds[1002]), .feature_above(feature_aboves[1002]), .feature_below(feature_belows[1002]), .scan_win_std_dev(scan_win_std_dev[1002]), .feature_accum(feature_accums[1002]));
  accum_calculator ac1003(.scan_win(scan_win1003), .rectangle1_x(rectangle1_xs[1003]), .rectangle1_y(rectangle1_ys[1003]), .rectangle1_width(rectangle1_widths[1003]), .rectangle1_height(rectangle1_heights[1003]), .rectangle1_weight(rectangle1_weights[1003]), .rectangle2_x(rectangle2_xs[1003]), .rectangle2_y(rectangle2_ys[1003]), .rectangle2_width(rectangle2_widths[1003]), .rectangle2_height(rectangle2_heights[1003]), .rectangle2_weight(rectangle2_weights[1003]), .rectangle3_x(rectangle3_xs[1003]), .rectangle3_y(rectangle3_ys[1003]), .rectangle3_width(rectangle3_widths[1003]), .rectangle3_height(rectangle3_heights[1003]), .rectangle3_weight(rectangle3_weights[1003]), .feature_threshold(feature_thresholds[1003]), .feature_above(feature_aboves[1003]), .feature_below(feature_belows[1003]), .scan_win_std_dev(scan_win_std_dev[1003]), .feature_accum(feature_accums[1003]));
  accum_calculator ac1004(.scan_win(scan_win1004), .rectangle1_x(rectangle1_xs[1004]), .rectangle1_y(rectangle1_ys[1004]), .rectangle1_width(rectangle1_widths[1004]), .rectangle1_height(rectangle1_heights[1004]), .rectangle1_weight(rectangle1_weights[1004]), .rectangle2_x(rectangle2_xs[1004]), .rectangle2_y(rectangle2_ys[1004]), .rectangle2_width(rectangle2_widths[1004]), .rectangle2_height(rectangle2_heights[1004]), .rectangle2_weight(rectangle2_weights[1004]), .rectangle3_x(rectangle3_xs[1004]), .rectangle3_y(rectangle3_ys[1004]), .rectangle3_width(rectangle3_widths[1004]), .rectangle3_height(rectangle3_heights[1004]), .rectangle3_weight(rectangle3_weights[1004]), .feature_threshold(feature_thresholds[1004]), .feature_above(feature_aboves[1004]), .feature_below(feature_belows[1004]), .scan_win_std_dev(scan_win_std_dev[1004]), .feature_accum(feature_accums[1004]));
  accum_calculator ac1005(.scan_win(scan_win1005), .rectangle1_x(rectangle1_xs[1005]), .rectangle1_y(rectangle1_ys[1005]), .rectangle1_width(rectangle1_widths[1005]), .rectangle1_height(rectangle1_heights[1005]), .rectangle1_weight(rectangle1_weights[1005]), .rectangle2_x(rectangle2_xs[1005]), .rectangle2_y(rectangle2_ys[1005]), .rectangle2_width(rectangle2_widths[1005]), .rectangle2_height(rectangle2_heights[1005]), .rectangle2_weight(rectangle2_weights[1005]), .rectangle3_x(rectangle3_xs[1005]), .rectangle3_y(rectangle3_ys[1005]), .rectangle3_width(rectangle3_widths[1005]), .rectangle3_height(rectangle3_heights[1005]), .rectangle3_weight(rectangle3_weights[1005]), .feature_threshold(feature_thresholds[1005]), .feature_above(feature_aboves[1005]), .feature_below(feature_belows[1005]), .scan_win_std_dev(scan_win_std_dev[1005]), .feature_accum(feature_accums[1005]));
  accum_calculator ac1006(.scan_win(scan_win1006), .rectangle1_x(rectangle1_xs[1006]), .rectangle1_y(rectangle1_ys[1006]), .rectangle1_width(rectangle1_widths[1006]), .rectangle1_height(rectangle1_heights[1006]), .rectangle1_weight(rectangle1_weights[1006]), .rectangle2_x(rectangle2_xs[1006]), .rectangle2_y(rectangle2_ys[1006]), .rectangle2_width(rectangle2_widths[1006]), .rectangle2_height(rectangle2_heights[1006]), .rectangle2_weight(rectangle2_weights[1006]), .rectangle3_x(rectangle3_xs[1006]), .rectangle3_y(rectangle3_ys[1006]), .rectangle3_width(rectangle3_widths[1006]), .rectangle3_height(rectangle3_heights[1006]), .rectangle3_weight(rectangle3_weights[1006]), .feature_threshold(feature_thresholds[1006]), .feature_above(feature_aboves[1006]), .feature_below(feature_belows[1006]), .scan_win_std_dev(scan_win_std_dev[1006]), .feature_accum(feature_accums[1006]));
  accum_calculator ac1007(.scan_win(scan_win1007), .rectangle1_x(rectangle1_xs[1007]), .rectangle1_y(rectangle1_ys[1007]), .rectangle1_width(rectangle1_widths[1007]), .rectangle1_height(rectangle1_heights[1007]), .rectangle1_weight(rectangle1_weights[1007]), .rectangle2_x(rectangle2_xs[1007]), .rectangle2_y(rectangle2_ys[1007]), .rectangle2_width(rectangle2_widths[1007]), .rectangle2_height(rectangle2_heights[1007]), .rectangle2_weight(rectangle2_weights[1007]), .rectangle3_x(rectangle3_xs[1007]), .rectangle3_y(rectangle3_ys[1007]), .rectangle3_width(rectangle3_widths[1007]), .rectangle3_height(rectangle3_heights[1007]), .rectangle3_weight(rectangle3_weights[1007]), .feature_threshold(feature_thresholds[1007]), .feature_above(feature_aboves[1007]), .feature_below(feature_belows[1007]), .scan_win_std_dev(scan_win_std_dev[1007]), .feature_accum(feature_accums[1007]));
  accum_calculator ac1008(.scan_win(scan_win1008), .rectangle1_x(rectangle1_xs[1008]), .rectangle1_y(rectangle1_ys[1008]), .rectangle1_width(rectangle1_widths[1008]), .rectangle1_height(rectangle1_heights[1008]), .rectangle1_weight(rectangle1_weights[1008]), .rectangle2_x(rectangle2_xs[1008]), .rectangle2_y(rectangle2_ys[1008]), .rectangle2_width(rectangle2_widths[1008]), .rectangle2_height(rectangle2_heights[1008]), .rectangle2_weight(rectangle2_weights[1008]), .rectangle3_x(rectangle3_xs[1008]), .rectangle3_y(rectangle3_ys[1008]), .rectangle3_width(rectangle3_widths[1008]), .rectangle3_height(rectangle3_heights[1008]), .rectangle3_weight(rectangle3_weights[1008]), .feature_threshold(feature_thresholds[1008]), .feature_above(feature_aboves[1008]), .feature_below(feature_belows[1008]), .scan_win_std_dev(scan_win_std_dev[1008]), .feature_accum(feature_accums[1008]));
  accum_calculator ac1009(.scan_win(scan_win1009), .rectangle1_x(rectangle1_xs[1009]), .rectangle1_y(rectangle1_ys[1009]), .rectangle1_width(rectangle1_widths[1009]), .rectangle1_height(rectangle1_heights[1009]), .rectangle1_weight(rectangle1_weights[1009]), .rectangle2_x(rectangle2_xs[1009]), .rectangle2_y(rectangle2_ys[1009]), .rectangle2_width(rectangle2_widths[1009]), .rectangle2_height(rectangle2_heights[1009]), .rectangle2_weight(rectangle2_weights[1009]), .rectangle3_x(rectangle3_xs[1009]), .rectangle3_y(rectangle3_ys[1009]), .rectangle3_width(rectangle3_widths[1009]), .rectangle3_height(rectangle3_heights[1009]), .rectangle3_weight(rectangle3_weights[1009]), .feature_threshold(feature_thresholds[1009]), .feature_above(feature_aboves[1009]), .feature_below(feature_belows[1009]), .scan_win_std_dev(scan_win_std_dev[1009]), .feature_accum(feature_accums[1009]));
  accum_calculator ac1010(.scan_win(scan_win1010), .rectangle1_x(rectangle1_xs[1010]), .rectangle1_y(rectangle1_ys[1010]), .rectangle1_width(rectangle1_widths[1010]), .rectangle1_height(rectangle1_heights[1010]), .rectangle1_weight(rectangle1_weights[1010]), .rectangle2_x(rectangle2_xs[1010]), .rectangle2_y(rectangle2_ys[1010]), .rectangle2_width(rectangle2_widths[1010]), .rectangle2_height(rectangle2_heights[1010]), .rectangle2_weight(rectangle2_weights[1010]), .rectangle3_x(rectangle3_xs[1010]), .rectangle3_y(rectangle3_ys[1010]), .rectangle3_width(rectangle3_widths[1010]), .rectangle3_height(rectangle3_heights[1010]), .rectangle3_weight(rectangle3_weights[1010]), .feature_threshold(feature_thresholds[1010]), .feature_above(feature_aboves[1010]), .feature_below(feature_belows[1010]), .scan_win_std_dev(scan_win_std_dev[1010]), .feature_accum(feature_accums[1010]));
  accum_calculator ac1011(.scan_win(scan_win1011), .rectangle1_x(rectangle1_xs[1011]), .rectangle1_y(rectangle1_ys[1011]), .rectangle1_width(rectangle1_widths[1011]), .rectangle1_height(rectangle1_heights[1011]), .rectangle1_weight(rectangle1_weights[1011]), .rectangle2_x(rectangle2_xs[1011]), .rectangle2_y(rectangle2_ys[1011]), .rectangle2_width(rectangle2_widths[1011]), .rectangle2_height(rectangle2_heights[1011]), .rectangle2_weight(rectangle2_weights[1011]), .rectangle3_x(rectangle3_xs[1011]), .rectangle3_y(rectangle3_ys[1011]), .rectangle3_width(rectangle3_widths[1011]), .rectangle3_height(rectangle3_heights[1011]), .rectangle3_weight(rectangle3_weights[1011]), .feature_threshold(feature_thresholds[1011]), .feature_above(feature_aboves[1011]), .feature_below(feature_belows[1011]), .scan_win_std_dev(scan_win_std_dev[1011]), .feature_accum(feature_accums[1011]));
  accum_calculator ac1012(.scan_win(scan_win1012), .rectangle1_x(rectangle1_xs[1012]), .rectangle1_y(rectangle1_ys[1012]), .rectangle1_width(rectangle1_widths[1012]), .rectangle1_height(rectangle1_heights[1012]), .rectangle1_weight(rectangle1_weights[1012]), .rectangle2_x(rectangle2_xs[1012]), .rectangle2_y(rectangle2_ys[1012]), .rectangle2_width(rectangle2_widths[1012]), .rectangle2_height(rectangle2_heights[1012]), .rectangle2_weight(rectangle2_weights[1012]), .rectangle3_x(rectangle3_xs[1012]), .rectangle3_y(rectangle3_ys[1012]), .rectangle3_width(rectangle3_widths[1012]), .rectangle3_height(rectangle3_heights[1012]), .rectangle3_weight(rectangle3_weights[1012]), .feature_threshold(feature_thresholds[1012]), .feature_above(feature_aboves[1012]), .feature_below(feature_belows[1012]), .scan_win_std_dev(scan_win_std_dev[1012]), .feature_accum(feature_accums[1012]));
  accum_calculator ac1013(.scan_win(scan_win1013), .rectangle1_x(rectangle1_xs[1013]), .rectangle1_y(rectangle1_ys[1013]), .rectangle1_width(rectangle1_widths[1013]), .rectangle1_height(rectangle1_heights[1013]), .rectangle1_weight(rectangle1_weights[1013]), .rectangle2_x(rectangle2_xs[1013]), .rectangle2_y(rectangle2_ys[1013]), .rectangle2_width(rectangle2_widths[1013]), .rectangle2_height(rectangle2_heights[1013]), .rectangle2_weight(rectangle2_weights[1013]), .rectangle3_x(rectangle3_xs[1013]), .rectangle3_y(rectangle3_ys[1013]), .rectangle3_width(rectangle3_widths[1013]), .rectangle3_height(rectangle3_heights[1013]), .rectangle3_weight(rectangle3_weights[1013]), .feature_threshold(feature_thresholds[1013]), .feature_above(feature_aboves[1013]), .feature_below(feature_belows[1013]), .scan_win_std_dev(scan_win_std_dev[1013]), .feature_accum(feature_accums[1013]));
  accum_calculator ac1014(.scan_win(scan_win1014), .rectangle1_x(rectangle1_xs[1014]), .rectangle1_y(rectangle1_ys[1014]), .rectangle1_width(rectangle1_widths[1014]), .rectangle1_height(rectangle1_heights[1014]), .rectangle1_weight(rectangle1_weights[1014]), .rectangle2_x(rectangle2_xs[1014]), .rectangle2_y(rectangle2_ys[1014]), .rectangle2_width(rectangle2_widths[1014]), .rectangle2_height(rectangle2_heights[1014]), .rectangle2_weight(rectangle2_weights[1014]), .rectangle3_x(rectangle3_xs[1014]), .rectangle3_y(rectangle3_ys[1014]), .rectangle3_width(rectangle3_widths[1014]), .rectangle3_height(rectangle3_heights[1014]), .rectangle3_weight(rectangle3_weights[1014]), .feature_threshold(feature_thresholds[1014]), .feature_above(feature_aboves[1014]), .feature_below(feature_belows[1014]), .scan_win_std_dev(scan_win_std_dev[1014]), .feature_accum(feature_accums[1014]));
  accum_calculator ac1015(.scan_win(scan_win1015), .rectangle1_x(rectangle1_xs[1015]), .rectangle1_y(rectangle1_ys[1015]), .rectangle1_width(rectangle1_widths[1015]), .rectangle1_height(rectangle1_heights[1015]), .rectangle1_weight(rectangle1_weights[1015]), .rectangle2_x(rectangle2_xs[1015]), .rectangle2_y(rectangle2_ys[1015]), .rectangle2_width(rectangle2_widths[1015]), .rectangle2_height(rectangle2_heights[1015]), .rectangle2_weight(rectangle2_weights[1015]), .rectangle3_x(rectangle3_xs[1015]), .rectangle3_y(rectangle3_ys[1015]), .rectangle3_width(rectangle3_widths[1015]), .rectangle3_height(rectangle3_heights[1015]), .rectangle3_weight(rectangle3_weights[1015]), .feature_threshold(feature_thresholds[1015]), .feature_above(feature_aboves[1015]), .feature_below(feature_belows[1015]), .scan_win_std_dev(scan_win_std_dev[1015]), .feature_accum(feature_accums[1015]));
  accum_calculator ac1016(.scan_win(scan_win1016), .rectangle1_x(rectangle1_xs[1016]), .rectangle1_y(rectangle1_ys[1016]), .rectangle1_width(rectangle1_widths[1016]), .rectangle1_height(rectangle1_heights[1016]), .rectangle1_weight(rectangle1_weights[1016]), .rectangle2_x(rectangle2_xs[1016]), .rectangle2_y(rectangle2_ys[1016]), .rectangle2_width(rectangle2_widths[1016]), .rectangle2_height(rectangle2_heights[1016]), .rectangle2_weight(rectangle2_weights[1016]), .rectangle3_x(rectangle3_xs[1016]), .rectangle3_y(rectangle3_ys[1016]), .rectangle3_width(rectangle3_widths[1016]), .rectangle3_height(rectangle3_heights[1016]), .rectangle3_weight(rectangle3_weights[1016]), .feature_threshold(feature_thresholds[1016]), .feature_above(feature_aboves[1016]), .feature_below(feature_belows[1016]), .scan_win_std_dev(scan_win_std_dev[1016]), .feature_accum(feature_accums[1016]));
  accum_calculator ac1017(.scan_win(scan_win1017), .rectangle1_x(rectangle1_xs[1017]), .rectangle1_y(rectangle1_ys[1017]), .rectangle1_width(rectangle1_widths[1017]), .rectangle1_height(rectangle1_heights[1017]), .rectangle1_weight(rectangle1_weights[1017]), .rectangle2_x(rectangle2_xs[1017]), .rectangle2_y(rectangle2_ys[1017]), .rectangle2_width(rectangle2_widths[1017]), .rectangle2_height(rectangle2_heights[1017]), .rectangle2_weight(rectangle2_weights[1017]), .rectangle3_x(rectangle3_xs[1017]), .rectangle3_y(rectangle3_ys[1017]), .rectangle3_width(rectangle3_widths[1017]), .rectangle3_height(rectangle3_heights[1017]), .rectangle3_weight(rectangle3_weights[1017]), .feature_threshold(feature_thresholds[1017]), .feature_above(feature_aboves[1017]), .feature_below(feature_belows[1017]), .scan_win_std_dev(scan_win_std_dev[1017]), .feature_accum(feature_accums[1017]));
  accum_calculator ac1018(.scan_win(scan_win1018), .rectangle1_x(rectangle1_xs[1018]), .rectangle1_y(rectangle1_ys[1018]), .rectangle1_width(rectangle1_widths[1018]), .rectangle1_height(rectangle1_heights[1018]), .rectangle1_weight(rectangle1_weights[1018]), .rectangle2_x(rectangle2_xs[1018]), .rectangle2_y(rectangle2_ys[1018]), .rectangle2_width(rectangle2_widths[1018]), .rectangle2_height(rectangle2_heights[1018]), .rectangle2_weight(rectangle2_weights[1018]), .rectangle3_x(rectangle3_xs[1018]), .rectangle3_y(rectangle3_ys[1018]), .rectangle3_width(rectangle3_widths[1018]), .rectangle3_height(rectangle3_heights[1018]), .rectangle3_weight(rectangle3_weights[1018]), .feature_threshold(feature_thresholds[1018]), .feature_above(feature_aboves[1018]), .feature_below(feature_belows[1018]), .scan_win_std_dev(scan_win_std_dev[1018]), .feature_accum(feature_accums[1018]));
  accum_calculator ac1019(.scan_win(scan_win1019), .rectangle1_x(rectangle1_xs[1019]), .rectangle1_y(rectangle1_ys[1019]), .rectangle1_width(rectangle1_widths[1019]), .rectangle1_height(rectangle1_heights[1019]), .rectangle1_weight(rectangle1_weights[1019]), .rectangle2_x(rectangle2_xs[1019]), .rectangle2_y(rectangle2_ys[1019]), .rectangle2_width(rectangle2_widths[1019]), .rectangle2_height(rectangle2_heights[1019]), .rectangle2_weight(rectangle2_weights[1019]), .rectangle3_x(rectangle3_xs[1019]), .rectangle3_y(rectangle3_ys[1019]), .rectangle3_width(rectangle3_widths[1019]), .rectangle3_height(rectangle3_heights[1019]), .rectangle3_weight(rectangle3_weights[1019]), .feature_threshold(feature_thresholds[1019]), .feature_above(feature_aboves[1019]), .feature_below(feature_belows[1019]), .scan_win_std_dev(scan_win_std_dev[1019]), .feature_accum(feature_accums[1019]));
  accum_calculator ac1020(.scan_win(scan_win1020), .rectangle1_x(rectangle1_xs[1020]), .rectangle1_y(rectangle1_ys[1020]), .rectangle1_width(rectangle1_widths[1020]), .rectangle1_height(rectangle1_heights[1020]), .rectangle1_weight(rectangle1_weights[1020]), .rectangle2_x(rectangle2_xs[1020]), .rectangle2_y(rectangle2_ys[1020]), .rectangle2_width(rectangle2_widths[1020]), .rectangle2_height(rectangle2_heights[1020]), .rectangle2_weight(rectangle2_weights[1020]), .rectangle3_x(rectangle3_xs[1020]), .rectangle3_y(rectangle3_ys[1020]), .rectangle3_width(rectangle3_widths[1020]), .rectangle3_height(rectangle3_heights[1020]), .rectangle3_weight(rectangle3_weights[1020]), .feature_threshold(feature_thresholds[1020]), .feature_above(feature_aboves[1020]), .feature_below(feature_belows[1020]), .scan_win_std_dev(scan_win_std_dev[1020]), .feature_accum(feature_accums[1020]));
  accum_calculator ac1021(.scan_win(scan_win1021), .rectangle1_x(rectangle1_xs[1021]), .rectangle1_y(rectangle1_ys[1021]), .rectangle1_width(rectangle1_widths[1021]), .rectangle1_height(rectangle1_heights[1021]), .rectangle1_weight(rectangle1_weights[1021]), .rectangle2_x(rectangle2_xs[1021]), .rectangle2_y(rectangle2_ys[1021]), .rectangle2_width(rectangle2_widths[1021]), .rectangle2_height(rectangle2_heights[1021]), .rectangle2_weight(rectangle2_weights[1021]), .rectangle3_x(rectangle3_xs[1021]), .rectangle3_y(rectangle3_ys[1021]), .rectangle3_width(rectangle3_widths[1021]), .rectangle3_height(rectangle3_heights[1021]), .rectangle3_weight(rectangle3_weights[1021]), .feature_threshold(feature_thresholds[1021]), .feature_above(feature_aboves[1021]), .feature_below(feature_belows[1021]), .scan_win_std_dev(scan_win_std_dev[1021]), .feature_accum(feature_accums[1021]));
  accum_calculator ac1022(.scan_win(scan_win1022), .rectangle1_x(rectangle1_xs[1022]), .rectangle1_y(rectangle1_ys[1022]), .rectangle1_width(rectangle1_widths[1022]), .rectangle1_height(rectangle1_heights[1022]), .rectangle1_weight(rectangle1_weights[1022]), .rectangle2_x(rectangle2_xs[1022]), .rectangle2_y(rectangle2_ys[1022]), .rectangle2_width(rectangle2_widths[1022]), .rectangle2_height(rectangle2_heights[1022]), .rectangle2_weight(rectangle2_weights[1022]), .rectangle3_x(rectangle3_xs[1022]), .rectangle3_y(rectangle3_ys[1022]), .rectangle3_width(rectangle3_widths[1022]), .rectangle3_height(rectangle3_heights[1022]), .rectangle3_weight(rectangle3_weights[1022]), .feature_threshold(feature_thresholds[1022]), .feature_above(feature_aboves[1022]), .feature_below(feature_belows[1022]), .scan_win_std_dev(scan_win_std_dev[1022]), .feature_accum(feature_accums[1022]));
  accum_calculator ac1023(.scan_win(scan_win1023), .rectangle1_x(rectangle1_xs[1023]), .rectangle1_y(rectangle1_ys[1023]), .rectangle1_width(rectangle1_widths[1023]), .rectangle1_height(rectangle1_heights[1023]), .rectangle1_weight(rectangle1_weights[1023]), .rectangle2_x(rectangle2_xs[1023]), .rectangle2_y(rectangle2_ys[1023]), .rectangle2_width(rectangle2_widths[1023]), .rectangle2_height(rectangle2_heights[1023]), .rectangle2_weight(rectangle2_weights[1023]), .rectangle3_x(rectangle3_xs[1023]), .rectangle3_y(rectangle3_ys[1023]), .rectangle3_width(rectangle3_widths[1023]), .rectangle3_height(rectangle3_heights[1023]), .rectangle3_weight(rectangle3_weights[1023]), .feature_threshold(feature_thresholds[1023]), .feature_above(feature_aboves[1023]), .feature_below(feature_belows[1023]), .scan_win_std_dev(scan_win_std_dev[1023]), .feature_accum(feature_accums[1023]));
  accum_calculator ac1024(.scan_win(scan_win1024), .rectangle1_x(rectangle1_xs[1024]), .rectangle1_y(rectangle1_ys[1024]), .rectangle1_width(rectangle1_widths[1024]), .rectangle1_height(rectangle1_heights[1024]), .rectangle1_weight(rectangle1_weights[1024]), .rectangle2_x(rectangle2_xs[1024]), .rectangle2_y(rectangle2_ys[1024]), .rectangle2_width(rectangle2_widths[1024]), .rectangle2_height(rectangle2_heights[1024]), .rectangle2_weight(rectangle2_weights[1024]), .rectangle3_x(rectangle3_xs[1024]), .rectangle3_y(rectangle3_ys[1024]), .rectangle3_width(rectangle3_widths[1024]), .rectangle3_height(rectangle3_heights[1024]), .rectangle3_weight(rectangle3_weights[1024]), .feature_threshold(feature_thresholds[1024]), .feature_above(feature_aboves[1024]), .feature_below(feature_belows[1024]), .scan_win_std_dev(scan_win_std_dev[1024]), .feature_accum(feature_accums[1024]));
  accum_calculator ac1025(.scan_win(scan_win1025), .rectangle1_x(rectangle1_xs[1025]), .rectangle1_y(rectangle1_ys[1025]), .rectangle1_width(rectangle1_widths[1025]), .rectangle1_height(rectangle1_heights[1025]), .rectangle1_weight(rectangle1_weights[1025]), .rectangle2_x(rectangle2_xs[1025]), .rectangle2_y(rectangle2_ys[1025]), .rectangle2_width(rectangle2_widths[1025]), .rectangle2_height(rectangle2_heights[1025]), .rectangle2_weight(rectangle2_weights[1025]), .rectangle3_x(rectangle3_xs[1025]), .rectangle3_y(rectangle3_ys[1025]), .rectangle3_width(rectangle3_widths[1025]), .rectangle3_height(rectangle3_heights[1025]), .rectangle3_weight(rectangle3_weights[1025]), .feature_threshold(feature_thresholds[1025]), .feature_above(feature_aboves[1025]), .feature_below(feature_belows[1025]), .scan_win_std_dev(scan_win_std_dev[1025]), .feature_accum(feature_accums[1025]));
  accum_calculator ac1026(.scan_win(scan_win1026), .rectangle1_x(rectangle1_xs[1026]), .rectangle1_y(rectangle1_ys[1026]), .rectangle1_width(rectangle1_widths[1026]), .rectangle1_height(rectangle1_heights[1026]), .rectangle1_weight(rectangle1_weights[1026]), .rectangle2_x(rectangle2_xs[1026]), .rectangle2_y(rectangle2_ys[1026]), .rectangle2_width(rectangle2_widths[1026]), .rectangle2_height(rectangle2_heights[1026]), .rectangle2_weight(rectangle2_weights[1026]), .rectangle3_x(rectangle3_xs[1026]), .rectangle3_y(rectangle3_ys[1026]), .rectangle3_width(rectangle3_widths[1026]), .rectangle3_height(rectangle3_heights[1026]), .rectangle3_weight(rectangle3_weights[1026]), .feature_threshold(feature_thresholds[1026]), .feature_above(feature_aboves[1026]), .feature_below(feature_belows[1026]), .scan_win_std_dev(scan_win_std_dev[1026]), .feature_accum(feature_accums[1026]));
  accum_calculator ac1027(.scan_win(scan_win1027), .rectangle1_x(rectangle1_xs[1027]), .rectangle1_y(rectangle1_ys[1027]), .rectangle1_width(rectangle1_widths[1027]), .rectangle1_height(rectangle1_heights[1027]), .rectangle1_weight(rectangle1_weights[1027]), .rectangle2_x(rectangle2_xs[1027]), .rectangle2_y(rectangle2_ys[1027]), .rectangle2_width(rectangle2_widths[1027]), .rectangle2_height(rectangle2_heights[1027]), .rectangle2_weight(rectangle2_weights[1027]), .rectangle3_x(rectangle3_xs[1027]), .rectangle3_y(rectangle3_ys[1027]), .rectangle3_width(rectangle3_widths[1027]), .rectangle3_height(rectangle3_heights[1027]), .rectangle3_weight(rectangle3_weights[1027]), .feature_threshold(feature_thresholds[1027]), .feature_above(feature_aboves[1027]), .feature_below(feature_belows[1027]), .scan_win_std_dev(scan_win_std_dev[1027]), .feature_accum(feature_accums[1027]));
  accum_calculator ac1028(.scan_win(scan_win1028), .rectangle1_x(rectangle1_xs[1028]), .rectangle1_y(rectangle1_ys[1028]), .rectangle1_width(rectangle1_widths[1028]), .rectangle1_height(rectangle1_heights[1028]), .rectangle1_weight(rectangle1_weights[1028]), .rectangle2_x(rectangle2_xs[1028]), .rectangle2_y(rectangle2_ys[1028]), .rectangle2_width(rectangle2_widths[1028]), .rectangle2_height(rectangle2_heights[1028]), .rectangle2_weight(rectangle2_weights[1028]), .rectangle3_x(rectangle3_xs[1028]), .rectangle3_y(rectangle3_ys[1028]), .rectangle3_width(rectangle3_widths[1028]), .rectangle3_height(rectangle3_heights[1028]), .rectangle3_weight(rectangle3_weights[1028]), .feature_threshold(feature_thresholds[1028]), .feature_above(feature_aboves[1028]), .feature_below(feature_belows[1028]), .scan_win_std_dev(scan_win_std_dev[1028]), .feature_accum(feature_accums[1028]));
  accum_calculator ac1029(.scan_win(scan_win1029), .rectangle1_x(rectangle1_xs[1029]), .rectangle1_y(rectangle1_ys[1029]), .rectangle1_width(rectangle1_widths[1029]), .rectangle1_height(rectangle1_heights[1029]), .rectangle1_weight(rectangle1_weights[1029]), .rectangle2_x(rectangle2_xs[1029]), .rectangle2_y(rectangle2_ys[1029]), .rectangle2_width(rectangle2_widths[1029]), .rectangle2_height(rectangle2_heights[1029]), .rectangle2_weight(rectangle2_weights[1029]), .rectangle3_x(rectangle3_xs[1029]), .rectangle3_y(rectangle3_ys[1029]), .rectangle3_width(rectangle3_widths[1029]), .rectangle3_height(rectangle3_heights[1029]), .rectangle3_weight(rectangle3_weights[1029]), .feature_threshold(feature_thresholds[1029]), .feature_above(feature_aboves[1029]), .feature_below(feature_belows[1029]), .scan_win_std_dev(scan_win_std_dev[1029]), .feature_accum(feature_accums[1029]));
  accum_calculator ac1030(.scan_win(scan_win1030), .rectangle1_x(rectangle1_xs[1030]), .rectangle1_y(rectangle1_ys[1030]), .rectangle1_width(rectangle1_widths[1030]), .rectangle1_height(rectangle1_heights[1030]), .rectangle1_weight(rectangle1_weights[1030]), .rectangle2_x(rectangle2_xs[1030]), .rectangle2_y(rectangle2_ys[1030]), .rectangle2_width(rectangle2_widths[1030]), .rectangle2_height(rectangle2_heights[1030]), .rectangle2_weight(rectangle2_weights[1030]), .rectangle3_x(rectangle3_xs[1030]), .rectangle3_y(rectangle3_ys[1030]), .rectangle3_width(rectangle3_widths[1030]), .rectangle3_height(rectangle3_heights[1030]), .rectangle3_weight(rectangle3_weights[1030]), .feature_threshold(feature_thresholds[1030]), .feature_above(feature_aboves[1030]), .feature_below(feature_belows[1030]), .scan_win_std_dev(scan_win_std_dev[1030]), .feature_accum(feature_accums[1030]));
  accum_calculator ac1031(.scan_win(scan_win1031), .rectangle1_x(rectangle1_xs[1031]), .rectangle1_y(rectangle1_ys[1031]), .rectangle1_width(rectangle1_widths[1031]), .rectangle1_height(rectangle1_heights[1031]), .rectangle1_weight(rectangle1_weights[1031]), .rectangle2_x(rectangle2_xs[1031]), .rectangle2_y(rectangle2_ys[1031]), .rectangle2_width(rectangle2_widths[1031]), .rectangle2_height(rectangle2_heights[1031]), .rectangle2_weight(rectangle2_weights[1031]), .rectangle3_x(rectangle3_xs[1031]), .rectangle3_y(rectangle3_ys[1031]), .rectangle3_width(rectangle3_widths[1031]), .rectangle3_height(rectangle3_heights[1031]), .rectangle3_weight(rectangle3_weights[1031]), .feature_threshold(feature_thresholds[1031]), .feature_above(feature_aboves[1031]), .feature_below(feature_belows[1031]), .scan_win_std_dev(scan_win_std_dev[1031]), .feature_accum(feature_accums[1031]));
  accum_calculator ac1032(.scan_win(scan_win1032), .rectangle1_x(rectangle1_xs[1032]), .rectangle1_y(rectangle1_ys[1032]), .rectangle1_width(rectangle1_widths[1032]), .rectangle1_height(rectangle1_heights[1032]), .rectangle1_weight(rectangle1_weights[1032]), .rectangle2_x(rectangle2_xs[1032]), .rectangle2_y(rectangle2_ys[1032]), .rectangle2_width(rectangle2_widths[1032]), .rectangle2_height(rectangle2_heights[1032]), .rectangle2_weight(rectangle2_weights[1032]), .rectangle3_x(rectangle3_xs[1032]), .rectangle3_y(rectangle3_ys[1032]), .rectangle3_width(rectangle3_widths[1032]), .rectangle3_height(rectangle3_heights[1032]), .rectangle3_weight(rectangle3_weights[1032]), .feature_threshold(feature_thresholds[1032]), .feature_above(feature_aboves[1032]), .feature_below(feature_belows[1032]), .scan_win_std_dev(scan_win_std_dev[1032]), .feature_accum(feature_accums[1032]));
  accum_calculator ac1033(.scan_win(scan_win1033), .rectangle1_x(rectangle1_xs[1033]), .rectangle1_y(rectangle1_ys[1033]), .rectangle1_width(rectangle1_widths[1033]), .rectangle1_height(rectangle1_heights[1033]), .rectangle1_weight(rectangle1_weights[1033]), .rectangle2_x(rectangle2_xs[1033]), .rectangle2_y(rectangle2_ys[1033]), .rectangle2_width(rectangle2_widths[1033]), .rectangle2_height(rectangle2_heights[1033]), .rectangle2_weight(rectangle2_weights[1033]), .rectangle3_x(rectangle3_xs[1033]), .rectangle3_y(rectangle3_ys[1033]), .rectangle3_width(rectangle3_widths[1033]), .rectangle3_height(rectangle3_heights[1033]), .rectangle3_weight(rectangle3_weights[1033]), .feature_threshold(feature_thresholds[1033]), .feature_above(feature_aboves[1033]), .feature_below(feature_belows[1033]), .scan_win_std_dev(scan_win_std_dev[1033]), .feature_accum(feature_accums[1033]));
  accum_calculator ac1034(.scan_win(scan_win1034), .rectangle1_x(rectangle1_xs[1034]), .rectangle1_y(rectangle1_ys[1034]), .rectangle1_width(rectangle1_widths[1034]), .rectangle1_height(rectangle1_heights[1034]), .rectangle1_weight(rectangle1_weights[1034]), .rectangle2_x(rectangle2_xs[1034]), .rectangle2_y(rectangle2_ys[1034]), .rectangle2_width(rectangle2_widths[1034]), .rectangle2_height(rectangle2_heights[1034]), .rectangle2_weight(rectangle2_weights[1034]), .rectangle3_x(rectangle3_xs[1034]), .rectangle3_y(rectangle3_ys[1034]), .rectangle3_width(rectangle3_widths[1034]), .rectangle3_height(rectangle3_heights[1034]), .rectangle3_weight(rectangle3_weights[1034]), .feature_threshold(feature_thresholds[1034]), .feature_above(feature_aboves[1034]), .feature_below(feature_belows[1034]), .scan_win_std_dev(scan_win_std_dev[1034]), .feature_accum(feature_accums[1034]));
  accum_calculator ac1035(.scan_win(scan_win1035), .rectangle1_x(rectangle1_xs[1035]), .rectangle1_y(rectangle1_ys[1035]), .rectangle1_width(rectangle1_widths[1035]), .rectangle1_height(rectangle1_heights[1035]), .rectangle1_weight(rectangle1_weights[1035]), .rectangle2_x(rectangle2_xs[1035]), .rectangle2_y(rectangle2_ys[1035]), .rectangle2_width(rectangle2_widths[1035]), .rectangle2_height(rectangle2_heights[1035]), .rectangle2_weight(rectangle2_weights[1035]), .rectangle3_x(rectangle3_xs[1035]), .rectangle3_y(rectangle3_ys[1035]), .rectangle3_width(rectangle3_widths[1035]), .rectangle3_height(rectangle3_heights[1035]), .rectangle3_weight(rectangle3_weights[1035]), .feature_threshold(feature_thresholds[1035]), .feature_above(feature_aboves[1035]), .feature_below(feature_belows[1035]), .scan_win_std_dev(scan_win_std_dev[1035]), .feature_accum(feature_accums[1035]));
  accum_calculator ac1036(.scan_win(scan_win1036), .rectangle1_x(rectangle1_xs[1036]), .rectangle1_y(rectangle1_ys[1036]), .rectangle1_width(rectangle1_widths[1036]), .rectangle1_height(rectangle1_heights[1036]), .rectangle1_weight(rectangle1_weights[1036]), .rectangle2_x(rectangle2_xs[1036]), .rectangle2_y(rectangle2_ys[1036]), .rectangle2_width(rectangle2_widths[1036]), .rectangle2_height(rectangle2_heights[1036]), .rectangle2_weight(rectangle2_weights[1036]), .rectangle3_x(rectangle3_xs[1036]), .rectangle3_y(rectangle3_ys[1036]), .rectangle3_width(rectangle3_widths[1036]), .rectangle3_height(rectangle3_heights[1036]), .rectangle3_weight(rectangle3_weights[1036]), .feature_threshold(feature_thresholds[1036]), .feature_above(feature_aboves[1036]), .feature_below(feature_belows[1036]), .scan_win_std_dev(scan_win_std_dev[1036]), .feature_accum(feature_accums[1036]));
  accum_calculator ac1037(.scan_win(scan_win1037), .rectangle1_x(rectangle1_xs[1037]), .rectangle1_y(rectangle1_ys[1037]), .rectangle1_width(rectangle1_widths[1037]), .rectangle1_height(rectangle1_heights[1037]), .rectangle1_weight(rectangle1_weights[1037]), .rectangle2_x(rectangle2_xs[1037]), .rectangle2_y(rectangle2_ys[1037]), .rectangle2_width(rectangle2_widths[1037]), .rectangle2_height(rectangle2_heights[1037]), .rectangle2_weight(rectangle2_weights[1037]), .rectangle3_x(rectangle3_xs[1037]), .rectangle3_y(rectangle3_ys[1037]), .rectangle3_width(rectangle3_widths[1037]), .rectangle3_height(rectangle3_heights[1037]), .rectangle3_weight(rectangle3_weights[1037]), .feature_threshold(feature_thresholds[1037]), .feature_above(feature_aboves[1037]), .feature_below(feature_belows[1037]), .scan_win_std_dev(scan_win_std_dev[1037]), .feature_accum(feature_accums[1037]));
  accum_calculator ac1038(.scan_win(scan_win1038), .rectangle1_x(rectangle1_xs[1038]), .rectangle1_y(rectangle1_ys[1038]), .rectangle1_width(rectangle1_widths[1038]), .rectangle1_height(rectangle1_heights[1038]), .rectangle1_weight(rectangle1_weights[1038]), .rectangle2_x(rectangle2_xs[1038]), .rectangle2_y(rectangle2_ys[1038]), .rectangle2_width(rectangle2_widths[1038]), .rectangle2_height(rectangle2_heights[1038]), .rectangle2_weight(rectangle2_weights[1038]), .rectangle3_x(rectangle3_xs[1038]), .rectangle3_y(rectangle3_ys[1038]), .rectangle3_width(rectangle3_widths[1038]), .rectangle3_height(rectangle3_heights[1038]), .rectangle3_weight(rectangle3_weights[1038]), .feature_threshold(feature_thresholds[1038]), .feature_above(feature_aboves[1038]), .feature_below(feature_belows[1038]), .scan_win_std_dev(scan_win_std_dev[1038]), .feature_accum(feature_accums[1038]));
  accum_calculator ac1039(.scan_win(scan_win1039), .rectangle1_x(rectangle1_xs[1039]), .rectangle1_y(rectangle1_ys[1039]), .rectangle1_width(rectangle1_widths[1039]), .rectangle1_height(rectangle1_heights[1039]), .rectangle1_weight(rectangle1_weights[1039]), .rectangle2_x(rectangle2_xs[1039]), .rectangle2_y(rectangle2_ys[1039]), .rectangle2_width(rectangle2_widths[1039]), .rectangle2_height(rectangle2_heights[1039]), .rectangle2_weight(rectangle2_weights[1039]), .rectangle3_x(rectangle3_xs[1039]), .rectangle3_y(rectangle3_ys[1039]), .rectangle3_width(rectangle3_widths[1039]), .rectangle3_height(rectangle3_heights[1039]), .rectangle3_weight(rectangle3_weights[1039]), .feature_threshold(feature_thresholds[1039]), .feature_above(feature_aboves[1039]), .feature_below(feature_belows[1039]), .scan_win_std_dev(scan_win_std_dev[1039]), .feature_accum(feature_accums[1039]));
  accum_calculator ac1040(.scan_win(scan_win1040), .rectangle1_x(rectangle1_xs[1040]), .rectangle1_y(rectangle1_ys[1040]), .rectangle1_width(rectangle1_widths[1040]), .rectangle1_height(rectangle1_heights[1040]), .rectangle1_weight(rectangle1_weights[1040]), .rectangle2_x(rectangle2_xs[1040]), .rectangle2_y(rectangle2_ys[1040]), .rectangle2_width(rectangle2_widths[1040]), .rectangle2_height(rectangle2_heights[1040]), .rectangle2_weight(rectangle2_weights[1040]), .rectangle3_x(rectangle3_xs[1040]), .rectangle3_y(rectangle3_ys[1040]), .rectangle3_width(rectangle3_widths[1040]), .rectangle3_height(rectangle3_heights[1040]), .rectangle3_weight(rectangle3_weights[1040]), .feature_threshold(feature_thresholds[1040]), .feature_above(feature_aboves[1040]), .feature_below(feature_belows[1040]), .scan_win_std_dev(scan_win_std_dev[1040]), .feature_accum(feature_accums[1040]));
  accum_calculator ac1041(.scan_win(scan_win1041), .rectangle1_x(rectangle1_xs[1041]), .rectangle1_y(rectangle1_ys[1041]), .rectangle1_width(rectangle1_widths[1041]), .rectangle1_height(rectangle1_heights[1041]), .rectangle1_weight(rectangle1_weights[1041]), .rectangle2_x(rectangle2_xs[1041]), .rectangle2_y(rectangle2_ys[1041]), .rectangle2_width(rectangle2_widths[1041]), .rectangle2_height(rectangle2_heights[1041]), .rectangle2_weight(rectangle2_weights[1041]), .rectangle3_x(rectangle3_xs[1041]), .rectangle3_y(rectangle3_ys[1041]), .rectangle3_width(rectangle3_widths[1041]), .rectangle3_height(rectangle3_heights[1041]), .rectangle3_weight(rectangle3_weights[1041]), .feature_threshold(feature_thresholds[1041]), .feature_above(feature_aboves[1041]), .feature_below(feature_belows[1041]), .scan_win_std_dev(scan_win_std_dev[1041]), .feature_accum(feature_accums[1041]));
  accum_calculator ac1042(.scan_win(scan_win1042), .rectangle1_x(rectangle1_xs[1042]), .rectangle1_y(rectangle1_ys[1042]), .rectangle1_width(rectangle1_widths[1042]), .rectangle1_height(rectangle1_heights[1042]), .rectangle1_weight(rectangle1_weights[1042]), .rectangle2_x(rectangle2_xs[1042]), .rectangle2_y(rectangle2_ys[1042]), .rectangle2_width(rectangle2_widths[1042]), .rectangle2_height(rectangle2_heights[1042]), .rectangle2_weight(rectangle2_weights[1042]), .rectangle3_x(rectangle3_xs[1042]), .rectangle3_y(rectangle3_ys[1042]), .rectangle3_width(rectangle3_widths[1042]), .rectangle3_height(rectangle3_heights[1042]), .rectangle3_weight(rectangle3_weights[1042]), .feature_threshold(feature_thresholds[1042]), .feature_above(feature_aboves[1042]), .feature_below(feature_belows[1042]), .scan_win_std_dev(scan_win_std_dev[1042]), .feature_accum(feature_accums[1042]));
  accum_calculator ac1043(.scan_win(scan_win1043), .rectangle1_x(rectangle1_xs[1043]), .rectangle1_y(rectangle1_ys[1043]), .rectangle1_width(rectangle1_widths[1043]), .rectangle1_height(rectangle1_heights[1043]), .rectangle1_weight(rectangle1_weights[1043]), .rectangle2_x(rectangle2_xs[1043]), .rectangle2_y(rectangle2_ys[1043]), .rectangle2_width(rectangle2_widths[1043]), .rectangle2_height(rectangle2_heights[1043]), .rectangle2_weight(rectangle2_weights[1043]), .rectangle3_x(rectangle3_xs[1043]), .rectangle3_y(rectangle3_ys[1043]), .rectangle3_width(rectangle3_widths[1043]), .rectangle3_height(rectangle3_heights[1043]), .rectangle3_weight(rectangle3_weights[1043]), .feature_threshold(feature_thresholds[1043]), .feature_above(feature_aboves[1043]), .feature_below(feature_belows[1043]), .scan_win_std_dev(scan_win_std_dev[1043]), .feature_accum(feature_accums[1043]));
  accum_calculator ac1044(.scan_win(scan_win1044), .rectangle1_x(rectangle1_xs[1044]), .rectangle1_y(rectangle1_ys[1044]), .rectangle1_width(rectangle1_widths[1044]), .rectangle1_height(rectangle1_heights[1044]), .rectangle1_weight(rectangle1_weights[1044]), .rectangle2_x(rectangle2_xs[1044]), .rectangle2_y(rectangle2_ys[1044]), .rectangle2_width(rectangle2_widths[1044]), .rectangle2_height(rectangle2_heights[1044]), .rectangle2_weight(rectangle2_weights[1044]), .rectangle3_x(rectangle3_xs[1044]), .rectangle3_y(rectangle3_ys[1044]), .rectangle3_width(rectangle3_widths[1044]), .rectangle3_height(rectangle3_heights[1044]), .rectangle3_weight(rectangle3_weights[1044]), .feature_threshold(feature_thresholds[1044]), .feature_above(feature_aboves[1044]), .feature_below(feature_belows[1044]), .scan_win_std_dev(scan_win_std_dev[1044]), .feature_accum(feature_accums[1044]));
  accum_calculator ac1045(.scan_win(scan_win1045), .rectangle1_x(rectangle1_xs[1045]), .rectangle1_y(rectangle1_ys[1045]), .rectangle1_width(rectangle1_widths[1045]), .rectangle1_height(rectangle1_heights[1045]), .rectangle1_weight(rectangle1_weights[1045]), .rectangle2_x(rectangle2_xs[1045]), .rectangle2_y(rectangle2_ys[1045]), .rectangle2_width(rectangle2_widths[1045]), .rectangle2_height(rectangle2_heights[1045]), .rectangle2_weight(rectangle2_weights[1045]), .rectangle3_x(rectangle3_xs[1045]), .rectangle3_y(rectangle3_ys[1045]), .rectangle3_width(rectangle3_widths[1045]), .rectangle3_height(rectangle3_heights[1045]), .rectangle3_weight(rectangle3_weights[1045]), .feature_threshold(feature_thresholds[1045]), .feature_above(feature_aboves[1045]), .feature_below(feature_belows[1045]), .scan_win_std_dev(scan_win_std_dev[1045]), .feature_accum(feature_accums[1045]));
  accum_calculator ac1046(.scan_win(scan_win1046), .rectangle1_x(rectangle1_xs[1046]), .rectangle1_y(rectangle1_ys[1046]), .rectangle1_width(rectangle1_widths[1046]), .rectangle1_height(rectangle1_heights[1046]), .rectangle1_weight(rectangle1_weights[1046]), .rectangle2_x(rectangle2_xs[1046]), .rectangle2_y(rectangle2_ys[1046]), .rectangle2_width(rectangle2_widths[1046]), .rectangle2_height(rectangle2_heights[1046]), .rectangle2_weight(rectangle2_weights[1046]), .rectangle3_x(rectangle3_xs[1046]), .rectangle3_y(rectangle3_ys[1046]), .rectangle3_width(rectangle3_widths[1046]), .rectangle3_height(rectangle3_heights[1046]), .rectangle3_weight(rectangle3_weights[1046]), .feature_threshold(feature_thresholds[1046]), .feature_above(feature_aboves[1046]), .feature_below(feature_belows[1046]), .scan_win_std_dev(scan_win_std_dev[1046]), .feature_accum(feature_accums[1046]));
  accum_calculator ac1047(.scan_win(scan_win1047), .rectangle1_x(rectangle1_xs[1047]), .rectangle1_y(rectangle1_ys[1047]), .rectangle1_width(rectangle1_widths[1047]), .rectangle1_height(rectangle1_heights[1047]), .rectangle1_weight(rectangle1_weights[1047]), .rectangle2_x(rectangle2_xs[1047]), .rectangle2_y(rectangle2_ys[1047]), .rectangle2_width(rectangle2_widths[1047]), .rectangle2_height(rectangle2_heights[1047]), .rectangle2_weight(rectangle2_weights[1047]), .rectangle3_x(rectangle3_xs[1047]), .rectangle3_y(rectangle3_ys[1047]), .rectangle3_width(rectangle3_widths[1047]), .rectangle3_height(rectangle3_heights[1047]), .rectangle3_weight(rectangle3_weights[1047]), .feature_threshold(feature_thresholds[1047]), .feature_above(feature_aboves[1047]), .feature_below(feature_belows[1047]), .scan_win_std_dev(scan_win_std_dev[1047]), .feature_accum(feature_accums[1047]));
  accum_calculator ac1048(.scan_win(scan_win1048), .rectangle1_x(rectangle1_xs[1048]), .rectangle1_y(rectangle1_ys[1048]), .rectangle1_width(rectangle1_widths[1048]), .rectangle1_height(rectangle1_heights[1048]), .rectangle1_weight(rectangle1_weights[1048]), .rectangle2_x(rectangle2_xs[1048]), .rectangle2_y(rectangle2_ys[1048]), .rectangle2_width(rectangle2_widths[1048]), .rectangle2_height(rectangle2_heights[1048]), .rectangle2_weight(rectangle2_weights[1048]), .rectangle3_x(rectangle3_xs[1048]), .rectangle3_y(rectangle3_ys[1048]), .rectangle3_width(rectangle3_widths[1048]), .rectangle3_height(rectangle3_heights[1048]), .rectangle3_weight(rectangle3_weights[1048]), .feature_threshold(feature_thresholds[1048]), .feature_above(feature_aboves[1048]), .feature_below(feature_belows[1048]), .scan_win_std_dev(scan_win_std_dev[1048]), .feature_accum(feature_accums[1048]));
  accum_calculator ac1049(.scan_win(scan_win1049), .rectangle1_x(rectangle1_xs[1049]), .rectangle1_y(rectangle1_ys[1049]), .rectangle1_width(rectangle1_widths[1049]), .rectangle1_height(rectangle1_heights[1049]), .rectangle1_weight(rectangle1_weights[1049]), .rectangle2_x(rectangle2_xs[1049]), .rectangle2_y(rectangle2_ys[1049]), .rectangle2_width(rectangle2_widths[1049]), .rectangle2_height(rectangle2_heights[1049]), .rectangle2_weight(rectangle2_weights[1049]), .rectangle3_x(rectangle3_xs[1049]), .rectangle3_y(rectangle3_ys[1049]), .rectangle3_width(rectangle3_widths[1049]), .rectangle3_height(rectangle3_heights[1049]), .rectangle3_weight(rectangle3_weights[1049]), .feature_threshold(feature_thresholds[1049]), .feature_above(feature_aboves[1049]), .feature_below(feature_belows[1049]), .scan_win_std_dev(scan_win_std_dev[1049]), .feature_accum(feature_accums[1049]));
  accum_calculator ac1050(.scan_win(scan_win1050), .rectangle1_x(rectangle1_xs[1050]), .rectangle1_y(rectangle1_ys[1050]), .rectangle1_width(rectangle1_widths[1050]), .rectangle1_height(rectangle1_heights[1050]), .rectangle1_weight(rectangle1_weights[1050]), .rectangle2_x(rectangle2_xs[1050]), .rectangle2_y(rectangle2_ys[1050]), .rectangle2_width(rectangle2_widths[1050]), .rectangle2_height(rectangle2_heights[1050]), .rectangle2_weight(rectangle2_weights[1050]), .rectangle3_x(rectangle3_xs[1050]), .rectangle3_y(rectangle3_ys[1050]), .rectangle3_width(rectangle3_widths[1050]), .rectangle3_height(rectangle3_heights[1050]), .rectangle3_weight(rectangle3_weights[1050]), .feature_threshold(feature_thresholds[1050]), .feature_above(feature_aboves[1050]), .feature_below(feature_belows[1050]), .scan_win_std_dev(scan_win_std_dev[1050]), .feature_accum(feature_accums[1050]));
  accum_calculator ac1051(.scan_win(scan_win1051), .rectangle1_x(rectangle1_xs[1051]), .rectangle1_y(rectangle1_ys[1051]), .rectangle1_width(rectangle1_widths[1051]), .rectangle1_height(rectangle1_heights[1051]), .rectangle1_weight(rectangle1_weights[1051]), .rectangle2_x(rectangle2_xs[1051]), .rectangle2_y(rectangle2_ys[1051]), .rectangle2_width(rectangle2_widths[1051]), .rectangle2_height(rectangle2_heights[1051]), .rectangle2_weight(rectangle2_weights[1051]), .rectangle3_x(rectangle3_xs[1051]), .rectangle3_y(rectangle3_ys[1051]), .rectangle3_width(rectangle3_widths[1051]), .rectangle3_height(rectangle3_heights[1051]), .rectangle3_weight(rectangle3_weights[1051]), .feature_threshold(feature_thresholds[1051]), .feature_above(feature_aboves[1051]), .feature_below(feature_belows[1051]), .scan_win_std_dev(scan_win_std_dev[1051]), .feature_accum(feature_accums[1051]));
  accum_calculator ac1052(.scan_win(scan_win1052), .rectangle1_x(rectangle1_xs[1052]), .rectangle1_y(rectangle1_ys[1052]), .rectangle1_width(rectangle1_widths[1052]), .rectangle1_height(rectangle1_heights[1052]), .rectangle1_weight(rectangle1_weights[1052]), .rectangle2_x(rectangle2_xs[1052]), .rectangle2_y(rectangle2_ys[1052]), .rectangle2_width(rectangle2_widths[1052]), .rectangle2_height(rectangle2_heights[1052]), .rectangle2_weight(rectangle2_weights[1052]), .rectangle3_x(rectangle3_xs[1052]), .rectangle3_y(rectangle3_ys[1052]), .rectangle3_width(rectangle3_widths[1052]), .rectangle3_height(rectangle3_heights[1052]), .rectangle3_weight(rectangle3_weights[1052]), .feature_threshold(feature_thresholds[1052]), .feature_above(feature_aboves[1052]), .feature_below(feature_belows[1052]), .scan_win_std_dev(scan_win_std_dev[1052]), .feature_accum(feature_accums[1052]));
  accum_calculator ac1053(.scan_win(scan_win1053), .rectangle1_x(rectangle1_xs[1053]), .rectangle1_y(rectangle1_ys[1053]), .rectangle1_width(rectangle1_widths[1053]), .rectangle1_height(rectangle1_heights[1053]), .rectangle1_weight(rectangle1_weights[1053]), .rectangle2_x(rectangle2_xs[1053]), .rectangle2_y(rectangle2_ys[1053]), .rectangle2_width(rectangle2_widths[1053]), .rectangle2_height(rectangle2_heights[1053]), .rectangle2_weight(rectangle2_weights[1053]), .rectangle3_x(rectangle3_xs[1053]), .rectangle3_y(rectangle3_ys[1053]), .rectangle3_width(rectangle3_widths[1053]), .rectangle3_height(rectangle3_heights[1053]), .rectangle3_weight(rectangle3_weights[1053]), .feature_threshold(feature_thresholds[1053]), .feature_above(feature_aboves[1053]), .feature_below(feature_belows[1053]), .scan_win_std_dev(scan_win_std_dev[1053]), .feature_accum(feature_accums[1053]));
  accum_calculator ac1054(.scan_win(scan_win1054), .rectangle1_x(rectangle1_xs[1054]), .rectangle1_y(rectangle1_ys[1054]), .rectangle1_width(rectangle1_widths[1054]), .rectangle1_height(rectangle1_heights[1054]), .rectangle1_weight(rectangle1_weights[1054]), .rectangle2_x(rectangle2_xs[1054]), .rectangle2_y(rectangle2_ys[1054]), .rectangle2_width(rectangle2_widths[1054]), .rectangle2_height(rectangle2_heights[1054]), .rectangle2_weight(rectangle2_weights[1054]), .rectangle3_x(rectangle3_xs[1054]), .rectangle3_y(rectangle3_ys[1054]), .rectangle3_width(rectangle3_widths[1054]), .rectangle3_height(rectangle3_heights[1054]), .rectangle3_weight(rectangle3_weights[1054]), .feature_threshold(feature_thresholds[1054]), .feature_above(feature_aboves[1054]), .feature_below(feature_belows[1054]), .scan_win_std_dev(scan_win_std_dev[1054]), .feature_accum(feature_accums[1054]));
  accum_calculator ac1055(.scan_win(scan_win1055), .rectangle1_x(rectangle1_xs[1055]), .rectangle1_y(rectangle1_ys[1055]), .rectangle1_width(rectangle1_widths[1055]), .rectangle1_height(rectangle1_heights[1055]), .rectangle1_weight(rectangle1_weights[1055]), .rectangle2_x(rectangle2_xs[1055]), .rectangle2_y(rectangle2_ys[1055]), .rectangle2_width(rectangle2_widths[1055]), .rectangle2_height(rectangle2_heights[1055]), .rectangle2_weight(rectangle2_weights[1055]), .rectangle3_x(rectangle3_xs[1055]), .rectangle3_y(rectangle3_ys[1055]), .rectangle3_width(rectangle3_widths[1055]), .rectangle3_height(rectangle3_heights[1055]), .rectangle3_weight(rectangle3_weights[1055]), .feature_threshold(feature_thresholds[1055]), .feature_above(feature_aboves[1055]), .feature_below(feature_belows[1055]), .scan_win_std_dev(scan_win_std_dev[1055]), .feature_accum(feature_accums[1055]));
  accum_calculator ac1056(.scan_win(scan_win1056), .rectangle1_x(rectangle1_xs[1056]), .rectangle1_y(rectangle1_ys[1056]), .rectangle1_width(rectangle1_widths[1056]), .rectangle1_height(rectangle1_heights[1056]), .rectangle1_weight(rectangle1_weights[1056]), .rectangle2_x(rectangle2_xs[1056]), .rectangle2_y(rectangle2_ys[1056]), .rectangle2_width(rectangle2_widths[1056]), .rectangle2_height(rectangle2_heights[1056]), .rectangle2_weight(rectangle2_weights[1056]), .rectangle3_x(rectangle3_xs[1056]), .rectangle3_y(rectangle3_ys[1056]), .rectangle3_width(rectangle3_widths[1056]), .rectangle3_height(rectangle3_heights[1056]), .rectangle3_weight(rectangle3_weights[1056]), .feature_threshold(feature_thresholds[1056]), .feature_above(feature_aboves[1056]), .feature_below(feature_belows[1056]), .scan_win_std_dev(scan_win_std_dev[1056]), .feature_accum(feature_accums[1056]));
  accum_calculator ac1057(.scan_win(scan_win1057), .rectangle1_x(rectangle1_xs[1057]), .rectangle1_y(rectangle1_ys[1057]), .rectangle1_width(rectangle1_widths[1057]), .rectangle1_height(rectangle1_heights[1057]), .rectangle1_weight(rectangle1_weights[1057]), .rectangle2_x(rectangle2_xs[1057]), .rectangle2_y(rectangle2_ys[1057]), .rectangle2_width(rectangle2_widths[1057]), .rectangle2_height(rectangle2_heights[1057]), .rectangle2_weight(rectangle2_weights[1057]), .rectangle3_x(rectangle3_xs[1057]), .rectangle3_y(rectangle3_ys[1057]), .rectangle3_width(rectangle3_widths[1057]), .rectangle3_height(rectangle3_heights[1057]), .rectangle3_weight(rectangle3_weights[1057]), .feature_threshold(feature_thresholds[1057]), .feature_above(feature_aboves[1057]), .feature_below(feature_belows[1057]), .scan_win_std_dev(scan_win_std_dev[1057]), .feature_accum(feature_accums[1057]));
  accum_calculator ac1058(.scan_win(scan_win1058), .rectangle1_x(rectangle1_xs[1058]), .rectangle1_y(rectangle1_ys[1058]), .rectangle1_width(rectangle1_widths[1058]), .rectangle1_height(rectangle1_heights[1058]), .rectangle1_weight(rectangle1_weights[1058]), .rectangle2_x(rectangle2_xs[1058]), .rectangle2_y(rectangle2_ys[1058]), .rectangle2_width(rectangle2_widths[1058]), .rectangle2_height(rectangle2_heights[1058]), .rectangle2_weight(rectangle2_weights[1058]), .rectangle3_x(rectangle3_xs[1058]), .rectangle3_y(rectangle3_ys[1058]), .rectangle3_width(rectangle3_widths[1058]), .rectangle3_height(rectangle3_heights[1058]), .rectangle3_weight(rectangle3_weights[1058]), .feature_threshold(feature_thresholds[1058]), .feature_above(feature_aboves[1058]), .feature_below(feature_belows[1058]), .scan_win_std_dev(scan_win_std_dev[1058]), .feature_accum(feature_accums[1058]));
  accum_calculator ac1059(.scan_win(scan_win1059), .rectangle1_x(rectangle1_xs[1059]), .rectangle1_y(rectangle1_ys[1059]), .rectangle1_width(rectangle1_widths[1059]), .rectangle1_height(rectangle1_heights[1059]), .rectangle1_weight(rectangle1_weights[1059]), .rectangle2_x(rectangle2_xs[1059]), .rectangle2_y(rectangle2_ys[1059]), .rectangle2_width(rectangle2_widths[1059]), .rectangle2_height(rectangle2_heights[1059]), .rectangle2_weight(rectangle2_weights[1059]), .rectangle3_x(rectangle3_xs[1059]), .rectangle3_y(rectangle3_ys[1059]), .rectangle3_width(rectangle3_widths[1059]), .rectangle3_height(rectangle3_heights[1059]), .rectangle3_weight(rectangle3_weights[1059]), .feature_threshold(feature_thresholds[1059]), .feature_above(feature_aboves[1059]), .feature_below(feature_belows[1059]), .scan_win_std_dev(scan_win_std_dev[1059]), .feature_accum(feature_accums[1059]));
  accum_calculator ac1060(.scan_win(scan_win1060), .rectangle1_x(rectangle1_xs[1060]), .rectangle1_y(rectangle1_ys[1060]), .rectangle1_width(rectangle1_widths[1060]), .rectangle1_height(rectangle1_heights[1060]), .rectangle1_weight(rectangle1_weights[1060]), .rectangle2_x(rectangle2_xs[1060]), .rectangle2_y(rectangle2_ys[1060]), .rectangle2_width(rectangle2_widths[1060]), .rectangle2_height(rectangle2_heights[1060]), .rectangle2_weight(rectangle2_weights[1060]), .rectangle3_x(rectangle3_xs[1060]), .rectangle3_y(rectangle3_ys[1060]), .rectangle3_width(rectangle3_widths[1060]), .rectangle3_height(rectangle3_heights[1060]), .rectangle3_weight(rectangle3_weights[1060]), .feature_threshold(feature_thresholds[1060]), .feature_above(feature_aboves[1060]), .feature_below(feature_belows[1060]), .scan_win_std_dev(scan_win_std_dev[1060]), .feature_accum(feature_accums[1060]));
  accum_calculator ac1061(.scan_win(scan_win1061), .rectangle1_x(rectangle1_xs[1061]), .rectangle1_y(rectangle1_ys[1061]), .rectangle1_width(rectangle1_widths[1061]), .rectangle1_height(rectangle1_heights[1061]), .rectangle1_weight(rectangle1_weights[1061]), .rectangle2_x(rectangle2_xs[1061]), .rectangle2_y(rectangle2_ys[1061]), .rectangle2_width(rectangle2_widths[1061]), .rectangle2_height(rectangle2_heights[1061]), .rectangle2_weight(rectangle2_weights[1061]), .rectangle3_x(rectangle3_xs[1061]), .rectangle3_y(rectangle3_ys[1061]), .rectangle3_width(rectangle3_widths[1061]), .rectangle3_height(rectangle3_heights[1061]), .rectangle3_weight(rectangle3_weights[1061]), .feature_threshold(feature_thresholds[1061]), .feature_above(feature_aboves[1061]), .feature_below(feature_belows[1061]), .scan_win_std_dev(scan_win_std_dev[1061]), .feature_accum(feature_accums[1061]));
  accum_calculator ac1062(.scan_win(scan_win1062), .rectangle1_x(rectangle1_xs[1062]), .rectangle1_y(rectangle1_ys[1062]), .rectangle1_width(rectangle1_widths[1062]), .rectangle1_height(rectangle1_heights[1062]), .rectangle1_weight(rectangle1_weights[1062]), .rectangle2_x(rectangle2_xs[1062]), .rectangle2_y(rectangle2_ys[1062]), .rectangle2_width(rectangle2_widths[1062]), .rectangle2_height(rectangle2_heights[1062]), .rectangle2_weight(rectangle2_weights[1062]), .rectangle3_x(rectangle3_xs[1062]), .rectangle3_y(rectangle3_ys[1062]), .rectangle3_width(rectangle3_widths[1062]), .rectangle3_height(rectangle3_heights[1062]), .rectangle3_weight(rectangle3_weights[1062]), .feature_threshold(feature_thresholds[1062]), .feature_above(feature_aboves[1062]), .feature_below(feature_belows[1062]), .scan_win_std_dev(scan_win_std_dev[1062]), .feature_accum(feature_accums[1062]));
  accum_calculator ac1063(.scan_win(scan_win1063), .rectangle1_x(rectangle1_xs[1063]), .rectangle1_y(rectangle1_ys[1063]), .rectangle1_width(rectangle1_widths[1063]), .rectangle1_height(rectangle1_heights[1063]), .rectangle1_weight(rectangle1_weights[1063]), .rectangle2_x(rectangle2_xs[1063]), .rectangle2_y(rectangle2_ys[1063]), .rectangle2_width(rectangle2_widths[1063]), .rectangle2_height(rectangle2_heights[1063]), .rectangle2_weight(rectangle2_weights[1063]), .rectangle3_x(rectangle3_xs[1063]), .rectangle3_y(rectangle3_ys[1063]), .rectangle3_width(rectangle3_widths[1063]), .rectangle3_height(rectangle3_heights[1063]), .rectangle3_weight(rectangle3_weights[1063]), .feature_threshold(feature_thresholds[1063]), .feature_above(feature_aboves[1063]), .feature_below(feature_belows[1063]), .scan_win_std_dev(scan_win_std_dev[1063]), .feature_accum(feature_accums[1063]));
  accum_calculator ac1064(.scan_win(scan_win1064), .rectangle1_x(rectangle1_xs[1064]), .rectangle1_y(rectangle1_ys[1064]), .rectangle1_width(rectangle1_widths[1064]), .rectangle1_height(rectangle1_heights[1064]), .rectangle1_weight(rectangle1_weights[1064]), .rectangle2_x(rectangle2_xs[1064]), .rectangle2_y(rectangle2_ys[1064]), .rectangle2_width(rectangle2_widths[1064]), .rectangle2_height(rectangle2_heights[1064]), .rectangle2_weight(rectangle2_weights[1064]), .rectangle3_x(rectangle3_xs[1064]), .rectangle3_y(rectangle3_ys[1064]), .rectangle3_width(rectangle3_widths[1064]), .rectangle3_height(rectangle3_heights[1064]), .rectangle3_weight(rectangle3_weights[1064]), .feature_threshold(feature_thresholds[1064]), .feature_above(feature_aboves[1064]), .feature_below(feature_belows[1064]), .scan_win_std_dev(scan_win_std_dev[1064]), .feature_accum(feature_accums[1064]));
  accum_calculator ac1065(.scan_win(scan_win1065), .rectangle1_x(rectangle1_xs[1065]), .rectangle1_y(rectangle1_ys[1065]), .rectangle1_width(rectangle1_widths[1065]), .rectangle1_height(rectangle1_heights[1065]), .rectangle1_weight(rectangle1_weights[1065]), .rectangle2_x(rectangle2_xs[1065]), .rectangle2_y(rectangle2_ys[1065]), .rectangle2_width(rectangle2_widths[1065]), .rectangle2_height(rectangle2_heights[1065]), .rectangle2_weight(rectangle2_weights[1065]), .rectangle3_x(rectangle3_xs[1065]), .rectangle3_y(rectangle3_ys[1065]), .rectangle3_width(rectangle3_widths[1065]), .rectangle3_height(rectangle3_heights[1065]), .rectangle3_weight(rectangle3_weights[1065]), .feature_threshold(feature_thresholds[1065]), .feature_above(feature_aboves[1065]), .feature_below(feature_belows[1065]), .scan_win_std_dev(scan_win_std_dev[1065]), .feature_accum(feature_accums[1065]));
  accum_calculator ac1066(.scan_win(scan_win1066), .rectangle1_x(rectangle1_xs[1066]), .rectangle1_y(rectangle1_ys[1066]), .rectangle1_width(rectangle1_widths[1066]), .rectangle1_height(rectangle1_heights[1066]), .rectangle1_weight(rectangle1_weights[1066]), .rectangle2_x(rectangle2_xs[1066]), .rectangle2_y(rectangle2_ys[1066]), .rectangle2_width(rectangle2_widths[1066]), .rectangle2_height(rectangle2_heights[1066]), .rectangle2_weight(rectangle2_weights[1066]), .rectangle3_x(rectangle3_xs[1066]), .rectangle3_y(rectangle3_ys[1066]), .rectangle3_width(rectangle3_widths[1066]), .rectangle3_height(rectangle3_heights[1066]), .rectangle3_weight(rectangle3_weights[1066]), .feature_threshold(feature_thresholds[1066]), .feature_above(feature_aboves[1066]), .feature_below(feature_belows[1066]), .scan_win_std_dev(scan_win_std_dev[1066]), .feature_accum(feature_accums[1066]));
  accum_calculator ac1067(.scan_win(scan_win1067), .rectangle1_x(rectangle1_xs[1067]), .rectangle1_y(rectangle1_ys[1067]), .rectangle1_width(rectangle1_widths[1067]), .rectangle1_height(rectangle1_heights[1067]), .rectangle1_weight(rectangle1_weights[1067]), .rectangle2_x(rectangle2_xs[1067]), .rectangle2_y(rectangle2_ys[1067]), .rectangle2_width(rectangle2_widths[1067]), .rectangle2_height(rectangle2_heights[1067]), .rectangle2_weight(rectangle2_weights[1067]), .rectangle3_x(rectangle3_xs[1067]), .rectangle3_y(rectangle3_ys[1067]), .rectangle3_width(rectangle3_widths[1067]), .rectangle3_height(rectangle3_heights[1067]), .rectangle3_weight(rectangle3_weights[1067]), .feature_threshold(feature_thresholds[1067]), .feature_above(feature_aboves[1067]), .feature_below(feature_belows[1067]), .scan_win_std_dev(scan_win_std_dev[1067]), .feature_accum(feature_accums[1067]));
  accum_calculator ac1068(.scan_win(scan_win1068), .rectangle1_x(rectangle1_xs[1068]), .rectangle1_y(rectangle1_ys[1068]), .rectangle1_width(rectangle1_widths[1068]), .rectangle1_height(rectangle1_heights[1068]), .rectangle1_weight(rectangle1_weights[1068]), .rectangle2_x(rectangle2_xs[1068]), .rectangle2_y(rectangle2_ys[1068]), .rectangle2_width(rectangle2_widths[1068]), .rectangle2_height(rectangle2_heights[1068]), .rectangle2_weight(rectangle2_weights[1068]), .rectangle3_x(rectangle3_xs[1068]), .rectangle3_y(rectangle3_ys[1068]), .rectangle3_width(rectangle3_widths[1068]), .rectangle3_height(rectangle3_heights[1068]), .rectangle3_weight(rectangle3_weights[1068]), .feature_threshold(feature_thresholds[1068]), .feature_above(feature_aboves[1068]), .feature_below(feature_belows[1068]), .scan_win_std_dev(scan_win_std_dev[1068]), .feature_accum(feature_accums[1068]));
  accum_calculator ac1069(.scan_win(scan_win1069), .rectangle1_x(rectangle1_xs[1069]), .rectangle1_y(rectangle1_ys[1069]), .rectangle1_width(rectangle1_widths[1069]), .rectangle1_height(rectangle1_heights[1069]), .rectangle1_weight(rectangle1_weights[1069]), .rectangle2_x(rectangle2_xs[1069]), .rectangle2_y(rectangle2_ys[1069]), .rectangle2_width(rectangle2_widths[1069]), .rectangle2_height(rectangle2_heights[1069]), .rectangle2_weight(rectangle2_weights[1069]), .rectangle3_x(rectangle3_xs[1069]), .rectangle3_y(rectangle3_ys[1069]), .rectangle3_width(rectangle3_widths[1069]), .rectangle3_height(rectangle3_heights[1069]), .rectangle3_weight(rectangle3_weights[1069]), .feature_threshold(feature_thresholds[1069]), .feature_above(feature_aboves[1069]), .feature_below(feature_belows[1069]), .scan_win_std_dev(scan_win_std_dev[1069]), .feature_accum(feature_accums[1069]));
  accum_calculator ac1070(.scan_win(scan_win1070), .rectangle1_x(rectangle1_xs[1070]), .rectangle1_y(rectangle1_ys[1070]), .rectangle1_width(rectangle1_widths[1070]), .rectangle1_height(rectangle1_heights[1070]), .rectangle1_weight(rectangle1_weights[1070]), .rectangle2_x(rectangle2_xs[1070]), .rectangle2_y(rectangle2_ys[1070]), .rectangle2_width(rectangle2_widths[1070]), .rectangle2_height(rectangle2_heights[1070]), .rectangle2_weight(rectangle2_weights[1070]), .rectangle3_x(rectangle3_xs[1070]), .rectangle3_y(rectangle3_ys[1070]), .rectangle3_width(rectangle3_widths[1070]), .rectangle3_height(rectangle3_heights[1070]), .rectangle3_weight(rectangle3_weights[1070]), .feature_threshold(feature_thresholds[1070]), .feature_above(feature_aboves[1070]), .feature_below(feature_belows[1070]), .scan_win_std_dev(scan_win_std_dev[1070]), .feature_accum(feature_accums[1070]));
  accum_calculator ac1071(.scan_win(scan_win1071), .rectangle1_x(rectangle1_xs[1071]), .rectangle1_y(rectangle1_ys[1071]), .rectangle1_width(rectangle1_widths[1071]), .rectangle1_height(rectangle1_heights[1071]), .rectangle1_weight(rectangle1_weights[1071]), .rectangle2_x(rectangle2_xs[1071]), .rectangle2_y(rectangle2_ys[1071]), .rectangle2_width(rectangle2_widths[1071]), .rectangle2_height(rectangle2_heights[1071]), .rectangle2_weight(rectangle2_weights[1071]), .rectangle3_x(rectangle3_xs[1071]), .rectangle3_y(rectangle3_ys[1071]), .rectangle3_width(rectangle3_widths[1071]), .rectangle3_height(rectangle3_heights[1071]), .rectangle3_weight(rectangle3_weights[1071]), .feature_threshold(feature_thresholds[1071]), .feature_above(feature_aboves[1071]), .feature_below(feature_belows[1071]), .scan_win_std_dev(scan_win_std_dev[1071]), .feature_accum(feature_accums[1071]));
  accum_calculator ac1072(.scan_win(scan_win1072), .rectangle1_x(rectangle1_xs[1072]), .rectangle1_y(rectangle1_ys[1072]), .rectangle1_width(rectangle1_widths[1072]), .rectangle1_height(rectangle1_heights[1072]), .rectangle1_weight(rectangle1_weights[1072]), .rectangle2_x(rectangle2_xs[1072]), .rectangle2_y(rectangle2_ys[1072]), .rectangle2_width(rectangle2_widths[1072]), .rectangle2_height(rectangle2_heights[1072]), .rectangle2_weight(rectangle2_weights[1072]), .rectangle3_x(rectangle3_xs[1072]), .rectangle3_y(rectangle3_ys[1072]), .rectangle3_width(rectangle3_widths[1072]), .rectangle3_height(rectangle3_heights[1072]), .rectangle3_weight(rectangle3_weights[1072]), .feature_threshold(feature_thresholds[1072]), .feature_above(feature_aboves[1072]), .feature_below(feature_belows[1072]), .scan_win_std_dev(scan_win_std_dev[1072]), .feature_accum(feature_accums[1072]));
  accum_calculator ac1073(.scan_win(scan_win1073), .rectangle1_x(rectangle1_xs[1073]), .rectangle1_y(rectangle1_ys[1073]), .rectangle1_width(rectangle1_widths[1073]), .rectangle1_height(rectangle1_heights[1073]), .rectangle1_weight(rectangle1_weights[1073]), .rectangle2_x(rectangle2_xs[1073]), .rectangle2_y(rectangle2_ys[1073]), .rectangle2_width(rectangle2_widths[1073]), .rectangle2_height(rectangle2_heights[1073]), .rectangle2_weight(rectangle2_weights[1073]), .rectangle3_x(rectangle3_xs[1073]), .rectangle3_y(rectangle3_ys[1073]), .rectangle3_width(rectangle3_widths[1073]), .rectangle3_height(rectangle3_heights[1073]), .rectangle3_weight(rectangle3_weights[1073]), .feature_threshold(feature_thresholds[1073]), .feature_above(feature_aboves[1073]), .feature_below(feature_belows[1073]), .scan_win_std_dev(scan_win_std_dev[1073]), .feature_accum(feature_accums[1073]));
  accum_calculator ac1074(.scan_win(scan_win1074), .rectangle1_x(rectangle1_xs[1074]), .rectangle1_y(rectangle1_ys[1074]), .rectangle1_width(rectangle1_widths[1074]), .rectangle1_height(rectangle1_heights[1074]), .rectangle1_weight(rectangle1_weights[1074]), .rectangle2_x(rectangle2_xs[1074]), .rectangle2_y(rectangle2_ys[1074]), .rectangle2_width(rectangle2_widths[1074]), .rectangle2_height(rectangle2_heights[1074]), .rectangle2_weight(rectangle2_weights[1074]), .rectangle3_x(rectangle3_xs[1074]), .rectangle3_y(rectangle3_ys[1074]), .rectangle3_width(rectangle3_widths[1074]), .rectangle3_height(rectangle3_heights[1074]), .rectangle3_weight(rectangle3_weights[1074]), .feature_threshold(feature_thresholds[1074]), .feature_above(feature_aboves[1074]), .feature_below(feature_belows[1074]), .scan_win_std_dev(scan_win_std_dev[1074]), .feature_accum(feature_accums[1074]));
  accum_calculator ac1075(.scan_win(scan_win1075), .rectangle1_x(rectangle1_xs[1075]), .rectangle1_y(rectangle1_ys[1075]), .rectangle1_width(rectangle1_widths[1075]), .rectangle1_height(rectangle1_heights[1075]), .rectangle1_weight(rectangle1_weights[1075]), .rectangle2_x(rectangle2_xs[1075]), .rectangle2_y(rectangle2_ys[1075]), .rectangle2_width(rectangle2_widths[1075]), .rectangle2_height(rectangle2_heights[1075]), .rectangle2_weight(rectangle2_weights[1075]), .rectangle3_x(rectangle3_xs[1075]), .rectangle3_y(rectangle3_ys[1075]), .rectangle3_width(rectangle3_widths[1075]), .rectangle3_height(rectangle3_heights[1075]), .rectangle3_weight(rectangle3_weights[1075]), .feature_threshold(feature_thresholds[1075]), .feature_above(feature_aboves[1075]), .feature_below(feature_belows[1075]), .scan_win_std_dev(scan_win_std_dev[1075]), .feature_accum(feature_accums[1075]));
  accum_calculator ac1076(.scan_win(scan_win1076), .rectangle1_x(rectangle1_xs[1076]), .rectangle1_y(rectangle1_ys[1076]), .rectangle1_width(rectangle1_widths[1076]), .rectangle1_height(rectangle1_heights[1076]), .rectangle1_weight(rectangle1_weights[1076]), .rectangle2_x(rectangle2_xs[1076]), .rectangle2_y(rectangle2_ys[1076]), .rectangle2_width(rectangle2_widths[1076]), .rectangle2_height(rectangle2_heights[1076]), .rectangle2_weight(rectangle2_weights[1076]), .rectangle3_x(rectangle3_xs[1076]), .rectangle3_y(rectangle3_ys[1076]), .rectangle3_width(rectangle3_widths[1076]), .rectangle3_height(rectangle3_heights[1076]), .rectangle3_weight(rectangle3_weights[1076]), .feature_threshold(feature_thresholds[1076]), .feature_above(feature_aboves[1076]), .feature_below(feature_belows[1076]), .scan_win_std_dev(scan_win_std_dev[1076]), .feature_accum(feature_accums[1076]));
  accum_calculator ac1077(.scan_win(scan_win1077), .rectangle1_x(rectangle1_xs[1077]), .rectangle1_y(rectangle1_ys[1077]), .rectangle1_width(rectangle1_widths[1077]), .rectangle1_height(rectangle1_heights[1077]), .rectangle1_weight(rectangle1_weights[1077]), .rectangle2_x(rectangle2_xs[1077]), .rectangle2_y(rectangle2_ys[1077]), .rectangle2_width(rectangle2_widths[1077]), .rectangle2_height(rectangle2_heights[1077]), .rectangle2_weight(rectangle2_weights[1077]), .rectangle3_x(rectangle3_xs[1077]), .rectangle3_y(rectangle3_ys[1077]), .rectangle3_width(rectangle3_widths[1077]), .rectangle3_height(rectangle3_heights[1077]), .rectangle3_weight(rectangle3_weights[1077]), .feature_threshold(feature_thresholds[1077]), .feature_above(feature_aboves[1077]), .feature_below(feature_belows[1077]), .scan_win_std_dev(scan_win_std_dev[1077]), .feature_accum(feature_accums[1077]));
  accum_calculator ac1078(.scan_win(scan_win1078), .rectangle1_x(rectangle1_xs[1078]), .rectangle1_y(rectangle1_ys[1078]), .rectangle1_width(rectangle1_widths[1078]), .rectangle1_height(rectangle1_heights[1078]), .rectangle1_weight(rectangle1_weights[1078]), .rectangle2_x(rectangle2_xs[1078]), .rectangle2_y(rectangle2_ys[1078]), .rectangle2_width(rectangle2_widths[1078]), .rectangle2_height(rectangle2_heights[1078]), .rectangle2_weight(rectangle2_weights[1078]), .rectangle3_x(rectangle3_xs[1078]), .rectangle3_y(rectangle3_ys[1078]), .rectangle3_width(rectangle3_widths[1078]), .rectangle3_height(rectangle3_heights[1078]), .rectangle3_weight(rectangle3_weights[1078]), .feature_threshold(feature_thresholds[1078]), .feature_above(feature_aboves[1078]), .feature_below(feature_belows[1078]), .scan_win_std_dev(scan_win_std_dev[1078]), .feature_accum(feature_accums[1078]));
  accum_calculator ac1079(.scan_win(scan_win1079), .rectangle1_x(rectangle1_xs[1079]), .rectangle1_y(rectangle1_ys[1079]), .rectangle1_width(rectangle1_widths[1079]), .rectangle1_height(rectangle1_heights[1079]), .rectangle1_weight(rectangle1_weights[1079]), .rectangle2_x(rectangle2_xs[1079]), .rectangle2_y(rectangle2_ys[1079]), .rectangle2_width(rectangle2_widths[1079]), .rectangle2_height(rectangle2_heights[1079]), .rectangle2_weight(rectangle2_weights[1079]), .rectangle3_x(rectangle3_xs[1079]), .rectangle3_y(rectangle3_ys[1079]), .rectangle3_width(rectangle3_widths[1079]), .rectangle3_height(rectangle3_heights[1079]), .rectangle3_weight(rectangle3_weights[1079]), .feature_threshold(feature_thresholds[1079]), .feature_above(feature_aboves[1079]), .feature_below(feature_belows[1079]), .scan_win_std_dev(scan_win_std_dev[1079]), .feature_accum(feature_accums[1079]));
  accum_calculator ac1080(.scan_win(scan_win1080), .rectangle1_x(rectangle1_xs[1080]), .rectangle1_y(rectangle1_ys[1080]), .rectangle1_width(rectangle1_widths[1080]), .rectangle1_height(rectangle1_heights[1080]), .rectangle1_weight(rectangle1_weights[1080]), .rectangle2_x(rectangle2_xs[1080]), .rectangle2_y(rectangle2_ys[1080]), .rectangle2_width(rectangle2_widths[1080]), .rectangle2_height(rectangle2_heights[1080]), .rectangle2_weight(rectangle2_weights[1080]), .rectangle3_x(rectangle3_xs[1080]), .rectangle3_y(rectangle3_ys[1080]), .rectangle3_width(rectangle3_widths[1080]), .rectangle3_height(rectangle3_heights[1080]), .rectangle3_weight(rectangle3_weights[1080]), .feature_threshold(feature_thresholds[1080]), .feature_above(feature_aboves[1080]), .feature_below(feature_belows[1080]), .scan_win_std_dev(scan_win_std_dev[1080]), .feature_accum(feature_accums[1080]));
  accum_calculator ac1081(.scan_win(scan_win1081), .rectangle1_x(rectangle1_xs[1081]), .rectangle1_y(rectangle1_ys[1081]), .rectangle1_width(rectangle1_widths[1081]), .rectangle1_height(rectangle1_heights[1081]), .rectangle1_weight(rectangle1_weights[1081]), .rectangle2_x(rectangle2_xs[1081]), .rectangle2_y(rectangle2_ys[1081]), .rectangle2_width(rectangle2_widths[1081]), .rectangle2_height(rectangle2_heights[1081]), .rectangle2_weight(rectangle2_weights[1081]), .rectangle3_x(rectangle3_xs[1081]), .rectangle3_y(rectangle3_ys[1081]), .rectangle3_width(rectangle3_widths[1081]), .rectangle3_height(rectangle3_heights[1081]), .rectangle3_weight(rectangle3_weights[1081]), .feature_threshold(feature_thresholds[1081]), .feature_above(feature_aboves[1081]), .feature_below(feature_belows[1081]), .scan_win_std_dev(scan_win_std_dev[1081]), .feature_accum(feature_accums[1081]));
  accum_calculator ac1082(.scan_win(scan_win1082), .rectangle1_x(rectangle1_xs[1082]), .rectangle1_y(rectangle1_ys[1082]), .rectangle1_width(rectangle1_widths[1082]), .rectangle1_height(rectangle1_heights[1082]), .rectangle1_weight(rectangle1_weights[1082]), .rectangle2_x(rectangle2_xs[1082]), .rectangle2_y(rectangle2_ys[1082]), .rectangle2_width(rectangle2_widths[1082]), .rectangle2_height(rectangle2_heights[1082]), .rectangle2_weight(rectangle2_weights[1082]), .rectangle3_x(rectangle3_xs[1082]), .rectangle3_y(rectangle3_ys[1082]), .rectangle3_width(rectangle3_widths[1082]), .rectangle3_height(rectangle3_heights[1082]), .rectangle3_weight(rectangle3_weights[1082]), .feature_threshold(feature_thresholds[1082]), .feature_above(feature_aboves[1082]), .feature_below(feature_belows[1082]), .scan_win_std_dev(scan_win_std_dev[1082]), .feature_accum(feature_accums[1082]));
  accum_calculator ac1083(.scan_win(scan_win1083), .rectangle1_x(rectangle1_xs[1083]), .rectangle1_y(rectangle1_ys[1083]), .rectangle1_width(rectangle1_widths[1083]), .rectangle1_height(rectangle1_heights[1083]), .rectangle1_weight(rectangle1_weights[1083]), .rectangle2_x(rectangle2_xs[1083]), .rectangle2_y(rectangle2_ys[1083]), .rectangle2_width(rectangle2_widths[1083]), .rectangle2_height(rectangle2_heights[1083]), .rectangle2_weight(rectangle2_weights[1083]), .rectangle3_x(rectangle3_xs[1083]), .rectangle3_y(rectangle3_ys[1083]), .rectangle3_width(rectangle3_widths[1083]), .rectangle3_height(rectangle3_heights[1083]), .rectangle3_weight(rectangle3_weights[1083]), .feature_threshold(feature_thresholds[1083]), .feature_above(feature_aboves[1083]), .feature_below(feature_belows[1083]), .scan_win_std_dev(scan_win_std_dev[1083]), .feature_accum(feature_accums[1083]));
  accum_calculator ac1084(.scan_win(scan_win1084), .rectangle1_x(rectangle1_xs[1084]), .rectangle1_y(rectangle1_ys[1084]), .rectangle1_width(rectangle1_widths[1084]), .rectangle1_height(rectangle1_heights[1084]), .rectangle1_weight(rectangle1_weights[1084]), .rectangle2_x(rectangle2_xs[1084]), .rectangle2_y(rectangle2_ys[1084]), .rectangle2_width(rectangle2_widths[1084]), .rectangle2_height(rectangle2_heights[1084]), .rectangle2_weight(rectangle2_weights[1084]), .rectangle3_x(rectangle3_xs[1084]), .rectangle3_y(rectangle3_ys[1084]), .rectangle3_width(rectangle3_widths[1084]), .rectangle3_height(rectangle3_heights[1084]), .rectangle3_weight(rectangle3_weights[1084]), .feature_threshold(feature_thresholds[1084]), .feature_above(feature_aboves[1084]), .feature_below(feature_belows[1084]), .scan_win_std_dev(scan_win_std_dev[1084]), .feature_accum(feature_accums[1084]));
  accum_calculator ac1085(.scan_win(scan_win1085), .rectangle1_x(rectangle1_xs[1085]), .rectangle1_y(rectangle1_ys[1085]), .rectangle1_width(rectangle1_widths[1085]), .rectangle1_height(rectangle1_heights[1085]), .rectangle1_weight(rectangle1_weights[1085]), .rectangle2_x(rectangle2_xs[1085]), .rectangle2_y(rectangle2_ys[1085]), .rectangle2_width(rectangle2_widths[1085]), .rectangle2_height(rectangle2_heights[1085]), .rectangle2_weight(rectangle2_weights[1085]), .rectangle3_x(rectangle3_xs[1085]), .rectangle3_y(rectangle3_ys[1085]), .rectangle3_width(rectangle3_widths[1085]), .rectangle3_height(rectangle3_heights[1085]), .rectangle3_weight(rectangle3_weights[1085]), .feature_threshold(feature_thresholds[1085]), .feature_above(feature_aboves[1085]), .feature_below(feature_belows[1085]), .scan_win_std_dev(scan_win_std_dev[1085]), .feature_accum(feature_accums[1085]));
  accum_calculator ac1086(.scan_win(scan_win1086), .rectangle1_x(rectangle1_xs[1086]), .rectangle1_y(rectangle1_ys[1086]), .rectangle1_width(rectangle1_widths[1086]), .rectangle1_height(rectangle1_heights[1086]), .rectangle1_weight(rectangle1_weights[1086]), .rectangle2_x(rectangle2_xs[1086]), .rectangle2_y(rectangle2_ys[1086]), .rectangle2_width(rectangle2_widths[1086]), .rectangle2_height(rectangle2_heights[1086]), .rectangle2_weight(rectangle2_weights[1086]), .rectangle3_x(rectangle3_xs[1086]), .rectangle3_y(rectangle3_ys[1086]), .rectangle3_width(rectangle3_widths[1086]), .rectangle3_height(rectangle3_heights[1086]), .rectangle3_weight(rectangle3_weights[1086]), .feature_threshold(feature_thresholds[1086]), .feature_above(feature_aboves[1086]), .feature_below(feature_belows[1086]), .scan_win_std_dev(scan_win_std_dev[1086]), .feature_accum(feature_accums[1086]));
  accum_calculator ac1087(.scan_win(scan_win1087), .rectangle1_x(rectangle1_xs[1087]), .rectangle1_y(rectangle1_ys[1087]), .rectangle1_width(rectangle1_widths[1087]), .rectangle1_height(rectangle1_heights[1087]), .rectangle1_weight(rectangle1_weights[1087]), .rectangle2_x(rectangle2_xs[1087]), .rectangle2_y(rectangle2_ys[1087]), .rectangle2_width(rectangle2_widths[1087]), .rectangle2_height(rectangle2_heights[1087]), .rectangle2_weight(rectangle2_weights[1087]), .rectangle3_x(rectangle3_xs[1087]), .rectangle3_y(rectangle3_ys[1087]), .rectangle3_width(rectangle3_widths[1087]), .rectangle3_height(rectangle3_heights[1087]), .rectangle3_weight(rectangle3_weights[1087]), .feature_threshold(feature_thresholds[1087]), .feature_above(feature_aboves[1087]), .feature_below(feature_belows[1087]), .scan_win_std_dev(scan_win_std_dev[1087]), .feature_accum(feature_accums[1087]));
  accum_calculator ac1088(.scan_win(scan_win1088), .rectangle1_x(rectangle1_xs[1088]), .rectangle1_y(rectangle1_ys[1088]), .rectangle1_width(rectangle1_widths[1088]), .rectangle1_height(rectangle1_heights[1088]), .rectangle1_weight(rectangle1_weights[1088]), .rectangle2_x(rectangle2_xs[1088]), .rectangle2_y(rectangle2_ys[1088]), .rectangle2_width(rectangle2_widths[1088]), .rectangle2_height(rectangle2_heights[1088]), .rectangle2_weight(rectangle2_weights[1088]), .rectangle3_x(rectangle3_xs[1088]), .rectangle3_y(rectangle3_ys[1088]), .rectangle3_width(rectangle3_widths[1088]), .rectangle3_height(rectangle3_heights[1088]), .rectangle3_weight(rectangle3_weights[1088]), .feature_threshold(feature_thresholds[1088]), .feature_above(feature_aboves[1088]), .feature_below(feature_belows[1088]), .scan_win_std_dev(scan_win_std_dev[1088]), .feature_accum(feature_accums[1088]));
  accum_calculator ac1089(.scan_win(scan_win1089), .rectangle1_x(rectangle1_xs[1089]), .rectangle1_y(rectangle1_ys[1089]), .rectangle1_width(rectangle1_widths[1089]), .rectangle1_height(rectangle1_heights[1089]), .rectangle1_weight(rectangle1_weights[1089]), .rectangle2_x(rectangle2_xs[1089]), .rectangle2_y(rectangle2_ys[1089]), .rectangle2_width(rectangle2_widths[1089]), .rectangle2_height(rectangle2_heights[1089]), .rectangle2_weight(rectangle2_weights[1089]), .rectangle3_x(rectangle3_xs[1089]), .rectangle3_y(rectangle3_ys[1089]), .rectangle3_width(rectangle3_widths[1089]), .rectangle3_height(rectangle3_heights[1089]), .rectangle3_weight(rectangle3_weights[1089]), .feature_threshold(feature_thresholds[1089]), .feature_above(feature_aboves[1089]), .feature_below(feature_belows[1089]), .scan_win_std_dev(scan_win_std_dev[1089]), .feature_accum(feature_accums[1089]));
  accum_calculator ac1090(.scan_win(scan_win1090), .rectangle1_x(rectangle1_xs[1090]), .rectangle1_y(rectangle1_ys[1090]), .rectangle1_width(rectangle1_widths[1090]), .rectangle1_height(rectangle1_heights[1090]), .rectangle1_weight(rectangle1_weights[1090]), .rectangle2_x(rectangle2_xs[1090]), .rectangle2_y(rectangle2_ys[1090]), .rectangle2_width(rectangle2_widths[1090]), .rectangle2_height(rectangle2_heights[1090]), .rectangle2_weight(rectangle2_weights[1090]), .rectangle3_x(rectangle3_xs[1090]), .rectangle3_y(rectangle3_ys[1090]), .rectangle3_width(rectangle3_widths[1090]), .rectangle3_height(rectangle3_heights[1090]), .rectangle3_weight(rectangle3_weights[1090]), .feature_threshold(feature_thresholds[1090]), .feature_above(feature_aboves[1090]), .feature_below(feature_belows[1090]), .scan_win_std_dev(scan_win_std_dev[1090]), .feature_accum(feature_accums[1090]));
  accum_calculator ac1091(.scan_win(scan_win1091), .rectangle1_x(rectangle1_xs[1091]), .rectangle1_y(rectangle1_ys[1091]), .rectangle1_width(rectangle1_widths[1091]), .rectangle1_height(rectangle1_heights[1091]), .rectangle1_weight(rectangle1_weights[1091]), .rectangle2_x(rectangle2_xs[1091]), .rectangle2_y(rectangle2_ys[1091]), .rectangle2_width(rectangle2_widths[1091]), .rectangle2_height(rectangle2_heights[1091]), .rectangle2_weight(rectangle2_weights[1091]), .rectangle3_x(rectangle3_xs[1091]), .rectangle3_y(rectangle3_ys[1091]), .rectangle3_width(rectangle3_widths[1091]), .rectangle3_height(rectangle3_heights[1091]), .rectangle3_weight(rectangle3_weights[1091]), .feature_threshold(feature_thresholds[1091]), .feature_above(feature_aboves[1091]), .feature_below(feature_belows[1091]), .scan_win_std_dev(scan_win_std_dev[1091]), .feature_accum(feature_accums[1091]));
  accum_calculator ac1092(.scan_win(scan_win1092), .rectangle1_x(rectangle1_xs[1092]), .rectangle1_y(rectangle1_ys[1092]), .rectangle1_width(rectangle1_widths[1092]), .rectangle1_height(rectangle1_heights[1092]), .rectangle1_weight(rectangle1_weights[1092]), .rectangle2_x(rectangle2_xs[1092]), .rectangle2_y(rectangle2_ys[1092]), .rectangle2_width(rectangle2_widths[1092]), .rectangle2_height(rectangle2_heights[1092]), .rectangle2_weight(rectangle2_weights[1092]), .rectangle3_x(rectangle3_xs[1092]), .rectangle3_y(rectangle3_ys[1092]), .rectangle3_width(rectangle3_widths[1092]), .rectangle3_height(rectangle3_heights[1092]), .rectangle3_weight(rectangle3_weights[1092]), .feature_threshold(feature_thresholds[1092]), .feature_above(feature_aboves[1092]), .feature_below(feature_belows[1092]), .scan_win_std_dev(scan_win_std_dev[1092]), .feature_accum(feature_accums[1092]));
  accum_calculator ac1093(.scan_win(scan_win1093), .rectangle1_x(rectangle1_xs[1093]), .rectangle1_y(rectangle1_ys[1093]), .rectangle1_width(rectangle1_widths[1093]), .rectangle1_height(rectangle1_heights[1093]), .rectangle1_weight(rectangle1_weights[1093]), .rectangle2_x(rectangle2_xs[1093]), .rectangle2_y(rectangle2_ys[1093]), .rectangle2_width(rectangle2_widths[1093]), .rectangle2_height(rectangle2_heights[1093]), .rectangle2_weight(rectangle2_weights[1093]), .rectangle3_x(rectangle3_xs[1093]), .rectangle3_y(rectangle3_ys[1093]), .rectangle3_width(rectangle3_widths[1093]), .rectangle3_height(rectangle3_heights[1093]), .rectangle3_weight(rectangle3_weights[1093]), .feature_threshold(feature_thresholds[1093]), .feature_above(feature_aboves[1093]), .feature_below(feature_belows[1093]), .scan_win_std_dev(scan_win_std_dev[1093]), .feature_accum(feature_accums[1093]));
  accum_calculator ac1094(.scan_win(scan_win1094), .rectangle1_x(rectangle1_xs[1094]), .rectangle1_y(rectangle1_ys[1094]), .rectangle1_width(rectangle1_widths[1094]), .rectangle1_height(rectangle1_heights[1094]), .rectangle1_weight(rectangle1_weights[1094]), .rectangle2_x(rectangle2_xs[1094]), .rectangle2_y(rectangle2_ys[1094]), .rectangle2_width(rectangle2_widths[1094]), .rectangle2_height(rectangle2_heights[1094]), .rectangle2_weight(rectangle2_weights[1094]), .rectangle3_x(rectangle3_xs[1094]), .rectangle3_y(rectangle3_ys[1094]), .rectangle3_width(rectangle3_widths[1094]), .rectangle3_height(rectangle3_heights[1094]), .rectangle3_weight(rectangle3_weights[1094]), .feature_threshold(feature_thresholds[1094]), .feature_above(feature_aboves[1094]), .feature_below(feature_belows[1094]), .scan_win_std_dev(scan_win_std_dev[1094]), .feature_accum(feature_accums[1094]));
  accum_calculator ac1095(.scan_win(scan_win1095), .rectangle1_x(rectangle1_xs[1095]), .rectangle1_y(rectangle1_ys[1095]), .rectangle1_width(rectangle1_widths[1095]), .rectangle1_height(rectangle1_heights[1095]), .rectangle1_weight(rectangle1_weights[1095]), .rectangle2_x(rectangle2_xs[1095]), .rectangle2_y(rectangle2_ys[1095]), .rectangle2_width(rectangle2_widths[1095]), .rectangle2_height(rectangle2_heights[1095]), .rectangle2_weight(rectangle2_weights[1095]), .rectangle3_x(rectangle3_xs[1095]), .rectangle3_y(rectangle3_ys[1095]), .rectangle3_width(rectangle3_widths[1095]), .rectangle3_height(rectangle3_heights[1095]), .rectangle3_weight(rectangle3_weights[1095]), .feature_threshold(feature_thresholds[1095]), .feature_above(feature_aboves[1095]), .feature_below(feature_belows[1095]), .scan_win_std_dev(scan_win_std_dev[1095]), .feature_accum(feature_accums[1095]));
  accum_calculator ac1096(.scan_win(scan_win1096), .rectangle1_x(rectangle1_xs[1096]), .rectangle1_y(rectangle1_ys[1096]), .rectangle1_width(rectangle1_widths[1096]), .rectangle1_height(rectangle1_heights[1096]), .rectangle1_weight(rectangle1_weights[1096]), .rectangle2_x(rectangle2_xs[1096]), .rectangle2_y(rectangle2_ys[1096]), .rectangle2_width(rectangle2_widths[1096]), .rectangle2_height(rectangle2_heights[1096]), .rectangle2_weight(rectangle2_weights[1096]), .rectangle3_x(rectangle3_xs[1096]), .rectangle3_y(rectangle3_ys[1096]), .rectangle3_width(rectangle3_widths[1096]), .rectangle3_height(rectangle3_heights[1096]), .rectangle3_weight(rectangle3_weights[1096]), .feature_threshold(feature_thresholds[1096]), .feature_above(feature_aboves[1096]), .feature_below(feature_belows[1096]), .scan_win_std_dev(scan_win_std_dev[1096]), .feature_accum(feature_accums[1096]));
  accum_calculator ac1097(.scan_win(scan_win1097), .rectangle1_x(rectangle1_xs[1097]), .rectangle1_y(rectangle1_ys[1097]), .rectangle1_width(rectangle1_widths[1097]), .rectangle1_height(rectangle1_heights[1097]), .rectangle1_weight(rectangle1_weights[1097]), .rectangle2_x(rectangle2_xs[1097]), .rectangle2_y(rectangle2_ys[1097]), .rectangle2_width(rectangle2_widths[1097]), .rectangle2_height(rectangle2_heights[1097]), .rectangle2_weight(rectangle2_weights[1097]), .rectangle3_x(rectangle3_xs[1097]), .rectangle3_y(rectangle3_ys[1097]), .rectangle3_width(rectangle3_widths[1097]), .rectangle3_height(rectangle3_heights[1097]), .rectangle3_weight(rectangle3_weights[1097]), .feature_threshold(feature_thresholds[1097]), .feature_above(feature_aboves[1097]), .feature_below(feature_belows[1097]), .scan_win_std_dev(scan_win_std_dev[1097]), .feature_accum(feature_accums[1097]));
  accum_calculator ac1098(.scan_win(scan_win1098), .rectangle1_x(rectangle1_xs[1098]), .rectangle1_y(rectangle1_ys[1098]), .rectangle1_width(rectangle1_widths[1098]), .rectangle1_height(rectangle1_heights[1098]), .rectangle1_weight(rectangle1_weights[1098]), .rectangle2_x(rectangle2_xs[1098]), .rectangle2_y(rectangle2_ys[1098]), .rectangle2_width(rectangle2_widths[1098]), .rectangle2_height(rectangle2_heights[1098]), .rectangle2_weight(rectangle2_weights[1098]), .rectangle3_x(rectangle3_xs[1098]), .rectangle3_y(rectangle3_ys[1098]), .rectangle3_width(rectangle3_widths[1098]), .rectangle3_height(rectangle3_heights[1098]), .rectangle3_weight(rectangle3_weights[1098]), .feature_threshold(feature_thresholds[1098]), .feature_above(feature_aboves[1098]), .feature_below(feature_belows[1098]), .scan_win_std_dev(scan_win_std_dev[1098]), .feature_accum(feature_accums[1098]));
  accum_calculator ac1099(.scan_win(scan_win1099), .rectangle1_x(rectangle1_xs[1099]), .rectangle1_y(rectangle1_ys[1099]), .rectangle1_width(rectangle1_widths[1099]), .rectangle1_height(rectangle1_heights[1099]), .rectangle1_weight(rectangle1_weights[1099]), .rectangle2_x(rectangle2_xs[1099]), .rectangle2_y(rectangle2_ys[1099]), .rectangle2_width(rectangle2_widths[1099]), .rectangle2_height(rectangle2_heights[1099]), .rectangle2_weight(rectangle2_weights[1099]), .rectangle3_x(rectangle3_xs[1099]), .rectangle3_y(rectangle3_ys[1099]), .rectangle3_width(rectangle3_widths[1099]), .rectangle3_height(rectangle3_heights[1099]), .rectangle3_weight(rectangle3_weights[1099]), .feature_threshold(feature_thresholds[1099]), .feature_above(feature_aboves[1099]), .feature_below(feature_belows[1099]), .scan_win_std_dev(scan_win_std_dev[1099]), .feature_accum(feature_accums[1099]));
  accum_calculator ac1100(.scan_win(scan_win1100), .rectangle1_x(rectangle1_xs[1100]), .rectangle1_y(rectangle1_ys[1100]), .rectangle1_width(rectangle1_widths[1100]), .rectangle1_height(rectangle1_heights[1100]), .rectangle1_weight(rectangle1_weights[1100]), .rectangle2_x(rectangle2_xs[1100]), .rectangle2_y(rectangle2_ys[1100]), .rectangle2_width(rectangle2_widths[1100]), .rectangle2_height(rectangle2_heights[1100]), .rectangle2_weight(rectangle2_weights[1100]), .rectangle3_x(rectangle3_xs[1100]), .rectangle3_y(rectangle3_ys[1100]), .rectangle3_width(rectangle3_widths[1100]), .rectangle3_height(rectangle3_heights[1100]), .rectangle3_weight(rectangle3_weights[1100]), .feature_threshold(feature_thresholds[1100]), .feature_above(feature_aboves[1100]), .feature_below(feature_belows[1100]), .scan_win_std_dev(scan_win_std_dev[1100]), .feature_accum(feature_accums[1100]));
  accum_calculator ac1101(.scan_win(scan_win1101), .rectangle1_x(rectangle1_xs[1101]), .rectangle1_y(rectangle1_ys[1101]), .rectangle1_width(rectangle1_widths[1101]), .rectangle1_height(rectangle1_heights[1101]), .rectangle1_weight(rectangle1_weights[1101]), .rectangle2_x(rectangle2_xs[1101]), .rectangle2_y(rectangle2_ys[1101]), .rectangle2_width(rectangle2_widths[1101]), .rectangle2_height(rectangle2_heights[1101]), .rectangle2_weight(rectangle2_weights[1101]), .rectangle3_x(rectangle3_xs[1101]), .rectangle3_y(rectangle3_ys[1101]), .rectangle3_width(rectangle3_widths[1101]), .rectangle3_height(rectangle3_heights[1101]), .rectangle3_weight(rectangle3_weights[1101]), .feature_threshold(feature_thresholds[1101]), .feature_above(feature_aboves[1101]), .feature_below(feature_belows[1101]), .scan_win_std_dev(scan_win_std_dev[1101]), .feature_accum(feature_accums[1101]));
  accum_calculator ac1102(.scan_win(scan_win1102), .rectangle1_x(rectangle1_xs[1102]), .rectangle1_y(rectangle1_ys[1102]), .rectangle1_width(rectangle1_widths[1102]), .rectangle1_height(rectangle1_heights[1102]), .rectangle1_weight(rectangle1_weights[1102]), .rectangle2_x(rectangle2_xs[1102]), .rectangle2_y(rectangle2_ys[1102]), .rectangle2_width(rectangle2_widths[1102]), .rectangle2_height(rectangle2_heights[1102]), .rectangle2_weight(rectangle2_weights[1102]), .rectangle3_x(rectangle3_xs[1102]), .rectangle3_y(rectangle3_ys[1102]), .rectangle3_width(rectangle3_widths[1102]), .rectangle3_height(rectangle3_heights[1102]), .rectangle3_weight(rectangle3_weights[1102]), .feature_threshold(feature_thresholds[1102]), .feature_above(feature_aboves[1102]), .feature_below(feature_belows[1102]), .scan_win_std_dev(scan_win_std_dev[1102]), .feature_accum(feature_accums[1102]));
  accum_calculator ac1103(.scan_win(scan_win1103), .rectangle1_x(rectangle1_xs[1103]), .rectangle1_y(rectangle1_ys[1103]), .rectangle1_width(rectangle1_widths[1103]), .rectangle1_height(rectangle1_heights[1103]), .rectangle1_weight(rectangle1_weights[1103]), .rectangle2_x(rectangle2_xs[1103]), .rectangle2_y(rectangle2_ys[1103]), .rectangle2_width(rectangle2_widths[1103]), .rectangle2_height(rectangle2_heights[1103]), .rectangle2_weight(rectangle2_weights[1103]), .rectangle3_x(rectangle3_xs[1103]), .rectangle3_y(rectangle3_ys[1103]), .rectangle3_width(rectangle3_widths[1103]), .rectangle3_height(rectangle3_heights[1103]), .rectangle3_weight(rectangle3_weights[1103]), .feature_threshold(feature_thresholds[1103]), .feature_above(feature_aboves[1103]), .feature_below(feature_belows[1103]), .scan_win_std_dev(scan_win_std_dev[1103]), .feature_accum(feature_accums[1103]));
  accum_calculator ac1104(.scan_win(scan_win1104), .rectangle1_x(rectangle1_xs[1104]), .rectangle1_y(rectangle1_ys[1104]), .rectangle1_width(rectangle1_widths[1104]), .rectangle1_height(rectangle1_heights[1104]), .rectangle1_weight(rectangle1_weights[1104]), .rectangle2_x(rectangle2_xs[1104]), .rectangle2_y(rectangle2_ys[1104]), .rectangle2_width(rectangle2_widths[1104]), .rectangle2_height(rectangle2_heights[1104]), .rectangle2_weight(rectangle2_weights[1104]), .rectangle3_x(rectangle3_xs[1104]), .rectangle3_y(rectangle3_ys[1104]), .rectangle3_width(rectangle3_widths[1104]), .rectangle3_height(rectangle3_heights[1104]), .rectangle3_weight(rectangle3_weights[1104]), .feature_threshold(feature_thresholds[1104]), .feature_above(feature_aboves[1104]), .feature_below(feature_belows[1104]), .scan_win_std_dev(scan_win_std_dev[1104]), .feature_accum(feature_accums[1104]));
  accum_calculator ac1105(.scan_win(scan_win1105), .rectangle1_x(rectangle1_xs[1105]), .rectangle1_y(rectangle1_ys[1105]), .rectangle1_width(rectangle1_widths[1105]), .rectangle1_height(rectangle1_heights[1105]), .rectangle1_weight(rectangle1_weights[1105]), .rectangle2_x(rectangle2_xs[1105]), .rectangle2_y(rectangle2_ys[1105]), .rectangle2_width(rectangle2_widths[1105]), .rectangle2_height(rectangle2_heights[1105]), .rectangle2_weight(rectangle2_weights[1105]), .rectangle3_x(rectangle3_xs[1105]), .rectangle3_y(rectangle3_ys[1105]), .rectangle3_width(rectangle3_widths[1105]), .rectangle3_height(rectangle3_heights[1105]), .rectangle3_weight(rectangle3_weights[1105]), .feature_threshold(feature_thresholds[1105]), .feature_above(feature_aboves[1105]), .feature_below(feature_belows[1105]), .scan_win_std_dev(scan_win_std_dev[1105]), .feature_accum(feature_accums[1105]));
  accum_calculator ac1106(.scan_win(scan_win1106), .rectangle1_x(rectangle1_xs[1106]), .rectangle1_y(rectangle1_ys[1106]), .rectangle1_width(rectangle1_widths[1106]), .rectangle1_height(rectangle1_heights[1106]), .rectangle1_weight(rectangle1_weights[1106]), .rectangle2_x(rectangle2_xs[1106]), .rectangle2_y(rectangle2_ys[1106]), .rectangle2_width(rectangle2_widths[1106]), .rectangle2_height(rectangle2_heights[1106]), .rectangle2_weight(rectangle2_weights[1106]), .rectangle3_x(rectangle3_xs[1106]), .rectangle3_y(rectangle3_ys[1106]), .rectangle3_width(rectangle3_widths[1106]), .rectangle3_height(rectangle3_heights[1106]), .rectangle3_weight(rectangle3_weights[1106]), .feature_threshold(feature_thresholds[1106]), .feature_above(feature_aboves[1106]), .feature_below(feature_belows[1106]), .scan_win_std_dev(scan_win_std_dev[1106]), .feature_accum(feature_accums[1106]));
  accum_calculator ac1107(.scan_win(scan_win1107), .rectangle1_x(rectangle1_xs[1107]), .rectangle1_y(rectangle1_ys[1107]), .rectangle1_width(rectangle1_widths[1107]), .rectangle1_height(rectangle1_heights[1107]), .rectangle1_weight(rectangle1_weights[1107]), .rectangle2_x(rectangle2_xs[1107]), .rectangle2_y(rectangle2_ys[1107]), .rectangle2_width(rectangle2_widths[1107]), .rectangle2_height(rectangle2_heights[1107]), .rectangle2_weight(rectangle2_weights[1107]), .rectangle3_x(rectangle3_xs[1107]), .rectangle3_y(rectangle3_ys[1107]), .rectangle3_width(rectangle3_widths[1107]), .rectangle3_height(rectangle3_heights[1107]), .rectangle3_weight(rectangle3_weights[1107]), .feature_threshold(feature_thresholds[1107]), .feature_above(feature_aboves[1107]), .feature_below(feature_belows[1107]), .scan_win_std_dev(scan_win_std_dev[1107]), .feature_accum(feature_accums[1107]));
  accum_calculator ac1108(.scan_win(scan_win1108), .rectangle1_x(rectangle1_xs[1108]), .rectangle1_y(rectangle1_ys[1108]), .rectangle1_width(rectangle1_widths[1108]), .rectangle1_height(rectangle1_heights[1108]), .rectangle1_weight(rectangle1_weights[1108]), .rectangle2_x(rectangle2_xs[1108]), .rectangle2_y(rectangle2_ys[1108]), .rectangle2_width(rectangle2_widths[1108]), .rectangle2_height(rectangle2_heights[1108]), .rectangle2_weight(rectangle2_weights[1108]), .rectangle3_x(rectangle3_xs[1108]), .rectangle3_y(rectangle3_ys[1108]), .rectangle3_width(rectangle3_widths[1108]), .rectangle3_height(rectangle3_heights[1108]), .rectangle3_weight(rectangle3_weights[1108]), .feature_threshold(feature_thresholds[1108]), .feature_above(feature_aboves[1108]), .feature_below(feature_belows[1108]), .scan_win_std_dev(scan_win_std_dev[1108]), .feature_accum(feature_accums[1108]));
  accum_calculator ac1109(.scan_win(scan_win1109), .rectangle1_x(rectangle1_xs[1109]), .rectangle1_y(rectangle1_ys[1109]), .rectangle1_width(rectangle1_widths[1109]), .rectangle1_height(rectangle1_heights[1109]), .rectangle1_weight(rectangle1_weights[1109]), .rectangle2_x(rectangle2_xs[1109]), .rectangle2_y(rectangle2_ys[1109]), .rectangle2_width(rectangle2_widths[1109]), .rectangle2_height(rectangle2_heights[1109]), .rectangle2_weight(rectangle2_weights[1109]), .rectangle3_x(rectangle3_xs[1109]), .rectangle3_y(rectangle3_ys[1109]), .rectangle3_width(rectangle3_widths[1109]), .rectangle3_height(rectangle3_heights[1109]), .rectangle3_weight(rectangle3_weights[1109]), .feature_threshold(feature_thresholds[1109]), .feature_above(feature_aboves[1109]), .feature_below(feature_belows[1109]), .scan_win_std_dev(scan_win_std_dev[1109]), .feature_accum(feature_accums[1109]));
  accum_calculator ac1110(.scan_win(scan_win1110), .rectangle1_x(rectangle1_xs[1110]), .rectangle1_y(rectangle1_ys[1110]), .rectangle1_width(rectangle1_widths[1110]), .rectangle1_height(rectangle1_heights[1110]), .rectangle1_weight(rectangle1_weights[1110]), .rectangle2_x(rectangle2_xs[1110]), .rectangle2_y(rectangle2_ys[1110]), .rectangle2_width(rectangle2_widths[1110]), .rectangle2_height(rectangle2_heights[1110]), .rectangle2_weight(rectangle2_weights[1110]), .rectangle3_x(rectangle3_xs[1110]), .rectangle3_y(rectangle3_ys[1110]), .rectangle3_width(rectangle3_widths[1110]), .rectangle3_height(rectangle3_heights[1110]), .rectangle3_weight(rectangle3_weights[1110]), .feature_threshold(feature_thresholds[1110]), .feature_above(feature_aboves[1110]), .feature_below(feature_belows[1110]), .scan_win_std_dev(scan_win_std_dev[1110]), .feature_accum(feature_accums[1110]));
  accum_calculator ac1111(.scan_win(scan_win1111), .rectangle1_x(rectangle1_xs[1111]), .rectangle1_y(rectangle1_ys[1111]), .rectangle1_width(rectangle1_widths[1111]), .rectangle1_height(rectangle1_heights[1111]), .rectangle1_weight(rectangle1_weights[1111]), .rectangle2_x(rectangle2_xs[1111]), .rectangle2_y(rectangle2_ys[1111]), .rectangle2_width(rectangle2_widths[1111]), .rectangle2_height(rectangle2_heights[1111]), .rectangle2_weight(rectangle2_weights[1111]), .rectangle3_x(rectangle3_xs[1111]), .rectangle3_y(rectangle3_ys[1111]), .rectangle3_width(rectangle3_widths[1111]), .rectangle3_height(rectangle3_heights[1111]), .rectangle3_weight(rectangle3_weights[1111]), .feature_threshold(feature_thresholds[1111]), .feature_above(feature_aboves[1111]), .feature_below(feature_belows[1111]), .scan_win_std_dev(scan_win_std_dev[1111]), .feature_accum(feature_accums[1111]));
  accum_calculator ac1112(.scan_win(scan_win1112), .rectangle1_x(rectangle1_xs[1112]), .rectangle1_y(rectangle1_ys[1112]), .rectangle1_width(rectangle1_widths[1112]), .rectangle1_height(rectangle1_heights[1112]), .rectangle1_weight(rectangle1_weights[1112]), .rectangle2_x(rectangle2_xs[1112]), .rectangle2_y(rectangle2_ys[1112]), .rectangle2_width(rectangle2_widths[1112]), .rectangle2_height(rectangle2_heights[1112]), .rectangle2_weight(rectangle2_weights[1112]), .rectangle3_x(rectangle3_xs[1112]), .rectangle3_y(rectangle3_ys[1112]), .rectangle3_width(rectangle3_widths[1112]), .rectangle3_height(rectangle3_heights[1112]), .rectangle3_weight(rectangle3_weights[1112]), .feature_threshold(feature_thresholds[1112]), .feature_above(feature_aboves[1112]), .feature_below(feature_belows[1112]), .scan_win_std_dev(scan_win_std_dev[1112]), .feature_accum(feature_accums[1112]));
  accum_calculator ac1113(.scan_win(scan_win1113), .rectangle1_x(rectangle1_xs[1113]), .rectangle1_y(rectangle1_ys[1113]), .rectangle1_width(rectangle1_widths[1113]), .rectangle1_height(rectangle1_heights[1113]), .rectangle1_weight(rectangle1_weights[1113]), .rectangle2_x(rectangle2_xs[1113]), .rectangle2_y(rectangle2_ys[1113]), .rectangle2_width(rectangle2_widths[1113]), .rectangle2_height(rectangle2_heights[1113]), .rectangle2_weight(rectangle2_weights[1113]), .rectangle3_x(rectangle3_xs[1113]), .rectangle3_y(rectangle3_ys[1113]), .rectangle3_width(rectangle3_widths[1113]), .rectangle3_height(rectangle3_heights[1113]), .rectangle3_weight(rectangle3_weights[1113]), .feature_threshold(feature_thresholds[1113]), .feature_above(feature_aboves[1113]), .feature_below(feature_belows[1113]), .scan_win_std_dev(scan_win_std_dev[1113]), .feature_accum(feature_accums[1113]));
  accum_calculator ac1114(.scan_win(scan_win1114), .rectangle1_x(rectangle1_xs[1114]), .rectangle1_y(rectangle1_ys[1114]), .rectangle1_width(rectangle1_widths[1114]), .rectangle1_height(rectangle1_heights[1114]), .rectangle1_weight(rectangle1_weights[1114]), .rectangle2_x(rectangle2_xs[1114]), .rectangle2_y(rectangle2_ys[1114]), .rectangle2_width(rectangle2_widths[1114]), .rectangle2_height(rectangle2_heights[1114]), .rectangle2_weight(rectangle2_weights[1114]), .rectangle3_x(rectangle3_xs[1114]), .rectangle3_y(rectangle3_ys[1114]), .rectangle3_width(rectangle3_widths[1114]), .rectangle3_height(rectangle3_heights[1114]), .rectangle3_weight(rectangle3_weights[1114]), .feature_threshold(feature_thresholds[1114]), .feature_above(feature_aboves[1114]), .feature_below(feature_belows[1114]), .scan_win_std_dev(scan_win_std_dev[1114]), .feature_accum(feature_accums[1114]));
  accum_calculator ac1115(.scan_win(scan_win1115), .rectangle1_x(rectangle1_xs[1115]), .rectangle1_y(rectangle1_ys[1115]), .rectangle1_width(rectangle1_widths[1115]), .rectangle1_height(rectangle1_heights[1115]), .rectangle1_weight(rectangle1_weights[1115]), .rectangle2_x(rectangle2_xs[1115]), .rectangle2_y(rectangle2_ys[1115]), .rectangle2_width(rectangle2_widths[1115]), .rectangle2_height(rectangle2_heights[1115]), .rectangle2_weight(rectangle2_weights[1115]), .rectangle3_x(rectangle3_xs[1115]), .rectangle3_y(rectangle3_ys[1115]), .rectangle3_width(rectangle3_widths[1115]), .rectangle3_height(rectangle3_heights[1115]), .rectangle3_weight(rectangle3_weights[1115]), .feature_threshold(feature_thresholds[1115]), .feature_above(feature_aboves[1115]), .feature_below(feature_belows[1115]), .scan_win_std_dev(scan_win_std_dev[1115]), .feature_accum(feature_accums[1115]));
  accum_calculator ac1116(.scan_win(scan_win1116), .rectangle1_x(rectangle1_xs[1116]), .rectangle1_y(rectangle1_ys[1116]), .rectangle1_width(rectangle1_widths[1116]), .rectangle1_height(rectangle1_heights[1116]), .rectangle1_weight(rectangle1_weights[1116]), .rectangle2_x(rectangle2_xs[1116]), .rectangle2_y(rectangle2_ys[1116]), .rectangle2_width(rectangle2_widths[1116]), .rectangle2_height(rectangle2_heights[1116]), .rectangle2_weight(rectangle2_weights[1116]), .rectangle3_x(rectangle3_xs[1116]), .rectangle3_y(rectangle3_ys[1116]), .rectangle3_width(rectangle3_widths[1116]), .rectangle3_height(rectangle3_heights[1116]), .rectangle3_weight(rectangle3_weights[1116]), .feature_threshold(feature_thresholds[1116]), .feature_above(feature_aboves[1116]), .feature_below(feature_belows[1116]), .scan_win_std_dev(scan_win_std_dev[1116]), .feature_accum(feature_accums[1116]));
  accum_calculator ac1117(.scan_win(scan_win1117), .rectangle1_x(rectangle1_xs[1117]), .rectangle1_y(rectangle1_ys[1117]), .rectangle1_width(rectangle1_widths[1117]), .rectangle1_height(rectangle1_heights[1117]), .rectangle1_weight(rectangle1_weights[1117]), .rectangle2_x(rectangle2_xs[1117]), .rectangle2_y(rectangle2_ys[1117]), .rectangle2_width(rectangle2_widths[1117]), .rectangle2_height(rectangle2_heights[1117]), .rectangle2_weight(rectangle2_weights[1117]), .rectangle3_x(rectangle3_xs[1117]), .rectangle3_y(rectangle3_ys[1117]), .rectangle3_width(rectangle3_widths[1117]), .rectangle3_height(rectangle3_heights[1117]), .rectangle3_weight(rectangle3_weights[1117]), .feature_threshold(feature_thresholds[1117]), .feature_above(feature_aboves[1117]), .feature_below(feature_belows[1117]), .scan_win_std_dev(scan_win_std_dev[1117]), .feature_accum(feature_accums[1117]));
  accum_calculator ac1118(.scan_win(scan_win1118), .rectangle1_x(rectangle1_xs[1118]), .rectangle1_y(rectangle1_ys[1118]), .rectangle1_width(rectangle1_widths[1118]), .rectangle1_height(rectangle1_heights[1118]), .rectangle1_weight(rectangle1_weights[1118]), .rectangle2_x(rectangle2_xs[1118]), .rectangle2_y(rectangle2_ys[1118]), .rectangle2_width(rectangle2_widths[1118]), .rectangle2_height(rectangle2_heights[1118]), .rectangle2_weight(rectangle2_weights[1118]), .rectangle3_x(rectangle3_xs[1118]), .rectangle3_y(rectangle3_ys[1118]), .rectangle3_width(rectangle3_widths[1118]), .rectangle3_height(rectangle3_heights[1118]), .rectangle3_weight(rectangle3_weights[1118]), .feature_threshold(feature_thresholds[1118]), .feature_above(feature_aboves[1118]), .feature_below(feature_belows[1118]), .scan_win_std_dev(scan_win_std_dev[1118]), .feature_accum(feature_accums[1118]));
  accum_calculator ac1119(.scan_win(scan_win1119), .rectangle1_x(rectangle1_xs[1119]), .rectangle1_y(rectangle1_ys[1119]), .rectangle1_width(rectangle1_widths[1119]), .rectangle1_height(rectangle1_heights[1119]), .rectangle1_weight(rectangle1_weights[1119]), .rectangle2_x(rectangle2_xs[1119]), .rectangle2_y(rectangle2_ys[1119]), .rectangle2_width(rectangle2_widths[1119]), .rectangle2_height(rectangle2_heights[1119]), .rectangle2_weight(rectangle2_weights[1119]), .rectangle3_x(rectangle3_xs[1119]), .rectangle3_y(rectangle3_ys[1119]), .rectangle3_width(rectangle3_widths[1119]), .rectangle3_height(rectangle3_heights[1119]), .rectangle3_weight(rectangle3_weights[1119]), .feature_threshold(feature_thresholds[1119]), .feature_above(feature_aboves[1119]), .feature_below(feature_belows[1119]), .scan_win_std_dev(scan_win_std_dev[1119]), .feature_accum(feature_accums[1119]));
  accum_calculator ac1120(.scan_win(scan_win1120), .rectangle1_x(rectangle1_xs[1120]), .rectangle1_y(rectangle1_ys[1120]), .rectangle1_width(rectangle1_widths[1120]), .rectangle1_height(rectangle1_heights[1120]), .rectangle1_weight(rectangle1_weights[1120]), .rectangle2_x(rectangle2_xs[1120]), .rectangle2_y(rectangle2_ys[1120]), .rectangle2_width(rectangle2_widths[1120]), .rectangle2_height(rectangle2_heights[1120]), .rectangle2_weight(rectangle2_weights[1120]), .rectangle3_x(rectangle3_xs[1120]), .rectangle3_y(rectangle3_ys[1120]), .rectangle3_width(rectangle3_widths[1120]), .rectangle3_height(rectangle3_heights[1120]), .rectangle3_weight(rectangle3_weights[1120]), .feature_threshold(feature_thresholds[1120]), .feature_above(feature_aboves[1120]), .feature_below(feature_belows[1120]), .scan_win_std_dev(scan_win_std_dev[1120]), .feature_accum(feature_accums[1120]));
  accum_calculator ac1121(.scan_win(scan_win1121), .rectangle1_x(rectangle1_xs[1121]), .rectangle1_y(rectangle1_ys[1121]), .rectangle1_width(rectangle1_widths[1121]), .rectangle1_height(rectangle1_heights[1121]), .rectangle1_weight(rectangle1_weights[1121]), .rectangle2_x(rectangle2_xs[1121]), .rectangle2_y(rectangle2_ys[1121]), .rectangle2_width(rectangle2_widths[1121]), .rectangle2_height(rectangle2_heights[1121]), .rectangle2_weight(rectangle2_weights[1121]), .rectangle3_x(rectangle3_xs[1121]), .rectangle3_y(rectangle3_ys[1121]), .rectangle3_width(rectangle3_widths[1121]), .rectangle3_height(rectangle3_heights[1121]), .rectangle3_weight(rectangle3_weights[1121]), .feature_threshold(feature_thresholds[1121]), .feature_above(feature_aboves[1121]), .feature_below(feature_belows[1121]), .scan_win_std_dev(scan_win_std_dev[1121]), .feature_accum(feature_accums[1121]));
  accum_calculator ac1122(.scan_win(scan_win1122), .rectangle1_x(rectangle1_xs[1122]), .rectangle1_y(rectangle1_ys[1122]), .rectangle1_width(rectangle1_widths[1122]), .rectangle1_height(rectangle1_heights[1122]), .rectangle1_weight(rectangle1_weights[1122]), .rectangle2_x(rectangle2_xs[1122]), .rectangle2_y(rectangle2_ys[1122]), .rectangle2_width(rectangle2_widths[1122]), .rectangle2_height(rectangle2_heights[1122]), .rectangle2_weight(rectangle2_weights[1122]), .rectangle3_x(rectangle3_xs[1122]), .rectangle3_y(rectangle3_ys[1122]), .rectangle3_width(rectangle3_widths[1122]), .rectangle3_height(rectangle3_heights[1122]), .rectangle3_weight(rectangle3_weights[1122]), .feature_threshold(feature_thresholds[1122]), .feature_above(feature_aboves[1122]), .feature_below(feature_belows[1122]), .scan_win_std_dev(scan_win_std_dev[1122]), .feature_accum(feature_accums[1122]));
  accum_calculator ac1123(.scan_win(scan_win1123), .rectangle1_x(rectangle1_xs[1123]), .rectangle1_y(rectangle1_ys[1123]), .rectangle1_width(rectangle1_widths[1123]), .rectangle1_height(rectangle1_heights[1123]), .rectangle1_weight(rectangle1_weights[1123]), .rectangle2_x(rectangle2_xs[1123]), .rectangle2_y(rectangle2_ys[1123]), .rectangle2_width(rectangle2_widths[1123]), .rectangle2_height(rectangle2_heights[1123]), .rectangle2_weight(rectangle2_weights[1123]), .rectangle3_x(rectangle3_xs[1123]), .rectangle3_y(rectangle3_ys[1123]), .rectangle3_width(rectangle3_widths[1123]), .rectangle3_height(rectangle3_heights[1123]), .rectangle3_weight(rectangle3_weights[1123]), .feature_threshold(feature_thresholds[1123]), .feature_above(feature_aboves[1123]), .feature_below(feature_belows[1123]), .scan_win_std_dev(scan_win_std_dev[1123]), .feature_accum(feature_accums[1123]));
  accum_calculator ac1124(.scan_win(scan_win1124), .rectangle1_x(rectangle1_xs[1124]), .rectangle1_y(rectangle1_ys[1124]), .rectangle1_width(rectangle1_widths[1124]), .rectangle1_height(rectangle1_heights[1124]), .rectangle1_weight(rectangle1_weights[1124]), .rectangle2_x(rectangle2_xs[1124]), .rectangle2_y(rectangle2_ys[1124]), .rectangle2_width(rectangle2_widths[1124]), .rectangle2_height(rectangle2_heights[1124]), .rectangle2_weight(rectangle2_weights[1124]), .rectangle3_x(rectangle3_xs[1124]), .rectangle3_y(rectangle3_ys[1124]), .rectangle3_width(rectangle3_widths[1124]), .rectangle3_height(rectangle3_heights[1124]), .rectangle3_weight(rectangle3_weights[1124]), .feature_threshold(feature_thresholds[1124]), .feature_above(feature_aboves[1124]), .feature_below(feature_belows[1124]), .scan_win_std_dev(scan_win_std_dev[1124]), .feature_accum(feature_accums[1124]));
  accum_calculator ac1125(.scan_win(scan_win1125), .rectangle1_x(rectangle1_xs[1125]), .rectangle1_y(rectangle1_ys[1125]), .rectangle1_width(rectangle1_widths[1125]), .rectangle1_height(rectangle1_heights[1125]), .rectangle1_weight(rectangle1_weights[1125]), .rectangle2_x(rectangle2_xs[1125]), .rectangle2_y(rectangle2_ys[1125]), .rectangle2_width(rectangle2_widths[1125]), .rectangle2_height(rectangle2_heights[1125]), .rectangle2_weight(rectangle2_weights[1125]), .rectangle3_x(rectangle3_xs[1125]), .rectangle3_y(rectangle3_ys[1125]), .rectangle3_width(rectangle3_widths[1125]), .rectangle3_height(rectangle3_heights[1125]), .rectangle3_weight(rectangle3_weights[1125]), .feature_threshold(feature_thresholds[1125]), .feature_above(feature_aboves[1125]), .feature_below(feature_belows[1125]), .scan_win_std_dev(scan_win_std_dev[1125]), .feature_accum(feature_accums[1125]));
  accum_calculator ac1126(.scan_win(scan_win1126), .rectangle1_x(rectangle1_xs[1126]), .rectangle1_y(rectangle1_ys[1126]), .rectangle1_width(rectangle1_widths[1126]), .rectangle1_height(rectangle1_heights[1126]), .rectangle1_weight(rectangle1_weights[1126]), .rectangle2_x(rectangle2_xs[1126]), .rectangle2_y(rectangle2_ys[1126]), .rectangle2_width(rectangle2_widths[1126]), .rectangle2_height(rectangle2_heights[1126]), .rectangle2_weight(rectangle2_weights[1126]), .rectangle3_x(rectangle3_xs[1126]), .rectangle3_y(rectangle3_ys[1126]), .rectangle3_width(rectangle3_widths[1126]), .rectangle3_height(rectangle3_heights[1126]), .rectangle3_weight(rectangle3_weights[1126]), .feature_threshold(feature_thresholds[1126]), .feature_above(feature_aboves[1126]), .feature_below(feature_belows[1126]), .scan_win_std_dev(scan_win_std_dev[1126]), .feature_accum(feature_accums[1126]));
  accum_calculator ac1127(.scan_win(scan_win1127), .rectangle1_x(rectangle1_xs[1127]), .rectangle1_y(rectangle1_ys[1127]), .rectangle1_width(rectangle1_widths[1127]), .rectangle1_height(rectangle1_heights[1127]), .rectangle1_weight(rectangle1_weights[1127]), .rectangle2_x(rectangle2_xs[1127]), .rectangle2_y(rectangle2_ys[1127]), .rectangle2_width(rectangle2_widths[1127]), .rectangle2_height(rectangle2_heights[1127]), .rectangle2_weight(rectangle2_weights[1127]), .rectangle3_x(rectangle3_xs[1127]), .rectangle3_y(rectangle3_ys[1127]), .rectangle3_width(rectangle3_widths[1127]), .rectangle3_height(rectangle3_heights[1127]), .rectangle3_weight(rectangle3_weights[1127]), .feature_threshold(feature_thresholds[1127]), .feature_above(feature_aboves[1127]), .feature_below(feature_belows[1127]), .scan_win_std_dev(scan_win_std_dev[1127]), .feature_accum(feature_accums[1127]));
  accum_calculator ac1128(.scan_win(scan_win1128), .rectangle1_x(rectangle1_xs[1128]), .rectangle1_y(rectangle1_ys[1128]), .rectangle1_width(rectangle1_widths[1128]), .rectangle1_height(rectangle1_heights[1128]), .rectangle1_weight(rectangle1_weights[1128]), .rectangle2_x(rectangle2_xs[1128]), .rectangle2_y(rectangle2_ys[1128]), .rectangle2_width(rectangle2_widths[1128]), .rectangle2_height(rectangle2_heights[1128]), .rectangle2_weight(rectangle2_weights[1128]), .rectangle3_x(rectangle3_xs[1128]), .rectangle3_y(rectangle3_ys[1128]), .rectangle3_width(rectangle3_widths[1128]), .rectangle3_height(rectangle3_heights[1128]), .rectangle3_weight(rectangle3_weights[1128]), .feature_threshold(feature_thresholds[1128]), .feature_above(feature_aboves[1128]), .feature_below(feature_belows[1128]), .scan_win_std_dev(scan_win_std_dev[1128]), .feature_accum(feature_accums[1128]));
  accum_calculator ac1129(.scan_win(scan_win1129), .rectangle1_x(rectangle1_xs[1129]), .rectangle1_y(rectangle1_ys[1129]), .rectangle1_width(rectangle1_widths[1129]), .rectangle1_height(rectangle1_heights[1129]), .rectangle1_weight(rectangle1_weights[1129]), .rectangle2_x(rectangle2_xs[1129]), .rectangle2_y(rectangle2_ys[1129]), .rectangle2_width(rectangle2_widths[1129]), .rectangle2_height(rectangle2_heights[1129]), .rectangle2_weight(rectangle2_weights[1129]), .rectangle3_x(rectangle3_xs[1129]), .rectangle3_y(rectangle3_ys[1129]), .rectangle3_width(rectangle3_widths[1129]), .rectangle3_height(rectangle3_heights[1129]), .rectangle3_weight(rectangle3_weights[1129]), .feature_threshold(feature_thresholds[1129]), .feature_above(feature_aboves[1129]), .feature_below(feature_belows[1129]), .scan_win_std_dev(scan_win_std_dev[1129]), .feature_accum(feature_accums[1129]));
  accum_calculator ac1130(.scan_win(scan_win1130), .rectangle1_x(rectangle1_xs[1130]), .rectangle1_y(rectangle1_ys[1130]), .rectangle1_width(rectangle1_widths[1130]), .rectangle1_height(rectangle1_heights[1130]), .rectangle1_weight(rectangle1_weights[1130]), .rectangle2_x(rectangle2_xs[1130]), .rectangle2_y(rectangle2_ys[1130]), .rectangle2_width(rectangle2_widths[1130]), .rectangle2_height(rectangle2_heights[1130]), .rectangle2_weight(rectangle2_weights[1130]), .rectangle3_x(rectangle3_xs[1130]), .rectangle3_y(rectangle3_ys[1130]), .rectangle3_width(rectangle3_widths[1130]), .rectangle3_height(rectangle3_heights[1130]), .rectangle3_weight(rectangle3_weights[1130]), .feature_threshold(feature_thresholds[1130]), .feature_above(feature_aboves[1130]), .feature_below(feature_belows[1130]), .scan_win_std_dev(scan_win_std_dev[1130]), .feature_accum(feature_accums[1130]));
  accum_calculator ac1131(.scan_win(scan_win1131), .rectangle1_x(rectangle1_xs[1131]), .rectangle1_y(rectangle1_ys[1131]), .rectangle1_width(rectangle1_widths[1131]), .rectangle1_height(rectangle1_heights[1131]), .rectangle1_weight(rectangle1_weights[1131]), .rectangle2_x(rectangle2_xs[1131]), .rectangle2_y(rectangle2_ys[1131]), .rectangle2_width(rectangle2_widths[1131]), .rectangle2_height(rectangle2_heights[1131]), .rectangle2_weight(rectangle2_weights[1131]), .rectangle3_x(rectangle3_xs[1131]), .rectangle3_y(rectangle3_ys[1131]), .rectangle3_width(rectangle3_widths[1131]), .rectangle3_height(rectangle3_heights[1131]), .rectangle3_weight(rectangle3_weights[1131]), .feature_threshold(feature_thresholds[1131]), .feature_above(feature_aboves[1131]), .feature_below(feature_belows[1131]), .scan_win_std_dev(scan_win_std_dev[1131]), .feature_accum(feature_accums[1131]));
  accum_calculator ac1132(.scan_win(scan_win1132), .rectangle1_x(rectangle1_xs[1132]), .rectangle1_y(rectangle1_ys[1132]), .rectangle1_width(rectangle1_widths[1132]), .rectangle1_height(rectangle1_heights[1132]), .rectangle1_weight(rectangle1_weights[1132]), .rectangle2_x(rectangle2_xs[1132]), .rectangle2_y(rectangle2_ys[1132]), .rectangle2_width(rectangle2_widths[1132]), .rectangle2_height(rectangle2_heights[1132]), .rectangle2_weight(rectangle2_weights[1132]), .rectangle3_x(rectangle3_xs[1132]), .rectangle3_y(rectangle3_ys[1132]), .rectangle3_width(rectangle3_widths[1132]), .rectangle3_height(rectangle3_heights[1132]), .rectangle3_weight(rectangle3_weights[1132]), .feature_threshold(feature_thresholds[1132]), .feature_above(feature_aboves[1132]), .feature_below(feature_belows[1132]), .scan_win_std_dev(scan_win_std_dev[1132]), .feature_accum(feature_accums[1132]));
  accum_calculator ac1133(.scan_win(scan_win1133), .rectangle1_x(rectangle1_xs[1133]), .rectangle1_y(rectangle1_ys[1133]), .rectangle1_width(rectangle1_widths[1133]), .rectangle1_height(rectangle1_heights[1133]), .rectangle1_weight(rectangle1_weights[1133]), .rectangle2_x(rectangle2_xs[1133]), .rectangle2_y(rectangle2_ys[1133]), .rectangle2_width(rectangle2_widths[1133]), .rectangle2_height(rectangle2_heights[1133]), .rectangle2_weight(rectangle2_weights[1133]), .rectangle3_x(rectangle3_xs[1133]), .rectangle3_y(rectangle3_ys[1133]), .rectangle3_width(rectangle3_widths[1133]), .rectangle3_height(rectangle3_heights[1133]), .rectangle3_weight(rectangle3_weights[1133]), .feature_threshold(feature_thresholds[1133]), .feature_above(feature_aboves[1133]), .feature_below(feature_belows[1133]), .scan_win_std_dev(scan_win_std_dev[1133]), .feature_accum(feature_accums[1133]));
  accum_calculator ac1134(.scan_win(scan_win1134), .rectangle1_x(rectangle1_xs[1134]), .rectangle1_y(rectangle1_ys[1134]), .rectangle1_width(rectangle1_widths[1134]), .rectangle1_height(rectangle1_heights[1134]), .rectangle1_weight(rectangle1_weights[1134]), .rectangle2_x(rectangle2_xs[1134]), .rectangle2_y(rectangle2_ys[1134]), .rectangle2_width(rectangle2_widths[1134]), .rectangle2_height(rectangle2_heights[1134]), .rectangle2_weight(rectangle2_weights[1134]), .rectangle3_x(rectangle3_xs[1134]), .rectangle3_y(rectangle3_ys[1134]), .rectangle3_width(rectangle3_widths[1134]), .rectangle3_height(rectangle3_heights[1134]), .rectangle3_weight(rectangle3_weights[1134]), .feature_threshold(feature_thresholds[1134]), .feature_above(feature_aboves[1134]), .feature_below(feature_belows[1134]), .scan_win_std_dev(scan_win_std_dev[1134]), .feature_accum(feature_accums[1134]));
  accum_calculator ac1135(.scan_win(scan_win1135), .rectangle1_x(rectangle1_xs[1135]), .rectangle1_y(rectangle1_ys[1135]), .rectangle1_width(rectangle1_widths[1135]), .rectangle1_height(rectangle1_heights[1135]), .rectangle1_weight(rectangle1_weights[1135]), .rectangle2_x(rectangle2_xs[1135]), .rectangle2_y(rectangle2_ys[1135]), .rectangle2_width(rectangle2_widths[1135]), .rectangle2_height(rectangle2_heights[1135]), .rectangle2_weight(rectangle2_weights[1135]), .rectangle3_x(rectangle3_xs[1135]), .rectangle3_y(rectangle3_ys[1135]), .rectangle3_width(rectangle3_widths[1135]), .rectangle3_height(rectangle3_heights[1135]), .rectangle3_weight(rectangle3_weights[1135]), .feature_threshold(feature_thresholds[1135]), .feature_above(feature_aboves[1135]), .feature_below(feature_belows[1135]), .scan_win_std_dev(scan_win_std_dev[1135]), .feature_accum(feature_accums[1135]));
  accum_calculator ac1136(.scan_win(scan_win1136), .rectangle1_x(rectangle1_xs[1136]), .rectangle1_y(rectangle1_ys[1136]), .rectangle1_width(rectangle1_widths[1136]), .rectangle1_height(rectangle1_heights[1136]), .rectangle1_weight(rectangle1_weights[1136]), .rectangle2_x(rectangle2_xs[1136]), .rectangle2_y(rectangle2_ys[1136]), .rectangle2_width(rectangle2_widths[1136]), .rectangle2_height(rectangle2_heights[1136]), .rectangle2_weight(rectangle2_weights[1136]), .rectangle3_x(rectangle3_xs[1136]), .rectangle3_y(rectangle3_ys[1136]), .rectangle3_width(rectangle3_widths[1136]), .rectangle3_height(rectangle3_heights[1136]), .rectangle3_weight(rectangle3_weights[1136]), .feature_threshold(feature_thresholds[1136]), .feature_above(feature_aboves[1136]), .feature_below(feature_belows[1136]), .scan_win_std_dev(scan_win_std_dev[1136]), .feature_accum(feature_accums[1136]));
  accum_calculator ac1137(.scan_win(scan_win1137), .rectangle1_x(rectangle1_xs[1137]), .rectangle1_y(rectangle1_ys[1137]), .rectangle1_width(rectangle1_widths[1137]), .rectangle1_height(rectangle1_heights[1137]), .rectangle1_weight(rectangle1_weights[1137]), .rectangle2_x(rectangle2_xs[1137]), .rectangle2_y(rectangle2_ys[1137]), .rectangle2_width(rectangle2_widths[1137]), .rectangle2_height(rectangle2_heights[1137]), .rectangle2_weight(rectangle2_weights[1137]), .rectangle3_x(rectangle3_xs[1137]), .rectangle3_y(rectangle3_ys[1137]), .rectangle3_width(rectangle3_widths[1137]), .rectangle3_height(rectangle3_heights[1137]), .rectangle3_weight(rectangle3_weights[1137]), .feature_threshold(feature_thresholds[1137]), .feature_above(feature_aboves[1137]), .feature_below(feature_belows[1137]), .scan_win_std_dev(scan_win_std_dev[1137]), .feature_accum(feature_accums[1137]));
  accum_calculator ac1138(.scan_win(scan_win1138), .rectangle1_x(rectangle1_xs[1138]), .rectangle1_y(rectangle1_ys[1138]), .rectangle1_width(rectangle1_widths[1138]), .rectangle1_height(rectangle1_heights[1138]), .rectangle1_weight(rectangle1_weights[1138]), .rectangle2_x(rectangle2_xs[1138]), .rectangle2_y(rectangle2_ys[1138]), .rectangle2_width(rectangle2_widths[1138]), .rectangle2_height(rectangle2_heights[1138]), .rectangle2_weight(rectangle2_weights[1138]), .rectangle3_x(rectangle3_xs[1138]), .rectangle3_y(rectangle3_ys[1138]), .rectangle3_width(rectangle3_widths[1138]), .rectangle3_height(rectangle3_heights[1138]), .rectangle3_weight(rectangle3_weights[1138]), .feature_threshold(feature_thresholds[1138]), .feature_above(feature_aboves[1138]), .feature_below(feature_belows[1138]), .scan_win_std_dev(scan_win_std_dev[1138]), .feature_accum(feature_accums[1138]));
  accum_calculator ac1139(.scan_win(scan_win1139), .rectangle1_x(rectangle1_xs[1139]), .rectangle1_y(rectangle1_ys[1139]), .rectangle1_width(rectangle1_widths[1139]), .rectangle1_height(rectangle1_heights[1139]), .rectangle1_weight(rectangle1_weights[1139]), .rectangle2_x(rectangle2_xs[1139]), .rectangle2_y(rectangle2_ys[1139]), .rectangle2_width(rectangle2_widths[1139]), .rectangle2_height(rectangle2_heights[1139]), .rectangle2_weight(rectangle2_weights[1139]), .rectangle3_x(rectangle3_xs[1139]), .rectangle3_y(rectangle3_ys[1139]), .rectangle3_width(rectangle3_widths[1139]), .rectangle3_height(rectangle3_heights[1139]), .rectangle3_weight(rectangle3_weights[1139]), .feature_threshold(feature_thresholds[1139]), .feature_above(feature_aboves[1139]), .feature_below(feature_belows[1139]), .scan_win_std_dev(scan_win_std_dev[1139]), .feature_accum(feature_accums[1139]));
  accum_calculator ac1140(.scan_win(scan_win1140), .rectangle1_x(rectangle1_xs[1140]), .rectangle1_y(rectangle1_ys[1140]), .rectangle1_width(rectangle1_widths[1140]), .rectangle1_height(rectangle1_heights[1140]), .rectangle1_weight(rectangle1_weights[1140]), .rectangle2_x(rectangle2_xs[1140]), .rectangle2_y(rectangle2_ys[1140]), .rectangle2_width(rectangle2_widths[1140]), .rectangle2_height(rectangle2_heights[1140]), .rectangle2_weight(rectangle2_weights[1140]), .rectangle3_x(rectangle3_xs[1140]), .rectangle3_y(rectangle3_ys[1140]), .rectangle3_width(rectangle3_widths[1140]), .rectangle3_height(rectangle3_heights[1140]), .rectangle3_weight(rectangle3_weights[1140]), .feature_threshold(feature_thresholds[1140]), .feature_above(feature_aboves[1140]), .feature_below(feature_belows[1140]), .scan_win_std_dev(scan_win_std_dev[1140]), .feature_accum(feature_accums[1140]));
  accum_calculator ac1141(.scan_win(scan_win1141), .rectangle1_x(rectangle1_xs[1141]), .rectangle1_y(rectangle1_ys[1141]), .rectangle1_width(rectangle1_widths[1141]), .rectangle1_height(rectangle1_heights[1141]), .rectangle1_weight(rectangle1_weights[1141]), .rectangle2_x(rectangle2_xs[1141]), .rectangle2_y(rectangle2_ys[1141]), .rectangle2_width(rectangle2_widths[1141]), .rectangle2_height(rectangle2_heights[1141]), .rectangle2_weight(rectangle2_weights[1141]), .rectangle3_x(rectangle3_xs[1141]), .rectangle3_y(rectangle3_ys[1141]), .rectangle3_width(rectangle3_widths[1141]), .rectangle3_height(rectangle3_heights[1141]), .rectangle3_weight(rectangle3_weights[1141]), .feature_threshold(feature_thresholds[1141]), .feature_above(feature_aboves[1141]), .feature_below(feature_belows[1141]), .scan_win_std_dev(scan_win_std_dev[1141]), .feature_accum(feature_accums[1141]));
  accum_calculator ac1142(.scan_win(scan_win1142), .rectangle1_x(rectangle1_xs[1142]), .rectangle1_y(rectangle1_ys[1142]), .rectangle1_width(rectangle1_widths[1142]), .rectangle1_height(rectangle1_heights[1142]), .rectangle1_weight(rectangle1_weights[1142]), .rectangle2_x(rectangle2_xs[1142]), .rectangle2_y(rectangle2_ys[1142]), .rectangle2_width(rectangle2_widths[1142]), .rectangle2_height(rectangle2_heights[1142]), .rectangle2_weight(rectangle2_weights[1142]), .rectangle3_x(rectangle3_xs[1142]), .rectangle3_y(rectangle3_ys[1142]), .rectangle3_width(rectangle3_widths[1142]), .rectangle3_height(rectangle3_heights[1142]), .rectangle3_weight(rectangle3_weights[1142]), .feature_threshold(feature_thresholds[1142]), .feature_above(feature_aboves[1142]), .feature_below(feature_belows[1142]), .scan_win_std_dev(scan_win_std_dev[1142]), .feature_accum(feature_accums[1142]));
  accum_calculator ac1143(.scan_win(scan_win1143), .rectangle1_x(rectangle1_xs[1143]), .rectangle1_y(rectangle1_ys[1143]), .rectangle1_width(rectangle1_widths[1143]), .rectangle1_height(rectangle1_heights[1143]), .rectangle1_weight(rectangle1_weights[1143]), .rectangle2_x(rectangle2_xs[1143]), .rectangle2_y(rectangle2_ys[1143]), .rectangle2_width(rectangle2_widths[1143]), .rectangle2_height(rectangle2_heights[1143]), .rectangle2_weight(rectangle2_weights[1143]), .rectangle3_x(rectangle3_xs[1143]), .rectangle3_y(rectangle3_ys[1143]), .rectangle3_width(rectangle3_widths[1143]), .rectangle3_height(rectangle3_heights[1143]), .rectangle3_weight(rectangle3_weights[1143]), .feature_threshold(feature_thresholds[1143]), .feature_above(feature_aboves[1143]), .feature_below(feature_belows[1143]), .scan_win_std_dev(scan_win_std_dev[1143]), .feature_accum(feature_accums[1143]));
  accum_calculator ac1144(.scan_win(scan_win1144), .rectangle1_x(rectangle1_xs[1144]), .rectangle1_y(rectangle1_ys[1144]), .rectangle1_width(rectangle1_widths[1144]), .rectangle1_height(rectangle1_heights[1144]), .rectangle1_weight(rectangle1_weights[1144]), .rectangle2_x(rectangle2_xs[1144]), .rectangle2_y(rectangle2_ys[1144]), .rectangle2_width(rectangle2_widths[1144]), .rectangle2_height(rectangle2_heights[1144]), .rectangle2_weight(rectangle2_weights[1144]), .rectangle3_x(rectangle3_xs[1144]), .rectangle3_y(rectangle3_ys[1144]), .rectangle3_width(rectangle3_widths[1144]), .rectangle3_height(rectangle3_heights[1144]), .rectangle3_weight(rectangle3_weights[1144]), .feature_threshold(feature_thresholds[1144]), .feature_above(feature_aboves[1144]), .feature_below(feature_belows[1144]), .scan_win_std_dev(scan_win_std_dev[1144]), .feature_accum(feature_accums[1144]));
  accum_calculator ac1145(.scan_win(scan_win1145), .rectangle1_x(rectangle1_xs[1145]), .rectangle1_y(rectangle1_ys[1145]), .rectangle1_width(rectangle1_widths[1145]), .rectangle1_height(rectangle1_heights[1145]), .rectangle1_weight(rectangle1_weights[1145]), .rectangle2_x(rectangle2_xs[1145]), .rectangle2_y(rectangle2_ys[1145]), .rectangle2_width(rectangle2_widths[1145]), .rectangle2_height(rectangle2_heights[1145]), .rectangle2_weight(rectangle2_weights[1145]), .rectangle3_x(rectangle3_xs[1145]), .rectangle3_y(rectangle3_ys[1145]), .rectangle3_width(rectangle3_widths[1145]), .rectangle3_height(rectangle3_heights[1145]), .rectangle3_weight(rectangle3_weights[1145]), .feature_threshold(feature_thresholds[1145]), .feature_above(feature_aboves[1145]), .feature_below(feature_belows[1145]), .scan_win_std_dev(scan_win_std_dev[1145]), .feature_accum(feature_accums[1145]));
  accum_calculator ac1146(.scan_win(scan_win1146), .rectangle1_x(rectangle1_xs[1146]), .rectangle1_y(rectangle1_ys[1146]), .rectangle1_width(rectangle1_widths[1146]), .rectangle1_height(rectangle1_heights[1146]), .rectangle1_weight(rectangle1_weights[1146]), .rectangle2_x(rectangle2_xs[1146]), .rectangle2_y(rectangle2_ys[1146]), .rectangle2_width(rectangle2_widths[1146]), .rectangle2_height(rectangle2_heights[1146]), .rectangle2_weight(rectangle2_weights[1146]), .rectangle3_x(rectangle3_xs[1146]), .rectangle3_y(rectangle3_ys[1146]), .rectangle3_width(rectangle3_widths[1146]), .rectangle3_height(rectangle3_heights[1146]), .rectangle3_weight(rectangle3_weights[1146]), .feature_threshold(feature_thresholds[1146]), .feature_above(feature_aboves[1146]), .feature_below(feature_belows[1146]), .scan_win_std_dev(scan_win_std_dev[1146]), .feature_accum(feature_accums[1146]));
  accum_calculator ac1147(.scan_win(scan_win1147), .rectangle1_x(rectangle1_xs[1147]), .rectangle1_y(rectangle1_ys[1147]), .rectangle1_width(rectangle1_widths[1147]), .rectangle1_height(rectangle1_heights[1147]), .rectangle1_weight(rectangle1_weights[1147]), .rectangle2_x(rectangle2_xs[1147]), .rectangle2_y(rectangle2_ys[1147]), .rectangle2_width(rectangle2_widths[1147]), .rectangle2_height(rectangle2_heights[1147]), .rectangle2_weight(rectangle2_weights[1147]), .rectangle3_x(rectangle3_xs[1147]), .rectangle3_y(rectangle3_ys[1147]), .rectangle3_width(rectangle3_widths[1147]), .rectangle3_height(rectangle3_heights[1147]), .rectangle3_weight(rectangle3_weights[1147]), .feature_threshold(feature_thresholds[1147]), .feature_above(feature_aboves[1147]), .feature_below(feature_belows[1147]), .scan_win_std_dev(scan_win_std_dev[1147]), .feature_accum(feature_accums[1147]));
  accum_calculator ac1148(.scan_win(scan_win1148), .rectangle1_x(rectangle1_xs[1148]), .rectangle1_y(rectangle1_ys[1148]), .rectangle1_width(rectangle1_widths[1148]), .rectangle1_height(rectangle1_heights[1148]), .rectangle1_weight(rectangle1_weights[1148]), .rectangle2_x(rectangle2_xs[1148]), .rectangle2_y(rectangle2_ys[1148]), .rectangle2_width(rectangle2_widths[1148]), .rectangle2_height(rectangle2_heights[1148]), .rectangle2_weight(rectangle2_weights[1148]), .rectangle3_x(rectangle3_xs[1148]), .rectangle3_y(rectangle3_ys[1148]), .rectangle3_width(rectangle3_widths[1148]), .rectangle3_height(rectangle3_heights[1148]), .rectangle3_weight(rectangle3_weights[1148]), .feature_threshold(feature_thresholds[1148]), .feature_above(feature_aboves[1148]), .feature_below(feature_belows[1148]), .scan_win_std_dev(scan_win_std_dev[1148]), .feature_accum(feature_accums[1148]));
  accum_calculator ac1149(.scan_win(scan_win1149), .rectangle1_x(rectangle1_xs[1149]), .rectangle1_y(rectangle1_ys[1149]), .rectangle1_width(rectangle1_widths[1149]), .rectangle1_height(rectangle1_heights[1149]), .rectangle1_weight(rectangle1_weights[1149]), .rectangle2_x(rectangle2_xs[1149]), .rectangle2_y(rectangle2_ys[1149]), .rectangle2_width(rectangle2_widths[1149]), .rectangle2_height(rectangle2_heights[1149]), .rectangle2_weight(rectangle2_weights[1149]), .rectangle3_x(rectangle3_xs[1149]), .rectangle3_y(rectangle3_ys[1149]), .rectangle3_width(rectangle3_widths[1149]), .rectangle3_height(rectangle3_heights[1149]), .rectangle3_weight(rectangle3_weights[1149]), .feature_threshold(feature_thresholds[1149]), .feature_above(feature_aboves[1149]), .feature_below(feature_belows[1149]), .scan_win_std_dev(scan_win_std_dev[1149]), .feature_accum(feature_accums[1149]));
  accum_calculator ac1150(.scan_win(scan_win1150), .rectangle1_x(rectangle1_xs[1150]), .rectangle1_y(rectangle1_ys[1150]), .rectangle1_width(rectangle1_widths[1150]), .rectangle1_height(rectangle1_heights[1150]), .rectangle1_weight(rectangle1_weights[1150]), .rectangle2_x(rectangle2_xs[1150]), .rectangle2_y(rectangle2_ys[1150]), .rectangle2_width(rectangle2_widths[1150]), .rectangle2_height(rectangle2_heights[1150]), .rectangle2_weight(rectangle2_weights[1150]), .rectangle3_x(rectangle3_xs[1150]), .rectangle3_y(rectangle3_ys[1150]), .rectangle3_width(rectangle3_widths[1150]), .rectangle3_height(rectangle3_heights[1150]), .rectangle3_weight(rectangle3_weights[1150]), .feature_threshold(feature_thresholds[1150]), .feature_above(feature_aboves[1150]), .feature_below(feature_belows[1150]), .scan_win_std_dev(scan_win_std_dev[1150]), .feature_accum(feature_accums[1150]));
  accum_calculator ac1151(.scan_win(scan_win1151), .rectangle1_x(rectangle1_xs[1151]), .rectangle1_y(rectangle1_ys[1151]), .rectangle1_width(rectangle1_widths[1151]), .rectangle1_height(rectangle1_heights[1151]), .rectangle1_weight(rectangle1_weights[1151]), .rectangle2_x(rectangle2_xs[1151]), .rectangle2_y(rectangle2_ys[1151]), .rectangle2_width(rectangle2_widths[1151]), .rectangle2_height(rectangle2_heights[1151]), .rectangle2_weight(rectangle2_weights[1151]), .rectangle3_x(rectangle3_xs[1151]), .rectangle3_y(rectangle3_ys[1151]), .rectangle3_width(rectangle3_widths[1151]), .rectangle3_height(rectangle3_heights[1151]), .rectangle3_weight(rectangle3_weights[1151]), .feature_threshold(feature_thresholds[1151]), .feature_above(feature_aboves[1151]), .feature_below(feature_belows[1151]), .scan_win_std_dev(scan_win_std_dev[1151]), .feature_accum(feature_accums[1151]));
  accum_calculator ac1152(.scan_win(scan_win1152), .rectangle1_x(rectangle1_xs[1152]), .rectangle1_y(rectangle1_ys[1152]), .rectangle1_width(rectangle1_widths[1152]), .rectangle1_height(rectangle1_heights[1152]), .rectangle1_weight(rectangle1_weights[1152]), .rectangle2_x(rectangle2_xs[1152]), .rectangle2_y(rectangle2_ys[1152]), .rectangle2_width(rectangle2_widths[1152]), .rectangle2_height(rectangle2_heights[1152]), .rectangle2_weight(rectangle2_weights[1152]), .rectangle3_x(rectangle3_xs[1152]), .rectangle3_y(rectangle3_ys[1152]), .rectangle3_width(rectangle3_widths[1152]), .rectangle3_height(rectangle3_heights[1152]), .rectangle3_weight(rectangle3_weights[1152]), .feature_threshold(feature_thresholds[1152]), .feature_above(feature_aboves[1152]), .feature_below(feature_belows[1152]), .scan_win_std_dev(scan_win_std_dev[1152]), .feature_accum(feature_accums[1152]));
  accum_calculator ac1153(.scan_win(scan_win1153), .rectangle1_x(rectangle1_xs[1153]), .rectangle1_y(rectangle1_ys[1153]), .rectangle1_width(rectangle1_widths[1153]), .rectangle1_height(rectangle1_heights[1153]), .rectangle1_weight(rectangle1_weights[1153]), .rectangle2_x(rectangle2_xs[1153]), .rectangle2_y(rectangle2_ys[1153]), .rectangle2_width(rectangle2_widths[1153]), .rectangle2_height(rectangle2_heights[1153]), .rectangle2_weight(rectangle2_weights[1153]), .rectangle3_x(rectangle3_xs[1153]), .rectangle3_y(rectangle3_ys[1153]), .rectangle3_width(rectangle3_widths[1153]), .rectangle3_height(rectangle3_heights[1153]), .rectangle3_weight(rectangle3_weights[1153]), .feature_threshold(feature_thresholds[1153]), .feature_above(feature_aboves[1153]), .feature_below(feature_belows[1153]), .scan_win_std_dev(scan_win_std_dev[1153]), .feature_accum(feature_accums[1153]));
  accum_calculator ac1154(.scan_win(scan_win1154), .rectangle1_x(rectangle1_xs[1154]), .rectangle1_y(rectangle1_ys[1154]), .rectangle1_width(rectangle1_widths[1154]), .rectangle1_height(rectangle1_heights[1154]), .rectangle1_weight(rectangle1_weights[1154]), .rectangle2_x(rectangle2_xs[1154]), .rectangle2_y(rectangle2_ys[1154]), .rectangle2_width(rectangle2_widths[1154]), .rectangle2_height(rectangle2_heights[1154]), .rectangle2_weight(rectangle2_weights[1154]), .rectangle3_x(rectangle3_xs[1154]), .rectangle3_y(rectangle3_ys[1154]), .rectangle3_width(rectangle3_widths[1154]), .rectangle3_height(rectangle3_heights[1154]), .rectangle3_weight(rectangle3_weights[1154]), .feature_threshold(feature_thresholds[1154]), .feature_above(feature_aboves[1154]), .feature_below(feature_belows[1154]), .scan_win_std_dev(scan_win_std_dev[1154]), .feature_accum(feature_accums[1154]));
  accum_calculator ac1155(.scan_win(scan_win1155), .rectangle1_x(rectangle1_xs[1155]), .rectangle1_y(rectangle1_ys[1155]), .rectangle1_width(rectangle1_widths[1155]), .rectangle1_height(rectangle1_heights[1155]), .rectangle1_weight(rectangle1_weights[1155]), .rectangle2_x(rectangle2_xs[1155]), .rectangle2_y(rectangle2_ys[1155]), .rectangle2_width(rectangle2_widths[1155]), .rectangle2_height(rectangle2_heights[1155]), .rectangle2_weight(rectangle2_weights[1155]), .rectangle3_x(rectangle3_xs[1155]), .rectangle3_y(rectangle3_ys[1155]), .rectangle3_width(rectangle3_widths[1155]), .rectangle3_height(rectangle3_heights[1155]), .rectangle3_weight(rectangle3_weights[1155]), .feature_threshold(feature_thresholds[1155]), .feature_above(feature_aboves[1155]), .feature_below(feature_belows[1155]), .scan_win_std_dev(scan_win_std_dev[1155]), .feature_accum(feature_accums[1155]));
  accum_calculator ac1156(.scan_win(scan_win1156), .rectangle1_x(rectangle1_xs[1156]), .rectangle1_y(rectangle1_ys[1156]), .rectangle1_width(rectangle1_widths[1156]), .rectangle1_height(rectangle1_heights[1156]), .rectangle1_weight(rectangle1_weights[1156]), .rectangle2_x(rectangle2_xs[1156]), .rectangle2_y(rectangle2_ys[1156]), .rectangle2_width(rectangle2_widths[1156]), .rectangle2_height(rectangle2_heights[1156]), .rectangle2_weight(rectangle2_weights[1156]), .rectangle3_x(rectangle3_xs[1156]), .rectangle3_y(rectangle3_ys[1156]), .rectangle3_width(rectangle3_widths[1156]), .rectangle3_height(rectangle3_heights[1156]), .rectangle3_weight(rectangle3_weights[1156]), .feature_threshold(feature_thresholds[1156]), .feature_above(feature_aboves[1156]), .feature_below(feature_belows[1156]), .scan_win_std_dev(scan_win_std_dev[1156]), .feature_accum(feature_accums[1156]));
  accum_calculator ac1157(.scan_win(scan_win1157), .rectangle1_x(rectangle1_xs[1157]), .rectangle1_y(rectangle1_ys[1157]), .rectangle1_width(rectangle1_widths[1157]), .rectangle1_height(rectangle1_heights[1157]), .rectangle1_weight(rectangle1_weights[1157]), .rectangle2_x(rectangle2_xs[1157]), .rectangle2_y(rectangle2_ys[1157]), .rectangle2_width(rectangle2_widths[1157]), .rectangle2_height(rectangle2_heights[1157]), .rectangle2_weight(rectangle2_weights[1157]), .rectangle3_x(rectangle3_xs[1157]), .rectangle3_y(rectangle3_ys[1157]), .rectangle3_width(rectangle3_widths[1157]), .rectangle3_height(rectangle3_heights[1157]), .rectangle3_weight(rectangle3_weights[1157]), .feature_threshold(feature_thresholds[1157]), .feature_above(feature_aboves[1157]), .feature_below(feature_belows[1157]), .scan_win_std_dev(scan_win_std_dev[1157]), .feature_accum(feature_accums[1157]));
  accum_calculator ac1158(.scan_win(scan_win1158), .rectangle1_x(rectangle1_xs[1158]), .rectangle1_y(rectangle1_ys[1158]), .rectangle1_width(rectangle1_widths[1158]), .rectangle1_height(rectangle1_heights[1158]), .rectangle1_weight(rectangle1_weights[1158]), .rectangle2_x(rectangle2_xs[1158]), .rectangle2_y(rectangle2_ys[1158]), .rectangle2_width(rectangle2_widths[1158]), .rectangle2_height(rectangle2_heights[1158]), .rectangle2_weight(rectangle2_weights[1158]), .rectangle3_x(rectangle3_xs[1158]), .rectangle3_y(rectangle3_ys[1158]), .rectangle3_width(rectangle3_widths[1158]), .rectangle3_height(rectangle3_heights[1158]), .rectangle3_weight(rectangle3_weights[1158]), .feature_threshold(feature_thresholds[1158]), .feature_above(feature_aboves[1158]), .feature_below(feature_belows[1158]), .scan_win_std_dev(scan_win_std_dev[1158]), .feature_accum(feature_accums[1158]));
  accum_calculator ac1159(.scan_win(scan_win1159), .rectangle1_x(rectangle1_xs[1159]), .rectangle1_y(rectangle1_ys[1159]), .rectangle1_width(rectangle1_widths[1159]), .rectangle1_height(rectangle1_heights[1159]), .rectangle1_weight(rectangle1_weights[1159]), .rectangle2_x(rectangle2_xs[1159]), .rectangle2_y(rectangle2_ys[1159]), .rectangle2_width(rectangle2_widths[1159]), .rectangle2_height(rectangle2_heights[1159]), .rectangle2_weight(rectangle2_weights[1159]), .rectangle3_x(rectangle3_xs[1159]), .rectangle3_y(rectangle3_ys[1159]), .rectangle3_width(rectangle3_widths[1159]), .rectangle3_height(rectangle3_heights[1159]), .rectangle3_weight(rectangle3_weights[1159]), .feature_threshold(feature_thresholds[1159]), .feature_above(feature_aboves[1159]), .feature_below(feature_belows[1159]), .scan_win_std_dev(scan_win_std_dev[1159]), .feature_accum(feature_accums[1159]));
  accum_calculator ac1160(.scan_win(scan_win1160), .rectangle1_x(rectangle1_xs[1160]), .rectangle1_y(rectangle1_ys[1160]), .rectangle1_width(rectangle1_widths[1160]), .rectangle1_height(rectangle1_heights[1160]), .rectangle1_weight(rectangle1_weights[1160]), .rectangle2_x(rectangle2_xs[1160]), .rectangle2_y(rectangle2_ys[1160]), .rectangle2_width(rectangle2_widths[1160]), .rectangle2_height(rectangle2_heights[1160]), .rectangle2_weight(rectangle2_weights[1160]), .rectangle3_x(rectangle3_xs[1160]), .rectangle3_y(rectangle3_ys[1160]), .rectangle3_width(rectangle3_widths[1160]), .rectangle3_height(rectangle3_heights[1160]), .rectangle3_weight(rectangle3_weights[1160]), .feature_threshold(feature_thresholds[1160]), .feature_above(feature_aboves[1160]), .feature_below(feature_belows[1160]), .scan_win_std_dev(scan_win_std_dev[1160]), .feature_accum(feature_accums[1160]));
  accum_calculator ac1161(.scan_win(scan_win1161), .rectangle1_x(rectangle1_xs[1161]), .rectangle1_y(rectangle1_ys[1161]), .rectangle1_width(rectangle1_widths[1161]), .rectangle1_height(rectangle1_heights[1161]), .rectangle1_weight(rectangle1_weights[1161]), .rectangle2_x(rectangle2_xs[1161]), .rectangle2_y(rectangle2_ys[1161]), .rectangle2_width(rectangle2_widths[1161]), .rectangle2_height(rectangle2_heights[1161]), .rectangle2_weight(rectangle2_weights[1161]), .rectangle3_x(rectangle3_xs[1161]), .rectangle3_y(rectangle3_ys[1161]), .rectangle3_width(rectangle3_widths[1161]), .rectangle3_height(rectangle3_heights[1161]), .rectangle3_weight(rectangle3_weights[1161]), .feature_threshold(feature_thresholds[1161]), .feature_above(feature_aboves[1161]), .feature_below(feature_belows[1161]), .scan_win_std_dev(scan_win_std_dev[1161]), .feature_accum(feature_accums[1161]));
  accum_calculator ac1162(.scan_win(scan_win1162), .rectangle1_x(rectangle1_xs[1162]), .rectangle1_y(rectangle1_ys[1162]), .rectangle1_width(rectangle1_widths[1162]), .rectangle1_height(rectangle1_heights[1162]), .rectangle1_weight(rectangle1_weights[1162]), .rectangle2_x(rectangle2_xs[1162]), .rectangle2_y(rectangle2_ys[1162]), .rectangle2_width(rectangle2_widths[1162]), .rectangle2_height(rectangle2_heights[1162]), .rectangle2_weight(rectangle2_weights[1162]), .rectangle3_x(rectangle3_xs[1162]), .rectangle3_y(rectangle3_ys[1162]), .rectangle3_width(rectangle3_widths[1162]), .rectangle3_height(rectangle3_heights[1162]), .rectangle3_weight(rectangle3_weights[1162]), .feature_threshold(feature_thresholds[1162]), .feature_above(feature_aboves[1162]), .feature_below(feature_belows[1162]), .scan_win_std_dev(scan_win_std_dev[1162]), .feature_accum(feature_accums[1162]));
  accum_calculator ac1163(.scan_win(scan_win1163), .rectangle1_x(rectangle1_xs[1163]), .rectangle1_y(rectangle1_ys[1163]), .rectangle1_width(rectangle1_widths[1163]), .rectangle1_height(rectangle1_heights[1163]), .rectangle1_weight(rectangle1_weights[1163]), .rectangle2_x(rectangle2_xs[1163]), .rectangle2_y(rectangle2_ys[1163]), .rectangle2_width(rectangle2_widths[1163]), .rectangle2_height(rectangle2_heights[1163]), .rectangle2_weight(rectangle2_weights[1163]), .rectangle3_x(rectangle3_xs[1163]), .rectangle3_y(rectangle3_ys[1163]), .rectangle3_width(rectangle3_widths[1163]), .rectangle3_height(rectangle3_heights[1163]), .rectangle3_weight(rectangle3_weights[1163]), .feature_threshold(feature_thresholds[1163]), .feature_above(feature_aboves[1163]), .feature_below(feature_belows[1163]), .scan_win_std_dev(scan_win_std_dev[1163]), .feature_accum(feature_accums[1163]));
  accum_calculator ac1164(.scan_win(scan_win1164), .rectangle1_x(rectangle1_xs[1164]), .rectangle1_y(rectangle1_ys[1164]), .rectangle1_width(rectangle1_widths[1164]), .rectangle1_height(rectangle1_heights[1164]), .rectangle1_weight(rectangle1_weights[1164]), .rectangle2_x(rectangle2_xs[1164]), .rectangle2_y(rectangle2_ys[1164]), .rectangle2_width(rectangle2_widths[1164]), .rectangle2_height(rectangle2_heights[1164]), .rectangle2_weight(rectangle2_weights[1164]), .rectangle3_x(rectangle3_xs[1164]), .rectangle3_y(rectangle3_ys[1164]), .rectangle3_width(rectangle3_widths[1164]), .rectangle3_height(rectangle3_heights[1164]), .rectangle3_weight(rectangle3_weights[1164]), .feature_threshold(feature_thresholds[1164]), .feature_above(feature_aboves[1164]), .feature_below(feature_belows[1164]), .scan_win_std_dev(scan_win_std_dev[1164]), .feature_accum(feature_accums[1164]));
  accum_calculator ac1165(.scan_win(scan_win1165), .rectangle1_x(rectangle1_xs[1165]), .rectangle1_y(rectangle1_ys[1165]), .rectangle1_width(rectangle1_widths[1165]), .rectangle1_height(rectangle1_heights[1165]), .rectangle1_weight(rectangle1_weights[1165]), .rectangle2_x(rectangle2_xs[1165]), .rectangle2_y(rectangle2_ys[1165]), .rectangle2_width(rectangle2_widths[1165]), .rectangle2_height(rectangle2_heights[1165]), .rectangle2_weight(rectangle2_weights[1165]), .rectangle3_x(rectangle3_xs[1165]), .rectangle3_y(rectangle3_ys[1165]), .rectangle3_width(rectangle3_widths[1165]), .rectangle3_height(rectangle3_heights[1165]), .rectangle3_weight(rectangle3_weights[1165]), .feature_threshold(feature_thresholds[1165]), .feature_above(feature_aboves[1165]), .feature_below(feature_belows[1165]), .scan_win_std_dev(scan_win_std_dev[1165]), .feature_accum(feature_accums[1165]));
  accum_calculator ac1166(.scan_win(scan_win1166), .rectangle1_x(rectangle1_xs[1166]), .rectangle1_y(rectangle1_ys[1166]), .rectangle1_width(rectangle1_widths[1166]), .rectangle1_height(rectangle1_heights[1166]), .rectangle1_weight(rectangle1_weights[1166]), .rectangle2_x(rectangle2_xs[1166]), .rectangle2_y(rectangle2_ys[1166]), .rectangle2_width(rectangle2_widths[1166]), .rectangle2_height(rectangle2_heights[1166]), .rectangle2_weight(rectangle2_weights[1166]), .rectangle3_x(rectangle3_xs[1166]), .rectangle3_y(rectangle3_ys[1166]), .rectangle3_width(rectangle3_widths[1166]), .rectangle3_height(rectangle3_heights[1166]), .rectangle3_weight(rectangle3_weights[1166]), .feature_threshold(feature_thresholds[1166]), .feature_above(feature_aboves[1166]), .feature_below(feature_belows[1166]), .scan_win_std_dev(scan_win_std_dev[1166]), .feature_accum(feature_accums[1166]));
  accum_calculator ac1167(.scan_win(scan_win1167), .rectangle1_x(rectangle1_xs[1167]), .rectangle1_y(rectangle1_ys[1167]), .rectangle1_width(rectangle1_widths[1167]), .rectangle1_height(rectangle1_heights[1167]), .rectangle1_weight(rectangle1_weights[1167]), .rectangle2_x(rectangle2_xs[1167]), .rectangle2_y(rectangle2_ys[1167]), .rectangle2_width(rectangle2_widths[1167]), .rectangle2_height(rectangle2_heights[1167]), .rectangle2_weight(rectangle2_weights[1167]), .rectangle3_x(rectangle3_xs[1167]), .rectangle3_y(rectangle3_ys[1167]), .rectangle3_width(rectangle3_widths[1167]), .rectangle3_height(rectangle3_heights[1167]), .rectangle3_weight(rectangle3_weights[1167]), .feature_threshold(feature_thresholds[1167]), .feature_above(feature_aboves[1167]), .feature_below(feature_belows[1167]), .scan_win_std_dev(scan_win_std_dev[1167]), .feature_accum(feature_accums[1167]));
  accum_calculator ac1168(.scan_win(scan_win1168), .rectangle1_x(rectangle1_xs[1168]), .rectangle1_y(rectangle1_ys[1168]), .rectangle1_width(rectangle1_widths[1168]), .rectangle1_height(rectangle1_heights[1168]), .rectangle1_weight(rectangle1_weights[1168]), .rectangle2_x(rectangle2_xs[1168]), .rectangle2_y(rectangle2_ys[1168]), .rectangle2_width(rectangle2_widths[1168]), .rectangle2_height(rectangle2_heights[1168]), .rectangle2_weight(rectangle2_weights[1168]), .rectangle3_x(rectangle3_xs[1168]), .rectangle3_y(rectangle3_ys[1168]), .rectangle3_width(rectangle3_widths[1168]), .rectangle3_height(rectangle3_heights[1168]), .rectangle3_weight(rectangle3_weights[1168]), .feature_threshold(feature_thresholds[1168]), .feature_above(feature_aboves[1168]), .feature_below(feature_belows[1168]), .scan_win_std_dev(scan_win_std_dev[1168]), .feature_accum(feature_accums[1168]));
  accum_calculator ac1169(.scan_win(scan_win1169), .rectangle1_x(rectangle1_xs[1169]), .rectangle1_y(rectangle1_ys[1169]), .rectangle1_width(rectangle1_widths[1169]), .rectangle1_height(rectangle1_heights[1169]), .rectangle1_weight(rectangle1_weights[1169]), .rectangle2_x(rectangle2_xs[1169]), .rectangle2_y(rectangle2_ys[1169]), .rectangle2_width(rectangle2_widths[1169]), .rectangle2_height(rectangle2_heights[1169]), .rectangle2_weight(rectangle2_weights[1169]), .rectangle3_x(rectangle3_xs[1169]), .rectangle3_y(rectangle3_ys[1169]), .rectangle3_width(rectangle3_widths[1169]), .rectangle3_height(rectangle3_heights[1169]), .rectangle3_weight(rectangle3_weights[1169]), .feature_threshold(feature_thresholds[1169]), .feature_above(feature_aboves[1169]), .feature_below(feature_belows[1169]), .scan_win_std_dev(scan_win_std_dev[1169]), .feature_accum(feature_accums[1169]));
  accum_calculator ac1170(.scan_win(scan_win1170), .rectangle1_x(rectangle1_xs[1170]), .rectangle1_y(rectangle1_ys[1170]), .rectangle1_width(rectangle1_widths[1170]), .rectangle1_height(rectangle1_heights[1170]), .rectangle1_weight(rectangle1_weights[1170]), .rectangle2_x(rectangle2_xs[1170]), .rectangle2_y(rectangle2_ys[1170]), .rectangle2_width(rectangle2_widths[1170]), .rectangle2_height(rectangle2_heights[1170]), .rectangle2_weight(rectangle2_weights[1170]), .rectangle3_x(rectangle3_xs[1170]), .rectangle3_y(rectangle3_ys[1170]), .rectangle3_width(rectangle3_widths[1170]), .rectangle3_height(rectangle3_heights[1170]), .rectangle3_weight(rectangle3_weights[1170]), .feature_threshold(feature_thresholds[1170]), .feature_above(feature_aboves[1170]), .feature_below(feature_belows[1170]), .scan_win_std_dev(scan_win_std_dev[1170]), .feature_accum(feature_accums[1170]));
  accum_calculator ac1171(.scan_win(scan_win1171), .rectangle1_x(rectangle1_xs[1171]), .rectangle1_y(rectangle1_ys[1171]), .rectangle1_width(rectangle1_widths[1171]), .rectangle1_height(rectangle1_heights[1171]), .rectangle1_weight(rectangle1_weights[1171]), .rectangle2_x(rectangle2_xs[1171]), .rectangle2_y(rectangle2_ys[1171]), .rectangle2_width(rectangle2_widths[1171]), .rectangle2_height(rectangle2_heights[1171]), .rectangle2_weight(rectangle2_weights[1171]), .rectangle3_x(rectangle3_xs[1171]), .rectangle3_y(rectangle3_ys[1171]), .rectangle3_width(rectangle3_widths[1171]), .rectangle3_height(rectangle3_heights[1171]), .rectangle3_weight(rectangle3_weights[1171]), .feature_threshold(feature_thresholds[1171]), .feature_above(feature_aboves[1171]), .feature_below(feature_belows[1171]), .scan_win_std_dev(scan_win_std_dev[1171]), .feature_accum(feature_accums[1171]));
  accum_calculator ac1172(.scan_win(scan_win1172), .rectangle1_x(rectangle1_xs[1172]), .rectangle1_y(rectangle1_ys[1172]), .rectangle1_width(rectangle1_widths[1172]), .rectangle1_height(rectangle1_heights[1172]), .rectangle1_weight(rectangle1_weights[1172]), .rectangle2_x(rectangle2_xs[1172]), .rectangle2_y(rectangle2_ys[1172]), .rectangle2_width(rectangle2_widths[1172]), .rectangle2_height(rectangle2_heights[1172]), .rectangle2_weight(rectangle2_weights[1172]), .rectangle3_x(rectangle3_xs[1172]), .rectangle3_y(rectangle3_ys[1172]), .rectangle3_width(rectangle3_widths[1172]), .rectangle3_height(rectangle3_heights[1172]), .rectangle3_weight(rectangle3_weights[1172]), .feature_threshold(feature_thresholds[1172]), .feature_above(feature_aboves[1172]), .feature_below(feature_belows[1172]), .scan_win_std_dev(scan_win_std_dev[1172]), .feature_accum(feature_accums[1172]));
  accum_calculator ac1173(.scan_win(scan_win1173), .rectangle1_x(rectangle1_xs[1173]), .rectangle1_y(rectangle1_ys[1173]), .rectangle1_width(rectangle1_widths[1173]), .rectangle1_height(rectangle1_heights[1173]), .rectangle1_weight(rectangle1_weights[1173]), .rectangle2_x(rectangle2_xs[1173]), .rectangle2_y(rectangle2_ys[1173]), .rectangle2_width(rectangle2_widths[1173]), .rectangle2_height(rectangle2_heights[1173]), .rectangle2_weight(rectangle2_weights[1173]), .rectangle3_x(rectangle3_xs[1173]), .rectangle3_y(rectangle3_ys[1173]), .rectangle3_width(rectangle3_widths[1173]), .rectangle3_height(rectangle3_heights[1173]), .rectangle3_weight(rectangle3_weights[1173]), .feature_threshold(feature_thresholds[1173]), .feature_above(feature_aboves[1173]), .feature_below(feature_belows[1173]), .scan_win_std_dev(scan_win_std_dev[1173]), .feature_accum(feature_accums[1173]));
  accum_calculator ac1174(.scan_win(scan_win1174), .rectangle1_x(rectangle1_xs[1174]), .rectangle1_y(rectangle1_ys[1174]), .rectangle1_width(rectangle1_widths[1174]), .rectangle1_height(rectangle1_heights[1174]), .rectangle1_weight(rectangle1_weights[1174]), .rectangle2_x(rectangle2_xs[1174]), .rectangle2_y(rectangle2_ys[1174]), .rectangle2_width(rectangle2_widths[1174]), .rectangle2_height(rectangle2_heights[1174]), .rectangle2_weight(rectangle2_weights[1174]), .rectangle3_x(rectangle3_xs[1174]), .rectangle3_y(rectangle3_ys[1174]), .rectangle3_width(rectangle3_widths[1174]), .rectangle3_height(rectangle3_heights[1174]), .rectangle3_weight(rectangle3_weights[1174]), .feature_threshold(feature_thresholds[1174]), .feature_above(feature_aboves[1174]), .feature_below(feature_belows[1174]), .scan_win_std_dev(scan_win_std_dev[1174]), .feature_accum(feature_accums[1174]));
  accum_calculator ac1175(.scan_win(scan_win1175), .rectangle1_x(rectangle1_xs[1175]), .rectangle1_y(rectangle1_ys[1175]), .rectangle1_width(rectangle1_widths[1175]), .rectangle1_height(rectangle1_heights[1175]), .rectangle1_weight(rectangle1_weights[1175]), .rectangle2_x(rectangle2_xs[1175]), .rectangle2_y(rectangle2_ys[1175]), .rectangle2_width(rectangle2_widths[1175]), .rectangle2_height(rectangle2_heights[1175]), .rectangle2_weight(rectangle2_weights[1175]), .rectangle3_x(rectangle3_xs[1175]), .rectangle3_y(rectangle3_ys[1175]), .rectangle3_width(rectangle3_widths[1175]), .rectangle3_height(rectangle3_heights[1175]), .rectangle3_weight(rectangle3_weights[1175]), .feature_threshold(feature_thresholds[1175]), .feature_above(feature_aboves[1175]), .feature_below(feature_belows[1175]), .scan_win_std_dev(scan_win_std_dev[1175]), .feature_accum(feature_accums[1175]));
  accum_calculator ac1176(.scan_win(scan_win1176), .rectangle1_x(rectangle1_xs[1176]), .rectangle1_y(rectangle1_ys[1176]), .rectangle1_width(rectangle1_widths[1176]), .rectangle1_height(rectangle1_heights[1176]), .rectangle1_weight(rectangle1_weights[1176]), .rectangle2_x(rectangle2_xs[1176]), .rectangle2_y(rectangle2_ys[1176]), .rectangle2_width(rectangle2_widths[1176]), .rectangle2_height(rectangle2_heights[1176]), .rectangle2_weight(rectangle2_weights[1176]), .rectangle3_x(rectangle3_xs[1176]), .rectangle3_y(rectangle3_ys[1176]), .rectangle3_width(rectangle3_widths[1176]), .rectangle3_height(rectangle3_heights[1176]), .rectangle3_weight(rectangle3_weights[1176]), .feature_threshold(feature_thresholds[1176]), .feature_above(feature_aboves[1176]), .feature_below(feature_belows[1176]), .scan_win_std_dev(scan_win_std_dev[1176]), .feature_accum(feature_accums[1176]));
  accum_calculator ac1177(.scan_win(scan_win1177), .rectangle1_x(rectangle1_xs[1177]), .rectangle1_y(rectangle1_ys[1177]), .rectangle1_width(rectangle1_widths[1177]), .rectangle1_height(rectangle1_heights[1177]), .rectangle1_weight(rectangle1_weights[1177]), .rectangle2_x(rectangle2_xs[1177]), .rectangle2_y(rectangle2_ys[1177]), .rectangle2_width(rectangle2_widths[1177]), .rectangle2_height(rectangle2_heights[1177]), .rectangle2_weight(rectangle2_weights[1177]), .rectangle3_x(rectangle3_xs[1177]), .rectangle3_y(rectangle3_ys[1177]), .rectangle3_width(rectangle3_widths[1177]), .rectangle3_height(rectangle3_heights[1177]), .rectangle3_weight(rectangle3_weights[1177]), .feature_threshold(feature_thresholds[1177]), .feature_above(feature_aboves[1177]), .feature_below(feature_belows[1177]), .scan_win_std_dev(scan_win_std_dev[1177]), .feature_accum(feature_accums[1177]));
  accum_calculator ac1178(.scan_win(scan_win1178), .rectangle1_x(rectangle1_xs[1178]), .rectangle1_y(rectangle1_ys[1178]), .rectangle1_width(rectangle1_widths[1178]), .rectangle1_height(rectangle1_heights[1178]), .rectangle1_weight(rectangle1_weights[1178]), .rectangle2_x(rectangle2_xs[1178]), .rectangle2_y(rectangle2_ys[1178]), .rectangle2_width(rectangle2_widths[1178]), .rectangle2_height(rectangle2_heights[1178]), .rectangle2_weight(rectangle2_weights[1178]), .rectangle3_x(rectangle3_xs[1178]), .rectangle3_y(rectangle3_ys[1178]), .rectangle3_width(rectangle3_widths[1178]), .rectangle3_height(rectangle3_heights[1178]), .rectangle3_weight(rectangle3_weights[1178]), .feature_threshold(feature_thresholds[1178]), .feature_above(feature_aboves[1178]), .feature_below(feature_belows[1178]), .scan_win_std_dev(scan_win_std_dev[1178]), .feature_accum(feature_accums[1178]));
  accum_calculator ac1179(.scan_win(scan_win1179), .rectangle1_x(rectangle1_xs[1179]), .rectangle1_y(rectangle1_ys[1179]), .rectangle1_width(rectangle1_widths[1179]), .rectangle1_height(rectangle1_heights[1179]), .rectangle1_weight(rectangle1_weights[1179]), .rectangle2_x(rectangle2_xs[1179]), .rectangle2_y(rectangle2_ys[1179]), .rectangle2_width(rectangle2_widths[1179]), .rectangle2_height(rectangle2_heights[1179]), .rectangle2_weight(rectangle2_weights[1179]), .rectangle3_x(rectangle3_xs[1179]), .rectangle3_y(rectangle3_ys[1179]), .rectangle3_width(rectangle3_widths[1179]), .rectangle3_height(rectangle3_heights[1179]), .rectangle3_weight(rectangle3_weights[1179]), .feature_threshold(feature_thresholds[1179]), .feature_above(feature_aboves[1179]), .feature_below(feature_belows[1179]), .scan_win_std_dev(scan_win_std_dev[1179]), .feature_accum(feature_accums[1179]));
  accum_calculator ac1180(.scan_win(scan_win1180), .rectangle1_x(rectangle1_xs[1180]), .rectangle1_y(rectangle1_ys[1180]), .rectangle1_width(rectangle1_widths[1180]), .rectangle1_height(rectangle1_heights[1180]), .rectangle1_weight(rectangle1_weights[1180]), .rectangle2_x(rectangle2_xs[1180]), .rectangle2_y(rectangle2_ys[1180]), .rectangle2_width(rectangle2_widths[1180]), .rectangle2_height(rectangle2_heights[1180]), .rectangle2_weight(rectangle2_weights[1180]), .rectangle3_x(rectangle3_xs[1180]), .rectangle3_y(rectangle3_ys[1180]), .rectangle3_width(rectangle3_widths[1180]), .rectangle3_height(rectangle3_heights[1180]), .rectangle3_weight(rectangle3_weights[1180]), .feature_threshold(feature_thresholds[1180]), .feature_above(feature_aboves[1180]), .feature_below(feature_belows[1180]), .scan_win_std_dev(scan_win_std_dev[1180]), .feature_accum(feature_accums[1180]));
  accum_calculator ac1181(.scan_win(scan_win1181), .rectangle1_x(rectangle1_xs[1181]), .rectangle1_y(rectangle1_ys[1181]), .rectangle1_width(rectangle1_widths[1181]), .rectangle1_height(rectangle1_heights[1181]), .rectangle1_weight(rectangle1_weights[1181]), .rectangle2_x(rectangle2_xs[1181]), .rectangle2_y(rectangle2_ys[1181]), .rectangle2_width(rectangle2_widths[1181]), .rectangle2_height(rectangle2_heights[1181]), .rectangle2_weight(rectangle2_weights[1181]), .rectangle3_x(rectangle3_xs[1181]), .rectangle3_y(rectangle3_ys[1181]), .rectangle3_width(rectangle3_widths[1181]), .rectangle3_height(rectangle3_heights[1181]), .rectangle3_weight(rectangle3_weights[1181]), .feature_threshold(feature_thresholds[1181]), .feature_above(feature_aboves[1181]), .feature_below(feature_belows[1181]), .scan_win_std_dev(scan_win_std_dev[1181]), .feature_accum(feature_accums[1181]));
  accum_calculator ac1182(.scan_win(scan_win1182), .rectangle1_x(rectangle1_xs[1182]), .rectangle1_y(rectangle1_ys[1182]), .rectangle1_width(rectangle1_widths[1182]), .rectangle1_height(rectangle1_heights[1182]), .rectangle1_weight(rectangle1_weights[1182]), .rectangle2_x(rectangle2_xs[1182]), .rectangle2_y(rectangle2_ys[1182]), .rectangle2_width(rectangle2_widths[1182]), .rectangle2_height(rectangle2_heights[1182]), .rectangle2_weight(rectangle2_weights[1182]), .rectangle3_x(rectangle3_xs[1182]), .rectangle3_y(rectangle3_ys[1182]), .rectangle3_width(rectangle3_widths[1182]), .rectangle3_height(rectangle3_heights[1182]), .rectangle3_weight(rectangle3_weights[1182]), .feature_threshold(feature_thresholds[1182]), .feature_above(feature_aboves[1182]), .feature_below(feature_belows[1182]), .scan_win_std_dev(scan_win_std_dev[1182]), .feature_accum(feature_accums[1182]));
  accum_calculator ac1183(.scan_win(scan_win1183), .rectangle1_x(rectangle1_xs[1183]), .rectangle1_y(rectangle1_ys[1183]), .rectangle1_width(rectangle1_widths[1183]), .rectangle1_height(rectangle1_heights[1183]), .rectangle1_weight(rectangle1_weights[1183]), .rectangle2_x(rectangle2_xs[1183]), .rectangle2_y(rectangle2_ys[1183]), .rectangle2_width(rectangle2_widths[1183]), .rectangle2_height(rectangle2_heights[1183]), .rectangle2_weight(rectangle2_weights[1183]), .rectangle3_x(rectangle3_xs[1183]), .rectangle3_y(rectangle3_ys[1183]), .rectangle3_width(rectangle3_widths[1183]), .rectangle3_height(rectangle3_heights[1183]), .rectangle3_weight(rectangle3_weights[1183]), .feature_threshold(feature_thresholds[1183]), .feature_above(feature_aboves[1183]), .feature_below(feature_belows[1183]), .scan_win_std_dev(scan_win_std_dev[1183]), .feature_accum(feature_accums[1183]));
  accum_calculator ac1184(.scan_win(scan_win1184), .rectangle1_x(rectangle1_xs[1184]), .rectangle1_y(rectangle1_ys[1184]), .rectangle1_width(rectangle1_widths[1184]), .rectangle1_height(rectangle1_heights[1184]), .rectangle1_weight(rectangle1_weights[1184]), .rectangle2_x(rectangle2_xs[1184]), .rectangle2_y(rectangle2_ys[1184]), .rectangle2_width(rectangle2_widths[1184]), .rectangle2_height(rectangle2_heights[1184]), .rectangle2_weight(rectangle2_weights[1184]), .rectangle3_x(rectangle3_xs[1184]), .rectangle3_y(rectangle3_ys[1184]), .rectangle3_width(rectangle3_widths[1184]), .rectangle3_height(rectangle3_heights[1184]), .rectangle3_weight(rectangle3_weights[1184]), .feature_threshold(feature_thresholds[1184]), .feature_above(feature_aboves[1184]), .feature_below(feature_belows[1184]), .scan_win_std_dev(scan_win_std_dev[1184]), .feature_accum(feature_accums[1184]));
  accum_calculator ac1185(.scan_win(scan_win1185), .rectangle1_x(rectangle1_xs[1185]), .rectangle1_y(rectangle1_ys[1185]), .rectangle1_width(rectangle1_widths[1185]), .rectangle1_height(rectangle1_heights[1185]), .rectangle1_weight(rectangle1_weights[1185]), .rectangle2_x(rectangle2_xs[1185]), .rectangle2_y(rectangle2_ys[1185]), .rectangle2_width(rectangle2_widths[1185]), .rectangle2_height(rectangle2_heights[1185]), .rectangle2_weight(rectangle2_weights[1185]), .rectangle3_x(rectangle3_xs[1185]), .rectangle3_y(rectangle3_ys[1185]), .rectangle3_width(rectangle3_widths[1185]), .rectangle3_height(rectangle3_heights[1185]), .rectangle3_weight(rectangle3_weights[1185]), .feature_threshold(feature_thresholds[1185]), .feature_above(feature_aboves[1185]), .feature_below(feature_belows[1185]), .scan_win_std_dev(scan_win_std_dev[1185]), .feature_accum(feature_accums[1185]));
  accum_calculator ac1186(.scan_win(scan_win1186), .rectangle1_x(rectangle1_xs[1186]), .rectangle1_y(rectangle1_ys[1186]), .rectangle1_width(rectangle1_widths[1186]), .rectangle1_height(rectangle1_heights[1186]), .rectangle1_weight(rectangle1_weights[1186]), .rectangle2_x(rectangle2_xs[1186]), .rectangle2_y(rectangle2_ys[1186]), .rectangle2_width(rectangle2_widths[1186]), .rectangle2_height(rectangle2_heights[1186]), .rectangle2_weight(rectangle2_weights[1186]), .rectangle3_x(rectangle3_xs[1186]), .rectangle3_y(rectangle3_ys[1186]), .rectangle3_width(rectangle3_widths[1186]), .rectangle3_height(rectangle3_heights[1186]), .rectangle3_weight(rectangle3_weights[1186]), .feature_threshold(feature_thresholds[1186]), .feature_above(feature_aboves[1186]), .feature_below(feature_belows[1186]), .scan_win_std_dev(scan_win_std_dev[1186]), .feature_accum(feature_accums[1186]));
  accum_calculator ac1187(.scan_win(scan_win1187), .rectangle1_x(rectangle1_xs[1187]), .rectangle1_y(rectangle1_ys[1187]), .rectangle1_width(rectangle1_widths[1187]), .rectangle1_height(rectangle1_heights[1187]), .rectangle1_weight(rectangle1_weights[1187]), .rectangle2_x(rectangle2_xs[1187]), .rectangle2_y(rectangle2_ys[1187]), .rectangle2_width(rectangle2_widths[1187]), .rectangle2_height(rectangle2_heights[1187]), .rectangle2_weight(rectangle2_weights[1187]), .rectangle3_x(rectangle3_xs[1187]), .rectangle3_y(rectangle3_ys[1187]), .rectangle3_width(rectangle3_widths[1187]), .rectangle3_height(rectangle3_heights[1187]), .rectangle3_weight(rectangle3_weights[1187]), .feature_threshold(feature_thresholds[1187]), .feature_above(feature_aboves[1187]), .feature_below(feature_belows[1187]), .scan_win_std_dev(scan_win_std_dev[1187]), .feature_accum(feature_accums[1187]));
  accum_calculator ac1188(.scan_win(scan_win1188), .rectangle1_x(rectangle1_xs[1188]), .rectangle1_y(rectangle1_ys[1188]), .rectangle1_width(rectangle1_widths[1188]), .rectangle1_height(rectangle1_heights[1188]), .rectangle1_weight(rectangle1_weights[1188]), .rectangle2_x(rectangle2_xs[1188]), .rectangle2_y(rectangle2_ys[1188]), .rectangle2_width(rectangle2_widths[1188]), .rectangle2_height(rectangle2_heights[1188]), .rectangle2_weight(rectangle2_weights[1188]), .rectangle3_x(rectangle3_xs[1188]), .rectangle3_y(rectangle3_ys[1188]), .rectangle3_width(rectangle3_widths[1188]), .rectangle3_height(rectangle3_heights[1188]), .rectangle3_weight(rectangle3_weights[1188]), .feature_threshold(feature_thresholds[1188]), .feature_above(feature_aboves[1188]), .feature_below(feature_belows[1188]), .scan_win_std_dev(scan_win_std_dev[1188]), .feature_accum(feature_accums[1188]));
  accum_calculator ac1189(.scan_win(scan_win1189), .rectangle1_x(rectangle1_xs[1189]), .rectangle1_y(rectangle1_ys[1189]), .rectangle1_width(rectangle1_widths[1189]), .rectangle1_height(rectangle1_heights[1189]), .rectangle1_weight(rectangle1_weights[1189]), .rectangle2_x(rectangle2_xs[1189]), .rectangle2_y(rectangle2_ys[1189]), .rectangle2_width(rectangle2_widths[1189]), .rectangle2_height(rectangle2_heights[1189]), .rectangle2_weight(rectangle2_weights[1189]), .rectangle3_x(rectangle3_xs[1189]), .rectangle3_y(rectangle3_ys[1189]), .rectangle3_width(rectangle3_widths[1189]), .rectangle3_height(rectangle3_heights[1189]), .rectangle3_weight(rectangle3_weights[1189]), .feature_threshold(feature_thresholds[1189]), .feature_above(feature_aboves[1189]), .feature_below(feature_belows[1189]), .scan_win_std_dev(scan_win_std_dev[1189]), .feature_accum(feature_accums[1189]));
  accum_calculator ac1190(.scan_win(scan_win1190), .rectangle1_x(rectangle1_xs[1190]), .rectangle1_y(rectangle1_ys[1190]), .rectangle1_width(rectangle1_widths[1190]), .rectangle1_height(rectangle1_heights[1190]), .rectangle1_weight(rectangle1_weights[1190]), .rectangle2_x(rectangle2_xs[1190]), .rectangle2_y(rectangle2_ys[1190]), .rectangle2_width(rectangle2_widths[1190]), .rectangle2_height(rectangle2_heights[1190]), .rectangle2_weight(rectangle2_weights[1190]), .rectangle3_x(rectangle3_xs[1190]), .rectangle3_y(rectangle3_ys[1190]), .rectangle3_width(rectangle3_widths[1190]), .rectangle3_height(rectangle3_heights[1190]), .rectangle3_weight(rectangle3_weights[1190]), .feature_threshold(feature_thresholds[1190]), .feature_above(feature_aboves[1190]), .feature_below(feature_belows[1190]), .scan_win_std_dev(scan_win_std_dev[1190]), .feature_accum(feature_accums[1190]));
  accum_calculator ac1191(.scan_win(scan_win1191), .rectangle1_x(rectangle1_xs[1191]), .rectangle1_y(rectangle1_ys[1191]), .rectangle1_width(rectangle1_widths[1191]), .rectangle1_height(rectangle1_heights[1191]), .rectangle1_weight(rectangle1_weights[1191]), .rectangle2_x(rectangle2_xs[1191]), .rectangle2_y(rectangle2_ys[1191]), .rectangle2_width(rectangle2_widths[1191]), .rectangle2_height(rectangle2_heights[1191]), .rectangle2_weight(rectangle2_weights[1191]), .rectangle3_x(rectangle3_xs[1191]), .rectangle3_y(rectangle3_ys[1191]), .rectangle3_width(rectangle3_widths[1191]), .rectangle3_height(rectangle3_heights[1191]), .rectangle3_weight(rectangle3_weights[1191]), .feature_threshold(feature_thresholds[1191]), .feature_above(feature_aboves[1191]), .feature_below(feature_belows[1191]), .scan_win_std_dev(scan_win_std_dev[1191]), .feature_accum(feature_accums[1191]));
  accum_calculator ac1192(.scan_win(scan_win1192), .rectangle1_x(rectangle1_xs[1192]), .rectangle1_y(rectangle1_ys[1192]), .rectangle1_width(rectangle1_widths[1192]), .rectangle1_height(rectangle1_heights[1192]), .rectangle1_weight(rectangle1_weights[1192]), .rectangle2_x(rectangle2_xs[1192]), .rectangle2_y(rectangle2_ys[1192]), .rectangle2_width(rectangle2_widths[1192]), .rectangle2_height(rectangle2_heights[1192]), .rectangle2_weight(rectangle2_weights[1192]), .rectangle3_x(rectangle3_xs[1192]), .rectangle3_y(rectangle3_ys[1192]), .rectangle3_width(rectangle3_widths[1192]), .rectangle3_height(rectangle3_heights[1192]), .rectangle3_weight(rectangle3_weights[1192]), .feature_threshold(feature_thresholds[1192]), .feature_above(feature_aboves[1192]), .feature_below(feature_belows[1192]), .scan_win_std_dev(scan_win_std_dev[1192]), .feature_accum(feature_accums[1192]));
  accum_calculator ac1193(.scan_win(scan_win1193), .rectangle1_x(rectangle1_xs[1193]), .rectangle1_y(rectangle1_ys[1193]), .rectangle1_width(rectangle1_widths[1193]), .rectangle1_height(rectangle1_heights[1193]), .rectangle1_weight(rectangle1_weights[1193]), .rectangle2_x(rectangle2_xs[1193]), .rectangle2_y(rectangle2_ys[1193]), .rectangle2_width(rectangle2_widths[1193]), .rectangle2_height(rectangle2_heights[1193]), .rectangle2_weight(rectangle2_weights[1193]), .rectangle3_x(rectangle3_xs[1193]), .rectangle3_y(rectangle3_ys[1193]), .rectangle3_width(rectangle3_widths[1193]), .rectangle3_height(rectangle3_heights[1193]), .rectangle3_weight(rectangle3_weights[1193]), .feature_threshold(feature_thresholds[1193]), .feature_above(feature_aboves[1193]), .feature_below(feature_belows[1193]), .scan_win_std_dev(scan_win_std_dev[1193]), .feature_accum(feature_accums[1193]));
  accum_calculator ac1194(.scan_win(scan_win1194), .rectangle1_x(rectangle1_xs[1194]), .rectangle1_y(rectangle1_ys[1194]), .rectangle1_width(rectangle1_widths[1194]), .rectangle1_height(rectangle1_heights[1194]), .rectangle1_weight(rectangle1_weights[1194]), .rectangle2_x(rectangle2_xs[1194]), .rectangle2_y(rectangle2_ys[1194]), .rectangle2_width(rectangle2_widths[1194]), .rectangle2_height(rectangle2_heights[1194]), .rectangle2_weight(rectangle2_weights[1194]), .rectangle3_x(rectangle3_xs[1194]), .rectangle3_y(rectangle3_ys[1194]), .rectangle3_width(rectangle3_widths[1194]), .rectangle3_height(rectangle3_heights[1194]), .rectangle3_weight(rectangle3_weights[1194]), .feature_threshold(feature_thresholds[1194]), .feature_above(feature_aboves[1194]), .feature_below(feature_belows[1194]), .scan_win_std_dev(scan_win_std_dev[1194]), .feature_accum(feature_accums[1194]));
  accum_calculator ac1195(.scan_win(scan_win1195), .rectangle1_x(rectangle1_xs[1195]), .rectangle1_y(rectangle1_ys[1195]), .rectangle1_width(rectangle1_widths[1195]), .rectangle1_height(rectangle1_heights[1195]), .rectangle1_weight(rectangle1_weights[1195]), .rectangle2_x(rectangle2_xs[1195]), .rectangle2_y(rectangle2_ys[1195]), .rectangle2_width(rectangle2_widths[1195]), .rectangle2_height(rectangle2_heights[1195]), .rectangle2_weight(rectangle2_weights[1195]), .rectangle3_x(rectangle3_xs[1195]), .rectangle3_y(rectangle3_ys[1195]), .rectangle3_width(rectangle3_widths[1195]), .rectangle3_height(rectangle3_heights[1195]), .rectangle3_weight(rectangle3_weights[1195]), .feature_threshold(feature_thresholds[1195]), .feature_above(feature_aboves[1195]), .feature_below(feature_belows[1195]), .scan_win_std_dev(scan_win_std_dev[1195]), .feature_accum(feature_accums[1195]));
  accum_calculator ac1196(.scan_win(scan_win1196), .rectangle1_x(rectangle1_xs[1196]), .rectangle1_y(rectangle1_ys[1196]), .rectangle1_width(rectangle1_widths[1196]), .rectangle1_height(rectangle1_heights[1196]), .rectangle1_weight(rectangle1_weights[1196]), .rectangle2_x(rectangle2_xs[1196]), .rectangle2_y(rectangle2_ys[1196]), .rectangle2_width(rectangle2_widths[1196]), .rectangle2_height(rectangle2_heights[1196]), .rectangle2_weight(rectangle2_weights[1196]), .rectangle3_x(rectangle3_xs[1196]), .rectangle3_y(rectangle3_ys[1196]), .rectangle3_width(rectangle3_widths[1196]), .rectangle3_height(rectangle3_heights[1196]), .rectangle3_weight(rectangle3_weights[1196]), .feature_threshold(feature_thresholds[1196]), .feature_above(feature_aboves[1196]), .feature_below(feature_belows[1196]), .scan_win_std_dev(scan_win_std_dev[1196]), .feature_accum(feature_accums[1196]));
  accum_calculator ac1197(.scan_win(scan_win1197), .rectangle1_x(rectangle1_xs[1197]), .rectangle1_y(rectangle1_ys[1197]), .rectangle1_width(rectangle1_widths[1197]), .rectangle1_height(rectangle1_heights[1197]), .rectangle1_weight(rectangle1_weights[1197]), .rectangle2_x(rectangle2_xs[1197]), .rectangle2_y(rectangle2_ys[1197]), .rectangle2_width(rectangle2_widths[1197]), .rectangle2_height(rectangle2_heights[1197]), .rectangle2_weight(rectangle2_weights[1197]), .rectangle3_x(rectangle3_xs[1197]), .rectangle3_y(rectangle3_ys[1197]), .rectangle3_width(rectangle3_widths[1197]), .rectangle3_height(rectangle3_heights[1197]), .rectangle3_weight(rectangle3_weights[1197]), .feature_threshold(feature_thresholds[1197]), .feature_above(feature_aboves[1197]), .feature_below(feature_belows[1197]), .scan_win_std_dev(scan_win_std_dev[1197]), .feature_accum(feature_accums[1197]));
  accum_calculator ac1198(.scan_win(scan_win1198), .rectangle1_x(rectangle1_xs[1198]), .rectangle1_y(rectangle1_ys[1198]), .rectangle1_width(rectangle1_widths[1198]), .rectangle1_height(rectangle1_heights[1198]), .rectangle1_weight(rectangle1_weights[1198]), .rectangle2_x(rectangle2_xs[1198]), .rectangle2_y(rectangle2_ys[1198]), .rectangle2_width(rectangle2_widths[1198]), .rectangle2_height(rectangle2_heights[1198]), .rectangle2_weight(rectangle2_weights[1198]), .rectangle3_x(rectangle3_xs[1198]), .rectangle3_y(rectangle3_ys[1198]), .rectangle3_width(rectangle3_widths[1198]), .rectangle3_height(rectangle3_heights[1198]), .rectangle3_weight(rectangle3_weights[1198]), .feature_threshold(feature_thresholds[1198]), .feature_above(feature_aboves[1198]), .feature_below(feature_belows[1198]), .scan_win_std_dev(scan_win_std_dev[1198]), .feature_accum(feature_accums[1198]));
  accum_calculator ac1199(.scan_win(scan_win1199), .rectangle1_x(rectangle1_xs[1199]), .rectangle1_y(rectangle1_ys[1199]), .rectangle1_width(rectangle1_widths[1199]), .rectangle1_height(rectangle1_heights[1199]), .rectangle1_weight(rectangle1_weights[1199]), .rectangle2_x(rectangle2_xs[1199]), .rectangle2_y(rectangle2_ys[1199]), .rectangle2_width(rectangle2_widths[1199]), .rectangle2_height(rectangle2_heights[1199]), .rectangle2_weight(rectangle2_weights[1199]), .rectangle3_x(rectangle3_xs[1199]), .rectangle3_y(rectangle3_ys[1199]), .rectangle3_width(rectangle3_widths[1199]), .rectangle3_height(rectangle3_heights[1199]), .rectangle3_weight(rectangle3_weights[1199]), .feature_threshold(feature_thresholds[1199]), .feature_above(feature_aboves[1199]), .feature_below(feature_belows[1199]), .scan_win_std_dev(scan_win_std_dev[1199]), .feature_accum(feature_accums[1199]));
  accum_calculator ac1200(.scan_win(scan_win1200), .rectangle1_x(rectangle1_xs[1200]), .rectangle1_y(rectangle1_ys[1200]), .rectangle1_width(rectangle1_widths[1200]), .rectangle1_height(rectangle1_heights[1200]), .rectangle1_weight(rectangle1_weights[1200]), .rectangle2_x(rectangle2_xs[1200]), .rectangle2_y(rectangle2_ys[1200]), .rectangle2_width(rectangle2_widths[1200]), .rectangle2_height(rectangle2_heights[1200]), .rectangle2_weight(rectangle2_weights[1200]), .rectangle3_x(rectangle3_xs[1200]), .rectangle3_y(rectangle3_ys[1200]), .rectangle3_width(rectangle3_widths[1200]), .rectangle3_height(rectangle3_heights[1200]), .rectangle3_weight(rectangle3_weights[1200]), .feature_threshold(feature_thresholds[1200]), .feature_above(feature_aboves[1200]), .feature_below(feature_belows[1200]), .scan_win_std_dev(scan_win_std_dev[1200]), .feature_accum(feature_accums[1200]));
  accum_calculator ac1201(.scan_win(scan_win1201), .rectangle1_x(rectangle1_xs[1201]), .rectangle1_y(rectangle1_ys[1201]), .rectangle1_width(rectangle1_widths[1201]), .rectangle1_height(rectangle1_heights[1201]), .rectangle1_weight(rectangle1_weights[1201]), .rectangle2_x(rectangle2_xs[1201]), .rectangle2_y(rectangle2_ys[1201]), .rectangle2_width(rectangle2_widths[1201]), .rectangle2_height(rectangle2_heights[1201]), .rectangle2_weight(rectangle2_weights[1201]), .rectangle3_x(rectangle3_xs[1201]), .rectangle3_y(rectangle3_ys[1201]), .rectangle3_width(rectangle3_widths[1201]), .rectangle3_height(rectangle3_heights[1201]), .rectangle3_weight(rectangle3_weights[1201]), .feature_threshold(feature_thresholds[1201]), .feature_above(feature_aboves[1201]), .feature_below(feature_belows[1201]), .scan_win_std_dev(scan_win_std_dev[1201]), .feature_accum(feature_accums[1201]));
  accum_calculator ac1202(.scan_win(scan_win1202), .rectangle1_x(rectangle1_xs[1202]), .rectangle1_y(rectangle1_ys[1202]), .rectangle1_width(rectangle1_widths[1202]), .rectangle1_height(rectangle1_heights[1202]), .rectangle1_weight(rectangle1_weights[1202]), .rectangle2_x(rectangle2_xs[1202]), .rectangle2_y(rectangle2_ys[1202]), .rectangle2_width(rectangle2_widths[1202]), .rectangle2_height(rectangle2_heights[1202]), .rectangle2_weight(rectangle2_weights[1202]), .rectangle3_x(rectangle3_xs[1202]), .rectangle3_y(rectangle3_ys[1202]), .rectangle3_width(rectangle3_widths[1202]), .rectangle3_height(rectangle3_heights[1202]), .rectangle3_weight(rectangle3_weights[1202]), .feature_threshold(feature_thresholds[1202]), .feature_above(feature_aboves[1202]), .feature_below(feature_belows[1202]), .scan_win_std_dev(scan_win_std_dev[1202]), .feature_accum(feature_accums[1202]));
  accum_calculator ac1203(.scan_win(scan_win1203), .rectangle1_x(rectangle1_xs[1203]), .rectangle1_y(rectangle1_ys[1203]), .rectangle1_width(rectangle1_widths[1203]), .rectangle1_height(rectangle1_heights[1203]), .rectangle1_weight(rectangle1_weights[1203]), .rectangle2_x(rectangle2_xs[1203]), .rectangle2_y(rectangle2_ys[1203]), .rectangle2_width(rectangle2_widths[1203]), .rectangle2_height(rectangle2_heights[1203]), .rectangle2_weight(rectangle2_weights[1203]), .rectangle3_x(rectangle3_xs[1203]), .rectangle3_y(rectangle3_ys[1203]), .rectangle3_width(rectangle3_widths[1203]), .rectangle3_height(rectangle3_heights[1203]), .rectangle3_weight(rectangle3_weights[1203]), .feature_threshold(feature_thresholds[1203]), .feature_above(feature_aboves[1203]), .feature_below(feature_belows[1203]), .scan_win_std_dev(scan_win_std_dev[1203]), .feature_accum(feature_accums[1203]));
  accum_calculator ac1204(.scan_win(scan_win1204), .rectangle1_x(rectangle1_xs[1204]), .rectangle1_y(rectangle1_ys[1204]), .rectangle1_width(rectangle1_widths[1204]), .rectangle1_height(rectangle1_heights[1204]), .rectangle1_weight(rectangle1_weights[1204]), .rectangle2_x(rectangle2_xs[1204]), .rectangle2_y(rectangle2_ys[1204]), .rectangle2_width(rectangle2_widths[1204]), .rectangle2_height(rectangle2_heights[1204]), .rectangle2_weight(rectangle2_weights[1204]), .rectangle3_x(rectangle3_xs[1204]), .rectangle3_y(rectangle3_ys[1204]), .rectangle3_width(rectangle3_widths[1204]), .rectangle3_height(rectangle3_heights[1204]), .rectangle3_weight(rectangle3_weights[1204]), .feature_threshold(feature_thresholds[1204]), .feature_above(feature_aboves[1204]), .feature_below(feature_belows[1204]), .scan_win_std_dev(scan_win_std_dev[1204]), .feature_accum(feature_accums[1204]));
  accum_calculator ac1205(.scan_win(scan_win1205), .rectangle1_x(rectangle1_xs[1205]), .rectangle1_y(rectangle1_ys[1205]), .rectangle1_width(rectangle1_widths[1205]), .rectangle1_height(rectangle1_heights[1205]), .rectangle1_weight(rectangle1_weights[1205]), .rectangle2_x(rectangle2_xs[1205]), .rectangle2_y(rectangle2_ys[1205]), .rectangle2_width(rectangle2_widths[1205]), .rectangle2_height(rectangle2_heights[1205]), .rectangle2_weight(rectangle2_weights[1205]), .rectangle3_x(rectangle3_xs[1205]), .rectangle3_y(rectangle3_ys[1205]), .rectangle3_width(rectangle3_widths[1205]), .rectangle3_height(rectangle3_heights[1205]), .rectangle3_weight(rectangle3_weights[1205]), .feature_threshold(feature_thresholds[1205]), .feature_above(feature_aboves[1205]), .feature_below(feature_belows[1205]), .scan_win_std_dev(scan_win_std_dev[1205]), .feature_accum(feature_accums[1205]));
  accum_calculator ac1206(.scan_win(scan_win1206), .rectangle1_x(rectangle1_xs[1206]), .rectangle1_y(rectangle1_ys[1206]), .rectangle1_width(rectangle1_widths[1206]), .rectangle1_height(rectangle1_heights[1206]), .rectangle1_weight(rectangle1_weights[1206]), .rectangle2_x(rectangle2_xs[1206]), .rectangle2_y(rectangle2_ys[1206]), .rectangle2_width(rectangle2_widths[1206]), .rectangle2_height(rectangle2_heights[1206]), .rectangle2_weight(rectangle2_weights[1206]), .rectangle3_x(rectangle3_xs[1206]), .rectangle3_y(rectangle3_ys[1206]), .rectangle3_width(rectangle3_widths[1206]), .rectangle3_height(rectangle3_heights[1206]), .rectangle3_weight(rectangle3_weights[1206]), .feature_threshold(feature_thresholds[1206]), .feature_above(feature_aboves[1206]), .feature_below(feature_belows[1206]), .scan_win_std_dev(scan_win_std_dev[1206]), .feature_accum(feature_accums[1206]));
  accum_calculator ac1207(.scan_win(scan_win1207), .rectangle1_x(rectangle1_xs[1207]), .rectangle1_y(rectangle1_ys[1207]), .rectangle1_width(rectangle1_widths[1207]), .rectangle1_height(rectangle1_heights[1207]), .rectangle1_weight(rectangle1_weights[1207]), .rectangle2_x(rectangle2_xs[1207]), .rectangle2_y(rectangle2_ys[1207]), .rectangle2_width(rectangle2_widths[1207]), .rectangle2_height(rectangle2_heights[1207]), .rectangle2_weight(rectangle2_weights[1207]), .rectangle3_x(rectangle3_xs[1207]), .rectangle3_y(rectangle3_ys[1207]), .rectangle3_width(rectangle3_widths[1207]), .rectangle3_height(rectangle3_heights[1207]), .rectangle3_weight(rectangle3_weights[1207]), .feature_threshold(feature_thresholds[1207]), .feature_above(feature_aboves[1207]), .feature_below(feature_belows[1207]), .scan_win_std_dev(scan_win_std_dev[1207]), .feature_accum(feature_accums[1207]));
  accum_calculator ac1208(.scan_win(scan_win1208), .rectangle1_x(rectangle1_xs[1208]), .rectangle1_y(rectangle1_ys[1208]), .rectangle1_width(rectangle1_widths[1208]), .rectangle1_height(rectangle1_heights[1208]), .rectangle1_weight(rectangle1_weights[1208]), .rectangle2_x(rectangle2_xs[1208]), .rectangle2_y(rectangle2_ys[1208]), .rectangle2_width(rectangle2_widths[1208]), .rectangle2_height(rectangle2_heights[1208]), .rectangle2_weight(rectangle2_weights[1208]), .rectangle3_x(rectangle3_xs[1208]), .rectangle3_y(rectangle3_ys[1208]), .rectangle3_width(rectangle3_widths[1208]), .rectangle3_height(rectangle3_heights[1208]), .rectangle3_weight(rectangle3_weights[1208]), .feature_threshold(feature_thresholds[1208]), .feature_above(feature_aboves[1208]), .feature_below(feature_belows[1208]), .scan_win_std_dev(scan_win_std_dev[1208]), .feature_accum(feature_accums[1208]));
  accum_calculator ac1209(.scan_win(scan_win1209), .rectangle1_x(rectangle1_xs[1209]), .rectangle1_y(rectangle1_ys[1209]), .rectangle1_width(rectangle1_widths[1209]), .rectangle1_height(rectangle1_heights[1209]), .rectangle1_weight(rectangle1_weights[1209]), .rectangle2_x(rectangle2_xs[1209]), .rectangle2_y(rectangle2_ys[1209]), .rectangle2_width(rectangle2_widths[1209]), .rectangle2_height(rectangle2_heights[1209]), .rectangle2_weight(rectangle2_weights[1209]), .rectangle3_x(rectangle3_xs[1209]), .rectangle3_y(rectangle3_ys[1209]), .rectangle3_width(rectangle3_widths[1209]), .rectangle3_height(rectangle3_heights[1209]), .rectangle3_weight(rectangle3_weights[1209]), .feature_threshold(feature_thresholds[1209]), .feature_above(feature_aboves[1209]), .feature_below(feature_belows[1209]), .scan_win_std_dev(scan_win_std_dev[1209]), .feature_accum(feature_accums[1209]));
  accum_calculator ac1210(.scan_win(scan_win1210), .rectangle1_x(rectangle1_xs[1210]), .rectangle1_y(rectangle1_ys[1210]), .rectangle1_width(rectangle1_widths[1210]), .rectangle1_height(rectangle1_heights[1210]), .rectangle1_weight(rectangle1_weights[1210]), .rectangle2_x(rectangle2_xs[1210]), .rectangle2_y(rectangle2_ys[1210]), .rectangle2_width(rectangle2_widths[1210]), .rectangle2_height(rectangle2_heights[1210]), .rectangle2_weight(rectangle2_weights[1210]), .rectangle3_x(rectangle3_xs[1210]), .rectangle3_y(rectangle3_ys[1210]), .rectangle3_width(rectangle3_widths[1210]), .rectangle3_height(rectangle3_heights[1210]), .rectangle3_weight(rectangle3_weights[1210]), .feature_threshold(feature_thresholds[1210]), .feature_above(feature_aboves[1210]), .feature_below(feature_belows[1210]), .scan_win_std_dev(scan_win_std_dev[1210]), .feature_accum(feature_accums[1210]));
  accum_calculator ac1211(.scan_win(scan_win1211), .rectangle1_x(rectangle1_xs[1211]), .rectangle1_y(rectangle1_ys[1211]), .rectangle1_width(rectangle1_widths[1211]), .rectangle1_height(rectangle1_heights[1211]), .rectangle1_weight(rectangle1_weights[1211]), .rectangle2_x(rectangle2_xs[1211]), .rectangle2_y(rectangle2_ys[1211]), .rectangle2_width(rectangle2_widths[1211]), .rectangle2_height(rectangle2_heights[1211]), .rectangle2_weight(rectangle2_weights[1211]), .rectangle3_x(rectangle3_xs[1211]), .rectangle3_y(rectangle3_ys[1211]), .rectangle3_width(rectangle3_widths[1211]), .rectangle3_height(rectangle3_heights[1211]), .rectangle3_weight(rectangle3_weights[1211]), .feature_threshold(feature_thresholds[1211]), .feature_above(feature_aboves[1211]), .feature_below(feature_belows[1211]), .scan_win_std_dev(scan_win_std_dev[1211]), .feature_accum(feature_accums[1211]));
  accum_calculator ac1212(.scan_win(scan_win1212), .rectangle1_x(rectangle1_xs[1212]), .rectangle1_y(rectangle1_ys[1212]), .rectangle1_width(rectangle1_widths[1212]), .rectangle1_height(rectangle1_heights[1212]), .rectangle1_weight(rectangle1_weights[1212]), .rectangle2_x(rectangle2_xs[1212]), .rectangle2_y(rectangle2_ys[1212]), .rectangle2_width(rectangle2_widths[1212]), .rectangle2_height(rectangle2_heights[1212]), .rectangle2_weight(rectangle2_weights[1212]), .rectangle3_x(rectangle3_xs[1212]), .rectangle3_y(rectangle3_ys[1212]), .rectangle3_width(rectangle3_widths[1212]), .rectangle3_height(rectangle3_heights[1212]), .rectangle3_weight(rectangle3_weights[1212]), .feature_threshold(feature_thresholds[1212]), .feature_above(feature_aboves[1212]), .feature_below(feature_belows[1212]), .scan_win_std_dev(scan_win_std_dev[1212]), .feature_accum(feature_accums[1212]));
  accum_calculator ac1213(.scan_win(scan_win1213), .rectangle1_x(rectangle1_xs[1213]), .rectangle1_y(rectangle1_ys[1213]), .rectangle1_width(rectangle1_widths[1213]), .rectangle1_height(rectangle1_heights[1213]), .rectangle1_weight(rectangle1_weights[1213]), .rectangle2_x(rectangle2_xs[1213]), .rectangle2_y(rectangle2_ys[1213]), .rectangle2_width(rectangle2_widths[1213]), .rectangle2_height(rectangle2_heights[1213]), .rectangle2_weight(rectangle2_weights[1213]), .rectangle3_x(rectangle3_xs[1213]), .rectangle3_y(rectangle3_ys[1213]), .rectangle3_width(rectangle3_widths[1213]), .rectangle3_height(rectangle3_heights[1213]), .rectangle3_weight(rectangle3_weights[1213]), .feature_threshold(feature_thresholds[1213]), .feature_above(feature_aboves[1213]), .feature_below(feature_belows[1213]), .scan_win_std_dev(scan_win_std_dev[1213]), .feature_accum(feature_accums[1213]));
  accum_calculator ac1214(.scan_win(scan_win1214), .rectangle1_x(rectangle1_xs[1214]), .rectangle1_y(rectangle1_ys[1214]), .rectangle1_width(rectangle1_widths[1214]), .rectangle1_height(rectangle1_heights[1214]), .rectangle1_weight(rectangle1_weights[1214]), .rectangle2_x(rectangle2_xs[1214]), .rectangle2_y(rectangle2_ys[1214]), .rectangle2_width(rectangle2_widths[1214]), .rectangle2_height(rectangle2_heights[1214]), .rectangle2_weight(rectangle2_weights[1214]), .rectangle3_x(rectangle3_xs[1214]), .rectangle3_y(rectangle3_ys[1214]), .rectangle3_width(rectangle3_widths[1214]), .rectangle3_height(rectangle3_heights[1214]), .rectangle3_weight(rectangle3_weights[1214]), .feature_threshold(feature_thresholds[1214]), .feature_above(feature_aboves[1214]), .feature_below(feature_belows[1214]), .scan_win_std_dev(scan_win_std_dev[1214]), .feature_accum(feature_accums[1214]));
  accum_calculator ac1215(.scan_win(scan_win1215), .rectangle1_x(rectangle1_xs[1215]), .rectangle1_y(rectangle1_ys[1215]), .rectangle1_width(rectangle1_widths[1215]), .rectangle1_height(rectangle1_heights[1215]), .rectangle1_weight(rectangle1_weights[1215]), .rectangle2_x(rectangle2_xs[1215]), .rectangle2_y(rectangle2_ys[1215]), .rectangle2_width(rectangle2_widths[1215]), .rectangle2_height(rectangle2_heights[1215]), .rectangle2_weight(rectangle2_weights[1215]), .rectangle3_x(rectangle3_xs[1215]), .rectangle3_y(rectangle3_ys[1215]), .rectangle3_width(rectangle3_widths[1215]), .rectangle3_height(rectangle3_heights[1215]), .rectangle3_weight(rectangle3_weights[1215]), .feature_threshold(feature_thresholds[1215]), .feature_above(feature_aboves[1215]), .feature_below(feature_belows[1215]), .scan_win_std_dev(scan_win_std_dev[1215]), .feature_accum(feature_accums[1215]));
  accum_calculator ac1216(.scan_win(scan_win1216), .rectangle1_x(rectangle1_xs[1216]), .rectangle1_y(rectangle1_ys[1216]), .rectangle1_width(rectangle1_widths[1216]), .rectangle1_height(rectangle1_heights[1216]), .rectangle1_weight(rectangle1_weights[1216]), .rectangle2_x(rectangle2_xs[1216]), .rectangle2_y(rectangle2_ys[1216]), .rectangle2_width(rectangle2_widths[1216]), .rectangle2_height(rectangle2_heights[1216]), .rectangle2_weight(rectangle2_weights[1216]), .rectangle3_x(rectangle3_xs[1216]), .rectangle3_y(rectangle3_ys[1216]), .rectangle3_width(rectangle3_widths[1216]), .rectangle3_height(rectangle3_heights[1216]), .rectangle3_weight(rectangle3_weights[1216]), .feature_threshold(feature_thresholds[1216]), .feature_above(feature_aboves[1216]), .feature_below(feature_belows[1216]), .scan_win_std_dev(scan_win_std_dev[1216]), .feature_accum(feature_accums[1216]));
  accum_calculator ac1217(.scan_win(scan_win1217), .rectangle1_x(rectangle1_xs[1217]), .rectangle1_y(rectangle1_ys[1217]), .rectangle1_width(rectangle1_widths[1217]), .rectangle1_height(rectangle1_heights[1217]), .rectangle1_weight(rectangle1_weights[1217]), .rectangle2_x(rectangle2_xs[1217]), .rectangle2_y(rectangle2_ys[1217]), .rectangle2_width(rectangle2_widths[1217]), .rectangle2_height(rectangle2_heights[1217]), .rectangle2_weight(rectangle2_weights[1217]), .rectangle3_x(rectangle3_xs[1217]), .rectangle3_y(rectangle3_ys[1217]), .rectangle3_width(rectangle3_widths[1217]), .rectangle3_height(rectangle3_heights[1217]), .rectangle3_weight(rectangle3_weights[1217]), .feature_threshold(feature_thresholds[1217]), .feature_above(feature_aboves[1217]), .feature_below(feature_belows[1217]), .scan_win_std_dev(scan_win_std_dev[1217]), .feature_accum(feature_accums[1217]));
  accum_calculator ac1218(.scan_win(scan_win1218), .rectangle1_x(rectangle1_xs[1218]), .rectangle1_y(rectangle1_ys[1218]), .rectangle1_width(rectangle1_widths[1218]), .rectangle1_height(rectangle1_heights[1218]), .rectangle1_weight(rectangle1_weights[1218]), .rectangle2_x(rectangle2_xs[1218]), .rectangle2_y(rectangle2_ys[1218]), .rectangle2_width(rectangle2_widths[1218]), .rectangle2_height(rectangle2_heights[1218]), .rectangle2_weight(rectangle2_weights[1218]), .rectangle3_x(rectangle3_xs[1218]), .rectangle3_y(rectangle3_ys[1218]), .rectangle3_width(rectangle3_widths[1218]), .rectangle3_height(rectangle3_heights[1218]), .rectangle3_weight(rectangle3_weights[1218]), .feature_threshold(feature_thresholds[1218]), .feature_above(feature_aboves[1218]), .feature_below(feature_belows[1218]), .scan_win_std_dev(scan_win_std_dev[1218]), .feature_accum(feature_accums[1218]));
  accum_calculator ac1219(.scan_win(scan_win1219), .rectangle1_x(rectangle1_xs[1219]), .rectangle1_y(rectangle1_ys[1219]), .rectangle1_width(rectangle1_widths[1219]), .rectangle1_height(rectangle1_heights[1219]), .rectangle1_weight(rectangle1_weights[1219]), .rectangle2_x(rectangle2_xs[1219]), .rectangle2_y(rectangle2_ys[1219]), .rectangle2_width(rectangle2_widths[1219]), .rectangle2_height(rectangle2_heights[1219]), .rectangle2_weight(rectangle2_weights[1219]), .rectangle3_x(rectangle3_xs[1219]), .rectangle3_y(rectangle3_ys[1219]), .rectangle3_width(rectangle3_widths[1219]), .rectangle3_height(rectangle3_heights[1219]), .rectangle3_weight(rectangle3_weights[1219]), .feature_threshold(feature_thresholds[1219]), .feature_above(feature_aboves[1219]), .feature_below(feature_belows[1219]), .scan_win_std_dev(scan_win_std_dev[1219]), .feature_accum(feature_accums[1219]));
  accum_calculator ac1220(.scan_win(scan_win1220), .rectangle1_x(rectangle1_xs[1220]), .rectangle1_y(rectangle1_ys[1220]), .rectangle1_width(rectangle1_widths[1220]), .rectangle1_height(rectangle1_heights[1220]), .rectangle1_weight(rectangle1_weights[1220]), .rectangle2_x(rectangle2_xs[1220]), .rectangle2_y(rectangle2_ys[1220]), .rectangle2_width(rectangle2_widths[1220]), .rectangle2_height(rectangle2_heights[1220]), .rectangle2_weight(rectangle2_weights[1220]), .rectangle3_x(rectangle3_xs[1220]), .rectangle3_y(rectangle3_ys[1220]), .rectangle3_width(rectangle3_widths[1220]), .rectangle3_height(rectangle3_heights[1220]), .rectangle3_weight(rectangle3_weights[1220]), .feature_threshold(feature_thresholds[1220]), .feature_above(feature_aboves[1220]), .feature_below(feature_belows[1220]), .scan_win_std_dev(scan_win_std_dev[1220]), .feature_accum(feature_accums[1220]));
  accum_calculator ac1221(.scan_win(scan_win1221), .rectangle1_x(rectangle1_xs[1221]), .rectangle1_y(rectangle1_ys[1221]), .rectangle1_width(rectangle1_widths[1221]), .rectangle1_height(rectangle1_heights[1221]), .rectangle1_weight(rectangle1_weights[1221]), .rectangle2_x(rectangle2_xs[1221]), .rectangle2_y(rectangle2_ys[1221]), .rectangle2_width(rectangle2_widths[1221]), .rectangle2_height(rectangle2_heights[1221]), .rectangle2_weight(rectangle2_weights[1221]), .rectangle3_x(rectangle3_xs[1221]), .rectangle3_y(rectangle3_ys[1221]), .rectangle3_width(rectangle3_widths[1221]), .rectangle3_height(rectangle3_heights[1221]), .rectangle3_weight(rectangle3_weights[1221]), .feature_threshold(feature_thresholds[1221]), .feature_above(feature_aboves[1221]), .feature_below(feature_belows[1221]), .scan_win_std_dev(scan_win_std_dev[1221]), .feature_accum(feature_accums[1221]));
  accum_calculator ac1222(.scan_win(scan_win1222), .rectangle1_x(rectangle1_xs[1222]), .rectangle1_y(rectangle1_ys[1222]), .rectangle1_width(rectangle1_widths[1222]), .rectangle1_height(rectangle1_heights[1222]), .rectangle1_weight(rectangle1_weights[1222]), .rectangle2_x(rectangle2_xs[1222]), .rectangle2_y(rectangle2_ys[1222]), .rectangle2_width(rectangle2_widths[1222]), .rectangle2_height(rectangle2_heights[1222]), .rectangle2_weight(rectangle2_weights[1222]), .rectangle3_x(rectangle3_xs[1222]), .rectangle3_y(rectangle3_ys[1222]), .rectangle3_width(rectangle3_widths[1222]), .rectangle3_height(rectangle3_heights[1222]), .rectangle3_weight(rectangle3_weights[1222]), .feature_threshold(feature_thresholds[1222]), .feature_above(feature_aboves[1222]), .feature_below(feature_belows[1222]), .scan_win_std_dev(scan_win_std_dev[1222]), .feature_accum(feature_accums[1222]));
  accum_calculator ac1223(.scan_win(scan_win1223), .rectangle1_x(rectangle1_xs[1223]), .rectangle1_y(rectangle1_ys[1223]), .rectangle1_width(rectangle1_widths[1223]), .rectangle1_height(rectangle1_heights[1223]), .rectangle1_weight(rectangle1_weights[1223]), .rectangle2_x(rectangle2_xs[1223]), .rectangle2_y(rectangle2_ys[1223]), .rectangle2_width(rectangle2_widths[1223]), .rectangle2_height(rectangle2_heights[1223]), .rectangle2_weight(rectangle2_weights[1223]), .rectangle3_x(rectangle3_xs[1223]), .rectangle3_y(rectangle3_ys[1223]), .rectangle3_width(rectangle3_widths[1223]), .rectangle3_height(rectangle3_heights[1223]), .rectangle3_weight(rectangle3_weights[1223]), .feature_threshold(feature_thresholds[1223]), .feature_above(feature_aboves[1223]), .feature_below(feature_belows[1223]), .scan_win_std_dev(scan_win_std_dev[1223]), .feature_accum(feature_accums[1223]));
  accum_calculator ac1224(.scan_win(scan_win1224), .rectangle1_x(rectangle1_xs[1224]), .rectangle1_y(rectangle1_ys[1224]), .rectangle1_width(rectangle1_widths[1224]), .rectangle1_height(rectangle1_heights[1224]), .rectangle1_weight(rectangle1_weights[1224]), .rectangle2_x(rectangle2_xs[1224]), .rectangle2_y(rectangle2_ys[1224]), .rectangle2_width(rectangle2_widths[1224]), .rectangle2_height(rectangle2_heights[1224]), .rectangle2_weight(rectangle2_weights[1224]), .rectangle3_x(rectangle3_xs[1224]), .rectangle3_y(rectangle3_ys[1224]), .rectangle3_width(rectangle3_widths[1224]), .rectangle3_height(rectangle3_heights[1224]), .rectangle3_weight(rectangle3_weights[1224]), .feature_threshold(feature_thresholds[1224]), .feature_above(feature_aboves[1224]), .feature_below(feature_belows[1224]), .scan_win_std_dev(scan_win_std_dev[1224]), .feature_accum(feature_accums[1224]));
  accum_calculator ac1225(.scan_win(scan_win1225), .rectangle1_x(rectangle1_xs[1225]), .rectangle1_y(rectangle1_ys[1225]), .rectangle1_width(rectangle1_widths[1225]), .rectangle1_height(rectangle1_heights[1225]), .rectangle1_weight(rectangle1_weights[1225]), .rectangle2_x(rectangle2_xs[1225]), .rectangle2_y(rectangle2_ys[1225]), .rectangle2_width(rectangle2_widths[1225]), .rectangle2_height(rectangle2_heights[1225]), .rectangle2_weight(rectangle2_weights[1225]), .rectangle3_x(rectangle3_xs[1225]), .rectangle3_y(rectangle3_ys[1225]), .rectangle3_width(rectangle3_widths[1225]), .rectangle3_height(rectangle3_heights[1225]), .rectangle3_weight(rectangle3_weights[1225]), .feature_threshold(feature_thresholds[1225]), .feature_above(feature_aboves[1225]), .feature_below(feature_belows[1225]), .scan_win_std_dev(scan_win_std_dev[1225]), .feature_accum(feature_accums[1225]));
  accum_calculator ac1226(.scan_win(scan_win1226), .rectangle1_x(rectangle1_xs[1226]), .rectangle1_y(rectangle1_ys[1226]), .rectangle1_width(rectangle1_widths[1226]), .rectangle1_height(rectangle1_heights[1226]), .rectangle1_weight(rectangle1_weights[1226]), .rectangle2_x(rectangle2_xs[1226]), .rectangle2_y(rectangle2_ys[1226]), .rectangle2_width(rectangle2_widths[1226]), .rectangle2_height(rectangle2_heights[1226]), .rectangle2_weight(rectangle2_weights[1226]), .rectangle3_x(rectangle3_xs[1226]), .rectangle3_y(rectangle3_ys[1226]), .rectangle3_width(rectangle3_widths[1226]), .rectangle3_height(rectangle3_heights[1226]), .rectangle3_weight(rectangle3_weights[1226]), .feature_threshold(feature_thresholds[1226]), .feature_above(feature_aboves[1226]), .feature_below(feature_belows[1226]), .scan_win_std_dev(scan_win_std_dev[1226]), .feature_accum(feature_accums[1226]));
  accum_calculator ac1227(.scan_win(scan_win1227), .rectangle1_x(rectangle1_xs[1227]), .rectangle1_y(rectangle1_ys[1227]), .rectangle1_width(rectangle1_widths[1227]), .rectangle1_height(rectangle1_heights[1227]), .rectangle1_weight(rectangle1_weights[1227]), .rectangle2_x(rectangle2_xs[1227]), .rectangle2_y(rectangle2_ys[1227]), .rectangle2_width(rectangle2_widths[1227]), .rectangle2_height(rectangle2_heights[1227]), .rectangle2_weight(rectangle2_weights[1227]), .rectangle3_x(rectangle3_xs[1227]), .rectangle3_y(rectangle3_ys[1227]), .rectangle3_width(rectangle3_widths[1227]), .rectangle3_height(rectangle3_heights[1227]), .rectangle3_weight(rectangle3_weights[1227]), .feature_threshold(feature_thresholds[1227]), .feature_above(feature_aboves[1227]), .feature_below(feature_belows[1227]), .scan_win_std_dev(scan_win_std_dev[1227]), .feature_accum(feature_accums[1227]));
  accum_calculator ac1228(.scan_win(scan_win1228), .rectangle1_x(rectangle1_xs[1228]), .rectangle1_y(rectangle1_ys[1228]), .rectangle1_width(rectangle1_widths[1228]), .rectangle1_height(rectangle1_heights[1228]), .rectangle1_weight(rectangle1_weights[1228]), .rectangle2_x(rectangle2_xs[1228]), .rectangle2_y(rectangle2_ys[1228]), .rectangle2_width(rectangle2_widths[1228]), .rectangle2_height(rectangle2_heights[1228]), .rectangle2_weight(rectangle2_weights[1228]), .rectangle3_x(rectangle3_xs[1228]), .rectangle3_y(rectangle3_ys[1228]), .rectangle3_width(rectangle3_widths[1228]), .rectangle3_height(rectangle3_heights[1228]), .rectangle3_weight(rectangle3_weights[1228]), .feature_threshold(feature_thresholds[1228]), .feature_above(feature_aboves[1228]), .feature_below(feature_belows[1228]), .scan_win_std_dev(scan_win_std_dev[1228]), .feature_accum(feature_accums[1228]));
  accum_calculator ac1229(.scan_win(scan_win1229), .rectangle1_x(rectangle1_xs[1229]), .rectangle1_y(rectangle1_ys[1229]), .rectangle1_width(rectangle1_widths[1229]), .rectangle1_height(rectangle1_heights[1229]), .rectangle1_weight(rectangle1_weights[1229]), .rectangle2_x(rectangle2_xs[1229]), .rectangle2_y(rectangle2_ys[1229]), .rectangle2_width(rectangle2_widths[1229]), .rectangle2_height(rectangle2_heights[1229]), .rectangle2_weight(rectangle2_weights[1229]), .rectangle3_x(rectangle3_xs[1229]), .rectangle3_y(rectangle3_ys[1229]), .rectangle3_width(rectangle3_widths[1229]), .rectangle3_height(rectangle3_heights[1229]), .rectangle3_weight(rectangle3_weights[1229]), .feature_threshold(feature_thresholds[1229]), .feature_above(feature_aboves[1229]), .feature_below(feature_belows[1229]), .scan_win_std_dev(scan_win_std_dev[1229]), .feature_accum(feature_accums[1229]));
  accum_calculator ac1230(.scan_win(scan_win1230), .rectangle1_x(rectangle1_xs[1230]), .rectangle1_y(rectangle1_ys[1230]), .rectangle1_width(rectangle1_widths[1230]), .rectangle1_height(rectangle1_heights[1230]), .rectangle1_weight(rectangle1_weights[1230]), .rectangle2_x(rectangle2_xs[1230]), .rectangle2_y(rectangle2_ys[1230]), .rectangle2_width(rectangle2_widths[1230]), .rectangle2_height(rectangle2_heights[1230]), .rectangle2_weight(rectangle2_weights[1230]), .rectangle3_x(rectangle3_xs[1230]), .rectangle3_y(rectangle3_ys[1230]), .rectangle3_width(rectangle3_widths[1230]), .rectangle3_height(rectangle3_heights[1230]), .rectangle3_weight(rectangle3_weights[1230]), .feature_threshold(feature_thresholds[1230]), .feature_above(feature_aboves[1230]), .feature_below(feature_belows[1230]), .scan_win_std_dev(scan_win_std_dev[1230]), .feature_accum(feature_accums[1230]));
  accum_calculator ac1231(.scan_win(scan_win1231), .rectangle1_x(rectangle1_xs[1231]), .rectangle1_y(rectangle1_ys[1231]), .rectangle1_width(rectangle1_widths[1231]), .rectangle1_height(rectangle1_heights[1231]), .rectangle1_weight(rectangle1_weights[1231]), .rectangle2_x(rectangle2_xs[1231]), .rectangle2_y(rectangle2_ys[1231]), .rectangle2_width(rectangle2_widths[1231]), .rectangle2_height(rectangle2_heights[1231]), .rectangle2_weight(rectangle2_weights[1231]), .rectangle3_x(rectangle3_xs[1231]), .rectangle3_y(rectangle3_ys[1231]), .rectangle3_width(rectangle3_widths[1231]), .rectangle3_height(rectangle3_heights[1231]), .rectangle3_weight(rectangle3_weights[1231]), .feature_threshold(feature_thresholds[1231]), .feature_above(feature_aboves[1231]), .feature_below(feature_belows[1231]), .scan_win_std_dev(scan_win_std_dev[1231]), .feature_accum(feature_accums[1231]));
  accum_calculator ac1232(.scan_win(scan_win1232), .rectangle1_x(rectangle1_xs[1232]), .rectangle1_y(rectangle1_ys[1232]), .rectangle1_width(rectangle1_widths[1232]), .rectangle1_height(rectangle1_heights[1232]), .rectangle1_weight(rectangle1_weights[1232]), .rectangle2_x(rectangle2_xs[1232]), .rectangle2_y(rectangle2_ys[1232]), .rectangle2_width(rectangle2_widths[1232]), .rectangle2_height(rectangle2_heights[1232]), .rectangle2_weight(rectangle2_weights[1232]), .rectangle3_x(rectangle3_xs[1232]), .rectangle3_y(rectangle3_ys[1232]), .rectangle3_width(rectangle3_widths[1232]), .rectangle3_height(rectangle3_heights[1232]), .rectangle3_weight(rectangle3_weights[1232]), .feature_threshold(feature_thresholds[1232]), .feature_above(feature_aboves[1232]), .feature_below(feature_belows[1232]), .scan_win_std_dev(scan_win_std_dev[1232]), .feature_accum(feature_accums[1232]));
  accum_calculator ac1233(.scan_win(scan_win1233), .rectangle1_x(rectangle1_xs[1233]), .rectangle1_y(rectangle1_ys[1233]), .rectangle1_width(rectangle1_widths[1233]), .rectangle1_height(rectangle1_heights[1233]), .rectangle1_weight(rectangle1_weights[1233]), .rectangle2_x(rectangle2_xs[1233]), .rectangle2_y(rectangle2_ys[1233]), .rectangle2_width(rectangle2_widths[1233]), .rectangle2_height(rectangle2_heights[1233]), .rectangle2_weight(rectangle2_weights[1233]), .rectangle3_x(rectangle3_xs[1233]), .rectangle3_y(rectangle3_ys[1233]), .rectangle3_width(rectangle3_widths[1233]), .rectangle3_height(rectangle3_heights[1233]), .rectangle3_weight(rectangle3_weights[1233]), .feature_threshold(feature_thresholds[1233]), .feature_above(feature_aboves[1233]), .feature_below(feature_belows[1233]), .scan_win_std_dev(scan_win_std_dev[1233]), .feature_accum(feature_accums[1233]));
  accum_calculator ac1234(.scan_win(scan_win1234), .rectangle1_x(rectangle1_xs[1234]), .rectangle1_y(rectangle1_ys[1234]), .rectangle1_width(rectangle1_widths[1234]), .rectangle1_height(rectangle1_heights[1234]), .rectangle1_weight(rectangle1_weights[1234]), .rectangle2_x(rectangle2_xs[1234]), .rectangle2_y(rectangle2_ys[1234]), .rectangle2_width(rectangle2_widths[1234]), .rectangle2_height(rectangle2_heights[1234]), .rectangle2_weight(rectangle2_weights[1234]), .rectangle3_x(rectangle3_xs[1234]), .rectangle3_y(rectangle3_ys[1234]), .rectangle3_width(rectangle3_widths[1234]), .rectangle3_height(rectangle3_heights[1234]), .rectangle3_weight(rectangle3_weights[1234]), .feature_threshold(feature_thresholds[1234]), .feature_above(feature_aboves[1234]), .feature_below(feature_belows[1234]), .scan_win_std_dev(scan_win_std_dev[1234]), .feature_accum(feature_accums[1234]));
  accum_calculator ac1235(.scan_win(scan_win1235), .rectangle1_x(rectangle1_xs[1235]), .rectangle1_y(rectangle1_ys[1235]), .rectangle1_width(rectangle1_widths[1235]), .rectangle1_height(rectangle1_heights[1235]), .rectangle1_weight(rectangle1_weights[1235]), .rectangle2_x(rectangle2_xs[1235]), .rectangle2_y(rectangle2_ys[1235]), .rectangle2_width(rectangle2_widths[1235]), .rectangle2_height(rectangle2_heights[1235]), .rectangle2_weight(rectangle2_weights[1235]), .rectangle3_x(rectangle3_xs[1235]), .rectangle3_y(rectangle3_ys[1235]), .rectangle3_width(rectangle3_widths[1235]), .rectangle3_height(rectangle3_heights[1235]), .rectangle3_weight(rectangle3_weights[1235]), .feature_threshold(feature_thresholds[1235]), .feature_above(feature_aboves[1235]), .feature_below(feature_belows[1235]), .scan_win_std_dev(scan_win_std_dev[1235]), .feature_accum(feature_accums[1235]));
  accum_calculator ac1236(.scan_win(scan_win1236), .rectangle1_x(rectangle1_xs[1236]), .rectangle1_y(rectangle1_ys[1236]), .rectangle1_width(rectangle1_widths[1236]), .rectangle1_height(rectangle1_heights[1236]), .rectangle1_weight(rectangle1_weights[1236]), .rectangle2_x(rectangle2_xs[1236]), .rectangle2_y(rectangle2_ys[1236]), .rectangle2_width(rectangle2_widths[1236]), .rectangle2_height(rectangle2_heights[1236]), .rectangle2_weight(rectangle2_weights[1236]), .rectangle3_x(rectangle3_xs[1236]), .rectangle3_y(rectangle3_ys[1236]), .rectangle3_width(rectangle3_widths[1236]), .rectangle3_height(rectangle3_heights[1236]), .rectangle3_weight(rectangle3_weights[1236]), .feature_threshold(feature_thresholds[1236]), .feature_above(feature_aboves[1236]), .feature_below(feature_belows[1236]), .scan_win_std_dev(scan_win_std_dev[1236]), .feature_accum(feature_accums[1236]));
  accum_calculator ac1237(.scan_win(scan_win1237), .rectangle1_x(rectangle1_xs[1237]), .rectangle1_y(rectangle1_ys[1237]), .rectangle1_width(rectangle1_widths[1237]), .rectangle1_height(rectangle1_heights[1237]), .rectangle1_weight(rectangle1_weights[1237]), .rectangle2_x(rectangle2_xs[1237]), .rectangle2_y(rectangle2_ys[1237]), .rectangle2_width(rectangle2_widths[1237]), .rectangle2_height(rectangle2_heights[1237]), .rectangle2_weight(rectangle2_weights[1237]), .rectangle3_x(rectangle3_xs[1237]), .rectangle3_y(rectangle3_ys[1237]), .rectangle3_width(rectangle3_widths[1237]), .rectangle3_height(rectangle3_heights[1237]), .rectangle3_weight(rectangle3_weights[1237]), .feature_threshold(feature_thresholds[1237]), .feature_above(feature_aboves[1237]), .feature_below(feature_belows[1237]), .scan_win_std_dev(scan_win_std_dev[1237]), .feature_accum(feature_accums[1237]));
  accum_calculator ac1238(.scan_win(scan_win1238), .rectangle1_x(rectangle1_xs[1238]), .rectangle1_y(rectangle1_ys[1238]), .rectangle1_width(rectangle1_widths[1238]), .rectangle1_height(rectangle1_heights[1238]), .rectangle1_weight(rectangle1_weights[1238]), .rectangle2_x(rectangle2_xs[1238]), .rectangle2_y(rectangle2_ys[1238]), .rectangle2_width(rectangle2_widths[1238]), .rectangle2_height(rectangle2_heights[1238]), .rectangle2_weight(rectangle2_weights[1238]), .rectangle3_x(rectangle3_xs[1238]), .rectangle3_y(rectangle3_ys[1238]), .rectangle3_width(rectangle3_widths[1238]), .rectangle3_height(rectangle3_heights[1238]), .rectangle3_weight(rectangle3_weights[1238]), .feature_threshold(feature_thresholds[1238]), .feature_above(feature_aboves[1238]), .feature_below(feature_belows[1238]), .scan_win_std_dev(scan_win_std_dev[1238]), .feature_accum(feature_accums[1238]));
  accum_calculator ac1239(.scan_win(scan_win1239), .rectangle1_x(rectangle1_xs[1239]), .rectangle1_y(rectangle1_ys[1239]), .rectangle1_width(rectangle1_widths[1239]), .rectangle1_height(rectangle1_heights[1239]), .rectangle1_weight(rectangle1_weights[1239]), .rectangle2_x(rectangle2_xs[1239]), .rectangle2_y(rectangle2_ys[1239]), .rectangle2_width(rectangle2_widths[1239]), .rectangle2_height(rectangle2_heights[1239]), .rectangle2_weight(rectangle2_weights[1239]), .rectangle3_x(rectangle3_xs[1239]), .rectangle3_y(rectangle3_ys[1239]), .rectangle3_width(rectangle3_widths[1239]), .rectangle3_height(rectangle3_heights[1239]), .rectangle3_weight(rectangle3_weights[1239]), .feature_threshold(feature_thresholds[1239]), .feature_above(feature_aboves[1239]), .feature_below(feature_belows[1239]), .scan_win_std_dev(scan_win_std_dev[1239]), .feature_accum(feature_accums[1239]));
  accum_calculator ac1240(.scan_win(scan_win1240), .rectangle1_x(rectangle1_xs[1240]), .rectangle1_y(rectangle1_ys[1240]), .rectangle1_width(rectangle1_widths[1240]), .rectangle1_height(rectangle1_heights[1240]), .rectangle1_weight(rectangle1_weights[1240]), .rectangle2_x(rectangle2_xs[1240]), .rectangle2_y(rectangle2_ys[1240]), .rectangle2_width(rectangle2_widths[1240]), .rectangle2_height(rectangle2_heights[1240]), .rectangle2_weight(rectangle2_weights[1240]), .rectangle3_x(rectangle3_xs[1240]), .rectangle3_y(rectangle3_ys[1240]), .rectangle3_width(rectangle3_widths[1240]), .rectangle3_height(rectangle3_heights[1240]), .rectangle3_weight(rectangle3_weights[1240]), .feature_threshold(feature_thresholds[1240]), .feature_above(feature_aboves[1240]), .feature_below(feature_belows[1240]), .scan_win_std_dev(scan_win_std_dev[1240]), .feature_accum(feature_accums[1240]));
  accum_calculator ac1241(.scan_win(scan_win1241), .rectangle1_x(rectangle1_xs[1241]), .rectangle1_y(rectangle1_ys[1241]), .rectangle1_width(rectangle1_widths[1241]), .rectangle1_height(rectangle1_heights[1241]), .rectangle1_weight(rectangle1_weights[1241]), .rectangle2_x(rectangle2_xs[1241]), .rectangle2_y(rectangle2_ys[1241]), .rectangle2_width(rectangle2_widths[1241]), .rectangle2_height(rectangle2_heights[1241]), .rectangle2_weight(rectangle2_weights[1241]), .rectangle3_x(rectangle3_xs[1241]), .rectangle3_y(rectangle3_ys[1241]), .rectangle3_width(rectangle3_widths[1241]), .rectangle3_height(rectangle3_heights[1241]), .rectangle3_weight(rectangle3_weights[1241]), .feature_threshold(feature_thresholds[1241]), .feature_above(feature_aboves[1241]), .feature_below(feature_belows[1241]), .scan_win_std_dev(scan_win_std_dev[1241]), .feature_accum(feature_accums[1241]));
  accum_calculator ac1242(.scan_win(scan_win1242), .rectangle1_x(rectangle1_xs[1242]), .rectangle1_y(rectangle1_ys[1242]), .rectangle1_width(rectangle1_widths[1242]), .rectangle1_height(rectangle1_heights[1242]), .rectangle1_weight(rectangle1_weights[1242]), .rectangle2_x(rectangle2_xs[1242]), .rectangle2_y(rectangle2_ys[1242]), .rectangle2_width(rectangle2_widths[1242]), .rectangle2_height(rectangle2_heights[1242]), .rectangle2_weight(rectangle2_weights[1242]), .rectangle3_x(rectangle3_xs[1242]), .rectangle3_y(rectangle3_ys[1242]), .rectangle3_width(rectangle3_widths[1242]), .rectangle3_height(rectangle3_heights[1242]), .rectangle3_weight(rectangle3_weights[1242]), .feature_threshold(feature_thresholds[1242]), .feature_above(feature_aboves[1242]), .feature_below(feature_belows[1242]), .scan_win_std_dev(scan_win_std_dev[1242]), .feature_accum(feature_accums[1242]));
  accum_calculator ac1243(.scan_win(scan_win1243), .rectangle1_x(rectangle1_xs[1243]), .rectangle1_y(rectangle1_ys[1243]), .rectangle1_width(rectangle1_widths[1243]), .rectangle1_height(rectangle1_heights[1243]), .rectangle1_weight(rectangle1_weights[1243]), .rectangle2_x(rectangle2_xs[1243]), .rectangle2_y(rectangle2_ys[1243]), .rectangle2_width(rectangle2_widths[1243]), .rectangle2_height(rectangle2_heights[1243]), .rectangle2_weight(rectangle2_weights[1243]), .rectangle3_x(rectangle3_xs[1243]), .rectangle3_y(rectangle3_ys[1243]), .rectangle3_width(rectangle3_widths[1243]), .rectangle3_height(rectangle3_heights[1243]), .rectangle3_weight(rectangle3_weights[1243]), .feature_threshold(feature_thresholds[1243]), .feature_above(feature_aboves[1243]), .feature_below(feature_belows[1243]), .scan_win_std_dev(scan_win_std_dev[1243]), .feature_accum(feature_accums[1243]));
  accum_calculator ac1244(.scan_win(scan_win1244), .rectangle1_x(rectangle1_xs[1244]), .rectangle1_y(rectangle1_ys[1244]), .rectangle1_width(rectangle1_widths[1244]), .rectangle1_height(rectangle1_heights[1244]), .rectangle1_weight(rectangle1_weights[1244]), .rectangle2_x(rectangle2_xs[1244]), .rectangle2_y(rectangle2_ys[1244]), .rectangle2_width(rectangle2_widths[1244]), .rectangle2_height(rectangle2_heights[1244]), .rectangle2_weight(rectangle2_weights[1244]), .rectangle3_x(rectangle3_xs[1244]), .rectangle3_y(rectangle3_ys[1244]), .rectangle3_width(rectangle3_widths[1244]), .rectangle3_height(rectangle3_heights[1244]), .rectangle3_weight(rectangle3_weights[1244]), .feature_threshold(feature_thresholds[1244]), .feature_above(feature_aboves[1244]), .feature_below(feature_belows[1244]), .scan_win_std_dev(scan_win_std_dev[1244]), .feature_accum(feature_accums[1244]));
  accum_calculator ac1245(.scan_win(scan_win1245), .rectangle1_x(rectangle1_xs[1245]), .rectangle1_y(rectangle1_ys[1245]), .rectangle1_width(rectangle1_widths[1245]), .rectangle1_height(rectangle1_heights[1245]), .rectangle1_weight(rectangle1_weights[1245]), .rectangle2_x(rectangle2_xs[1245]), .rectangle2_y(rectangle2_ys[1245]), .rectangle2_width(rectangle2_widths[1245]), .rectangle2_height(rectangle2_heights[1245]), .rectangle2_weight(rectangle2_weights[1245]), .rectangle3_x(rectangle3_xs[1245]), .rectangle3_y(rectangle3_ys[1245]), .rectangle3_width(rectangle3_widths[1245]), .rectangle3_height(rectangle3_heights[1245]), .rectangle3_weight(rectangle3_weights[1245]), .feature_threshold(feature_thresholds[1245]), .feature_above(feature_aboves[1245]), .feature_below(feature_belows[1245]), .scan_win_std_dev(scan_win_std_dev[1245]), .feature_accum(feature_accums[1245]));
  accum_calculator ac1246(.scan_win(scan_win1246), .rectangle1_x(rectangle1_xs[1246]), .rectangle1_y(rectangle1_ys[1246]), .rectangle1_width(rectangle1_widths[1246]), .rectangle1_height(rectangle1_heights[1246]), .rectangle1_weight(rectangle1_weights[1246]), .rectangle2_x(rectangle2_xs[1246]), .rectangle2_y(rectangle2_ys[1246]), .rectangle2_width(rectangle2_widths[1246]), .rectangle2_height(rectangle2_heights[1246]), .rectangle2_weight(rectangle2_weights[1246]), .rectangle3_x(rectangle3_xs[1246]), .rectangle3_y(rectangle3_ys[1246]), .rectangle3_width(rectangle3_widths[1246]), .rectangle3_height(rectangle3_heights[1246]), .rectangle3_weight(rectangle3_weights[1246]), .feature_threshold(feature_thresholds[1246]), .feature_above(feature_aboves[1246]), .feature_below(feature_belows[1246]), .scan_win_std_dev(scan_win_std_dev[1246]), .feature_accum(feature_accums[1246]));
  accum_calculator ac1247(.scan_win(scan_win1247), .rectangle1_x(rectangle1_xs[1247]), .rectangle1_y(rectangle1_ys[1247]), .rectangle1_width(rectangle1_widths[1247]), .rectangle1_height(rectangle1_heights[1247]), .rectangle1_weight(rectangle1_weights[1247]), .rectangle2_x(rectangle2_xs[1247]), .rectangle2_y(rectangle2_ys[1247]), .rectangle2_width(rectangle2_widths[1247]), .rectangle2_height(rectangle2_heights[1247]), .rectangle2_weight(rectangle2_weights[1247]), .rectangle3_x(rectangle3_xs[1247]), .rectangle3_y(rectangle3_ys[1247]), .rectangle3_width(rectangle3_widths[1247]), .rectangle3_height(rectangle3_heights[1247]), .rectangle3_weight(rectangle3_weights[1247]), .feature_threshold(feature_thresholds[1247]), .feature_above(feature_aboves[1247]), .feature_below(feature_belows[1247]), .scan_win_std_dev(scan_win_std_dev[1247]), .feature_accum(feature_accums[1247]));
  accum_calculator ac1248(.scan_win(scan_win1248), .rectangle1_x(rectangle1_xs[1248]), .rectangle1_y(rectangle1_ys[1248]), .rectangle1_width(rectangle1_widths[1248]), .rectangle1_height(rectangle1_heights[1248]), .rectangle1_weight(rectangle1_weights[1248]), .rectangle2_x(rectangle2_xs[1248]), .rectangle2_y(rectangle2_ys[1248]), .rectangle2_width(rectangle2_widths[1248]), .rectangle2_height(rectangle2_heights[1248]), .rectangle2_weight(rectangle2_weights[1248]), .rectangle3_x(rectangle3_xs[1248]), .rectangle3_y(rectangle3_ys[1248]), .rectangle3_width(rectangle3_widths[1248]), .rectangle3_height(rectangle3_heights[1248]), .rectangle3_weight(rectangle3_weights[1248]), .feature_threshold(feature_thresholds[1248]), .feature_above(feature_aboves[1248]), .feature_below(feature_belows[1248]), .scan_win_std_dev(scan_win_std_dev[1248]), .feature_accum(feature_accums[1248]));
  accum_calculator ac1249(.scan_win(scan_win1249), .rectangle1_x(rectangle1_xs[1249]), .rectangle1_y(rectangle1_ys[1249]), .rectangle1_width(rectangle1_widths[1249]), .rectangle1_height(rectangle1_heights[1249]), .rectangle1_weight(rectangle1_weights[1249]), .rectangle2_x(rectangle2_xs[1249]), .rectangle2_y(rectangle2_ys[1249]), .rectangle2_width(rectangle2_widths[1249]), .rectangle2_height(rectangle2_heights[1249]), .rectangle2_weight(rectangle2_weights[1249]), .rectangle3_x(rectangle3_xs[1249]), .rectangle3_y(rectangle3_ys[1249]), .rectangle3_width(rectangle3_widths[1249]), .rectangle3_height(rectangle3_heights[1249]), .rectangle3_weight(rectangle3_weights[1249]), .feature_threshold(feature_thresholds[1249]), .feature_above(feature_aboves[1249]), .feature_below(feature_belows[1249]), .scan_win_std_dev(scan_win_std_dev[1249]), .feature_accum(feature_accums[1249]));
  accum_calculator ac1250(.scan_win(scan_win1250), .rectangle1_x(rectangle1_xs[1250]), .rectangle1_y(rectangle1_ys[1250]), .rectangle1_width(rectangle1_widths[1250]), .rectangle1_height(rectangle1_heights[1250]), .rectangle1_weight(rectangle1_weights[1250]), .rectangle2_x(rectangle2_xs[1250]), .rectangle2_y(rectangle2_ys[1250]), .rectangle2_width(rectangle2_widths[1250]), .rectangle2_height(rectangle2_heights[1250]), .rectangle2_weight(rectangle2_weights[1250]), .rectangle3_x(rectangle3_xs[1250]), .rectangle3_y(rectangle3_ys[1250]), .rectangle3_width(rectangle3_widths[1250]), .rectangle3_height(rectangle3_heights[1250]), .rectangle3_weight(rectangle3_weights[1250]), .feature_threshold(feature_thresholds[1250]), .feature_above(feature_aboves[1250]), .feature_below(feature_belows[1250]), .scan_win_std_dev(scan_win_std_dev[1250]), .feature_accum(feature_accums[1250]));
  accum_calculator ac1251(.scan_win(scan_win1251), .rectangle1_x(rectangle1_xs[1251]), .rectangle1_y(rectangle1_ys[1251]), .rectangle1_width(rectangle1_widths[1251]), .rectangle1_height(rectangle1_heights[1251]), .rectangle1_weight(rectangle1_weights[1251]), .rectangle2_x(rectangle2_xs[1251]), .rectangle2_y(rectangle2_ys[1251]), .rectangle2_width(rectangle2_widths[1251]), .rectangle2_height(rectangle2_heights[1251]), .rectangle2_weight(rectangle2_weights[1251]), .rectangle3_x(rectangle3_xs[1251]), .rectangle3_y(rectangle3_ys[1251]), .rectangle3_width(rectangle3_widths[1251]), .rectangle3_height(rectangle3_heights[1251]), .rectangle3_weight(rectangle3_weights[1251]), .feature_threshold(feature_thresholds[1251]), .feature_above(feature_aboves[1251]), .feature_below(feature_belows[1251]), .scan_win_std_dev(scan_win_std_dev[1251]), .feature_accum(feature_accums[1251]));
  accum_calculator ac1252(.scan_win(scan_win1252), .rectangle1_x(rectangle1_xs[1252]), .rectangle1_y(rectangle1_ys[1252]), .rectangle1_width(rectangle1_widths[1252]), .rectangle1_height(rectangle1_heights[1252]), .rectangle1_weight(rectangle1_weights[1252]), .rectangle2_x(rectangle2_xs[1252]), .rectangle2_y(rectangle2_ys[1252]), .rectangle2_width(rectangle2_widths[1252]), .rectangle2_height(rectangle2_heights[1252]), .rectangle2_weight(rectangle2_weights[1252]), .rectangle3_x(rectangle3_xs[1252]), .rectangle3_y(rectangle3_ys[1252]), .rectangle3_width(rectangle3_widths[1252]), .rectangle3_height(rectangle3_heights[1252]), .rectangle3_weight(rectangle3_weights[1252]), .feature_threshold(feature_thresholds[1252]), .feature_above(feature_aboves[1252]), .feature_below(feature_belows[1252]), .scan_win_std_dev(scan_win_std_dev[1252]), .feature_accum(feature_accums[1252]));
  accum_calculator ac1253(.scan_win(scan_win1253), .rectangle1_x(rectangle1_xs[1253]), .rectangle1_y(rectangle1_ys[1253]), .rectangle1_width(rectangle1_widths[1253]), .rectangle1_height(rectangle1_heights[1253]), .rectangle1_weight(rectangle1_weights[1253]), .rectangle2_x(rectangle2_xs[1253]), .rectangle2_y(rectangle2_ys[1253]), .rectangle2_width(rectangle2_widths[1253]), .rectangle2_height(rectangle2_heights[1253]), .rectangle2_weight(rectangle2_weights[1253]), .rectangle3_x(rectangle3_xs[1253]), .rectangle3_y(rectangle3_ys[1253]), .rectangle3_width(rectangle3_widths[1253]), .rectangle3_height(rectangle3_heights[1253]), .rectangle3_weight(rectangle3_weights[1253]), .feature_threshold(feature_thresholds[1253]), .feature_above(feature_aboves[1253]), .feature_below(feature_belows[1253]), .scan_win_std_dev(scan_win_std_dev[1253]), .feature_accum(feature_accums[1253]));
  accum_calculator ac1254(.scan_win(scan_win1254), .rectangle1_x(rectangle1_xs[1254]), .rectangle1_y(rectangle1_ys[1254]), .rectangle1_width(rectangle1_widths[1254]), .rectangle1_height(rectangle1_heights[1254]), .rectangle1_weight(rectangle1_weights[1254]), .rectangle2_x(rectangle2_xs[1254]), .rectangle2_y(rectangle2_ys[1254]), .rectangle2_width(rectangle2_widths[1254]), .rectangle2_height(rectangle2_heights[1254]), .rectangle2_weight(rectangle2_weights[1254]), .rectangle3_x(rectangle3_xs[1254]), .rectangle3_y(rectangle3_ys[1254]), .rectangle3_width(rectangle3_widths[1254]), .rectangle3_height(rectangle3_heights[1254]), .rectangle3_weight(rectangle3_weights[1254]), .feature_threshold(feature_thresholds[1254]), .feature_above(feature_aboves[1254]), .feature_below(feature_belows[1254]), .scan_win_std_dev(scan_win_std_dev[1254]), .feature_accum(feature_accums[1254]));
  accum_calculator ac1255(.scan_win(scan_win1255), .rectangle1_x(rectangle1_xs[1255]), .rectangle1_y(rectangle1_ys[1255]), .rectangle1_width(rectangle1_widths[1255]), .rectangle1_height(rectangle1_heights[1255]), .rectangle1_weight(rectangle1_weights[1255]), .rectangle2_x(rectangle2_xs[1255]), .rectangle2_y(rectangle2_ys[1255]), .rectangle2_width(rectangle2_widths[1255]), .rectangle2_height(rectangle2_heights[1255]), .rectangle2_weight(rectangle2_weights[1255]), .rectangle3_x(rectangle3_xs[1255]), .rectangle3_y(rectangle3_ys[1255]), .rectangle3_width(rectangle3_widths[1255]), .rectangle3_height(rectangle3_heights[1255]), .rectangle3_weight(rectangle3_weights[1255]), .feature_threshold(feature_thresholds[1255]), .feature_above(feature_aboves[1255]), .feature_below(feature_belows[1255]), .scan_win_std_dev(scan_win_std_dev[1255]), .feature_accum(feature_accums[1255]));
  accum_calculator ac1256(.scan_win(scan_win1256), .rectangle1_x(rectangle1_xs[1256]), .rectangle1_y(rectangle1_ys[1256]), .rectangle1_width(rectangle1_widths[1256]), .rectangle1_height(rectangle1_heights[1256]), .rectangle1_weight(rectangle1_weights[1256]), .rectangle2_x(rectangle2_xs[1256]), .rectangle2_y(rectangle2_ys[1256]), .rectangle2_width(rectangle2_widths[1256]), .rectangle2_height(rectangle2_heights[1256]), .rectangle2_weight(rectangle2_weights[1256]), .rectangle3_x(rectangle3_xs[1256]), .rectangle3_y(rectangle3_ys[1256]), .rectangle3_width(rectangle3_widths[1256]), .rectangle3_height(rectangle3_heights[1256]), .rectangle3_weight(rectangle3_weights[1256]), .feature_threshold(feature_thresholds[1256]), .feature_above(feature_aboves[1256]), .feature_below(feature_belows[1256]), .scan_win_std_dev(scan_win_std_dev[1256]), .feature_accum(feature_accums[1256]));
  accum_calculator ac1257(.scan_win(scan_win1257), .rectangle1_x(rectangle1_xs[1257]), .rectangle1_y(rectangle1_ys[1257]), .rectangle1_width(rectangle1_widths[1257]), .rectangle1_height(rectangle1_heights[1257]), .rectangle1_weight(rectangle1_weights[1257]), .rectangle2_x(rectangle2_xs[1257]), .rectangle2_y(rectangle2_ys[1257]), .rectangle2_width(rectangle2_widths[1257]), .rectangle2_height(rectangle2_heights[1257]), .rectangle2_weight(rectangle2_weights[1257]), .rectangle3_x(rectangle3_xs[1257]), .rectangle3_y(rectangle3_ys[1257]), .rectangle3_width(rectangle3_widths[1257]), .rectangle3_height(rectangle3_heights[1257]), .rectangle3_weight(rectangle3_weights[1257]), .feature_threshold(feature_thresholds[1257]), .feature_above(feature_aboves[1257]), .feature_below(feature_belows[1257]), .scan_win_std_dev(scan_win_std_dev[1257]), .feature_accum(feature_accums[1257]));
  accum_calculator ac1258(.scan_win(scan_win1258), .rectangle1_x(rectangle1_xs[1258]), .rectangle1_y(rectangle1_ys[1258]), .rectangle1_width(rectangle1_widths[1258]), .rectangle1_height(rectangle1_heights[1258]), .rectangle1_weight(rectangle1_weights[1258]), .rectangle2_x(rectangle2_xs[1258]), .rectangle2_y(rectangle2_ys[1258]), .rectangle2_width(rectangle2_widths[1258]), .rectangle2_height(rectangle2_heights[1258]), .rectangle2_weight(rectangle2_weights[1258]), .rectangle3_x(rectangle3_xs[1258]), .rectangle3_y(rectangle3_ys[1258]), .rectangle3_width(rectangle3_widths[1258]), .rectangle3_height(rectangle3_heights[1258]), .rectangle3_weight(rectangle3_weights[1258]), .feature_threshold(feature_thresholds[1258]), .feature_above(feature_aboves[1258]), .feature_below(feature_belows[1258]), .scan_win_std_dev(scan_win_std_dev[1258]), .feature_accum(feature_accums[1258]));
  accum_calculator ac1259(.scan_win(scan_win1259), .rectangle1_x(rectangle1_xs[1259]), .rectangle1_y(rectangle1_ys[1259]), .rectangle1_width(rectangle1_widths[1259]), .rectangle1_height(rectangle1_heights[1259]), .rectangle1_weight(rectangle1_weights[1259]), .rectangle2_x(rectangle2_xs[1259]), .rectangle2_y(rectangle2_ys[1259]), .rectangle2_width(rectangle2_widths[1259]), .rectangle2_height(rectangle2_heights[1259]), .rectangle2_weight(rectangle2_weights[1259]), .rectangle3_x(rectangle3_xs[1259]), .rectangle3_y(rectangle3_ys[1259]), .rectangle3_width(rectangle3_widths[1259]), .rectangle3_height(rectangle3_heights[1259]), .rectangle3_weight(rectangle3_weights[1259]), .feature_threshold(feature_thresholds[1259]), .feature_above(feature_aboves[1259]), .feature_below(feature_belows[1259]), .scan_win_std_dev(scan_win_std_dev[1259]), .feature_accum(feature_accums[1259]));
  accum_calculator ac1260(.scan_win(scan_win1260), .rectangle1_x(rectangle1_xs[1260]), .rectangle1_y(rectangle1_ys[1260]), .rectangle1_width(rectangle1_widths[1260]), .rectangle1_height(rectangle1_heights[1260]), .rectangle1_weight(rectangle1_weights[1260]), .rectangle2_x(rectangle2_xs[1260]), .rectangle2_y(rectangle2_ys[1260]), .rectangle2_width(rectangle2_widths[1260]), .rectangle2_height(rectangle2_heights[1260]), .rectangle2_weight(rectangle2_weights[1260]), .rectangle3_x(rectangle3_xs[1260]), .rectangle3_y(rectangle3_ys[1260]), .rectangle3_width(rectangle3_widths[1260]), .rectangle3_height(rectangle3_heights[1260]), .rectangle3_weight(rectangle3_weights[1260]), .feature_threshold(feature_thresholds[1260]), .feature_above(feature_aboves[1260]), .feature_below(feature_belows[1260]), .scan_win_std_dev(scan_win_std_dev[1260]), .feature_accum(feature_accums[1260]));
  accum_calculator ac1261(.scan_win(scan_win1261), .rectangle1_x(rectangle1_xs[1261]), .rectangle1_y(rectangle1_ys[1261]), .rectangle1_width(rectangle1_widths[1261]), .rectangle1_height(rectangle1_heights[1261]), .rectangle1_weight(rectangle1_weights[1261]), .rectangle2_x(rectangle2_xs[1261]), .rectangle2_y(rectangle2_ys[1261]), .rectangle2_width(rectangle2_widths[1261]), .rectangle2_height(rectangle2_heights[1261]), .rectangle2_weight(rectangle2_weights[1261]), .rectangle3_x(rectangle3_xs[1261]), .rectangle3_y(rectangle3_ys[1261]), .rectangle3_width(rectangle3_widths[1261]), .rectangle3_height(rectangle3_heights[1261]), .rectangle3_weight(rectangle3_weights[1261]), .feature_threshold(feature_thresholds[1261]), .feature_above(feature_aboves[1261]), .feature_below(feature_belows[1261]), .scan_win_std_dev(scan_win_std_dev[1261]), .feature_accum(feature_accums[1261]));
  accum_calculator ac1262(.scan_win(scan_win1262), .rectangle1_x(rectangle1_xs[1262]), .rectangle1_y(rectangle1_ys[1262]), .rectangle1_width(rectangle1_widths[1262]), .rectangle1_height(rectangle1_heights[1262]), .rectangle1_weight(rectangle1_weights[1262]), .rectangle2_x(rectangle2_xs[1262]), .rectangle2_y(rectangle2_ys[1262]), .rectangle2_width(rectangle2_widths[1262]), .rectangle2_height(rectangle2_heights[1262]), .rectangle2_weight(rectangle2_weights[1262]), .rectangle3_x(rectangle3_xs[1262]), .rectangle3_y(rectangle3_ys[1262]), .rectangle3_width(rectangle3_widths[1262]), .rectangle3_height(rectangle3_heights[1262]), .rectangle3_weight(rectangle3_weights[1262]), .feature_threshold(feature_thresholds[1262]), .feature_above(feature_aboves[1262]), .feature_below(feature_belows[1262]), .scan_win_std_dev(scan_win_std_dev[1262]), .feature_accum(feature_accums[1262]));
  accum_calculator ac1263(.scan_win(scan_win1263), .rectangle1_x(rectangle1_xs[1263]), .rectangle1_y(rectangle1_ys[1263]), .rectangle1_width(rectangle1_widths[1263]), .rectangle1_height(rectangle1_heights[1263]), .rectangle1_weight(rectangle1_weights[1263]), .rectangle2_x(rectangle2_xs[1263]), .rectangle2_y(rectangle2_ys[1263]), .rectangle2_width(rectangle2_widths[1263]), .rectangle2_height(rectangle2_heights[1263]), .rectangle2_weight(rectangle2_weights[1263]), .rectangle3_x(rectangle3_xs[1263]), .rectangle3_y(rectangle3_ys[1263]), .rectangle3_width(rectangle3_widths[1263]), .rectangle3_height(rectangle3_heights[1263]), .rectangle3_weight(rectangle3_weights[1263]), .feature_threshold(feature_thresholds[1263]), .feature_above(feature_aboves[1263]), .feature_below(feature_belows[1263]), .scan_win_std_dev(scan_win_std_dev[1263]), .feature_accum(feature_accums[1263]));
  accum_calculator ac1264(.scan_win(scan_win1264), .rectangle1_x(rectangle1_xs[1264]), .rectangle1_y(rectangle1_ys[1264]), .rectangle1_width(rectangle1_widths[1264]), .rectangle1_height(rectangle1_heights[1264]), .rectangle1_weight(rectangle1_weights[1264]), .rectangle2_x(rectangle2_xs[1264]), .rectangle2_y(rectangle2_ys[1264]), .rectangle2_width(rectangle2_widths[1264]), .rectangle2_height(rectangle2_heights[1264]), .rectangle2_weight(rectangle2_weights[1264]), .rectangle3_x(rectangle3_xs[1264]), .rectangle3_y(rectangle3_ys[1264]), .rectangle3_width(rectangle3_widths[1264]), .rectangle3_height(rectangle3_heights[1264]), .rectangle3_weight(rectangle3_weights[1264]), .feature_threshold(feature_thresholds[1264]), .feature_above(feature_aboves[1264]), .feature_below(feature_belows[1264]), .scan_win_std_dev(scan_win_std_dev[1264]), .feature_accum(feature_accums[1264]));
  accum_calculator ac1265(.scan_win(scan_win1265), .rectangle1_x(rectangle1_xs[1265]), .rectangle1_y(rectangle1_ys[1265]), .rectangle1_width(rectangle1_widths[1265]), .rectangle1_height(rectangle1_heights[1265]), .rectangle1_weight(rectangle1_weights[1265]), .rectangle2_x(rectangle2_xs[1265]), .rectangle2_y(rectangle2_ys[1265]), .rectangle2_width(rectangle2_widths[1265]), .rectangle2_height(rectangle2_heights[1265]), .rectangle2_weight(rectangle2_weights[1265]), .rectangle3_x(rectangle3_xs[1265]), .rectangle3_y(rectangle3_ys[1265]), .rectangle3_width(rectangle3_widths[1265]), .rectangle3_height(rectangle3_heights[1265]), .rectangle3_weight(rectangle3_weights[1265]), .feature_threshold(feature_thresholds[1265]), .feature_above(feature_aboves[1265]), .feature_below(feature_belows[1265]), .scan_win_std_dev(scan_win_std_dev[1265]), .feature_accum(feature_accums[1265]));
  accum_calculator ac1266(.scan_win(scan_win1266), .rectangle1_x(rectangle1_xs[1266]), .rectangle1_y(rectangle1_ys[1266]), .rectangle1_width(rectangle1_widths[1266]), .rectangle1_height(rectangle1_heights[1266]), .rectangle1_weight(rectangle1_weights[1266]), .rectangle2_x(rectangle2_xs[1266]), .rectangle2_y(rectangle2_ys[1266]), .rectangle2_width(rectangle2_widths[1266]), .rectangle2_height(rectangle2_heights[1266]), .rectangle2_weight(rectangle2_weights[1266]), .rectangle3_x(rectangle3_xs[1266]), .rectangle3_y(rectangle3_ys[1266]), .rectangle3_width(rectangle3_widths[1266]), .rectangle3_height(rectangle3_heights[1266]), .rectangle3_weight(rectangle3_weights[1266]), .feature_threshold(feature_thresholds[1266]), .feature_above(feature_aboves[1266]), .feature_below(feature_belows[1266]), .scan_win_std_dev(scan_win_std_dev[1266]), .feature_accum(feature_accums[1266]));
  accum_calculator ac1267(.scan_win(scan_win1267), .rectangle1_x(rectangle1_xs[1267]), .rectangle1_y(rectangle1_ys[1267]), .rectangle1_width(rectangle1_widths[1267]), .rectangle1_height(rectangle1_heights[1267]), .rectangle1_weight(rectangle1_weights[1267]), .rectangle2_x(rectangle2_xs[1267]), .rectangle2_y(rectangle2_ys[1267]), .rectangle2_width(rectangle2_widths[1267]), .rectangle2_height(rectangle2_heights[1267]), .rectangle2_weight(rectangle2_weights[1267]), .rectangle3_x(rectangle3_xs[1267]), .rectangle3_y(rectangle3_ys[1267]), .rectangle3_width(rectangle3_widths[1267]), .rectangle3_height(rectangle3_heights[1267]), .rectangle3_weight(rectangle3_weights[1267]), .feature_threshold(feature_thresholds[1267]), .feature_above(feature_aboves[1267]), .feature_below(feature_belows[1267]), .scan_win_std_dev(scan_win_std_dev[1267]), .feature_accum(feature_accums[1267]));
  accum_calculator ac1268(.scan_win(scan_win1268), .rectangle1_x(rectangle1_xs[1268]), .rectangle1_y(rectangle1_ys[1268]), .rectangle1_width(rectangle1_widths[1268]), .rectangle1_height(rectangle1_heights[1268]), .rectangle1_weight(rectangle1_weights[1268]), .rectangle2_x(rectangle2_xs[1268]), .rectangle2_y(rectangle2_ys[1268]), .rectangle2_width(rectangle2_widths[1268]), .rectangle2_height(rectangle2_heights[1268]), .rectangle2_weight(rectangle2_weights[1268]), .rectangle3_x(rectangle3_xs[1268]), .rectangle3_y(rectangle3_ys[1268]), .rectangle3_width(rectangle3_widths[1268]), .rectangle3_height(rectangle3_heights[1268]), .rectangle3_weight(rectangle3_weights[1268]), .feature_threshold(feature_thresholds[1268]), .feature_above(feature_aboves[1268]), .feature_below(feature_belows[1268]), .scan_win_std_dev(scan_win_std_dev[1268]), .feature_accum(feature_accums[1268]));
  accum_calculator ac1269(.scan_win(scan_win1269), .rectangle1_x(rectangle1_xs[1269]), .rectangle1_y(rectangle1_ys[1269]), .rectangle1_width(rectangle1_widths[1269]), .rectangle1_height(rectangle1_heights[1269]), .rectangle1_weight(rectangle1_weights[1269]), .rectangle2_x(rectangle2_xs[1269]), .rectangle2_y(rectangle2_ys[1269]), .rectangle2_width(rectangle2_widths[1269]), .rectangle2_height(rectangle2_heights[1269]), .rectangle2_weight(rectangle2_weights[1269]), .rectangle3_x(rectangle3_xs[1269]), .rectangle3_y(rectangle3_ys[1269]), .rectangle3_width(rectangle3_widths[1269]), .rectangle3_height(rectangle3_heights[1269]), .rectangle3_weight(rectangle3_weights[1269]), .feature_threshold(feature_thresholds[1269]), .feature_above(feature_aboves[1269]), .feature_below(feature_belows[1269]), .scan_win_std_dev(scan_win_std_dev[1269]), .feature_accum(feature_accums[1269]));
  accum_calculator ac1270(.scan_win(scan_win1270), .rectangle1_x(rectangle1_xs[1270]), .rectangle1_y(rectangle1_ys[1270]), .rectangle1_width(rectangle1_widths[1270]), .rectangle1_height(rectangle1_heights[1270]), .rectangle1_weight(rectangle1_weights[1270]), .rectangle2_x(rectangle2_xs[1270]), .rectangle2_y(rectangle2_ys[1270]), .rectangle2_width(rectangle2_widths[1270]), .rectangle2_height(rectangle2_heights[1270]), .rectangle2_weight(rectangle2_weights[1270]), .rectangle3_x(rectangle3_xs[1270]), .rectangle3_y(rectangle3_ys[1270]), .rectangle3_width(rectangle3_widths[1270]), .rectangle3_height(rectangle3_heights[1270]), .rectangle3_weight(rectangle3_weights[1270]), .feature_threshold(feature_thresholds[1270]), .feature_above(feature_aboves[1270]), .feature_below(feature_belows[1270]), .scan_win_std_dev(scan_win_std_dev[1270]), .feature_accum(feature_accums[1270]));
  accum_calculator ac1271(.scan_win(scan_win1271), .rectangle1_x(rectangle1_xs[1271]), .rectangle1_y(rectangle1_ys[1271]), .rectangle1_width(rectangle1_widths[1271]), .rectangle1_height(rectangle1_heights[1271]), .rectangle1_weight(rectangle1_weights[1271]), .rectangle2_x(rectangle2_xs[1271]), .rectangle2_y(rectangle2_ys[1271]), .rectangle2_width(rectangle2_widths[1271]), .rectangle2_height(rectangle2_heights[1271]), .rectangle2_weight(rectangle2_weights[1271]), .rectangle3_x(rectangle3_xs[1271]), .rectangle3_y(rectangle3_ys[1271]), .rectangle3_width(rectangle3_widths[1271]), .rectangle3_height(rectangle3_heights[1271]), .rectangle3_weight(rectangle3_weights[1271]), .feature_threshold(feature_thresholds[1271]), .feature_above(feature_aboves[1271]), .feature_below(feature_belows[1271]), .scan_win_std_dev(scan_win_std_dev[1271]), .feature_accum(feature_accums[1271]));
  accum_calculator ac1272(.scan_win(scan_win1272), .rectangle1_x(rectangle1_xs[1272]), .rectangle1_y(rectangle1_ys[1272]), .rectangle1_width(rectangle1_widths[1272]), .rectangle1_height(rectangle1_heights[1272]), .rectangle1_weight(rectangle1_weights[1272]), .rectangle2_x(rectangle2_xs[1272]), .rectangle2_y(rectangle2_ys[1272]), .rectangle2_width(rectangle2_widths[1272]), .rectangle2_height(rectangle2_heights[1272]), .rectangle2_weight(rectangle2_weights[1272]), .rectangle3_x(rectangle3_xs[1272]), .rectangle3_y(rectangle3_ys[1272]), .rectangle3_width(rectangle3_widths[1272]), .rectangle3_height(rectangle3_heights[1272]), .rectangle3_weight(rectangle3_weights[1272]), .feature_threshold(feature_thresholds[1272]), .feature_above(feature_aboves[1272]), .feature_below(feature_belows[1272]), .scan_win_std_dev(scan_win_std_dev[1272]), .feature_accum(feature_accums[1272]));
  accum_calculator ac1273(.scan_win(scan_win1273), .rectangle1_x(rectangle1_xs[1273]), .rectangle1_y(rectangle1_ys[1273]), .rectangle1_width(rectangle1_widths[1273]), .rectangle1_height(rectangle1_heights[1273]), .rectangle1_weight(rectangle1_weights[1273]), .rectangle2_x(rectangle2_xs[1273]), .rectangle2_y(rectangle2_ys[1273]), .rectangle2_width(rectangle2_widths[1273]), .rectangle2_height(rectangle2_heights[1273]), .rectangle2_weight(rectangle2_weights[1273]), .rectangle3_x(rectangle3_xs[1273]), .rectangle3_y(rectangle3_ys[1273]), .rectangle3_width(rectangle3_widths[1273]), .rectangle3_height(rectangle3_heights[1273]), .rectangle3_weight(rectangle3_weights[1273]), .feature_threshold(feature_thresholds[1273]), .feature_above(feature_aboves[1273]), .feature_below(feature_belows[1273]), .scan_win_std_dev(scan_win_std_dev[1273]), .feature_accum(feature_accums[1273]));
  accum_calculator ac1274(.scan_win(scan_win1274), .rectangle1_x(rectangle1_xs[1274]), .rectangle1_y(rectangle1_ys[1274]), .rectangle1_width(rectangle1_widths[1274]), .rectangle1_height(rectangle1_heights[1274]), .rectangle1_weight(rectangle1_weights[1274]), .rectangle2_x(rectangle2_xs[1274]), .rectangle2_y(rectangle2_ys[1274]), .rectangle2_width(rectangle2_widths[1274]), .rectangle2_height(rectangle2_heights[1274]), .rectangle2_weight(rectangle2_weights[1274]), .rectangle3_x(rectangle3_xs[1274]), .rectangle3_y(rectangle3_ys[1274]), .rectangle3_width(rectangle3_widths[1274]), .rectangle3_height(rectangle3_heights[1274]), .rectangle3_weight(rectangle3_weights[1274]), .feature_threshold(feature_thresholds[1274]), .feature_above(feature_aboves[1274]), .feature_below(feature_belows[1274]), .scan_win_std_dev(scan_win_std_dev[1274]), .feature_accum(feature_accums[1274]));
  accum_calculator ac1275(.scan_win(scan_win1275), .rectangle1_x(rectangle1_xs[1275]), .rectangle1_y(rectangle1_ys[1275]), .rectangle1_width(rectangle1_widths[1275]), .rectangle1_height(rectangle1_heights[1275]), .rectangle1_weight(rectangle1_weights[1275]), .rectangle2_x(rectangle2_xs[1275]), .rectangle2_y(rectangle2_ys[1275]), .rectangle2_width(rectangle2_widths[1275]), .rectangle2_height(rectangle2_heights[1275]), .rectangle2_weight(rectangle2_weights[1275]), .rectangle3_x(rectangle3_xs[1275]), .rectangle3_y(rectangle3_ys[1275]), .rectangle3_width(rectangle3_widths[1275]), .rectangle3_height(rectangle3_heights[1275]), .rectangle3_weight(rectangle3_weights[1275]), .feature_threshold(feature_thresholds[1275]), .feature_above(feature_aboves[1275]), .feature_below(feature_belows[1275]), .scan_win_std_dev(scan_win_std_dev[1275]), .feature_accum(feature_accums[1275]));
  accum_calculator ac1276(.scan_win(scan_win1276), .rectangle1_x(rectangle1_xs[1276]), .rectangle1_y(rectangle1_ys[1276]), .rectangle1_width(rectangle1_widths[1276]), .rectangle1_height(rectangle1_heights[1276]), .rectangle1_weight(rectangle1_weights[1276]), .rectangle2_x(rectangle2_xs[1276]), .rectangle2_y(rectangle2_ys[1276]), .rectangle2_width(rectangle2_widths[1276]), .rectangle2_height(rectangle2_heights[1276]), .rectangle2_weight(rectangle2_weights[1276]), .rectangle3_x(rectangle3_xs[1276]), .rectangle3_y(rectangle3_ys[1276]), .rectangle3_width(rectangle3_widths[1276]), .rectangle3_height(rectangle3_heights[1276]), .rectangle3_weight(rectangle3_weights[1276]), .feature_threshold(feature_thresholds[1276]), .feature_above(feature_aboves[1276]), .feature_below(feature_belows[1276]), .scan_win_std_dev(scan_win_std_dev[1276]), .feature_accum(feature_accums[1276]));
  accum_calculator ac1277(.scan_win(scan_win1277), .rectangle1_x(rectangle1_xs[1277]), .rectangle1_y(rectangle1_ys[1277]), .rectangle1_width(rectangle1_widths[1277]), .rectangle1_height(rectangle1_heights[1277]), .rectangle1_weight(rectangle1_weights[1277]), .rectangle2_x(rectangle2_xs[1277]), .rectangle2_y(rectangle2_ys[1277]), .rectangle2_width(rectangle2_widths[1277]), .rectangle2_height(rectangle2_heights[1277]), .rectangle2_weight(rectangle2_weights[1277]), .rectangle3_x(rectangle3_xs[1277]), .rectangle3_y(rectangle3_ys[1277]), .rectangle3_width(rectangle3_widths[1277]), .rectangle3_height(rectangle3_heights[1277]), .rectangle3_weight(rectangle3_weights[1277]), .feature_threshold(feature_thresholds[1277]), .feature_above(feature_aboves[1277]), .feature_below(feature_belows[1277]), .scan_win_std_dev(scan_win_std_dev[1277]), .feature_accum(feature_accums[1277]));
  accum_calculator ac1278(.scan_win(scan_win1278), .rectangle1_x(rectangle1_xs[1278]), .rectangle1_y(rectangle1_ys[1278]), .rectangle1_width(rectangle1_widths[1278]), .rectangle1_height(rectangle1_heights[1278]), .rectangle1_weight(rectangle1_weights[1278]), .rectangle2_x(rectangle2_xs[1278]), .rectangle2_y(rectangle2_ys[1278]), .rectangle2_width(rectangle2_widths[1278]), .rectangle2_height(rectangle2_heights[1278]), .rectangle2_weight(rectangle2_weights[1278]), .rectangle3_x(rectangle3_xs[1278]), .rectangle3_y(rectangle3_ys[1278]), .rectangle3_width(rectangle3_widths[1278]), .rectangle3_height(rectangle3_heights[1278]), .rectangle3_weight(rectangle3_weights[1278]), .feature_threshold(feature_thresholds[1278]), .feature_above(feature_aboves[1278]), .feature_below(feature_belows[1278]), .scan_win_std_dev(scan_win_std_dev[1278]), .feature_accum(feature_accums[1278]));
  accum_calculator ac1279(.scan_win(scan_win1279), .rectangle1_x(rectangle1_xs[1279]), .rectangle1_y(rectangle1_ys[1279]), .rectangle1_width(rectangle1_widths[1279]), .rectangle1_height(rectangle1_heights[1279]), .rectangle1_weight(rectangle1_weights[1279]), .rectangle2_x(rectangle2_xs[1279]), .rectangle2_y(rectangle2_ys[1279]), .rectangle2_width(rectangle2_widths[1279]), .rectangle2_height(rectangle2_heights[1279]), .rectangle2_weight(rectangle2_weights[1279]), .rectangle3_x(rectangle3_xs[1279]), .rectangle3_y(rectangle3_ys[1279]), .rectangle3_width(rectangle3_widths[1279]), .rectangle3_height(rectangle3_heights[1279]), .rectangle3_weight(rectangle3_weights[1279]), .feature_threshold(feature_thresholds[1279]), .feature_above(feature_aboves[1279]), .feature_below(feature_belows[1279]), .scan_win_std_dev(scan_win_std_dev[1279]), .feature_accum(feature_accums[1279]));
  accum_calculator ac1280(.scan_win(scan_win1280), .rectangle1_x(rectangle1_xs[1280]), .rectangle1_y(rectangle1_ys[1280]), .rectangle1_width(rectangle1_widths[1280]), .rectangle1_height(rectangle1_heights[1280]), .rectangle1_weight(rectangle1_weights[1280]), .rectangle2_x(rectangle2_xs[1280]), .rectangle2_y(rectangle2_ys[1280]), .rectangle2_width(rectangle2_widths[1280]), .rectangle2_height(rectangle2_heights[1280]), .rectangle2_weight(rectangle2_weights[1280]), .rectangle3_x(rectangle3_xs[1280]), .rectangle3_y(rectangle3_ys[1280]), .rectangle3_width(rectangle3_widths[1280]), .rectangle3_height(rectangle3_heights[1280]), .rectangle3_weight(rectangle3_weights[1280]), .feature_threshold(feature_thresholds[1280]), .feature_above(feature_aboves[1280]), .feature_below(feature_belows[1280]), .scan_win_std_dev(scan_win_std_dev[1280]), .feature_accum(feature_accums[1280]));
  accum_calculator ac1281(.scan_win(scan_win1281), .rectangle1_x(rectangle1_xs[1281]), .rectangle1_y(rectangle1_ys[1281]), .rectangle1_width(rectangle1_widths[1281]), .rectangle1_height(rectangle1_heights[1281]), .rectangle1_weight(rectangle1_weights[1281]), .rectangle2_x(rectangle2_xs[1281]), .rectangle2_y(rectangle2_ys[1281]), .rectangle2_width(rectangle2_widths[1281]), .rectangle2_height(rectangle2_heights[1281]), .rectangle2_weight(rectangle2_weights[1281]), .rectangle3_x(rectangle3_xs[1281]), .rectangle3_y(rectangle3_ys[1281]), .rectangle3_width(rectangle3_widths[1281]), .rectangle3_height(rectangle3_heights[1281]), .rectangle3_weight(rectangle3_weights[1281]), .feature_threshold(feature_thresholds[1281]), .feature_above(feature_aboves[1281]), .feature_below(feature_belows[1281]), .scan_win_std_dev(scan_win_std_dev[1281]), .feature_accum(feature_accums[1281]));
  accum_calculator ac1282(.scan_win(scan_win1282), .rectangle1_x(rectangle1_xs[1282]), .rectangle1_y(rectangle1_ys[1282]), .rectangle1_width(rectangle1_widths[1282]), .rectangle1_height(rectangle1_heights[1282]), .rectangle1_weight(rectangle1_weights[1282]), .rectangle2_x(rectangle2_xs[1282]), .rectangle2_y(rectangle2_ys[1282]), .rectangle2_width(rectangle2_widths[1282]), .rectangle2_height(rectangle2_heights[1282]), .rectangle2_weight(rectangle2_weights[1282]), .rectangle3_x(rectangle3_xs[1282]), .rectangle3_y(rectangle3_ys[1282]), .rectangle3_width(rectangle3_widths[1282]), .rectangle3_height(rectangle3_heights[1282]), .rectangle3_weight(rectangle3_weights[1282]), .feature_threshold(feature_thresholds[1282]), .feature_above(feature_aboves[1282]), .feature_below(feature_belows[1282]), .scan_win_std_dev(scan_win_std_dev[1282]), .feature_accum(feature_accums[1282]));
  accum_calculator ac1283(.scan_win(scan_win1283), .rectangle1_x(rectangle1_xs[1283]), .rectangle1_y(rectangle1_ys[1283]), .rectangle1_width(rectangle1_widths[1283]), .rectangle1_height(rectangle1_heights[1283]), .rectangle1_weight(rectangle1_weights[1283]), .rectangle2_x(rectangle2_xs[1283]), .rectangle2_y(rectangle2_ys[1283]), .rectangle2_width(rectangle2_widths[1283]), .rectangle2_height(rectangle2_heights[1283]), .rectangle2_weight(rectangle2_weights[1283]), .rectangle3_x(rectangle3_xs[1283]), .rectangle3_y(rectangle3_ys[1283]), .rectangle3_width(rectangle3_widths[1283]), .rectangle3_height(rectangle3_heights[1283]), .rectangle3_weight(rectangle3_weights[1283]), .feature_threshold(feature_thresholds[1283]), .feature_above(feature_aboves[1283]), .feature_below(feature_belows[1283]), .scan_win_std_dev(scan_win_std_dev[1283]), .feature_accum(feature_accums[1283]));
  accum_calculator ac1284(.scan_win(scan_win1284), .rectangle1_x(rectangle1_xs[1284]), .rectangle1_y(rectangle1_ys[1284]), .rectangle1_width(rectangle1_widths[1284]), .rectangle1_height(rectangle1_heights[1284]), .rectangle1_weight(rectangle1_weights[1284]), .rectangle2_x(rectangle2_xs[1284]), .rectangle2_y(rectangle2_ys[1284]), .rectangle2_width(rectangle2_widths[1284]), .rectangle2_height(rectangle2_heights[1284]), .rectangle2_weight(rectangle2_weights[1284]), .rectangle3_x(rectangle3_xs[1284]), .rectangle3_y(rectangle3_ys[1284]), .rectangle3_width(rectangle3_widths[1284]), .rectangle3_height(rectangle3_heights[1284]), .rectangle3_weight(rectangle3_weights[1284]), .feature_threshold(feature_thresholds[1284]), .feature_above(feature_aboves[1284]), .feature_below(feature_belows[1284]), .scan_win_std_dev(scan_win_std_dev[1284]), .feature_accum(feature_accums[1284]));
  accum_calculator ac1285(.scan_win(scan_win1285), .rectangle1_x(rectangle1_xs[1285]), .rectangle1_y(rectangle1_ys[1285]), .rectangle1_width(rectangle1_widths[1285]), .rectangle1_height(rectangle1_heights[1285]), .rectangle1_weight(rectangle1_weights[1285]), .rectangle2_x(rectangle2_xs[1285]), .rectangle2_y(rectangle2_ys[1285]), .rectangle2_width(rectangle2_widths[1285]), .rectangle2_height(rectangle2_heights[1285]), .rectangle2_weight(rectangle2_weights[1285]), .rectangle3_x(rectangle3_xs[1285]), .rectangle3_y(rectangle3_ys[1285]), .rectangle3_width(rectangle3_widths[1285]), .rectangle3_height(rectangle3_heights[1285]), .rectangle3_weight(rectangle3_weights[1285]), .feature_threshold(feature_thresholds[1285]), .feature_above(feature_aboves[1285]), .feature_below(feature_belows[1285]), .scan_win_std_dev(scan_win_std_dev[1285]), .feature_accum(feature_accums[1285]));
  accum_calculator ac1286(.scan_win(scan_win1286), .rectangle1_x(rectangle1_xs[1286]), .rectangle1_y(rectangle1_ys[1286]), .rectangle1_width(rectangle1_widths[1286]), .rectangle1_height(rectangle1_heights[1286]), .rectangle1_weight(rectangle1_weights[1286]), .rectangle2_x(rectangle2_xs[1286]), .rectangle2_y(rectangle2_ys[1286]), .rectangle2_width(rectangle2_widths[1286]), .rectangle2_height(rectangle2_heights[1286]), .rectangle2_weight(rectangle2_weights[1286]), .rectangle3_x(rectangle3_xs[1286]), .rectangle3_y(rectangle3_ys[1286]), .rectangle3_width(rectangle3_widths[1286]), .rectangle3_height(rectangle3_heights[1286]), .rectangle3_weight(rectangle3_weights[1286]), .feature_threshold(feature_thresholds[1286]), .feature_above(feature_aboves[1286]), .feature_below(feature_belows[1286]), .scan_win_std_dev(scan_win_std_dev[1286]), .feature_accum(feature_accums[1286]));
  accum_calculator ac1287(.scan_win(scan_win1287), .rectangle1_x(rectangle1_xs[1287]), .rectangle1_y(rectangle1_ys[1287]), .rectangle1_width(rectangle1_widths[1287]), .rectangle1_height(rectangle1_heights[1287]), .rectangle1_weight(rectangle1_weights[1287]), .rectangle2_x(rectangle2_xs[1287]), .rectangle2_y(rectangle2_ys[1287]), .rectangle2_width(rectangle2_widths[1287]), .rectangle2_height(rectangle2_heights[1287]), .rectangle2_weight(rectangle2_weights[1287]), .rectangle3_x(rectangle3_xs[1287]), .rectangle3_y(rectangle3_ys[1287]), .rectangle3_width(rectangle3_widths[1287]), .rectangle3_height(rectangle3_heights[1287]), .rectangle3_weight(rectangle3_weights[1287]), .feature_threshold(feature_thresholds[1287]), .feature_above(feature_aboves[1287]), .feature_below(feature_belows[1287]), .scan_win_std_dev(scan_win_std_dev[1287]), .feature_accum(feature_accums[1287]));
  accum_calculator ac1288(.scan_win(scan_win1288), .rectangle1_x(rectangle1_xs[1288]), .rectangle1_y(rectangle1_ys[1288]), .rectangle1_width(rectangle1_widths[1288]), .rectangle1_height(rectangle1_heights[1288]), .rectangle1_weight(rectangle1_weights[1288]), .rectangle2_x(rectangle2_xs[1288]), .rectangle2_y(rectangle2_ys[1288]), .rectangle2_width(rectangle2_widths[1288]), .rectangle2_height(rectangle2_heights[1288]), .rectangle2_weight(rectangle2_weights[1288]), .rectangle3_x(rectangle3_xs[1288]), .rectangle3_y(rectangle3_ys[1288]), .rectangle3_width(rectangle3_widths[1288]), .rectangle3_height(rectangle3_heights[1288]), .rectangle3_weight(rectangle3_weights[1288]), .feature_threshold(feature_thresholds[1288]), .feature_above(feature_aboves[1288]), .feature_below(feature_belows[1288]), .scan_win_std_dev(scan_win_std_dev[1288]), .feature_accum(feature_accums[1288]));
  accum_calculator ac1289(.scan_win(scan_win1289), .rectangle1_x(rectangle1_xs[1289]), .rectangle1_y(rectangle1_ys[1289]), .rectangle1_width(rectangle1_widths[1289]), .rectangle1_height(rectangle1_heights[1289]), .rectangle1_weight(rectangle1_weights[1289]), .rectangle2_x(rectangle2_xs[1289]), .rectangle2_y(rectangle2_ys[1289]), .rectangle2_width(rectangle2_widths[1289]), .rectangle2_height(rectangle2_heights[1289]), .rectangle2_weight(rectangle2_weights[1289]), .rectangle3_x(rectangle3_xs[1289]), .rectangle3_y(rectangle3_ys[1289]), .rectangle3_width(rectangle3_widths[1289]), .rectangle3_height(rectangle3_heights[1289]), .rectangle3_weight(rectangle3_weights[1289]), .feature_threshold(feature_thresholds[1289]), .feature_above(feature_aboves[1289]), .feature_below(feature_belows[1289]), .scan_win_std_dev(scan_win_std_dev[1289]), .feature_accum(feature_accums[1289]));
  accum_calculator ac1290(.scan_win(scan_win1290), .rectangle1_x(rectangle1_xs[1290]), .rectangle1_y(rectangle1_ys[1290]), .rectangle1_width(rectangle1_widths[1290]), .rectangle1_height(rectangle1_heights[1290]), .rectangle1_weight(rectangle1_weights[1290]), .rectangle2_x(rectangle2_xs[1290]), .rectangle2_y(rectangle2_ys[1290]), .rectangle2_width(rectangle2_widths[1290]), .rectangle2_height(rectangle2_heights[1290]), .rectangle2_weight(rectangle2_weights[1290]), .rectangle3_x(rectangle3_xs[1290]), .rectangle3_y(rectangle3_ys[1290]), .rectangle3_width(rectangle3_widths[1290]), .rectangle3_height(rectangle3_heights[1290]), .rectangle3_weight(rectangle3_weights[1290]), .feature_threshold(feature_thresholds[1290]), .feature_above(feature_aboves[1290]), .feature_below(feature_belows[1290]), .scan_win_std_dev(scan_win_std_dev[1290]), .feature_accum(feature_accums[1290]));
  accum_calculator ac1291(.scan_win(scan_win1291), .rectangle1_x(rectangle1_xs[1291]), .rectangle1_y(rectangle1_ys[1291]), .rectangle1_width(rectangle1_widths[1291]), .rectangle1_height(rectangle1_heights[1291]), .rectangle1_weight(rectangle1_weights[1291]), .rectangle2_x(rectangle2_xs[1291]), .rectangle2_y(rectangle2_ys[1291]), .rectangle2_width(rectangle2_widths[1291]), .rectangle2_height(rectangle2_heights[1291]), .rectangle2_weight(rectangle2_weights[1291]), .rectangle3_x(rectangle3_xs[1291]), .rectangle3_y(rectangle3_ys[1291]), .rectangle3_width(rectangle3_widths[1291]), .rectangle3_height(rectangle3_heights[1291]), .rectangle3_weight(rectangle3_weights[1291]), .feature_threshold(feature_thresholds[1291]), .feature_above(feature_aboves[1291]), .feature_below(feature_belows[1291]), .scan_win_std_dev(scan_win_std_dev[1291]), .feature_accum(feature_accums[1291]));
  accum_calculator ac1292(.scan_win(scan_win1292), .rectangle1_x(rectangle1_xs[1292]), .rectangle1_y(rectangle1_ys[1292]), .rectangle1_width(rectangle1_widths[1292]), .rectangle1_height(rectangle1_heights[1292]), .rectangle1_weight(rectangle1_weights[1292]), .rectangle2_x(rectangle2_xs[1292]), .rectangle2_y(rectangle2_ys[1292]), .rectangle2_width(rectangle2_widths[1292]), .rectangle2_height(rectangle2_heights[1292]), .rectangle2_weight(rectangle2_weights[1292]), .rectangle3_x(rectangle3_xs[1292]), .rectangle3_y(rectangle3_ys[1292]), .rectangle3_width(rectangle3_widths[1292]), .rectangle3_height(rectangle3_heights[1292]), .rectangle3_weight(rectangle3_weights[1292]), .feature_threshold(feature_thresholds[1292]), .feature_above(feature_aboves[1292]), .feature_below(feature_belows[1292]), .scan_win_std_dev(scan_win_std_dev[1292]), .feature_accum(feature_accums[1292]));
  accum_calculator ac1293(.scan_win(scan_win1293), .rectangle1_x(rectangle1_xs[1293]), .rectangle1_y(rectangle1_ys[1293]), .rectangle1_width(rectangle1_widths[1293]), .rectangle1_height(rectangle1_heights[1293]), .rectangle1_weight(rectangle1_weights[1293]), .rectangle2_x(rectangle2_xs[1293]), .rectangle2_y(rectangle2_ys[1293]), .rectangle2_width(rectangle2_widths[1293]), .rectangle2_height(rectangle2_heights[1293]), .rectangle2_weight(rectangle2_weights[1293]), .rectangle3_x(rectangle3_xs[1293]), .rectangle3_y(rectangle3_ys[1293]), .rectangle3_width(rectangle3_widths[1293]), .rectangle3_height(rectangle3_heights[1293]), .rectangle3_weight(rectangle3_weights[1293]), .feature_threshold(feature_thresholds[1293]), .feature_above(feature_aboves[1293]), .feature_below(feature_belows[1293]), .scan_win_std_dev(scan_win_std_dev[1293]), .feature_accum(feature_accums[1293]));
  accum_calculator ac1294(.scan_win(scan_win1294), .rectangle1_x(rectangle1_xs[1294]), .rectangle1_y(rectangle1_ys[1294]), .rectangle1_width(rectangle1_widths[1294]), .rectangle1_height(rectangle1_heights[1294]), .rectangle1_weight(rectangle1_weights[1294]), .rectangle2_x(rectangle2_xs[1294]), .rectangle2_y(rectangle2_ys[1294]), .rectangle2_width(rectangle2_widths[1294]), .rectangle2_height(rectangle2_heights[1294]), .rectangle2_weight(rectangle2_weights[1294]), .rectangle3_x(rectangle3_xs[1294]), .rectangle3_y(rectangle3_ys[1294]), .rectangle3_width(rectangle3_widths[1294]), .rectangle3_height(rectangle3_heights[1294]), .rectangle3_weight(rectangle3_weights[1294]), .feature_threshold(feature_thresholds[1294]), .feature_above(feature_aboves[1294]), .feature_below(feature_belows[1294]), .scan_win_std_dev(scan_win_std_dev[1294]), .feature_accum(feature_accums[1294]));
  accum_calculator ac1295(.scan_win(scan_win1295), .rectangle1_x(rectangle1_xs[1295]), .rectangle1_y(rectangle1_ys[1295]), .rectangle1_width(rectangle1_widths[1295]), .rectangle1_height(rectangle1_heights[1295]), .rectangle1_weight(rectangle1_weights[1295]), .rectangle2_x(rectangle2_xs[1295]), .rectangle2_y(rectangle2_ys[1295]), .rectangle2_width(rectangle2_widths[1295]), .rectangle2_height(rectangle2_heights[1295]), .rectangle2_weight(rectangle2_weights[1295]), .rectangle3_x(rectangle3_xs[1295]), .rectangle3_y(rectangle3_ys[1295]), .rectangle3_width(rectangle3_widths[1295]), .rectangle3_height(rectangle3_heights[1295]), .rectangle3_weight(rectangle3_weights[1295]), .feature_threshold(feature_thresholds[1295]), .feature_above(feature_aboves[1295]), .feature_below(feature_belows[1295]), .scan_win_std_dev(scan_win_std_dev[1295]), .feature_accum(feature_accums[1295]));
  accum_calculator ac1296(.scan_win(scan_win1296), .rectangle1_x(rectangle1_xs[1296]), .rectangle1_y(rectangle1_ys[1296]), .rectangle1_width(rectangle1_widths[1296]), .rectangle1_height(rectangle1_heights[1296]), .rectangle1_weight(rectangle1_weights[1296]), .rectangle2_x(rectangle2_xs[1296]), .rectangle2_y(rectangle2_ys[1296]), .rectangle2_width(rectangle2_widths[1296]), .rectangle2_height(rectangle2_heights[1296]), .rectangle2_weight(rectangle2_weights[1296]), .rectangle3_x(rectangle3_xs[1296]), .rectangle3_y(rectangle3_ys[1296]), .rectangle3_width(rectangle3_widths[1296]), .rectangle3_height(rectangle3_heights[1296]), .rectangle3_weight(rectangle3_weights[1296]), .feature_threshold(feature_thresholds[1296]), .feature_above(feature_aboves[1296]), .feature_below(feature_belows[1296]), .scan_win_std_dev(scan_win_std_dev[1296]), .feature_accum(feature_accums[1296]));
  accum_calculator ac1297(.scan_win(scan_win1297), .rectangle1_x(rectangle1_xs[1297]), .rectangle1_y(rectangle1_ys[1297]), .rectangle1_width(rectangle1_widths[1297]), .rectangle1_height(rectangle1_heights[1297]), .rectangle1_weight(rectangle1_weights[1297]), .rectangle2_x(rectangle2_xs[1297]), .rectangle2_y(rectangle2_ys[1297]), .rectangle2_width(rectangle2_widths[1297]), .rectangle2_height(rectangle2_heights[1297]), .rectangle2_weight(rectangle2_weights[1297]), .rectangle3_x(rectangle3_xs[1297]), .rectangle3_y(rectangle3_ys[1297]), .rectangle3_width(rectangle3_widths[1297]), .rectangle3_height(rectangle3_heights[1297]), .rectangle3_weight(rectangle3_weights[1297]), .feature_threshold(feature_thresholds[1297]), .feature_above(feature_aboves[1297]), .feature_below(feature_belows[1297]), .scan_win_std_dev(scan_win_std_dev[1297]), .feature_accum(feature_accums[1297]));
  accum_calculator ac1298(.scan_win(scan_win1298), .rectangle1_x(rectangle1_xs[1298]), .rectangle1_y(rectangle1_ys[1298]), .rectangle1_width(rectangle1_widths[1298]), .rectangle1_height(rectangle1_heights[1298]), .rectangle1_weight(rectangle1_weights[1298]), .rectangle2_x(rectangle2_xs[1298]), .rectangle2_y(rectangle2_ys[1298]), .rectangle2_width(rectangle2_widths[1298]), .rectangle2_height(rectangle2_heights[1298]), .rectangle2_weight(rectangle2_weights[1298]), .rectangle3_x(rectangle3_xs[1298]), .rectangle3_y(rectangle3_ys[1298]), .rectangle3_width(rectangle3_widths[1298]), .rectangle3_height(rectangle3_heights[1298]), .rectangle3_weight(rectangle3_weights[1298]), .feature_threshold(feature_thresholds[1298]), .feature_above(feature_aboves[1298]), .feature_below(feature_belows[1298]), .scan_win_std_dev(scan_win_std_dev[1298]), .feature_accum(feature_accums[1298]));
  accum_calculator ac1299(.scan_win(scan_win1299), .rectangle1_x(rectangle1_xs[1299]), .rectangle1_y(rectangle1_ys[1299]), .rectangle1_width(rectangle1_widths[1299]), .rectangle1_height(rectangle1_heights[1299]), .rectangle1_weight(rectangle1_weights[1299]), .rectangle2_x(rectangle2_xs[1299]), .rectangle2_y(rectangle2_ys[1299]), .rectangle2_width(rectangle2_widths[1299]), .rectangle2_height(rectangle2_heights[1299]), .rectangle2_weight(rectangle2_weights[1299]), .rectangle3_x(rectangle3_xs[1299]), .rectangle3_y(rectangle3_ys[1299]), .rectangle3_width(rectangle3_widths[1299]), .rectangle3_height(rectangle3_heights[1299]), .rectangle3_weight(rectangle3_weights[1299]), .feature_threshold(feature_thresholds[1299]), .feature_above(feature_aboves[1299]), .feature_below(feature_belows[1299]), .scan_win_std_dev(scan_win_std_dev[1299]), .feature_accum(feature_accums[1299]));
  accum_calculator ac1300(.scan_win(scan_win1300), .rectangle1_x(rectangle1_xs[1300]), .rectangle1_y(rectangle1_ys[1300]), .rectangle1_width(rectangle1_widths[1300]), .rectangle1_height(rectangle1_heights[1300]), .rectangle1_weight(rectangle1_weights[1300]), .rectangle2_x(rectangle2_xs[1300]), .rectangle2_y(rectangle2_ys[1300]), .rectangle2_width(rectangle2_widths[1300]), .rectangle2_height(rectangle2_heights[1300]), .rectangle2_weight(rectangle2_weights[1300]), .rectangle3_x(rectangle3_xs[1300]), .rectangle3_y(rectangle3_ys[1300]), .rectangle3_width(rectangle3_widths[1300]), .rectangle3_height(rectangle3_heights[1300]), .rectangle3_weight(rectangle3_weights[1300]), .feature_threshold(feature_thresholds[1300]), .feature_above(feature_aboves[1300]), .feature_below(feature_belows[1300]), .scan_win_std_dev(scan_win_std_dev[1300]), .feature_accum(feature_accums[1300]));
  accum_calculator ac1301(.scan_win(scan_win1301), .rectangle1_x(rectangle1_xs[1301]), .rectangle1_y(rectangle1_ys[1301]), .rectangle1_width(rectangle1_widths[1301]), .rectangle1_height(rectangle1_heights[1301]), .rectangle1_weight(rectangle1_weights[1301]), .rectangle2_x(rectangle2_xs[1301]), .rectangle2_y(rectangle2_ys[1301]), .rectangle2_width(rectangle2_widths[1301]), .rectangle2_height(rectangle2_heights[1301]), .rectangle2_weight(rectangle2_weights[1301]), .rectangle3_x(rectangle3_xs[1301]), .rectangle3_y(rectangle3_ys[1301]), .rectangle3_width(rectangle3_widths[1301]), .rectangle3_height(rectangle3_heights[1301]), .rectangle3_weight(rectangle3_weights[1301]), .feature_threshold(feature_thresholds[1301]), .feature_above(feature_aboves[1301]), .feature_below(feature_belows[1301]), .scan_win_std_dev(scan_win_std_dev[1301]), .feature_accum(feature_accums[1301]));
  accum_calculator ac1302(.scan_win(scan_win1302), .rectangle1_x(rectangle1_xs[1302]), .rectangle1_y(rectangle1_ys[1302]), .rectangle1_width(rectangle1_widths[1302]), .rectangle1_height(rectangle1_heights[1302]), .rectangle1_weight(rectangle1_weights[1302]), .rectangle2_x(rectangle2_xs[1302]), .rectangle2_y(rectangle2_ys[1302]), .rectangle2_width(rectangle2_widths[1302]), .rectangle2_height(rectangle2_heights[1302]), .rectangle2_weight(rectangle2_weights[1302]), .rectangle3_x(rectangle3_xs[1302]), .rectangle3_y(rectangle3_ys[1302]), .rectangle3_width(rectangle3_widths[1302]), .rectangle3_height(rectangle3_heights[1302]), .rectangle3_weight(rectangle3_weights[1302]), .feature_threshold(feature_thresholds[1302]), .feature_above(feature_aboves[1302]), .feature_below(feature_belows[1302]), .scan_win_std_dev(scan_win_std_dev[1302]), .feature_accum(feature_accums[1302]));
  accum_calculator ac1303(.scan_win(scan_win1303), .rectangle1_x(rectangle1_xs[1303]), .rectangle1_y(rectangle1_ys[1303]), .rectangle1_width(rectangle1_widths[1303]), .rectangle1_height(rectangle1_heights[1303]), .rectangle1_weight(rectangle1_weights[1303]), .rectangle2_x(rectangle2_xs[1303]), .rectangle2_y(rectangle2_ys[1303]), .rectangle2_width(rectangle2_widths[1303]), .rectangle2_height(rectangle2_heights[1303]), .rectangle2_weight(rectangle2_weights[1303]), .rectangle3_x(rectangle3_xs[1303]), .rectangle3_y(rectangle3_ys[1303]), .rectangle3_width(rectangle3_widths[1303]), .rectangle3_height(rectangle3_heights[1303]), .rectangle3_weight(rectangle3_weights[1303]), .feature_threshold(feature_thresholds[1303]), .feature_above(feature_aboves[1303]), .feature_below(feature_belows[1303]), .scan_win_std_dev(scan_win_std_dev[1303]), .feature_accum(feature_accums[1303]));
  accum_calculator ac1304(.scan_win(scan_win1304), .rectangle1_x(rectangle1_xs[1304]), .rectangle1_y(rectangle1_ys[1304]), .rectangle1_width(rectangle1_widths[1304]), .rectangle1_height(rectangle1_heights[1304]), .rectangle1_weight(rectangle1_weights[1304]), .rectangle2_x(rectangle2_xs[1304]), .rectangle2_y(rectangle2_ys[1304]), .rectangle2_width(rectangle2_widths[1304]), .rectangle2_height(rectangle2_heights[1304]), .rectangle2_weight(rectangle2_weights[1304]), .rectangle3_x(rectangle3_xs[1304]), .rectangle3_y(rectangle3_ys[1304]), .rectangle3_width(rectangle3_widths[1304]), .rectangle3_height(rectangle3_heights[1304]), .rectangle3_weight(rectangle3_weights[1304]), .feature_threshold(feature_thresholds[1304]), .feature_above(feature_aboves[1304]), .feature_below(feature_belows[1304]), .scan_win_std_dev(scan_win_std_dev[1304]), .feature_accum(feature_accums[1304]));
  accum_calculator ac1305(.scan_win(scan_win1305), .rectangle1_x(rectangle1_xs[1305]), .rectangle1_y(rectangle1_ys[1305]), .rectangle1_width(rectangle1_widths[1305]), .rectangle1_height(rectangle1_heights[1305]), .rectangle1_weight(rectangle1_weights[1305]), .rectangle2_x(rectangle2_xs[1305]), .rectangle2_y(rectangle2_ys[1305]), .rectangle2_width(rectangle2_widths[1305]), .rectangle2_height(rectangle2_heights[1305]), .rectangle2_weight(rectangle2_weights[1305]), .rectangle3_x(rectangle3_xs[1305]), .rectangle3_y(rectangle3_ys[1305]), .rectangle3_width(rectangle3_widths[1305]), .rectangle3_height(rectangle3_heights[1305]), .rectangle3_weight(rectangle3_weights[1305]), .feature_threshold(feature_thresholds[1305]), .feature_above(feature_aboves[1305]), .feature_below(feature_belows[1305]), .scan_win_std_dev(scan_win_std_dev[1305]), .feature_accum(feature_accums[1305]));
  accum_calculator ac1306(.scan_win(scan_win1306), .rectangle1_x(rectangle1_xs[1306]), .rectangle1_y(rectangle1_ys[1306]), .rectangle1_width(rectangle1_widths[1306]), .rectangle1_height(rectangle1_heights[1306]), .rectangle1_weight(rectangle1_weights[1306]), .rectangle2_x(rectangle2_xs[1306]), .rectangle2_y(rectangle2_ys[1306]), .rectangle2_width(rectangle2_widths[1306]), .rectangle2_height(rectangle2_heights[1306]), .rectangle2_weight(rectangle2_weights[1306]), .rectangle3_x(rectangle3_xs[1306]), .rectangle3_y(rectangle3_ys[1306]), .rectangle3_width(rectangle3_widths[1306]), .rectangle3_height(rectangle3_heights[1306]), .rectangle3_weight(rectangle3_weights[1306]), .feature_threshold(feature_thresholds[1306]), .feature_above(feature_aboves[1306]), .feature_below(feature_belows[1306]), .scan_win_std_dev(scan_win_std_dev[1306]), .feature_accum(feature_accums[1306]));
  accum_calculator ac1307(.scan_win(scan_win1307), .rectangle1_x(rectangle1_xs[1307]), .rectangle1_y(rectangle1_ys[1307]), .rectangle1_width(rectangle1_widths[1307]), .rectangle1_height(rectangle1_heights[1307]), .rectangle1_weight(rectangle1_weights[1307]), .rectangle2_x(rectangle2_xs[1307]), .rectangle2_y(rectangle2_ys[1307]), .rectangle2_width(rectangle2_widths[1307]), .rectangle2_height(rectangle2_heights[1307]), .rectangle2_weight(rectangle2_weights[1307]), .rectangle3_x(rectangle3_xs[1307]), .rectangle3_y(rectangle3_ys[1307]), .rectangle3_width(rectangle3_widths[1307]), .rectangle3_height(rectangle3_heights[1307]), .rectangle3_weight(rectangle3_weights[1307]), .feature_threshold(feature_thresholds[1307]), .feature_above(feature_aboves[1307]), .feature_below(feature_belows[1307]), .scan_win_std_dev(scan_win_std_dev[1307]), .feature_accum(feature_accums[1307]));
  accum_calculator ac1308(.scan_win(scan_win1308), .rectangle1_x(rectangle1_xs[1308]), .rectangle1_y(rectangle1_ys[1308]), .rectangle1_width(rectangle1_widths[1308]), .rectangle1_height(rectangle1_heights[1308]), .rectangle1_weight(rectangle1_weights[1308]), .rectangle2_x(rectangle2_xs[1308]), .rectangle2_y(rectangle2_ys[1308]), .rectangle2_width(rectangle2_widths[1308]), .rectangle2_height(rectangle2_heights[1308]), .rectangle2_weight(rectangle2_weights[1308]), .rectangle3_x(rectangle3_xs[1308]), .rectangle3_y(rectangle3_ys[1308]), .rectangle3_width(rectangle3_widths[1308]), .rectangle3_height(rectangle3_heights[1308]), .rectangle3_weight(rectangle3_weights[1308]), .feature_threshold(feature_thresholds[1308]), .feature_above(feature_aboves[1308]), .feature_below(feature_belows[1308]), .scan_win_std_dev(scan_win_std_dev[1308]), .feature_accum(feature_accums[1308]));
  accum_calculator ac1309(.scan_win(scan_win1309), .rectangle1_x(rectangle1_xs[1309]), .rectangle1_y(rectangle1_ys[1309]), .rectangle1_width(rectangle1_widths[1309]), .rectangle1_height(rectangle1_heights[1309]), .rectangle1_weight(rectangle1_weights[1309]), .rectangle2_x(rectangle2_xs[1309]), .rectangle2_y(rectangle2_ys[1309]), .rectangle2_width(rectangle2_widths[1309]), .rectangle2_height(rectangle2_heights[1309]), .rectangle2_weight(rectangle2_weights[1309]), .rectangle3_x(rectangle3_xs[1309]), .rectangle3_y(rectangle3_ys[1309]), .rectangle3_width(rectangle3_widths[1309]), .rectangle3_height(rectangle3_heights[1309]), .rectangle3_weight(rectangle3_weights[1309]), .feature_threshold(feature_thresholds[1309]), .feature_above(feature_aboves[1309]), .feature_below(feature_belows[1309]), .scan_win_std_dev(scan_win_std_dev[1309]), .feature_accum(feature_accums[1309]));
  accum_calculator ac1310(.scan_win(scan_win1310), .rectangle1_x(rectangle1_xs[1310]), .rectangle1_y(rectangle1_ys[1310]), .rectangle1_width(rectangle1_widths[1310]), .rectangle1_height(rectangle1_heights[1310]), .rectangle1_weight(rectangle1_weights[1310]), .rectangle2_x(rectangle2_xs[1310]), .rectangle2_y(rectangle2_ys[1310]), .rectangle2_width(rectangle2_widths[1310]), .rectangle2_height(rectangle2_heights[1310]), .rectangle2_weight(rectangle2_weights[1310]), .rectangle3_x(rectangle3_xs[1310]), .rectangle3_y(rectangle3_ys[1310]), .rectangle3_width(rectangle3_widths[1310]), .rectangle3_height(rectangle3_heights[1310]), .rectangle3_weight(rectangle3_weights[1310]), .feature_threshold(feature_thresholds[1310]), .feature_above(feature_aboves[1310]), .feature_below(feature_belows[1310]), .scan_win_std_dev(scan_win_std_dev[1310]), .feature_accum(feature_accums[1310]));
  accum_calculator ac1311(.scan_win(scan_win1311), .rectangle1_x(rectangle1_xs[1311]), .rectangle1_y(rectangle1_ys[1311]), .rectangle1_width(rectangle1_widths[1311]), .rectangle1_height(rectangle1_heights[1311]), .rectangle1_weight(rectangle1_weights[1311]), .rectangle2_x(rectangle2_xs[1311]), .rectangle2_y(rectangle2_ys[1311]), .rectangle2_width(rectangle2_widths[1311]), .rectangle2_height(rectangle2_heights[1311]), .rectangle2_weight(rectangle2_weights[1311]), .rectangle3_x(rectangle3_xs[1311]), .rectangle3_y(rectangle3_ys[1311]), .rectangle3_width(rectangle3_widths[1311]), .rectangle3_height(rectangle3_heights[1311]), .rectangle3_weight(rectangle3_weights[1311]), .feature_threshold(feature_thresholds[1311]), .feature_above(feature_aboves[1311]), .feature_below(feature_belows[1311]), .scan_win_std_dev(scan_win_std_dev[1311]), .feature_accum(feature_accums[1311]));
  accum_calculator ac1312(.scan_win(scan_win1312), .rectangle1_x(rectangle1_xs[1312]), .rectangle1_y(rectangle1_ys[1312]), .rectangle1_width(rectangle1_widths[1312]), .rectangle1_height(rectangle1_heights[1312]), .rectangle1_weight(rectangle1_weights[1312]), .rectangle2_x(rectangle2_xs[1312]), .rectangle2_y(rectangle2_ys[1312]), .rectangle2_width(rectangle2_widths[1312]), .rectangle2_height(rectangle2_heights[1312]), .rectangle2_weight(rectangle2_weights[1312]), .rectangle3_x(rectangle3_xs[1312]), .rectangle3_y(rectangle3_ys[1312]), .rectangle3_width(rectangle3_widths[1312]), .rectangle3_height(rectangle3_heights[1312]), .rectangle3_weight(rectangle3_weights[1312]), .feature_threshold(feature_thresholds[1312]), .feature_above(feature_aboves[1312]), .feature_below(feature_belows[1312]), .scan_win_std_dev(scan_win_std_dev[1312]), .feature_accum(feature_accums[1312]));
  accum_calculator ac1313(.scan_win(scan_win1313), .rectangle1_x(rectangle1_xs[1313]), .rectangle1_y(rectangle1_ys[1313]), .rectangle1_width(rectangle1_widths[1313]), .rectangle1_height(rectangle1_heights[1313]), .rectangle1_weight(rectangle1_weights[1313]), .rectangle2_x(rectangle2_xs[1313]), .rectangle2_y(rectangle2_ys[1313]), .rectangle2_width(rectangle2_widths[1313]), .rectangle2_height(rectangle2_heights[1313]), .rectangle2_weight(rectangle2_weights[1313]), .rectangle3_x(rectangle3_xs[1313]), .rectangle3_y(rectangle3_ys[1313]), .rectangle3_width(rectangle3_widths[1313]), .rectangle3_height(rectangle3_heights[1313]), .rectangle3_weight(rectangle3_weights[1313]), .feature_threshold(feature_thresholds[1313]), .feature_above(feature_aboves[1313]), .feature_below(feature_belows[1313]), .scan_win_std_dev(scan_win_std_dev[1313]), .feature_accum(feature_accums[1313]));
  accum_calculator ac1314(.scan_win(scan_win1314), .rectangle1_x(rectangle1_xs[1314]), .rectangle1_y(rectangle1_ys[1314]), .rectangle1_width(rectangle1_widths[1314]), .rectangle1_height(rectangle1_heights[1314]), .rectangle1_weight(rectangle1_weights[1314]), .rectangle2_x(rectangle2_xs[1314]), .rectangle2_y(rectangle2_ys[1314]), .rectangle2_width(rectangle2_widths[1314]), .rectangle2_height(rectangle2_heights[1314]), .rectangle2_weight(rectangle2_weights[1314]), .rectangle3_x(rectangle3_xs[1314]), .rectangle3_y(rectangle3_ys[1314]), .rectangle3_width(rectangle3_widths[1314]), .rectangle3_height(rectangle3_heights[1314]), .rectangle3_weight(rectangle3_weights[1314]), .feature_threshold(feature_thresholds[1314]), .feature_above(feature_aboves[1314]), .feature_below(feature_belows[1314]), .scan_win_std_dev(scan_win_std_dev[1314]), .feature_accum(feature_accums[1314]));
  accum_calculator ac1315(.scan_win(scan_win1315), .rectangle1_x(rectangle1_xs[1315]), .rectangle1_y(rectangle1_ys[1315]), .rectangle1_width(rectangle1_widths[1315]), .rectangle1_height(rectangle1_heights[1315]), .rectangle1_weight(rectangle1_weights[1315]), .rectangle2_x(rectangle2_xs[1315]), .rectangle2_y(rectangle2_ys[1315]), .rectangle2_width(rectangle2_widths[1315]), .rectangle2_height(rectangle2_heights[1315]), .rectangle2_weight(rectangle2_weights[1315]), .rectangle3_x(rectangle3_xs[1315]), .rectangle3_y(rectangle3_ys[1315]), .rectangle3_width(rectangle3_widths[1315]), .rectangle3_height(rectangle3_heights[1315]), .rectangle3_weight(rectangle3_weights[1315]), .feature_threshold(feature_thresholds[1315]), .feature_above(feature_aboves[1315]), .feature_below(feature_belows[1315]), .scan_win_std_dev(scan_win_std_dev[1315]), .feature_accum(feature_accums[1315]));
  accum_calculator ac1316(.scan_win(scan_win1316), .rectangle1_x(rectangle1_xs[1316]), .rectangle1_y(rectangle1_ys[1316]), .rectangle1_width(rectangle1_widths[1316]), .rectangle1_height(rectangle1_heights[1316]), .rectangle1_weight(rectangle1_weights[1316]), .rectangle2_x(rectangle2_xs[1316]), .rectangle2_y(rectangle2_ys[1316]), .rectangle2_width(rectangle2_widths[1316]), .rectangle2_height(rectangle2_heights[1316]), .rectangle2_weight(rectangle2_weights[1316]), .rectangle3_x(rectangle3_xs[1316]), .rectangle3_y(rectangle3_ys[1316]), .rectangle3_width(rectangle3_widths[1316]), .rectangle3_height(rectangle3_heights[1316]), .rectangle3_weight(rectangle3_weights[1316]), .feature_threshold(feature_thresholds[1316]), .feature_above(feature_aboves[1316]), .feature_below(feature_belows[1316]), .scan_win_std_dev(scan_win_std_dev[1316]), .feature_accum(feature_accums[1316]));
  accum_calculator ac1317(.scan_win(scan_win1317), .rectangle1_x(rectangle1_xs[1317]), .rectangle1_y(rectangle1_ys[1317]), .rectangle1_width(rectangle1_widths[1317]), .rectangle1_height(rectangle1_heights[1317]), .rectangle1_weight(rectangle1_weights[1317]), .rectangle2_x(rectangle2_xs[1317]), .rectangle2_y(rectangle2_ys[1317]), .rectangle2_width(rectangle2_widths[1317]), .rectangle2_height(rectangle2_heights[1317]), .rectangle2_weight(rectangle2_weights[1317]), .rectangle3_x(rectangle3_xs[1317]), .rectangle3_y(rectangle3_ys[1317]), .rectangle3_width(rectangle3_widths[1317]), .rectangle3_height(rectangle3_heights[1317]), .rectangle3_weight(rectangle3_weights[1317]), .feature_threshold(feature_thresholds[1317]), .feature_above(feature_aboves[1317]), .feature_below(feature_belows[1317]), .scan_win_std_dev(scan_win_std_dev[1317]), .feature_accum(feature_accums[1317]));
  accum_calculator ac1318(.scan_win(scan_win1318), .rectangle1_x(rectangle1_xs[1318]), .rectangle1_y(rectangle1_ys[1318]), .rectangle1_width(rectangle1_widths[1318]), .rectangle1_height(rectangle1_heights[1318]), .rectangle1_weight(rectangle1_weights[1318]), .rectangle2_x(rectangle2_xs[1318]), .rectangle2_y(rectangle2_ys[1318]), .rectangle2_width(rectangle2_widths[1318]), .rectangle2_height(rectangle2_heights[1318]), .rectangle2_weight(rectangle2_weights[1318]), .rectangle3_x(rectangle3_xs[1318]), .rectangle3_y(rectangle3_ys[1318]), .rectangle3_width(rectangle3_widths[1318]), .rectangle3_height(rectangle3_heights[1318]), .rectangle3_weight(rectangle3_weights[1318]), .feature_threshold(feature_thresholds[1318]), .feature_above(feature_aboves[1318]), .feature_below(feature_belows[1318]), .scan_win_std_dev(scan_win_std_dev[1318]), .feature_accum(feature_accums[1318]));
  accum_calculator ac1319(.scan_win(scan_win1319), .rectangle1_x(rectangle1_xs[1319]), .rectangle1_y(rectangle1_ys[1319]), .rectangle1_width(rectangle1_widths[1319]), .rectangle1_height(rectangle1_heights[1319]), .rectangle1_weight(rectangle1_weights[1319]), .rectangle2_x(rectangle2_xs[1319]), .rectangle2_y(rectangle2_ys[1319]), .rectangle2_width(rectangle2_widths[1319]), .rectangle2_height(rectangle2_heights[1319]), .rectangle2_weight(rectangle2_weights[1319]), .rectangle3_x(rectangle3_xs[1319]), .rectangle3_y(rectangle3_ys[1319]), .rectangle3_width(rectangle3_widths[1319]), .rectangle3_height(rectangle3_heights[1319]), .rectangle3_weight(rectangle3_weights[1319]), .feature_threshold(feature_thresholds[1319]), .feature_above(feature_aboves[1319]), .feature_below(feature_belows[1319]), .scan_win_std_dev(scan_win_std_dev[1319]), .feature_accum(feature_accums[1319]));
  accum_calculator ac1320(.scan_win(scan_win1320), .rectangle1_x(rectangle1_xs[1320]), .rectangle1_y(rectangle1_ys[1320]), .rectangle1_width(rectangle1_widths[1320]), .rectangle1_height(rectangle1_heights[1320]), .rectangle1_weight(rectangle1_weights[1320]), .rectangle2_x(rectangle2_xs[1320]), .rectangle2_y(rectangle2_ys[1320]), .rectangle2_width(rectangle2_widths[1320]), .rectangle2_height(rectangle2_heights[1320]), .rectangle2_weight(rectangle2_weights[1320]), .rectangle3_x(rectangle3_xs[1320]), .rectangle3_y(rectangle3_ys[1320]), .rectangle3_width(rectangle3_widths[1320]), .rectangle3_height(rectangle3_heights[1320]), .rectangle3_weight(rectangle3_weights[1320]), .feature_threshold(feature_thresholds[1320]), .feature_above(feature_aboves[1320]), .feature_below(feature_belows[1320]), .scan_win_std_dev(scan_win_std_dev[1320]), .feature_accum(feature_accums[1320]));
  accum_calculator ac1321(.scan_win(scan_win1321), .rectangle1_x(rectangle1_xs[1321]), .rectangle1_y(rectangle1_ys[1321]), .rectangle1_width(rectangle1_widths[1321]), .rectangle1_height(rectangle1_heights[1321]), .rectangle1_weight(rectangle1_weights[1321]), .rectangle2_x(rectangle2_xs[1321]), .rectangle2_y(rectangle2_ys[1321]), .rectangle2_width(rectangle2_widths[1321]), .rectangle2_height(rectangle2_heights[1321]), .rectangle2_weight(rectangle2_weights[1321]), .rectangle3_x(rectangle3_xs[1321]), .rectangle3_y(rectangle3_ys[1321]), .rectangle3_width(rectangle3_widths[1321]), .rectangle3_height(rectangle3_heights[1321]), .rectangle3_weight(rectangle3_weights[1321]), .feature_threshold(feature_thresholds[1321]), .feature_above(feature_aboves[1321]), .feature_below(feature_belows[1321]), .scan_win_std_dev(scan_win_std_dev[1321]), .feature_accum(feature_accums[1321]));
  accum_calculator ac1322(.scan_win(scan_win1322), .rectangle1_x(rectangle1_xs[1322]), .rectangle1_y(rectangle1_ys[1322]), .rectangle1_width(rectangle1_widths[1322]), .rectangle1_height(rectangle1_heights[1322]), .rectangle1_weight(rectangle1_weights[1322]), .rectangle2_x(rectangle2_xs[1322]), .rectangle2_y(rectangle2_ys[1322]), .rectangle2_width(rectangle2_widths[1322]), .rectangle2_height(rectangle2_heights[1322]), .rectangle2_weight(rectangle2_weights[1322]), .rectangle3_x(rectangle3_xs[1322]), .rectangle3_y(rectangle3_ys[1322]), .rectangle3_width(rectangle3_widths[1322]), .rectangle3_height(rectangle3_heights[1322]), .rectangle3_weight(rectangle3_weights[1322]), .feature_threshold(feature_thresholds[1322]), .feature_above(feature_aboves[1322]), .feature_below(feature_belows[1322]), .scan_win_std_dev(scan_win_std_dev[1322]), .feature_accum(feature_accums[1322]));
  accum_calculator ac1323(.scan_win(scan_win1323), .rectangle1_x(rectangle1_xs[1323]), .rectangle1_y(rectangle1_ys[1323]), .rectangle1_width(rectangle1_widths[1323]), .rectangle1_height(rectangle1_heights[1323]), .rectangle1_weight(rectangle1_weights[1323]), .rectangle2_x(rectangle2_xs[1323]), .rectangle2_y(rectangle2_ys[1323]), .rectangle2_width(rectangle2_widths[1323]), .rectangle2_height(rectangle2_heights[1323]), .rectangle2_weight(rectangle2_weights[1323]), .rectangle3_x(rectangle3_xs[1323]), .rectangle3_y(rectangle3_ys[1323]), .rectangle3_width(rectangle3_widths[1323]), .rectangle3_height(rectangle3_heights[1323]), .rectangle3_weight(rectangle3_weights[1323]), .feature_threshold(feature_thresholds[1323]), .feature_above(feature_aboves[1323]), .feature_below(feature_belows[1323]), .scan_win_std_dev(scan_win_std_dev[1323]), .feature_accum(feature_accums[1323]));
  accum_calculator ac1324(.scan_win(scan_win1324), .rectangle1_x(rectangle1_xs[1324]), .rectangle1_y(rectangle1_ys[1324]), .rectangle1_width(rectangle1_widths[1324]), .rectangle1_height(rectangle1_heights[1324]), .rectangle1_weight(rectangle1_weights[1324]), .rectangle2_x(rectangle2_xs[1324]), .rectangle2_y(rectangle2_ys[1324]), .rectangle2_width(rectangle2_widths[1324]), .rectangle2_height(rectangle2_heights[1324]), .rectangle2_weight(rectangle2_weights[1324]), .rectangle3_x(rectangle3_xs[1324]), .rectangle3_y(rectangle3_ys[1324]), .rectangle3_width(rectangle3_widths[1324]), .rectangle3_height(rectangle3_heights[1324]), .rectangle3_weight(rectangle3_weights[1324]), .feature_threshold(feature_thresholds[1324]), .feature_above(feature_aboves[1324]), .feature_below(feature_belows[1324]), .scan_win_std_dev(scan_win_std_dev[1324]), .feature_accum(feature_accums[1324]));
  accum_calculator ac1325(.scan_win(scan_win1325), .rectangle1_x(rectangle1_xs[1325]), .rectangle1_y(rectangle1_ys[1325]), .rectangle1_width(rectangle1_widths[1325]), .rectangle1_height(rectangle1_heights[1325]), .rectangle1_weight(rectangle1_weights[1325]), .rectangle2_x(rectangle2_xs[1325]), .rectangle2_y(rectangle2_ys[1325]), .rectangle2_width(rectangle2_widths[1325]), .rectangle2_height(rectangle2_heights[1325]), .rectangle2_weight(rectangle2_weights[1325]), .rectangle3_x(rectangle3_xs[1325]), .rectangle3_y(rectangle3_ys[1325]), .rectangle3_width(rectangle3_widths[1325]), .rectangle3_height(rectangle3_heights[1325]), .rectangle3_weight(rectangle3_weights[1325]), .feature_threshold(feature_thresholds[1325]), .feature_above(feature_aboves[1325]), .feature_below(feature_belows[1325]), .scan_win_std_dev(scan_win_std_dev[1325]), .feature_accum(feature_accums[1325]));
  accum_calculator ac1326(.scan_win(scan_win1326), .rectangle1_x(rectangle1_xs[1326]), .rectangle1_y(rectangle1_ys[1326]), .rectangle1_width(rectangle1_widths[1326]), .rectangle1_height(rectangle1_heights[1326]), .rectangle1_weight(rectangle1_weights[1326]), .rectangle2_x(rectangle2_xs[1326]), .rectangle2_y(rectangle2_ys[1326]), .rectangle2_width(rectangle2_widths[1326]), .rectangle2_height(rectangle2_heights[1326]), .rectangle2_weight(rectangle2_weights[1326]), .rectangle3_x(rectangle3_xs[1326]), .rectangle3_y(rectangle3_ys[1326]), .rectangle3_width(rectangle3_widths[1326]), .rectangle3_height(rectangle3_heights[1326]), .rectangle3_weight(rectangle3_weights[1326]), .feature_threshold(feature_thresholds[1326]), .feature_above(feature_aboves[1326]), .feature_below(feature_belows[1326]), .scan_win_std_dev(scan_win_std_dev[1326]), .feature_accum(feature_accums[1326]));
  accum_calculator ac1327(.scan_win(scan_win1327), .rectangle1_x(rectangle1_xs[1327]), .rectangle1_y(rectangle1_ys[1327]), .rectangle1_width(rectangle1_widths[1327]), .rectangle1_height(rectangle1_heights[1327]), .rectangle1_weight(rectangle1_weights[1327]), .rectangle2_x(rectangle2_xs[1327]), .rectangle2_y(rectangle2_ys[1327]), .rectangle2_width(rectangle2_widths[1327]), .rectangle2_height(rectangle2_heights[1327]), .rectangle2_weight(rectangle2_weights[1327]), .rectangle3_x(rectangle3_xs[1327]), .rectangle3_y(rectangle3_ys[1327]), .rectangle3_width(rectangle3_widths[1327]), .rectangle3_height(rectangle3_heights[1327]), .rectangle3_weight(rectangle3_weights[1327]), .feature_threshold(feature_thresholds[1327]), .feature_above(feature_aboves[1327]), .feature_below(feature_belows[1327]), .scan_win_std_dev(scan_win_std_dev[1327]), .feature_accum(feature_accums[1327]));
  accum_calculator ac1328(.scan_win(scan_win1328), .rectangle1_x(rectangle1_xs[1328]), .rectangle1_y(rectangle1_ys[1328]), .rectangle1_width(rectangle1_widths[1328]), .rectangle1_height(rectangle1_heights[1328]), .rectangle1_weight(rectangle1_weights[1328]), .rectangle2_x(rectangle2_xs[1328]), .rectangle2_y(rectangle2_ys[1328]), .rectangle2_width(rectangle2_widths[1328]), .rectangle2_height(rectangle2_heights[1328]), .rectangle2_weight(rectangle2_weights[1328]), .rectangle3_x(rectangle3_xs[1328]), .rectangle3_y(rectangle3_ys[1328]), .rectangle3_width(rectangle3_widths[1328]), .rectangle3_height(rectangle3_heights[1328]), .rectangle3_weight(rectangle3_weights[1328]), .feature_threshold(feature_thresholds[1328]), .feature_above(feature_aboves[1328]), .feature_below(feature_belows[1328]), .scan_win_std_dev(scan_win_std_dev[1328]), .feature_accum(feature_accums[1328]));
  accum_calculator ac1329(.scan_win(scan_win1329), .rectangle1_x(rectangle1_xs[1329]), .rectangle1_y(rectangle1_ys[1329]), .rectangle1_width(rectangle1_widths[1329]), .rectangle1_height(rectangle1_heights[1329]), .rectangle1_weight(rectangle1_weights[1329]), .rectangle2_x(rectangle2_xs[1329]), .rectangle2_y(rectangle2_ys[1329]), .rectangle2_width(rectangle2_widths[1329]), .rectangle2_height(rectangle2_heights[1329]), .rectangle2_weight(rectangle2_weights[1329]), .rectangle3_x(rectangle3_xs[1329]), .rectangle3_y(rectangle3_ys[1329]), .rectangle3_width(rectangle3_widths[1329]), .rectangle3_height(rectangle3_heights[1329]), .rectangle3_weight(rectangle3_weights[1329]), .feature_threshold(feature_thresholds[1329]), .feature_above(feature_aboves[1329]), .feature_below(feature_belows[1329]), .scan_win_std_dev(scan_win_std_dev[1329]), .feature_accum(feature_accums[1329]));
  accum_calculator ac1330(.scan_win(scan_win1330), .rectangle1_x(rectangle1_xs[1330]), .rectangle1_y(rectangle1_ys[1330]), .rectangle1_width(rectangle1_widths[1330]), .rectangle1_height(rectangle1_heights[1330]), .rectangle1_weight(rectangle1_weights[1330]), .rectangle2_x(rectangle2_xs[1330]), .rectangle2_y(rectangle2_ys[1330]), .rectangle2_width(rectangle2_widths[1330]), .rectangle2_height(rectangle2_heights[1330]), .rectangle2_weight(rectangle2_weights[1330]), .rectangle3_x(rectangle3_xs[1330]), .rectangle3_y(rectangle3_ys[1330]), .rectangle3_width(rectangle3_widths[1330]), .rectangle3_height(rectangle3_heights[1330]), .rectangle3_weight(rectangle3_weights[1330]), .feature_threshold(feature_thresholds[1330]), .feature_above(feature_aboves[1330]), .feature_below(feature_belows[1330]), .scan_win_std_dev(scan_win_std_dev[1330]), .feature_accum(feature_accums[1330]));
  accum_calculator ac1331(.scan_win(scan_win1331), .rectangle1_x(rectangle1_xs[1331]), .rectangle1_y(rectangle1_ys[1331]), .rectangle1_width(rectangle1_widths[1331]), .rectangle1_height(rectangle1_heights[1331]), .rectangle1_weight(rectangle1_weights[1331]), .rectangle2_x(rectangle2_xs[1331]), .rectangle2_y(rectangle2_ys[1331]), .rectangle2_width(rectangle2_widths[1331]), .rectangle2_height(rectangle2_heights[1331]), .rectangle2_weight(rectangle2_weights[1331]), .rectangle3_x(rectangle3_xs[1331]), .rectangle3_y(rectangle3_ys[1331]), .rectangle3_width(rectangle3_widths[1331]), .rectangle3_height(rectangle3_heights[1331]), .rectangle3_weight(rectangle3_weights[1331]), .feature_threshold(feature_thresholds[1331]), .feature_above(feature_aboves[1331]), .feature_below(feature_belows[1331]), .scan_win_std_dev(scan_win_std_dev[1331]), .feature_accum(feature_accums[1331]));
  accum_calculator ac1332(.scan_win(scan_win1332), .rectangle1_x(rectangle1_xs[1332]), .rectangle1_y(rectangle1_ys[1332]), .rectangle1_width(rectangle1_widths[1332]), .rectangle1_height(rectangle1_heights[1332]), .rectangle1_weight(rectangle1_weights[1332]), .rectangle2_x(rectangle2_xs[1332]), .rectangle2_y(rectangle2_ys[1332]), .rectangle2_width(rectangle2_widths[1332]), .rectangle2_height(rectangle2_heights[1332]), .rectangle2_weight(rectangle2_weights[1332]), .rectangle3_x(rectangle3_xs[1332]), .rectangle3_y(rectangle3_ys[1332]), .rectangle3_width(rectangle3_widths[1332]), .rectangle3_height(rectangle3_heights[1332]), .rectangle3_weight(rectangle3_weights[1332]), .feature_threshold(feature_thresholds[1332]), .feature_above(feature_aboves[1332]), .feature_below(feature_belows[1332]), .scan_win_std_dev(scan_win_std_dev[1332]), .feature_accum(feature_accums[1332]));
  accum_calculator ac1333(.scan_win(scan_win1333), .rectangle1_x(rectangle1_xs[1333]), .rectangle1_y(rectangle1_ys[1333]), .rectangle1_width(rectangle1_widths[1333]), .rectangle1_height(rectangle1_heights[1333]), .rectangle1_weight(rectangle1_weights[1333]), .rectangle2_x(rectangle2_xs[1333]), .rectangle2_y(rectangle2_ys[1333]), .rectangle2_width(rectangle2_widths[1333]), .rectangle2_height(rectangle2_heights[1333]), .rectangle2_weight(rectangle2_weights[1333]), .rectangle3_x(rectangle3_xs[1333]), .rectangle3_y(rectangle3_ys[1333]), .rectangle3_width(rectangle3_widths[1333]), .rectangle3_height(rectangle3_heights[1333]), .rectangle3_weight(rectangle3_weights[1333]), .feature_threshold(feature_thresholds[1333]), .feature_above(feature_aboves[1333]), .feature_below(feature_belows[1333]), .scan_win_std_dev(scan_win_std_dev[1333]), .feature_accum(feature_accums[1333]));
  accum_calculator ac1334(.scan_win(scan_win1334), .rectangle1_x(rectangle1_xs[1334]), .rectangle1_y(rectangle1_ys[1334]), .rectangle1_width(rectangle1_widths[1334]), .rectangle1_height(rectangle1_heights[1334]), .rectangle1_weight(rectangle1_weights[1334]), .rectangle2_x(rectangle2_xs[1334]), .rectangle2_y(rectangle2_ys[1334]), .rectangle2_width(rectangle2_widths[1334]), .rectangle2_height(rectangle2_heights[1334]), .rectangle2_weight(rectangle2_weights[1334]), .rectangle3_x(rectangle3_xs[1334]), .rectangle3_y(rectangle3_ys[1334]), .rectangle3_width(rectangle3_widths[1334]), .rectangle3_height(rectangle3_heights[1334]), .rectangle3_weight(rectangle3_weights[1334]), .feature_threshold(feature_thresholds[1334]), .feature_above(feature_aboves[1334]), .feature_below(feature_belows[1334]), .scan_win_std_dev(scan_win_std_dev[1334]), .feature_accum(feature_accums[1334]));
  accum_calculator ac1335(.scan_win(scan_win1335), .rectangle1_x(rectangle1_xs[1335]), .rectangle1_y(rectangle1_ys[1335]), .rectangle1_width(rectangle1_widths[1335]), .rectangle1_height(rectangle1_heights[1335]), .rectangle1_weight(rectangle1_weights[1335]), .rectangle2_x(rectangle2_xs[1335]), .rectangle2_y(rectangle2_ys[1335]), .rectangle2_width(rectangle2_widths[1335]), .rectangle2_height(rectangle2_heights[1335]), .rectangle2_weight(rectangle2_weights[1335]), .rectangle3_x(rectangle3_xs[1335]), .rectangle3_y(rectangle3_ys[1335]), .rectangle3_width(rectangle3_widths[1335]), .rectangle3_height(rectangle3_heights[1335]), .rectangle3_weight(rectangle3_weights[1335]), .feature_threshold(feature_thresholds[1335]), .feature_above(feature_aboves[1335]), .feature_below(feature_belows[1335]), .scan_win_std_dev(scan_win_std_dev[1335]), .feature_accum(feature_accums[1335]));
  accum_calculator ac1336(.scan_win(scan_win1336), .rectangle1_x(rectangle1_xs[1336]), .rectangle1_y(rectangle1_ys[1336]), .rectangle1_width(rectangle1_widths[1336]), .rectangle1_height(rectangle1_heights[1336]), .rectangle1_weight(rectangle1_weights[1336]), .rectangle2_x(rectangle2_xs[1336]), .rectangle2_y(rectangle2_ys[1336]), .rectangle2_width(rectangle2_widths[1336]), .rectangle2_height(rectangle2_heights[1336]), .rectangle2_weight(rectangle2_weights[1336]), .rectangle3_x(rectangle3_xs[1336]), .rectangle3_y(rectangle3_ys[1336]), .rectangle3_width(rectangle3_widths[1336]), .rectangle3_height(rectangle3_heights[1336]), .rectangle3_weight(rectangle3_weights[1336]), .feature_threshold(feature_thresholds[1336]), .feature_above(feature_aboves[1336]), .feature_below(feature_belows[1336]), .scan_win_std_dev(scan_win_std_dev[1336]), .feature_accum(feature_accums[1336]));
  accum_calculator ac1337(.scan_win(scan_win1337), .rectangle1_x(rectangle1_xs[1337]), .rectangle1_y(rectangle1_ys[1337]), .rectangle1_width(rectangle1_widths[1337]), .rectangle1_height(rectangle1_heights[1337]), .rectangle1_weight(rectangle1_weights[1337]), .rectangle2_x(rectangle2_xs[1337]), .rectangle2_y(rectangle2_ys[1337]), .rectangle2_width(rectangle2_widths[1337]), .rectangle2_height(rectangle2_heights[1337]), .rectangle2_weight(rectangle2_weights[1337]), .rectangle3_x(rectangle3_xs[1337]), .rectangle3_y(rectangle3_ys[1337]), .rectangle3_width(rectangle3_widths[1337]), .rectangle3_height(rectangle3_heights[1337]), .rectangle3_weight(rectangle3_weights[1337]), .feature_threshold(feature_thresholds[1337]), .feature_above(feature_aboves[1337]), .feature_below(feature_belows[1337]), .scan_win_std_dev(scan_win_std_dev[1337]), .feature_accum(feature_accums[1337]));
  accum_calculator ac1338(.scan_win(scan_win1338), .rectangle1_x(rectangle1_xs[1338]), .rectangle1_y(rectangle1_ys[1338]), .rectangle1_width(rectangle1_widths[1338]), .rectangle1_height(rectangle1_heights[1338]), .rectangle1_weight(rectangle1_weights[1338]), .rectangle2_x(rectangle2_xs[1338]), .rectangle2_y(rectangle2_ys[1338]), .rectangle2_width(rectangle2_widths[1338]), .rectangle2_height(rectangle2_heights[1338]), .rectangle2_weight(rectangle2_weights[1338]), .rectangle3_x(rectangle3_xs[1338]), .rectangle3_y(rectangle3_ys[1338]), .rectangle3_width(rectangle3_widths[1338]), .rectangle3_height(rectangle3_heights[1338]), .rectangle3_weight(rectangle3_weights[1338]), .feature_threshold(feature_thresholds[1338]), .feature_above(feature_aboves[1338]), .feature_below(feature_belows[1338]), .scan_win_std_dev(scan_win_std_dev[1338]), .feature_accum(feature_accums[1338]));
  accum_calculator ac1339(.scan_win(scan_win1339), .rectangle1_x(rectangle1_xs[1339]), .rectangle1_y(rectangle1_ys[1339]), .rectangle1_width(rectangle1_widths[1339]), .rectangle1_height(rectangle1_heights[1339]), .rectangle1_weight(rectangle1_weights[1339]), .rectangle2_x(rectangle2_xs[1339]), .rectangle2_y(rectangle2_ys[1339]), .rectangle2_width(rectangle2_widths[1339]), .rectangle2_height(rectangle2_heights[1339]), .rectangle2_weight(rectangle2_weights[1339]), .rectangle3_x(rectangle3_xs[1339]), .rectangle3_y(rectangle3_ys[1339]), .rectangle3_width(rectangle3_widths[1339]), .rectangle3_height(rectangle3_heights[1339]), .rectangle3_weight(rectangle3_weights[1339]), .feature_threshold(feature_thresholds[1339]), .feature_above(feature_aboves[1339]), .feature_below(feature_belows[1339]), .scan_win_std_dev(scan_win_std_dev[1339]), .feature_accum(feature_accums[1339]));
  accum_calculator ac1340(.scan_win(scan_win1340), .rectangle1_x(rectangle1_xs[1340]), .rectangle1_y(rectangle1_ys[1340]), .rectangle1_width(rectangle1_widths[1340]), .rectangle1_height(rectangle1_heights[1340]), .rectangle1_weight(rectangle1_weights[1340]), .rectangle2_x(rectangle2_xs[1340]), .rectangle2_y(rectangle2_ys[1340]), .rectangle2_width(rectangle2_widths[1340]), .rectangle2_height(rectangle2_heights[1340]), .rectangle2_weight(rectangle2_weights[1340]), .rectangle3_x(rectangle3_xs[1340]), .rectangle3_y(rectangle3_ys[1340]), .rectangle3_width(rectangle3_widths[1340]), .rectangle3_height(rectangle3_heights[1340]), .rectangle3_weight(rectangle3_weights[1340]), .feature_threshold(feature_thresholds[1340]), .feature_above(feature_aboves[1340]), .feature_below(feature_belows[1340]), .scan_win_std_dev(scan_win_std_dev[1340]), .feature_accum(feature_accums[1340]));
  accum_calculator ac1341(.scan_win(scan_win1341), .rectangle1_x(rectangle1_xs[1341]), .rectangle1_y(rectangle1_ys[1341]), .rectangle1_width(rectangle1_widths[1341]), .rectangle1_height(rectangle1_heights[1341]), .rectangle1_weight(rectangle1_weights[1341]), .rectangle2_x(rectangle2_xs[1341]), .rectangle2_y(rectangle2_ys[1341]), .rectangle2_width(rectangle2_widths[1341]), .rectangle2_height(rectangle2_heights[1341]), .rectangle2_weight(rectangle2_weights[1341]), .rectangle3_x(rectangle3_xs[1341]), .rectangle3_y(rectangle3_ys[1341]), .rectangle3_width(rectangle3_widths[1341]), .rectangle3_height(rectangle3_heights[1341]), .rectangle3_weight(rectangle3_weights[1341]), .feature_threshold(feature_thresholds[1341]), .feature_above(feature_aboves[1341]), .feature_below(feature_belows[1341]), .scan_win_std_dev(scan_win_std_dev[1341]), .feature_accum(feature_accums[1341]));
  accum_calculator ac1342(.scan_win(scan_win1342), .rectangle1_x(rectangle1_xs[1342]), .rectangle1_y(rectangle1_ys[1342]), .rectangle1_width(rectangle1_widths[1342]), .rectangle1_height(rectangle1_heights[1342]), .rectangle1_weight(rectangle1_weights[1342]), .rectangle2_x(rectangle2_xs[1342]), .rectangle2_y(rectangle2_ys[1342]), .rectangle2_width(rectangle2_widths[1342]), .rectangle2_height(rectangle2_heights[1342]), .rectangle2_weight(rectangle2_weights[1342]), .rectangle3_x(rectangle3_xs[1342]), .rectangle3_y(rectangle3_ys[1342]), .rectangle3_width(rectangle3_widths[1342]), .rectangle3_height(rectangle3_heights[1342]), .rectangle3_weight(rectangle3_weights[1342]), .feature_threshold(feature_thresholds[1342]), .feature_above(feature_aboves[1342]), .feature_below(feature_belows[1342]), .scan_win_std_dev(scan_win_std_dev[1342]), .feature_accum(feature_accums[1342]));
  accum_calculator ac1343(.scan_win(scan_win1343), .rectangle1_x(rectangle1_xs[1343]), .rectangle1_y(rectangle1_ys[1343]), .rectangle1_width(rectangle1_widths[1343]), .rectangle1_height(rectangle1_heights[1343]), .rectangle1_weight(rectangle1_weights[1343]), .rectangle2_x(rectangle2_xs[1343]), .rectangle2_y(rectangle2_ys[1343]), .rectangle2_width(rectangle2_widths[1343]), .rectangle2_height(rectangle2_heights[1343]), .rectangle2_weight(rectangle2_weights[1343]), .rectangle3_x(rectangle3_xs[1343]), .rectangle3_y(rectangle3_ys[1343]), .rectangle3_width(rectangle3_widths[1343]), .rectangle3_height(rectangle3_heights[1343]), .rectangle3_weight(rectangle3_weights[1343]), .feature_threshold(feature_thresholds[1343]), .feature_above(feature_aboves[1343]), .feature_below(feature_belows[1343]), .scan_win_std_dev(scan_win_std_dev[1343]), .feature_accum(feature_accums[1343]));
  accum_calculator ac1344(.scan_win(scan_win1344), .rectangle1_x(rectangle1_xs[1344]), .rectangle1_y(rectangle1_ys[1344]), .rectangle1_width(rectangle1_widths[1344]), .rectangle1_height(rectangle1_heights[1344]), .rectangle1_weight(rectangle1_weights[1344]), .rectangle2_x(rectangle2_xs[1344]), .rectangle2_y(rectangle2_ys[1344]), .rectangle2_width(rectangle2_widths[1344]), .rectangle2_height(rectangle2_heights[1344]), .rectangle2_weight(rectangle2_weights[1344]), .rectangle3_x(rectangle3_xs[1344]), .rectangle3_y(rectangle3_ys[1344]), .rectangle3_width(rectangle3_widths[1344]), .rectangle3_height(rectangle3_heights[1344]), .rectangle3_weight(rectangle3_weights[1344]), .feature_threshold(feature_thresholds[1344]), .feature_above(feature_aboves[1344]), .feature_below(feature_belows[1344]), .scan_win_std_dev(scan_win_std_dev[1344]), .feature_accum(feature_accums[1344]));
  accum_calculator ac1345(.scan_win(scan_win1345), .rectangle1_x(rectangle1_xs[1345]), .rectangle1_y(rectangle1_ys[1345]), .rectangle1_width(rectangle1_widths[1345]), .rectangle1_height(rectangle1_heights[1345]), .rectangle1_weight(rectangle1_weights[1345]), .rectangle2_x(rectangle2_xs[1345]), .rectangle2_y(rectangle2_ys[1345]), .rectangle2_width(rectangle2_widths[1345]), .rectangle2_height(rectangle2_heights[1345]), .rectangle2_weight(rectangle2_weights[1345]), .rectangle3_x(rectangle3_xs[1345]), .rectangle3_y(rectangle3_ys[1345]), .rectangle3_width(rectangle3_widths[1345]), .rectangle3_height(rectangle3_heights[1345]), .rectangle3_weight(rectangle3_weights[1345]), .feature_threshold(feature_thresholds[1345]), .feature_above(feature_aboves[1345]), .feature_below(feature_belows[1345]), .scan_win_std_dev(scan_win_std_dev[1345]), .feature_accum(feature_accums[1345]));
  accum_calculator ac1346(.scan_win(scan_win1346), .rectangle1_x(rectangle1_xs[1346]), .rectangle1_y(rectangle1_ys[1346]), .rectangle1_width(rectangle1_widths[1346]), .rectangle1_height(rectangle1_heights[1346]), .rectangle1_weight(rectangle1_weights[1346]), .rectangle2_x(rectangle2_xs[1346]), .rectangle2_y(rectangle2_ys[1346]), .rectangle2_width(rectangle2_widths[1346]), .rectangle2_height(rectangle2_heights[1346]), .rectangle2_weight(rectangle2_weights[1346]), .rectangle3_x(rectangle3_xs[1346]), .rectangle3_y(rectangle3_ys[1346]), .rectangle3_width(rectangle3_widths[1346]), .rectangle3_height(rectangle3_heights[1346]), .rectangle3_weight(rectangle3_weights[1346]), .feature_threshold(feature_thresholds[1346]), .feature_above(feature_aboves[1346]), .feature_below(feature_belows[1346]), .scan_win_std_dev(scan_win_std_dev[1346]), .feature_accum(feature_accums[1346]));
  accum_calculator ac1347(.scan_win(scan_win1347), .rectangle1_x(rectangle1_xs[1347]), .rectangle1_y(rectangle1_ys[1347]), .rectangle1_width(rectangle1_widths[1347]), .rectangle1_height(rectangle1_heights[1347]), .rectangle1_weight(rectangle1_weights[1347]), .rectangle2_x(rectangle2_xs[1347]), .rectangle2_y(rectangle2_ys[1347]), .rectangle2_width(rectangle2_widths[1347]), .rectangle2_height(rectangle2_heights[1347]), .rectangle2_weight(rectangle2_weights[1347]), .rectangle3_x(rectangle3_xs[1347]), .rectangle3_y(rectangle3_ys[1347]), .rectangle3_width(rectangle3_widths[1347]), .rectangle3_height(rectangle3_heights[1347]), .rectangle3_weight(rectangle3_weights[1347]), .feature_threshold(feature_thresholds[1347]), .feature_above(feature_aboves[1347]), .feature_below(feature_belows[1347]), .scan_win_std_dev(scan_win_std_dev[1347]), .feature_accum(feature_accums[1347]));
  accum_calculator ac1348(.scan_win(scan_win1348), .rectangle1_x(rectangle1_xs[1348]), .rectangle1_y(rectangle1_ys[1348]), .rectangle1_width(rectangle1_widths[1348]), .rectangle1_height(rectangle1_heights[1348]), .rectangle1_weight(rectangle1_weights[1348]), .rectangle2_x(rectangle2_xs[1348]), .rectangle2_y(rectangle2_ys[1348]), .rectangle2_width(rectangle2_widths[1348]), .rectangle2_height(rectangle2_heights[1348]), .rectangle2_weight(rectangle2_weights[1348]), .rectangle3_x(rectangle3_xs[1348]), .rectangle3_y(rectangle3_ys[1348]), .rectangle3_width(rectangle3_widths[1348]), .rectangle3_height(rectangle3_heights[1348]), .rectangle3_weight(rectangle3_weights[1348]), .feature_threshold(feature_thresholds[1348]), .feature_above(feature_aboves[1348]), .feature_below(feature_belows[1348]), .scan_win_std_dev(scan_win_std_dev[1348]), .feature_accum(feature_accums[1348]));
  accum_calculator ac1349(.scan_win(scan_win1349), .rectangle1_x(rectangle1_xs[1349]), .rectangle1_y(rectangle1_ys[1349]), .rectangle1_width(rectangle1_widths[1349]), .rectangle1_height(rectangle1_heights[1349]), .rectangle1_weight(rectangle1_weights[1349]), .rectangle2_x(rectangle2_xs[1349]), .rectangle2_y(rectangle2_ys[1349]), .rectangle2_width(rectangle2_widths[1349]), .rectangle2_height(rectangle2_heights[1349]), .rectangle2_weight(rectangle2_weights[1349]), .rectangle3_x(rectangle3_xs[1349]), .rectangle3_y(rectangle3_ys[1349]), .rectangle3_width(rectangle3_widths[1349]), .rectangle3_height(rectangle3_heights[1349]), .rectangle3_weight(rectangle3_weights[1349]), .feature_threshold(feature_thresholds[1349]), .feature_above(feature_aboves[1349]), .feature_below(feature_belows[1349]), .scan_win_std_dev(scan_win_std_dev[1349]), .feature_accum(feature_accums[1349]));
  accum_calculator ac1350(.scan_win(scan_win1350), .rectangle1_x(rectangle1_xs[1350]), .rectangle1_y(rectangle1_ys[1350]), .rectangle1_width(rectangle1_widths[1350]), .rectangle1_height(rectangle1_heights[1350]), .rectangle1_weight(rectangle1_weights[1350]), .rectangle2_x(rectangle2_xs[1350]), .rectangle2_y(rectangle2_ys[1350]), .rectangle2_width(rectangle2_widths[1350]), .rectangle2_height(rectangle2_heights[1350]), .rectangle2_weight(rectangle2_weights[1350]), .rectangle3_x(rectangle3_xs[1350]), .rectangle3_y(rectangle3_ys[1350]), .rectangle3_width(rectangle3_widths[1350]), .rectangle3_height(rectangle3_heights[1350]), .rectangle3_weight(rectangle3_weights[1350]), .feature_threshold(feature_thresholds[1350]), .feature_above(feature_aboves[1350]), .feature_below(feature_belows[1350]), .scan_win_std_dev(scan_win_std_dev[1350]), .feature_accum(feature_accums[1350]));
  accum_calculator ac1351(.scan_win(scan_win1351), .rectangle1_x(rectangle1_xs[1351]), .rectangle1_y(rectangle1_ys[1351]), .rectangle1_width(rectangle1_widths[1351]), .rectangle1_height(rectangle1_heights[1351]), .rectangle1_weight(rectangle1_weights[1351]), .rectangle2_x(rectangle2_xs[1351]), .rectangle2_y(rectangle2_ys[1351]), .rectangle2_width(rectangle2_widths[1351]), .rectangle2_height(rectangle2_heights[1351]), .rectangle2_weight(rectangle2_weights[1351]), .rectangle3_x(rectangle3_xs[1351]), .rectangle3_y(rectangle3_ys[1351]), .rectangle3_width(rectangle3_widths[1351]), .rectangle3_height(rectangle3_heights[1351]), .rectangle3_weight(rectangle3_weights[1351]), .feature_threshold(feature_thresholds[1351]), .feature_above(feature_aboves[1351]), .feature_below(feature_belows[1351]), .scan_win_std_dev(scan_win_std_dev[1351]), .feature_accum(feature_accums[1351]));
  accum_calculator ac1352(.scan_win(scan_win1352), .rectangle1_x(rectangle1_xs[1352]), .rectangle1_y(rectangle1_ys[1352]), .rectangle1_width(rectangle1_widths[1352]), .rectangle1_height(rectangle1_heights[1352]), .rectangle1_weight(rectangle1_weights[1352]), .rectangle2_x(rectangle2_xs[1352]), .rectangle2_y(rectangle2_ys[1352]), .rectangle2_width(rectangle2_widths[1352]), .rectangle2_height(rectangle2_heights[1352]), .rectangle2_weight(rectangle2_weights[1352]), .rectangle3_x(rectangle3_xs[1352]), .rectangle3_y(rectangle3_ys[1352]), .rectangle3_width(rectangle3_widths[1352]), .rectangle3_height(rectangle3_heights[1352]), .rectangle3_weight(rectangle3_weights[1352]), .feature_threshold(feature_thresholds[1352]), .feature_above(feature_aboves[1352]), .feature_below(feature_belows[1352]), .scan_win_std_dev(scan_win_std_dev[1352]), .feature_accum(feature_accums[1352]));
  accum_calculator ac1353(.scan_win(scan_win1353), .rectangle1_x(rectangle1_xs[1353]), .rectangle1_y(rectangle1_ys[1353]), .rectangle1_width(rectangle1_widths[1353]), .rectangle1_height(rectangle1_heights[1353]), .rectangle1_weight(rectangle1_weights[1353]), .rectangle2_x(rectangle2_xs[1353]), .rectangle2_y(rectangle2_ys[1353]), .rectangle2_width(rectangle2_widths[1353]), .rectangle2_height(rectangle2_heights[1353]), .rectangle2_weight(rectangle2_weights[1353]), .rectangle3_x(rectangle3_xs[1353]), .rectangle3_y(rectangle3_ys[1353]), .rectangle3_width(rectangle3_widths[1353]), .rectangle3_height(rectangle3_heights[1353]), .rectangle3_weight(rectangle3_weights[1353]), .feature_threshold(feature_thresholds[1353]), .feature_above(feature_aboves[1353]), .feature_below(feature_belows[1353]), .scan_win_std_dev(scan_win_std_dev[1353]), .feature_accum(feature_accums[1353]));
  accum_calculator ac1354(.scan_win(scan_win1354), .rectangle1_x(rectangle1_xs[1354]), .rectangle1_y(rectangle1_ys[1354]), .rectangle1_width(rectangle1_widths[1354]), .rectangle1_height(rectangle1_heights[1354]), .rectangle1_weight(rectangle1_weights[1354]), .rectangle2_x(rectangle2_xs[1354]), .rectangle2_y(rectangle2_ys[1354]), .rectangle2_width(rectangle2_widths[1354]), .rectangle2_height(rectangle2_heights[1354]), .rectangle2_weight(rectangle2_weights[1354]), .rectangle3_x(rectangle3_xs[1354]), .rectangle3_y(rectangle3_ys[1354]), .rectangle3_width(rectangle3_widths[1354]), .rectangle3_height(rectangle3_heights[1354]), .rectangle3_weight(rectangle3_weights[1354]), .feature_threshold(feature_thresholds[1354]), .feature_above(feature_aboves[1354]), .feature_below(feature_belows[1354]), .scan_win_std_dev(scan_win_std_dev[1354]), .feature_accum(feature_accums[1354]));
  accum_calculator ac1355(.scan_win(scan_win1355), .rectangle1_x(rectangle1_xs[1355]), .rectangle1_y(rectangle1_ys[1355]), .rectangle1_width(rectangle1_widths[1355]), .rectangle1_height(rectangle1_heights[1355]), .rectangle1_weight(rectangle1_weights[1355]), .rectangle2_x(rectangle2_xs[1355]), .rectangle2_y(rectangle2_ys[1355]), .rectangle2_width(rectangle2_widths[1355]), .rectangle2_height(rectangle2_heights[1355]), .rectangle2_weight(rectangle2_weights[1355]), .rectangle3_x(rectangle3_xs[1355]), .rectangle3_y(rectangle3_ys[1355]), .rectangle3_width(rectangle3_widths[1355]), .rectangle3_height(rectangle3_heights[1355]), .rectangle3_weight(rectangle3_weights[1355]), .feature_threshold(feature_thresholds[1355]), .feature_above(feature_aboves[1355]), .feature_below(feature_belows[1355]), .scan_win_std_dev(scan_win_std_dev[1355]), .feature_accum(feature_accums[1355]));
  accum_calculator ac1356(.scan_win(scan_win1356), .rectangle1_x(rectangle1_xs[1356]), .rectangle1_y(rectangle1_ys[1356]), .rectangle1_width(rectangle1_widths[1356]), .rectangle1_height(rectangle1_heights[1356]), .rectangle1_weight(rectangle1_weights[1356]), .rectangle2_x(rectangle2_xs[1356]), .rectangle2_y(rectangle2_ys[1356]), .rectangle2_width(rectangle2_widths[1356]), .rectangle2_height(rectangle2_heights[1356]), .rectangle2_weight(rectangle2_weights[1356]), .rectangle3_x(rectangle3_xs[1356]), .rectangle3_y(rectangle3_ys[1356]), .rectangle3_width(rectangle3_widths[1356]), .rectangle3_height(rectangle3_heights[1356]), .rectangle3_weight(rectangle3_weights[1356]), .feature_threshold(feature_thresholds[1356]), .feature_above(feature_aboves[1356]), .feature_below(feature_belows[1356]), .scan_win_std_dev(scan_win_std_dev[1356]), .feature_accum(feature_accums[1356]));
  accum_calculator ac1357(.scan_win(scan_win1357), .rectangle1_x(rectangle1_xs[1357]), .rectangle1_y(rectangle1_ys[1357]), .rectangle1_width(rectangle1_widths[1357]), .rectangle1_height(rectangle1_heights[1357]), .rectangle1_weight(rectangle1_weights[1357]), .rectangle2_x(rectangle2_xs[1357]), .rectangle2_y(rectangle2_ys[1357]), .rectangle2_width(rectangle2_widths[1357]), .rectangle2_height(rectangle2_heights[1357]), .rectangle2_weight(rectangle2_weights[1357]), .rectangle3_x(rectangle3_xs[1357]), .rectangle3_y(rectangle3_ys[1357]), .rectangle3_width(rectangle3_widths[1357]), .rectangle3_height(rectangle3_heights[1357]), .rectangle3_weight(rectangle3_weights[1357]), .feature_threshold(feature_thresholds[1357]), .feature_above(feature_aboves[1357]), .feature_below(feature_belows[1357]), .scan_win_std_dev(scan_win_std_dev[1357]), .feature_accum(feature_accums[1357]));
  accum_calculator ac1358(.scan_win(scan_win1358), .rectangle1_x(rectangle1_xs[1358]), .rectangle1_y(rectangle1_ys[1358]), .rectangle1_width(rectangle1_widths[1358]), .rectangle1_height(rectangle1_heights[1358]), .rectangle1_weight(rectangle1_weights[1358]), .rectangle2_x(rectangle2_xs[1358]), .rectangle2_y(rectangle2_ys[1358]), .rectangle2_width(rectangle2_widths[1358]), .rectangle2_height(rectangle2_heights[1358]), .rectangle2_weight(rectangle2_weights[1358]), .rectangle3_x(rectangle3_xs[1358]), .rectangle3_y(rectangle3_ys[1358]), .rectangle3_width(rectangle3_widths[1358]), .rectangle3_height(rectangle3_heights[1358]), .rectangle3_weight(rectangle3_weights[1358]), .feature_threshold(feature_thresholds[1358]), .feature_above(feature_aboves[1358]), .feature_below(feature_belows[1358]), .scan_win_std_dev(scan_win_std_dev[1358]), .feature_accum(feature_accums[1358]));
  accum_calculator ac1359(.scan_win(scan_win1359), .rectangle1_x(rectangle1_xs[1359]), .rectangle1_y(rectangle1_ys[1359]), .rectangle1_width(rectangle1_widths[1359]), .rectangle1_height(rectangle1_heights[1359]), .rectangle1_weight(rectangle1_weights[1359]), .rectangle2_x(rectangle2_xs[1359]), .rectangle2_y(rectangle2_ys[1359]), .rectangle2_width(rectangle2_widths[1359]), .rectangle2_height(rectangle2_heights[1359]), .rectangle2_weight(rectangle2_weights[1359]), .rectangle3_x(rectangle3_xs[1359]), .rectangle3_y(rectangle3_ys[1359]), .rectangle3_width(rectangle3_widths[1359]), .rectangle3_height(rectangle3_heights[1359]), .rectangle3_weight(rectangle3_weights[1359]), .feature_threshold(feature_thresholds[1359]), .feature_above(feature_aboves[1359]), .feature_below(feature_belows[1359]), .scan_win_std_dev(scan_win_std_dev[1359]), .feature_accum(feature_accums[1359]));
  accum_calculator ac1360(.scan_win(scan_win1360), .rectangle1_x(rectangle1_xs[1360]), .rectangle1_y(rectangle1_ys[1360]), .rectangle1_width(rectangle1_widths[1360]), .rectangle1_height(rectangle1_heights[1360]), .rectangle1_weight(rectangle1_weights[1360]), .rectangle2_x(rectangle2_xs[1360]), .rectangle2_y(rectangle2_ys[1360]), .rectangle2_width(rectangle2_widths[1360]), .rectangle2_height(rectangle2_heights[1360]), .rectangle2_weight(rectangle2_weights[1360]), .rectangle3_x(rectangle3_xs[1360]), .rectangle3_y(rectangle3_ys[1360]), .rectangle3_width(rectangle3_widths[1360]), .rectangle3_height(rectangle3_heights[1360]), .rectangle3_weight(rectangle3_weights[1360]), .feature_threshold(feature_thresholds[1360]), .feature_above(feature_aboves[1360]), .feature_below(feature_belows[1360]), .scan_win_std_dev(scan_win_std_dev[1360]), .feature_accum(feature_accums[1360]));
  accum_calculator ac1361(.scan_win(scan_win1361), .rectangle1_x(rectangle1_xs[1361]), .rectangle1_y(rectangle1_ys[1361]), .rectangle1_width(rectangle1_widths[1361]), .rectangle1_height(rectangle1_heights[1361]), .rectangle1_weight(rectangle1_weights[1361]), .rectangle2_x(rectangle2_xs[1361]), .rectangle2_y(rectangle2_ys[1361]), .rectangle2_width(rectangle2_widths[1361]), .rectangle2_height(rectangle2_heights[1361]), .rectangle2_weight(rectangle2_weights[1361]), .rectangle3_x(rectangle3_xs[1361]), .rectangle3_y(rectangle3_ys[1361]), .rectangle3_width(rectangle3_widths[1361]), .rectangle3_height(rectangle3_heights[1361]), .rectangle3_weight(rectangle3_weights[1361]), .feature_threshold(feature_thresholds[1361]), .feature_above(feature_aboves[1361]), .feature_below(feature_belows[1361]), .scan_win_std_dev(scan_win_std_dev[1361]), .feature_accum(feature_accums[1361]));
  accum_calculator ac1362(.scan_win(scan_win1362), .rectangle1_x(rectangle1_xs[1362]), .rectangle1_y(rectangle1_ys[1362]), .rectangle1_width(rectangle1_widths[1362]), .rectangle1_height(rectangle1_heights[1362]), .rectangle1_weight(rectangle1_weights[1362]), .rectangle2_x(rectangle2_xs[1362]), .rectangle2_y(rectangle2_ys[1362]), .rectangle2_width(rectangle2_widths[1362]), .rectangle2_height(rectangle2_heights[1362]), .rectangle2_weight(rectangle2_weights[1362]), .rectangle3_x(rectangle3_xs[1362]), .rectangle3_y(rectangle3_ys[1362]), .rectangle3_width(rectangle3_widths[1362]), .rectangle3_height(rectangle3_heights[1362]), .rectangle3_weight(rectangle3_weights[1362]), .feature_threshold(feature_thresholds[1362]), .feature_above(feature_aboves[1362]), .feature_below(feature_belows[1362]), .scan_win_std_dev(scan_win_std_dev[1362]), .feature_accum(feature_accums[1362]));
  accum_calculator ac1363(.scan_win(scan_win1363), .rectangle1_x(rectangle1_xs[1363]), .rectangle1_y(rectangle1_ys[1363]), .rectangle1_width(rectangle1_widths[1363]), .rectangle1_height(rectangle1_heights[1363]), .rectangle1_weight(rectangle1_weights[1363]), .rectangle2_x(rectangle2_xs[1363]), .rectangle2_y(rectangle2_ys[1363]), .rectangle2_width(rectangle2_widths[1363]), .rectangle2_height(rectangle2_heights[1363]), .rectangle2_weight(rectangle2_weights[1363]), .rectangle3_x(rectangle3_xs[1363]), .rectangle3_y(rectangle3_ys[1363]), .rectangle3_width(rectangle3_widths[1363]), .rectangle3_height(rectangle3_heights[1363]), .rectangle3_weight(rectangle3_weights[1363]), .feature_threshold(feature_thresholds[1363]), .feature_above(feature_aboves[1363]), .feature_below(feature_belows[1363]), .scan_win_std_dev(scan_win_std_dev[1363]), .feature_accum(feature_accums[1363]));
  accum_calculator ac1364(.scan_win(scan_win1364), .rectangle1_x(rectangle1_xs[1364]), .rectangle1_y(rectangle1_ys[1364]), .rectangle1_width(rectangle1_widths[1364]), .rectangle1_height(rectangle1_heights[1364]), .rectangle1_weight(rectangle1_weights[1364]), .rectangle2_x(rectangle2_xs[1364]), .rectangle2_y(rectangle2_ys[1364]), .rectangle2_width(rectangle2_widths[1364]), .rectangle2_height(rectangle2_heights[1364]), .rectangle2_weight(rectangle2_weights[1364]), .rectangle3_x(rectangle3_xs[1364]), .rectangle3_y(rectangle3_ys[1364]), .rectangle3_width(rectangle3_widths[1364]), .rectangle3_height(rectangle3_heights[1364]), .rectangle3_weight(rectangle3_weights[1364]), .feature_threshold(feature_thresholds[1364]), .feature_above(feature_aboves[1364]), .feature_below(feature_belows[1364]), .scan_win_std_dev(scan_win_std_dev[1364]), .feature_accum(feature_accums[1364]));
  accum_calculator ac1365(.scan_win(scan_win1365), .rectangle1_x(rectangle1_xs[1365]), .rectangle1_y(rectangle1_ys[1365]), .rectangle1_width(rectangle1_widths[1365]), .rectangle1_height(rectangle1_heights[1365]), .rectangle1_weight(rectangle1_weights[1365]), .rectangle2_x(rectangle2_xs[1365]), .rectangle2_y(rectangle2_ys[1365]), .rectangle2_width(rectangle2_widths[1365]), .rectangle2_height(rectangle2_heights[1365]), .rectangle2_weight(rectangle2_weights[1365]), .rectangle3_x(rectangle3_xs[1365]), .rectangle3_y(rectangle3_ys[1365]), .rectangle3_width(rectangle3_widths[1365]), .rectangle3_height(rectangle3_heights[1365]), .rectangle3_weight(rectangle3_weights[1365]), .feature_threshold(feature_thresholds[1365]), .feature_above(feature_aboves[1365]), .feature_below(feature_belows[1365]), .scan_win_std_dev(scan_win_std_dev[1365]), .feature_accum(feature_accums[1365]));
  accum_calculator ac1366(.scan_win(scan_win1366), .rectangle1_x(rectangle1_xs[1366]), .rectangle1_y(rectangle1_ys[1366]), .rectangle1_width(rectangle1_widths[1366]), .rectangle1_height(rectangle1_heights[1366]), .rectangle1_weight(rectangle1_weights[1366]), .rectangle2_x(rectangle2_xs[1366]), .rectangle2_y(rectangle2_ys[1366]), .rectangle2_width(rectangle2_widths[1366]), .rectangle2_height(rectangle2_heights[1366]), .rectangle2_weight(rectangle2_weights[1366]), .rectangle3_x(rectangle3_xs[1366]), .rectangle3_y(rectangle3_ys[1366]), .rectangle3_width(rectangle3_widths[1366]), .rectangle3_height(rectangle3_heights[1366]), .rectangle3_weight(rectangle3_weights[1366]), .feature_threshold(feature_thresholds[1366]), .feature_above(feature_aboves[1366]), .feature_below(feature_belows[1366]), .scan_win_std_dev(scan_win_std_dev[1366]), .feature_accum(feature_accums[1366]));
  accum_calculator ac1367(.scan_win(scan_win1367), .rectangle1_x(rectangle1_xs[1367]), .rectangle1_y(rectangle1_ys[1367]), .rectangle1_width(rectangle1_widths[1367]), .rectangle1_height(rectangle1_heights[1367]), .rectangle1_weight(rectangle1_weights[1367]), .rectangle2_x(rectangle2_xs[1367]), .rectangle2_y(rectangle2_ys[1367]), .rectangle2_width(rectangle2_widths[1367]), .rectangle2_height(rectangle2_heights[1367]), .rectangle2_weight(rectangle2_weights[1367]), .rectangle3_x(rectangle3_xs[1367]), .rectangle3_y(rectangle3_ys[1367]), .rectangle3_width(rectangle3_widths[1367]), .rectangle3_height(rectangle3_heights[1367]), .rectangle3_weight(rectangle3_weights[1367]), .feature_threshold(feature_thresholds[1367]), .feature_above(feature_aboves[1367]), .feature_below(feature_belows[1367]), .scan_win_std_dev(scan_win_std_dev[1367]), .feature_accum(feature_accums[1367]));
  accum_calculator ac1368(.scan_win(scan_win1368), .rectangle1_x(rectangle1_xs[1368]), .rectangle1_y(rectangle1_ys[1368]), .rectangle1_width(rectangle1_widths[1368]), .rectangle1_height(rectangle1_heights[1368]), .rectangle1_weight(rectangle1_weights[1368]), .rectangle2_x(rectangle2_xs[1368]), .rectangle2_y(rectangle2_ys[1368]), .rectangle2_width(rectangle2_widths[1368]), .rectangle2_height(rectangle2_heights[1368]), .rectangle2_weight(rectangle2_weights[1368]), .rectangle3_x(rectangle3_xs[1368]), .rectangle3_y(rectangle3_ys[1368]), .rectangle3_width(rectangle3_widths[1368]), .rectangle3_height(rectangle3_heights[1368]), .rectangle3_weight(rectangle3_weights[1368]), .feature_threshold(feature_thresholds[1368]), .feature_above(feature_aboves[1368]), .feature_below(feature_belows[1368]), .scan_win_std_dev(scan_win_std_dev[1368]), .feature_accum(feature_accums[1368]));
  accum_calculator ac1369(.scan_win(scan_win1369), .rectangle1_x(rectangle1_xs[1369]), .rectangle1_y(rectangle1_ys[1369]), .rectangle1_width(rectangle1_widths[1369]), .rectangle1_height(rectangle1_heights[1369]), .rectangle1_weight(rectangle1_weights[1369]), .rectangle2_x(rectangle2_xs[1369]), .rectangle2_y(rectangle2_ys[1369]), .rectangle2_width(rectangle2_widths[1369]), .rectangle2_height(rectangle2_heights[1369]), .rectangle2_weight(rectangle2_weights[1369]), .rectangle3_x(rectangle3_xs[1369]), .rectangle3_y(rectangle3_ys[1369]), .rectangle3_width(rectangle3_widths[1369]), .rectangle3_height(rectangle3_heights[1369]), .rectangle3_weight(rectangle3_weights[1369]), .feature_threshold(feature_thresholds[1369]), .feature_above(feature_aboves[1369]), .feature_below(feature_belows[1369]), .scan_win_std_dev(scan_win_std_dev[1369]), .feature_accum(feature_accums[1369]));
  accum_calculator ac1370(.scan_win(scan_win1370), .rectangle1_x(rectangle1_xs[1370]), .rectangle1_y(rectangle1_ys[1370]), .rectangle1_width(rectangle1_widths[1370]), .rectangle1_height(rectangle1_heights[1370]), .rectangle1_weight(rectangle1_weights[1370]), .rectangle2_x(rectangle2_xs[1370]), .rectangle2_y(rectangle2_ys[1370]), .rectangle2_width(rectangle2_widths[1370]), .rectangle2_height(rectangle2_heights[1370]), .rectangle2_weight(rectangle2_weights[1370]), .rectangle3_x(rectangle3_xs[1370]), .rectangle3_y(rectangle3_ys[1370]), .rectangle3_width(rectangle3_widths[1370]), .rectangle3_height(rectangle3_heights[1370]), .rectangle3_weight(rectangle3_weights[1370]), .feature_threshold(feature_thresholds[1370]), .feature_above(feature_aboves[1370]), .feature_below(feature_belows[1370]), .scan_win_std_dev(scan_win_std_dev[1370]), .feature_accum(feature_accums[1370]));
  accum_calculator ac1371(.scan_win(scan_win1371), .rectangle1_x(rectangle1_xs[1371]), .rectangle1_y(rectangle1_ys[1371]), .rectangle1_width(rectangle1_widths[1371]), .rectangle1_height(rectangle1_heights[1371]), .rectangle1_weight(rectangle1_weights[1371]), .rectangle2_x(rectangle2_xs[1371]), .rectangle2_y(rectangle2_ys[1371]), .rectangle2_width(rectangle2_widths[1371]), .rectangle2_height(rectangle2_heights[1371]), .rectangle2_weight(rectangle2_weights[1371]), .rectangle3_x(rectangle3_xs[1371]), .rectangle3_y(rectangle3_ys[1371]), .rectangle3_width(rectangle3_widths[1371]), .rectangle3_height(rectangle3_heights[1371]), .rectangle3_weight(rectangle3_weights[1371]), .feature_threshold(feature_thresholds[1371]), .feature_above(feature_aboves[1371]), .feature_below(feature_belows[1371]), .scan_win_std_dev(scan_win_std_dev[1371]), .feature_accum(feature_accums[1371]));
  accum_calculator ac1372(.scan_win(scan_win1372), .rectangle1_x(rectangle1_xs[1372]), .rectangle1_y(rectangle1_ys[1372]), .rectangle1_width(rectangle1_widths[1372]), .rectangle1_height(rectangle1_heights[1372]), .rectangle1_weight(rectangle1_weights[1372]), .rectangle2_x(rectangle2_xs[1372]), .rectangle2_y(rectangle2_ys[1372]), .rectangle2_width(rectangle2_widths[1372]), .rectangle2_height(rectangle2_heights[1372]), .rectangle2_weight(rectangle2_weights[1372]), .rectangle3_x(rectangle3_xs[1372]), .rectangle3_y(rectangle3_ys[1372]), .rectangle3_width(rectangle3_widths[1372]), .rectangle3_height(rectangle3_heights[1372]), .rectangle3_weight(rectangle3_weights[1372]), .feature_threshold(feature_thresholds[1372]), .feature_above(feature_aboves[1372]), .feature_below(feature_belows[1372]), .scan_win_std_dev(scan_win_std_dev[1372]), .feature_accum(feature_accums[1372]));
  accum_calculator ac1373(.scan_win(scan_win1373), .rectangle1_x(rectangle1_xs[1373]), .rectangle1_y(rectangle1_ys[1373]), .rectangle1_width(rectangle1_widths[1373]), .rectangle1_height(rectangle1_heights[1373]), .rectangle1_weight(rectangle1_weights[1373]), .rectangle2_x(rectangle2_xs[1373]), .rectangle2_y(rectangle2_ys[1373]), .rectangle2_width(rectangle2_widths[1373]), .rectangle2_height(rectangle2_heights[1373]), .rectangle2_weight(rectangle2_weights[1373]), .rectangle3_x(rectangle3_xs[1373]), .rectangle3_y(rectangle3_ys[1373]), .rectangle3_width(rectangle3_widths[1373]), .rectangle3_height(rectangle3_heights[1373]), .rectangle3_weight(rectangle3_weights[1373]), .feature_threshold(feature_thresholds[1373]), .feature_above(feature_aboves[1373]), .feature_below(feature_belows[1373]), .scan_win_std_dev(scan_win_std_dev[1373]), .feature_accum(feature_accums[1373]));
  accum_calculator ac1374(.scan_win(scan_win1374), .rectangle1_x(rectangle1_xs[1374]), .rectangle1_y(rectangle1_ys[1374]), .rectangle1_width(rectangle1_widths[1374]), .rectangle1_height(rectangle1_heights[1374]), .rectangle1_weight(rectangle1_weights[1374]), .rectangle2_x(rectangle2_xs[1374]), .rectangle2_y(rectangle2_ys[1374]), .rectangle2_width(rectangle2_widths[1374]), .rectangle2_height(rectangle2_heights[1374]), .rectangle2_weight(rectangle2_weights[1374]), .rectangle3_x(rectangle3_xs[1374]), .rectangle3_y(rectangle3_ys[1374]), .rectangle3_width(rectangle3_widths[1374]), .rectangle3_height(rectangle3_heights[1374]), .rectangle3_weight(rectangle3_weights[1374]), .feature_threshold(feature_thresholds[1374]), .feature_above(feature_aboves[1374]), .feature_below(feature_belows[1374]), .scan_win_std_dev(scan_win_std_dev[1374]), .feature_accum(feature_accums[1374]));
  accum_calculator ac1375(.scan_win(scan_win1375), .rectangle1_x(rectangle1_xs[1375]), .rectangle1_y(rectangle1_ys[1375]), .rectangle1_width(rectangle1_widths[1375]), .rectangle1_height(rectangle1_heights[1375]), .rectangle1_weight(rectangle1_weights[1375]), .rectangle2_x(rectangle2_xs[1375]), .rectangle2_y(rectangle2_ys[1375]), .rectangle2_width(rectangle2_widths[1375]), .rectangle2_height(rectangle2_heights[1375]), .rectangle2_weight(rectangle2_weights[1375]), .rectangle3_x(rectangle3_xs[1375]), .rectangle3_y(rectangle3_ys[1375]), .rectangle3_width(rectangle3_widths[1375]), .rectangle3_height(rectangle3_heights[1375]), .rectangle3_weight(rectangle3_weights[1375]), .feature_threshold(feature_thresholds[1375]), .feature_above(feature_aboves[1375]), .feature_below(feature_belows[1375]), .scan_win_std_dev(scan_win_std_dev[1375]), .feature_accum(feature_accums[1375]));
  accum_calculator ac1376(.scan_win(scan_win1376), .rectangle1_x(rectangle1_xs[1376]), .rectangle1_y(rectangle1_ys[1376]), .rectangle1_width(rectangle1_widths[1376]), .rectangle1_height(rectangle1_heights[1376]), .rectangle1_weight(rectangle1_weights[1376]), .rectangle2_x(rectangle2_xs[1376]), .rectangle2_y(rectangle2_ys[1376]), .rectangle2_width(rectangle2_widths[1376]), .rectangle2_height(rectangle2_heights[1376]), .rectangle2_weight(rectangle2_weights[1376]), .rectangle3_x(rectangle3_xs[1376]), .rectangle3_y(rectangle3_ys[1376]), .rectangle3_width(rectangle3_widths[1376]), .rectangle3_height(rectangle3_heights[1376]), .rectangle3_weight(rectangle3_weights[1376]), .feature_threshold(feature_thresholds[1376]), .feature_above(feature_aboves[1376]), .feature_below(feature_belows[1376]), .scan_win_std_dev(scan_win_std_dev[1376]), .feature_accum(feature_accums[1376]));
  accum_calculator ac1377(.scan_win(scan_win1377), .rectangle1_x(rectangle1_xs[1377]), .rectangle1_y(rectangle1_ys[1377]), .rectangle1_width(rectangle1_widths[1377]), .rectangle1_height(rectangle1_heights[1377]), .rectangle1_weight(rectangle1_weights[1377]), .rectangle2_x(rectangle2_xs[1377]), .rectangle2_y(rectangle2_ys[1377]), .rectangle2_width(rectangle2_widths[1377]), .rectangle2_height(rectangle2_heights[1377]), .rectangle2_weight(rectangle2_weights[1377]), .rectangle3_x(rectangle3_xs[1377]), .rectangle3_y(rectangle3_ys[1377]), .rectangle3_width(rectangle3_widths[1377]), .rectangle3_height(rectangle3_heights[1377]), .rectangle3_weight(rectangle3_weights[1377]), .feature_threshold(feature_thresholds[1377]), .feature_above(feature_aboves[1377]), .feature_below(feature_belows[1377]), .scan_win_std_dev(scan_win_std_dev[1377]), .feature_accum(feature_accums[1377]));
  accum_calculator ac1378(.scan_win(scan_win1378), .rectangle1_x(rectangle1_xs[1378]), .rectangle1_y(rectangle1_ys[1378]), .rectangle1_width(rectangle1_widths[1378]), .rectangle1_height(rectangle1_heights[1378]), .rectangle1_weight(rectangle1_weights[1378]), .rectangle2_x(rectangle2_xs[1378]), .rectangle2_y(rectangle2_ys[1378]), .rectangle2_width(rectangle2_widths[1378]), .rectangle2_height(rectangle2_heights[1378]), .rectangle2_weight(rectangle2_weights[1378]), .rectangle3_x(rectangle3_xs[1378]), .rectangle3_y(rectangle3_ys[1378]), .rectangle3_width(rectangle3_widths[1378]), .rectangle3_height(rectangle3_heights[1378]), .rectangle3_weight(rectangle3_weights[1378]), .feature_threshold(feature_thresholds[1378]), .feature_above(feature_aboves[1378]), .feature_below(feature_belows[1378]), .scan_win_std_dev(scan_win_std_dev[1378]), .feature_accum(feature_accums[1378]));
  accum_calculator ac1379(.scan_win(scan_win1379), .rectangle1_x(rectangle1_xs[1379]), .rectangle1_y(rectangle1_ys[1379]), .rectangle1_width(rectangle1_widths[1379]), .rectangle1_height(rectangle1_heights[1379]), .rectangle1_weight(rectangle1_weights[1379]), .rectangle2_x(rectangle2_xs[1379]), .rectangle2_y(rectangle2_ys[1379]), .rectangle2_width(rectangle2_widths[1379]), .rectangle2_height(rectangle2_heights[1379]), .rectangle2_weight(rectangle2_weights[1379]), .rectangle3_x(rectangle3_xs[1379]), .rectangle3_y(rectangle3_ys[1379]), .rectangle3_width(rectangle3_widths[1379]), .rectangle3_height(rectangle3_heights[1379]), .rectangle3_weight(rectangle3_weights[1379]), .feature_threshold(feature_thresholds[1379]), .feature_above(feature_aboves[1379]), .feature_below(feature_belows[1379]), .scan_win_std_dev(scan_win_std_dev[1379]), .feature_accum(feature_accums[1379]));
  accum_calculator ac1380(.scan_win(scan_win1380), .rectangle1_x(rectangle1_xs[1380]), .rectangle1_y(rectangle1_ys[1380]), .rectangle1_width(rectangle1_widths[1380]), .rectangle1_height(rectangle1_heights[1380]), .rectangle1_weight(rectangle1_weights[1380]), .rectangle2_x(rectangle2_xs[1380]), .rectangle2_y(rectangle2_ys[1380]), .rectangle2_width(rectangle2_widths[1380]), .rectangle2_height(rectangle2_heights[1380]), .rectangle2_weight(rectangle2_weights[1380]), .rectangle3_x(rectangle3_xs[1380]), .rectangle3_y(rectangle3_ys[1380]), .rectangle3_width(rectangle3_widths[1380]), .rectangle3_height(rectangle3_heights[1380]), .rectangle3_weight(rectangle3_weights[1380]), .feature_threshold(feature_thresholds[1380]), .feature_above(feature_aboves[1380]), .feature_below(feature_belows[1380]), .scan_win_std_dev(scan_win_std_dev[1380]), .feature_accum(feature_accums[1380]));
  accum_calculator ac1381(.scan_win(scan_win1381), .rectangle1_x(rectangle1_xs[1381]), .rectangle1_y(rectangle1_ys[1381]), .rectangle1_width(rectangle1_widths[1381]), .rectangle1_height(rectangle1_heights[1381]), .rectangle1_weight(rectangle1_weights[1381]), .rectangle2_x(rectangle2_xs[1381]), .rectangle2_y(rectangle2_ys[1381]), .rectangle2_width(rectangle2_widths[1381]), .rectangle2_height(rectangle2_heights[1381]), .rectangle2_weight(rectangle2_weights[1381]), .rectangle3_x(rectangle3_xs[1381]), .rectangle3_y(rectangle3_ys[1381]), .rectangle3_width(rectangle3_widths[1381]), .rectangle3_height(rectangle3_heights[1381]), .rectangle3_weight(rectangle3_weights[1381]), .feature_threshold(feature_thresholds[1381]), .feature_above(feature_aboves[1381]), .feature_below(feature_belows[1381]), .scan_win_std_dev(scan_win_std_dev[1381]), .feature_accum(feature_accums[1381]));
  accum_calculator ac1382(.scan_win(scan_win1382), .rectangle1_x(rectangle1_xs[1382]), .rectangle1_y(rectangle1_ys[1382]), .rectangle1_width(rectangle1_widths[1382]), .rectangle1_height(rectangle1_heights[1382]), .rectangle1_weight(rectangle1_weights[1382]), .rectangle2_x(rectangle2_xs[1382]), .rectangle2_y(rectangle2_ys[1382]), .rectangle2_width(rectangle2_widths[1382]), .rectangle2_height(rectangle2_heights[1382]), .rectangle2_weight(rectangle2_weights[1382]), .rectangle3_x(rectangle3_xs[1382]), .rectangle3_y(rectangle3_ys[1382]), .rectangle3_width(rectangle3_widths[1382]), .rectangle3_height(rectangle3_heights[1382]), .rectangle3_weight(rectangle3_weights[1382]), .feature_threshold(feature_thresholds[1382]), .feature_above(feature_aboves[1382]), .feature_below(feature_belows[1382]), .scan_win_std_dev(scan_win_std_dev[1382]), .feature_accum(feature_accums[1382]));
  accum_calculator ac1383(.scan_win(scan_win1383), .rectangle1_x(rectangle1_xs[1383]), .rectangle1_y(rectangle1_ys[1383]), .rectangle1_width(rectangle1_widths[1383]), .rectangle1_height(rectangle1_heights[1383]), .rectangle1_weight(rectangle1_weights[1383]), .rectangle2_x(rectangle2_xs[1383]), .rectangle2_y(rectangle2_ys[1383]), .rectangle2_width(rectangle2_widths[1383]), .rectangle2_height(rectangle2_heights[1383]), .rectangle2_weight(rectangle2_weights[1383]), .rectangle3_x(rectangle3_xs[1383]), .rectangle3_y(rectangle3_ys[1383]), .rectangle3_width(rectangle3_widths[1383]), .rectangle3_height(rectangle3_heights[1383]), .rectangle3_weight(rectangle3_weights[1383]), .feature_threshold(feature_thresholds[1383]), .feature_above(feature_aboves[1383]), .feature_below(feature_belows[1383]), .scan_win_std_dev(scan_win_std_dev[1383]), .feature_accum(feature_accums[1383]));
  accum_calculator ac1384(.scan_win(scan_win1384), .rectangle1_x(rectangle1_xs[1384]), .rectangle1_y(rectangle1_ys[1384]), .rectangle1_width(rectangle1_widths[1384]), .rectangle1_height(rectangle1_heights[1384]), .rectangle1_weight(rectangle1_weights[1384]), .rectangle2_x(rectangle2_xs[1384]), .rectangle2_y(rectangle2_ys[1384]), .rectangle2_width(rectangle2_widths[1384]), .rectangle2_height(rectangle2_heights[1384]), .rectangle2_weight(rectangle2_weights[1384]), .rectangle3_x(rectangle3_xs[1384]), .rectangle3_y(rectangle3_ys[1384]), .rectangle3_width(rectangle3_widths[1384]), .rectangle3_height(rectangle3_heights[1384]), .rectangle3_weight(rectangle3_weights[1384]), .feature_threshold(feature_thresholds[1384]), .feature_above(feature_aboves[1384]), .feature_below(feature_belows[1384]), .scan_win_std_dev(scan_win_std_dev[1384]), .feature_accum(feature_accums[1384]));
  accum_calculator ac1385(.scan_win(scan_win1385), .rectangle1_x(rectangle1_xs[1385]), .rectangle1_y(rectangle1_ys[1385]), .rectangle1_width(rectangle1_widths[1385]), .rectangle1_height(rectangle1_heights[1385]), .rectangle1_weight(rectangle1_weights[1385]), .rectangle2_x(rectangle2_xs[1385]), .rectangle2_y(rectangle2_ys[1385]), .rectangle2_width(rectangle2_widths[1385]), .rectangle2_height(rectangle2_heights[1385]), .rectangle2_weight(rectangle2_weights[1385]), .rectangle3_x(rectangle3_xs[1385]), .rectangle3_y(rectangle3_ys[1385]), .rectangle3_width(rectangle3_widths[1385]), .rectangle3_height(rectangle3_heights[1385]), .rectangle3_weight(rectangle3_weights[1385]), .feature_threshold(feature_thresholds[1385]), .feature_above(feature_aboves[1385]), .feature_below(feature_belows[1385]), .scan_win_std_dev(scan_win_std_dev[1385]), .feature_accum(feature_accums[1385]));
  accum_calculator ac1386(.scan_win(scan_win1386), .rectangle1_x(rectangle1_xs[1386]), .rectangle1_y(rectangle1_ys[1386]), .rectangle1_width(rectangle1_widths[1386]), .rectangle1_height(rectangle1_heights[1386]), .rectangle1_weight(rectangle1_weights[1386]), .rectangle2_x(rectangle2_xs[1386]), .rectangle2_y(rectangle2_ys[1386]), .rectangle2_width(rectangle2_widths[1386]), .rectangle2_height(rectangle2_heights[1386]), .rectangle2_weight(rectangle2_weights[1386]), .rectangle3_x(rectangle3_xs[1386]), .rectangle3_y(rectangle3_ys[1386]), .rectangle3_width(rectangle3_widths[1386]), .rectangle3_height(rectangle3_heights[1386]), .rectangle3_weight(rectangle3_weights[1386]), .feature_threshold(feature_thresholds[1386]), .feature_above(feature_aboves[1386]), .feature_below(feature_belows[1386]), .scan_win_std_dev(scan_win_std_dev[1386]), .feature_accum(feature_accums[1386]));
  accum_calculator ac1387(.scan_win(scan_win1387), .rectangle1_x(rectangle1_xs[1387]), .rectangle1_y(rectangle1_ys[1387]), .rectangle1_width(rectangle1_widths[1387]), .rectangle1_height(rectangle1_heights[1387]), .rectangle1_weight(rectangle1_weights[1387]), .rectangle2_x(rectangle2_xs[1387]), .rectangle2_y(rectangle2_ys[1387]), .rectangle2_width(rectangle2_widths[1387]), .rectangle2_height(rectangle2_heights[1387]), .rectangle2_weight(rectangle2_weights[1387]), .rectangle3_x(rectangle3_xs[1387]), .rectangle3_y(rectangle3_ys[1387]), .rectangle3_width(rectangle3_widths[1387]), .rectangle3_height(rectangle3_heights[1387]), .rectangle3_weight(rectangle3_weights[1387]), .feature_threshold(feature_thresholds[1387]), .feature_above(feature_aboves[1387]), .feature_below(feature_belows[1387]), .scan_win_std_dev(scan_win_std_dev[1387]), .feature_accum(feature_accums[1387]));
  accum_calculator ac1388(.scan_win(scan_win1388), .rectangle1_x(rectangle1_xs[1388]), .rectangle1_y(rectangle1_ys[1388]), .rectangle1_width(rectangle1_widths[1388]), .rectangle1_height(rectangle1_heights[1388]), .rectangle1_weight(rectangle1_weights[1388]), .rectangle2_x(rectangle2_xs[1388]), .rectangle2_y(rectangle2_ys[1388]), .rectangle2_width(rectangle2_widths[1388]), .rectangle2_height(rectangle2_heights[1388]), .rectangle2_weight(rectangle2_weights[1388]), .rectangle3_x(rectangle3_xs[1388]), .rectangle3_y(rectangle3_ys[1388]), .rectangle3_width(rectangle3_widths[1388]), .rectangle3_height(rectangle3_heights[1388]), .rectangle3_weight(rectangle3_weights[1388]), .feature_threshold(feature_thresholds[1388]), .feature_above(feature_aboves[1388]), .feature_below(feature_belows[1388]), .scan_win_std_dev(scan_win_std_dev[1388]), .feature_accum(feature_accums[1388]));
  accum_calculator ac1389(.scan_win(scan_win1389), .rectangle1_x(rectangle1_xs[1389]), .rectangle1_y(rectangle1_ys[1389]), .rectangle1_width(rectangle1_widths[1389]), .rectangle1_height(rectangle1_heights[1389]), .rectangle1_weight(rectangle1_weights[1389]), .rectangle2_x(rectangle2_xs[1389]), .rectangle2_y(rectangle2_ys[1389]), .rectangle2_width(rectangle2_widths[1389]), .rectangle2_height(rectangle2_heights[1389]), .rectangle2_weight(rectangle2_weights[1389]), .rectangle3_x(rectangle3_xs[1389]), .rectangle3_y(rectangle3_ys[1389]), .rectangle3_width(rectangle3_widths[1389]), .rectangle3_height(rectangle3_heights[1389]), .rectangle3_weight(rectangle3_weights[1389]), .feature_threshold(feature_thresholds[1389]), .feature_above(feature_aboves[1389]), .feature_below(feature_belows[1389]), .scan_win_std_dev(scan_win_std_dev[1389]), .feature_accum(feature_accums[1389]));
  accum_calculator ac1390(.scan_win(scan_win1390), .rectangle1_x(rectangle1_xs[1390]), .rectangle1_y(rectangle1_ys[1390]), .rectangle1_width(rectangle1_widths[1390]), .rectangle1_height(rectangle1_heights[1390]), .rectangle1_weight(rectangle1_weights[1390]), .rectangle2_x(rectangle2_xs[1390]), .rectangle2_y(rectangle2_ys[1390]), .rectangle2_width(rectangle2_widths[1390]), .rectangle2_height(rectangle2_heights[1390]), .rectangle2_weight(rectangle2_weights[1390]), .rectangle3_x(rectangle3_xs[1390]), .rectangle3_y(rectangle3_ys[1390]), .rectangle3_width(rectangle3_widths[1390]), .rectangle3_height(rectangle3_heights[1390]), .rectangle3_weight(rectangle3_weights[1390]), .feature_threshold(feature_thresholds[1390]), .feature_above(feature_aboves[1390]), .feature_below(feature_belows[1390]), .scan_win_std_dev(scan_win_std_dev[1390]), .feature_accum(feature_accums[1390]));
  accum_calculator ac1391(.scan_win(scan_win1391), .rectangle1_x(rectangle1_xs[1391]), .rectangle1_y(rectangle1_ys[1391]), .rectangle1_width(rectangle1_widths[1391]), .rectangle1_height(rectangle1_heights[1391]), .rectangle1_weight(rectangle1_weights[1391]), .rectangle2_x(rectangle2_xs[1391]), .rectangle2_y(rectangle2_ys[1391]), .rectangle2_width(rectangle2_widths[1391]), .rectangle2_height(rectangle2_heights[1391]), .rectangle2_weight(rectangle2_weights[1391]), .rectangle3_x(rectangle3_xs[1391]), .rectangle3_y(rectangle3_ys[1391]), .rectangle3_width(rectangle3_widths[1391]), .rectangle3_height(rectangle3_heights[1391]), .rectangle3_weight(rectangle3_weights[1391]), .feature_threshold(feature_thresholds[1391]), .feature_above(feature_aboves[1391]), .feature_below(feature_belows[1391]), .scan_win_std_dev(scan_win_std_dev[1391]), .feature_accum(feature_accums[1391]));
  accum_calculator ac1392(.scan_win(scan_win1392), .rectangle1_x(rectangle1_xs[1392]), .rectangle1_y(rectangle1_ys[1392]), .rectangle1_width(rectangle1_widths[1392]), .rectangle1_height(rectangle1_heights[1392]), .rectangle1_weight(rectangle1_weights[1392]), .rectangle2_x(rectangle2_xs[1392]), .rectangle2_y(rectangle2_ys[1392]), .rectangle2_width(rectangle2_widths[1392]), .rectangle2_height(rectangle2_heights[1392]), .rectangle2_weight(rectangle2_weights[1392]), .rectangle3_x(rectangle3_xs[1392]), .rectangle3_y(rectangle3_ys[1392]), .rectangle3_width(rectangle3_widths[1392]), .rectangle3_height(rectangle3_heights[1392]), .rectangle3_weight(rectangle3_weights[1392]), .feature_threshold(feature_thresholds[1392]), .feature_above(feature_aboves[1392]), .feature_below(feature_belows[1392]), .scan_win_std_dev(scan_win_std_dev[1392]), .feature_accum(feature_accums[1392]));
  accum_calculator ac1393(.scan_win(scan_win1393), .rectangle1_x(rectangle1_xs[1393]), .rectangle1_y(rectangle1_ys[1393]), .rectangle1_width(rectangle1_widths[1393]), .rectangle1_height(rectangle1_heights[1393]), .rectangle1_weight(rectangle1_weights[1393]), .rectangle2_x(rectangle2_xs[1393]), .rectangle2_y(rectangle2_ys[1393]), .rectangle2_width(rectangle2_widths[1393]), .rectangle2_height(rectangle2_heights[1393]), .rectangle2_weight(rectangle2_weights[1393]), .rectangle3_x(rectangle3_xs[1393]), .rectangle3_y(rectangle3_ys[1393]), .rectangle3_width(rectangle3_widths[1393]), .rectangle3_height(rectangle3_heights[1393]), .rectangle3_weight(rectangle3_weights[1393]), .feature_threshold(feature_thresholds[1393]), .feature_above(feature_aboves[1393]), .feature_below(feature_belows[1393]), .scan_win_std_dev(scan_win_std_dev[1393]), .feature_accum(feature_accums[1393]));
  accum_calculator ac1394(.scan_win(scan_win1394), .rectangle1_x(rectangle1_xs[1394]), .rectangle1_y(rectangle1_ys[1394]), .rectangle1_width(rectangle1_widths[1394]), .rectangle1_height(rectangle1_heights[1394]), .rectangle1_weight(rectangle1_weights[1394]), .rectangle2_x(rectangle2_xs[1394]), .rectangle2_y(rectangle2_ys[1394]), .rectangle2_width(rectangle2_widths[1394]), .rectangle2_height(rectangle2_heights[1394]), .rectangle2_weight(rectangle2_weights[1394]), .rectangle3_x(rectangle3_xs[1394]), .rectangle3_y(rectangle3_ys[1394]), .rectangle3_width(rectangle3_widths[1394]), .rectangle3_height(rectangle3_heights[1394]), .rectangle3_weight(rectangle3_weights[1394]), .feature_threshold(feature_thresholds[1394]), .feature_above(feature_aboves[1394]), .feature_below(feature_belows[1394]), .scan_win_std_dev(scan_win_std_dev[1394]), .feature_accum(feature_accums[1394]));
  accum_calculator ac1395(.scan_win(scan_win1395), .rectangle1_x(rectangle1_xs[1395]), .rectangle1_y(rectangle1_ys[1395]), .rectangle1_width(rectangle1_widths[1395]), .rectangle1_height(rectangle1_heights[1395]), .rectangle1_weight(rectangle1_weights[1395]), .rectangle2_x(rectangle2_xs[1395]), .rectangle2_y(rectangle2_ys[1395]), .rectangle2_width(rectangle2_widths[1395]), .rectangle2_height(rectangle2_heights[1395]), .rectangle2_weight(rectangle2_weights[1395]), .rectangle3_x(rectangle3_xs[1395]), .rectangle3_y(rectangle3_ys[1395]), .rectangle3_width(rectangle3_widths[1395]), .rectangle3_height(rectangle3_heights[1395]), .rectangle3_weight(rectangle3_weights[1395]), .feature_threshold(feature_thresholds[1395]), .feature_above(feature_aboves[1395]), .feature_below(feature_belows[1395]), .scan_win_std_dev(scan_win_std_dev[1395]), .feature_accum(feature_accums[1395]));
  accum_calculator ac1396(.scan_win(scan_win1396), .rectangle1_x(rectangle1_xs[1396]), .rectangle1_y(rectangle1_ys[1396]), .rectangle1_width(rectangle1_widths[1396]), .rectangle1_height(rectangle1_heights[1396]), .rectangle1_weight(rectangle1_weights[1396]), .rectangle2_x(rectangle2_xs[1396]), .rectangle2_y(rectangle2_ys[1396]), .rectangle2_width(rectangle2_widths[1396]), .rectangle2_height(rectangle2_heights[1396]), .rectangle2_weight(rectangle2_weights[1396]), .rectangle3_x(rectangle3_xs[1396]), .rectangle3_y(rectangle3_ys[1396]), .rectangle3_width(rectangle3_widths[1396]), .rectangle3_height(rectangle3_heights[1396]), .rectangle3_weight(rectangle3_weights[1396]), .feature_threshold(feature_thresholds[1396]), .feature_above(feature_aboves[1396]), .feature_below(feature_belows[1396]), .scan_win_std_dev(scan_win_std_dev[1396]), .feature_accum(feature_accums[1396]));
  accum_calculator ac1397(.scan_win(scan_win1397), .rectangle1_x(rectangle1_xs[1397]), .rectangle1_y(rectangle1_ys[1397]), .rectangle1_width(rectangle1_widths[1397]), .rectangle1_height(rectangle1_heights[1397]), .rectangle1_weight(rectangle1_weights[1397]), .rectangle2_x(rectangle2_xs[1397]), .rectangle2_y(rectangle2_ys[1397]), .rectangle2_width(rectangle2_widths[1397]), .rectangle2_height(rectangle2_heights[1397]), .rectangle2_weight(rectangle2_weights[1397]), .rectangle3_x(rectangle3_xs[1397]), .rectangle3_y(rectangle3_ys[1397]), .rectangle3_width(rectangle3_widths[1397]), .rectangle3_height(rectangle3_heights[1397]), .rectangle3_weight(rectangle3_weights[1397]), .feature_threshold(feature_thresholds[1397]), .feature_above(feature_aboves[1397]), .feature_below(feature_belows[1397]), .scan_win_std_dev(scan_win_std_dev[1397]), .feature_accum(feature_accums[1397]));
  accum_calculator ac1398(.scan_win(scan_win1398), .rectangle1_x(rectangle1_xs[1398]), .rectangle1_y(rectangle1_ys[1398]), .rectangle1_width(rectangle1_widths[1398]), .rectangle1_height(rectangle1_heights[1398]), .rectangle1_weight(rectangle1_weights[1398]), .rectangle2_x(rectangle2_xs[1398]), .rectangle2_y(rectangle2_ys[1398]), .rectangle2_width(rectangle2_widths[1398]), .rectangle2_height(rectangle2_heights[1398]), .rectangle2_weight(rectangle2_weights[1398]), .rectangle3_x(rectangle3_xs[1398]), .rectangle3_y(rectangle3_ys[1398]), .rectangle3_width(rectangle3_widths[1398]), .rectangle3_height(rectangle3_heights[1398]), .rectangle3_weight(rectangle3_weights[1398]), .feature_threshold(feature_thresholds[1398]), .feature_above(feature_aboves[1398]), .feature_below(feature_belows[1398]), .scan_win_std_dev(scan_win_std_dev[1398]), .feature_accum(feature_accums[1398]));
  accum_calculator ac1399(.scan_win(scan_win1399), .rectangle1_x(rectangle1_xs[1399]), .rectangle1_y(rectangle1_ys[1399]), .rectangle1_width(rectangle1_widths[1399]), .rectangle1_height(rectangle1_heights[1399]), .rectangle1_weight(rectangle1_weights[1399]), .rectangle2_x(rectangle2_xs[1399]), .rectangle2_y(rectangle2_ys[1399]), .rectangle2_width(rectangle2_widths[1399]), .rectangle2_height(rectangle2_heights[1399]), .rectangle2_weight(rectangle2_weights[1399]), .rectangle3_x(rectangle3_xs[1399]), .rectangle3_y(rectangle3_ys[1399]), .rectangle3_width(rectangle3_widths[1399]), .rectangle3_height(rectangle3_heights[1399]), .rectangle3_weight(rectangle3_weights[1399]), .feature_threshold(feature_thresholds[1399]), .feature_above(feature_aboves[1399]), .feature_below(feature_belows[1399]), .scan_win_std_dev(scan_win_std_dev[1399]), .feature_accum(feature_accums[1399]));
  accum_calculator ac1400(.scan_win(scan_win1400), .rectangle1_x(rectangle1_xs[1400]), .rectangle1_y(rectangle1_ys[1400]), .rectangle1_width(rectangle1_widths[1400]), .rectangle1_height(rectangle1_heights[1400]), .rectangle1_weight(rectangle1_weights[1400]), .rectangle2_x(rectangle2_xs[1400]), .rectangle2_y(rectangle2_ys[1400]), .rectangle2_width(rectangle2_widths[1400]), .rectangle2_height(rectangle2_heights[1400]), .rectangle2_weight(rectangle2_weights[1400]), .rectangle3_x(rectangle3_xs[1400]), .rectangle3_y(rectangle3_ys[1400]), .rectangle3_width(rectangle3_widths[1400]), .rectangle3_height(rectangle3_heights[1400]), .rectangle3_weight(rectangle3_weights[1400]), .feature_threshold(feature_thresholds[1400]), .feature_above(feature_aboves[1400]), .feature_below(feature_belows[1400]), .scan_win_std_dev(scan_win_std_dev[1400]), .feature_accum(feature_accums[1400]));
  accum_calculator ac1401(.scan_win(scan_win1401), .rectangle1_x(rectangle1_xs[1401]), .rectangle1_y(rectangle1_ys[1401]), .rectangle1_width(rectangle1_widths[1401]), .rectangle1_height(rectangle1_heights[1401]), .rectangle1_weight(rectangle1_weights[1401]), .rectangle2_x(rectangle2_xs[1401]), .rectangle2_y(rectangle2_ys[1401]), .rectangle2_width(rectangle2_widths[1401]), .rectangle2_height(rectangle2_heights[1401]), .rectangle2_weight(rectangle2_weights[1401]), .rectangle3_x(rectangle3_xs[1401]), .rectangle3_y(rectangle3_ys[1401]), .rectangle3_width(rectangle3_widths[1401]), .rectangle3_height(rectangle3_heights[1401]), .rectangle3_weight(rectangle3_weights[1401]), .feature_threshold(feature_thresholds[1401]), .feature_above(feature_aboves[1401]), .feature_below(feature_belows[1401]), .scan_win_std_dev(scan_win_std_dev[1401]), .feature_accum(feature_accums[1401]));
  accum_calculator ac1402(.scan_win(scan_win1402), .rectangle1_x(rectangle1_xs[1402]), .rectangle1_y(rectangle1_ys[1402]), .rectangle1_width(rectangle1_widths[1402]), .rectangle1_height(rectangle1_heights[1402]), .rectangle1_weight(rectangle1_weights[1402]), .rectangle2_x(rectangle2_xs[1402]), .rectangle2_y(rectangle2_ys[1402]), .rectangle2_width(rectangle2_widths[1402]), .rectangle2_height(rectangle2_heights[1402]), .rectangle2_weight(rectangle2_weights[1402]), .rectangle3_x(rectangle3_xs[1402]), .rectangle3_y(rectangle3_ys[1402]), .rectangle3_width(rectangle3_widths[1402]), .rectangle3_height(rectangle3_heights[1402]), .rectangle3_weight(rectangle3_weights[1402]), .feature_threshold(feature_thresholds[1402]), .feature_above(feature_aboves[1402]), .feature_below(feature_belows[1402]), .scan_win_std_dev(scan_win_std_dev[1402]), .feature_accum(feature_accums[1402]));
  accum_calculator ac1403(.scan_win(scan_win1403), .rectangle1_x(rectangle1_xs[1403]), .rectangle1_y(rectangle1_ys[1403]), .rectangle1_width(rectangle1_widths[1403]), .rectangle1_height(rectangle1_heights[1403]), .rectangle1_weight(rectangle1_weights[1403]), .rectangle2_x(rectangle2_xs[1403]), .rectangle2_y(rectangle2_ys[1403]), .rectangle2_width(rectangle2_widths[1403]), .rectangle2_height(rectangle2_heights[1403]), .rectangle2_weight(rectangle2_weights[1403]), .rectangle3_x(rectangle3_xs[1403]), .rectangle3_y(rectangle3_ys[1403]), .rectangle3_width(rectangle3_widths[1403]), .rectangle3_height(rectangle3_heights[1403]), .rectangle3_weight(rectangle3_weights[1403]), .feature_threshold(feature_thresholds[1403]), .feature_above(feature_aboves[1403]), .feature_below(feature_belows[1403]), .scan_win_std_dev(scan_win_std_dev[1403]), .feature_accum(feature_accums[1403]));
  accum_calculator ac1404(.scan_win(scan_win1404), .rectangle1_x(rectangle1_xs[1404]), .rectangle1_y(rectangle1_ys[1404]), .rectangle1_width(rectangle1_widths[1404]), .rectangle1_height(rectangle1_heights[1404]), .rectangle1_weight(rectangle1_weights[1404]), .rectangle2_x(rectangle2_xs[1404]), .rectangle2_y(rectangle2_ys[1404]), .rectangle2_width(rectangle2_widths[1404]), .rectangle2_height(rectangle2_heights[1404]), .rectangle2_weight(rectangle2_weights[1404]), .rectangle3_x(rectangle3_xs[1404]), .rectangle3_y(rectangle3_ys[1404]), .rectangle3_width(rectangle3_widths[1404]), .rectangle3_height(rectangle3_heights[1404]), .rectangle3_weight(rectangle3_weights[1404]), .feature_threshold(feature_thresholds[1404]), .feature_above(feature_aboves[1404]), .feature_below(feature_belows[1404]), .scan_win_std_dev(scan_win_std_dev[1404]), .feature_accum(feature_accums[1404]));
  accum_calculator ac1405(.scan_win(scan_win1405), .rectangle1_x(rectangle1_xs[1405]), .rectangle1_y(rectangle1_ys[1405]), .rectangle1_width(rectangle1_widths[1405]), .rectangle1_height(rectangle1_heights[1405]), .rectangle1_weight(rectangle1_weights[1405]), .rectangle2_x(rectangle2_xs[1405]), .rectangle2_y(rectangle2_ys[1405]), .rectangle2_width(rectangle2_widths[1405]), .rectangle2_height(rectangle2_heights[1405]), .rectangle2_weight(rectangle2_weights[1405]), .rectangle3_x(rectangle3_xs[1405]), .rectangle3_y(rectangle3_ys[1405]), .rectangle3_width(rectangle3_widths[1405]), .rectangle3_height(rectangle3_heights[1405]), .rectangle3_weight(rectangle3_weights[1405]), .feature_threshold(feature_thresholds[1405]), .feature_above(feature_aboves[1405]), .feature_below(feature_belows[1405]), .scan_win_std_dev(scan_win_std_dev[1405]), .feature_accum(feature_accums[1405]));
  accum_calculator ac1406(.scan_win(scan_win1406), .rectangle1_x(rectangle1_xs[1406]), .rectangle1_y(rectangle1_ys[1406]), .rectangle1_width(rectangle1_widths[1406]), .rectangle1_height(rectangle1_heights[1406]), .rectangle1_weight(rectangle1_weights[1406]), .rectangle2_x(rectangle2_xs[1406]), .rectangle2_y(rectangle2_ys[1406]), .rectangle2_width(rectangle2_widths[1406]), .rectangle2_height(rectangle2_heights[1406]), .rectangle2_weight(rectangle2_weights[1406]), .rectangle3_x(rectangle3_xs[1406]), .rectangle3_y(rectangle3_ys[1406]), .rectangle3_width(rectangle3_widths[1406]), .rectangle3_height(rectangle3_heights[1406]), .rectangle3_weight(rectangle3_weights[1406]), .feature_threshold(feature_thresholds[1406]), .feature_above(feature_aboves[1406]), .feature_below(feature_belows[1406]), .scan_win_std_dev(scan_win_std_dev[1406]), .feature_accum(feature_accums[1406]));
  accum_calculator ac1407(.scan_win(scan_win1407), .rectangle1_x(rectangle1_xs[1407]), .rectangle1_y(rectangle1_ys[1407]), .rectangle1_width(rectangle1_widths[1407]), .rectangle1_height(rectangle1_heights[1407]), .rectangle1_weight(rectangle1_weights[1407]), .rectangle2_x(rectangle2_xs[1407]), .rectangle2_y(rectangle2_ys[1407]), .rectangle2_width(rectangle2_widths[1407]), .rectangle2_height(rectangle2_heights[1407]), .rectangle2_weight(rectangle2_weights[1407]), .rectangle3_x(rectangle3_xs[1407]), .rectangle3_y(rectangle3_ys[1407]), .rectangle3_width(rectangle3_widths[1407]), .rectangle3_height(rectangle3_heights[1407]), .rectangle3_weight(rectangle3_weights[1407]), .feature_threshold(feature_thresholds[1407]), .feature_above(feature_aboves[1407]), .feature_below(feature_belows[1407]), .scan_win_std_dev(scan_win_std_dev[1407]), .feature_accum(feature_accums[1407]));
  accum_calculator ac1408(.scan_win(scan_win1408), .rectangle1_x(rectangle1_xs[1408]), .rectangle1_y(rectangle1_ys[1408]), .rectangle1_width(rectangle1_widths[1408]), .rectangle1_height(rectangle1_heights[1408]), .rectangle1_weight(rectangle1_weights[1408]), .rectangle2_x(rectangle2_xs[1408]), .rectangle2_y(rectangle2_ys[1408]), .rectangle2_width(rectangle2_widths[1408]), .rectangle2_height(rectangle2_heights[1408]), .rectangle2_weight(rectangle2_weights[1408]), .rectangle3_x(rectangle3_xs[1408]), .rectangle3_y(rectangle3_ys[1408]), .rectangle3_width(rectangle3_widths[1408]), .rectangle3_height(rectangle3_heights[1408]), .rectangle3_weight(rectangle3_weights[1408]), .feature_threshold(feature_thresholds[1408]), .feature_above(feature_aboves[1408]), .feature_below(feature_belows[1408]), .scan_win_std_dev(scan_win_std_dev[1408]), .feature_accum(feature_accums[1408]));
  accum_calculator ac1409(.scan_win(scan_win1409), .rectangle1_x(rectangle1_xs[1409]), .rectangle1_y(rectangle1_ys[1409]), .rectangle1_width(rectangle1_widths[1409]), .rectangle1_height(rectangle1_heights[1409]), .rectangle1_weight(rectangle1_weights[1409]), .rectangle2_x(rectangle2_xs[1409]), .rectangle2_y(rectangle2_ys[1409]), .rectangle2_width(rectangle2_widths[1409]), .rectangle2_height(rectangle2_heights[1409]), .rectangle2_weight(rectangle2_weights[1409]), .rectangle3_x(rectangle3_xs[1409]), .rectangle3_y(rectangle3_ys[1409]), .rectangle3_width(rectangle3_widths[1409]), .rectangle3_height(rectangle3_heights[1409]), .rectangle3_weight(rectangle3_weights[1409]), .feature_threshold(feature_thresholds[1409]), .feature_above(feature_aboves[1409]), .feature_below(feature_belows[1409]), .scan_win_std_dev(scan_win_std_dev[1409]), .feature_accum(feature_accums[1409]));
  accum_calculator ac1410(.scan_win(scan_win1410), .rectangle1_x(rectangle1_xs[1410]), .rectangle1_y(rectangle1_ys[1410]), .rectangle1_width(rectangle1_widths[1410]), .rectangle1_height(rectangle1_heights[1410]), .rectangle1_weight(rectangle1_weights[1410]), .rectangle2_x(rectangle2_xs[1410]), .rectangle2_y(rectangle2_ys[1410]), .rectangle2_width(rectangle2_widths[1410]), .rectangle2_height(rectangle2_heights[1410]), .rectangle2_weight(rectangle2_weights[1410]), .rectangle3_x(rectangle3_xs[1410]), .rectangle3_y(rectangle3_ys[1410]), .rectangle3_width(rectangle3_widths[1410]), .rectangle3_height(rectangle3_heights[1410]), .rectangle3_weight(rectangle3_weights[1410]), .feature_threshold(feature_thresholds[1410]), .feature_above(feature_aboves[1410]), .feature_below(feature_belows[1410]), .scan_win_std_dev(scan_win_std_dev[1410]), .feature_accum(feature_accums[1410]));
  accum_calculator ac1411(.scan_win(scan_win1411), .rectangle1_x(rectangle1_xs[1411]), .rectangle1_y(rectangle1_ys[1411]), .rectangle1_width(rectangle1_widths[1411]), .rectangle1_height(rectangle1_heights[1411]), .rectangle1_weight(rectangle1_weights[1411]), .rectangle2_x(rectangle2_xs[1411]), .rectangle2_y(rectangle2_ys[1411]), .rectangle2_width(rectangle2_widths[1411]), .rectangle2_height(rectangle2_heights[1411]), .rectangle2_weight(rectangle2_weights[1411]), .rectangle3_x(rectangle3_xs[1411]), .rectangle3_y(rectangle3_ys[1411]), .rectangle3_width(rectangle3_widths[1411]), .rectangle3_height(rectangle3_heights[1411]), .rectangle3_weight(rectangle3_weights[1411]), .feature_threshold(feature_thresholds[1411]), .feature_above(feature_aboves[1411]), .feature_below(feature_belows[1411]), .scan_win_std_dev(scan_win_std_dev[1411]), .feature_accum(feature_accums[1411]));
  accum_calculator ac1412(.scan_win(scan_win1412), .rectangle1_x(rectangle1_xs[1412]), .rectangle1_y(rectangle1_ys[1412]), .rectangle1_width(rectangle1_widths[1412]), .rectangle1_height(rectangle1_heights[1412]), .rectangle1_weight(rectangle1_weights[1412]), .rectangle2_x(rectangle2_xs[1412]), .rectangle2_y(rectangle2_ys[1412]), .rectangle2_width(rectangle2_widths[1412]), .rectangle2_height(rectangle2_heights[1412]), .rectangle2_weight(rectangle2_weights[1412]), .rectangle3_x(rectangle3_xs[1412]), .rectangle3_y(rectangle3_ys[1412]), .rectangle3_width(rectangle3_widths[1412]), .rectangle3_height(rectangle3_heights[1412]), .rectangle3_weight(rectangle3_weights[1412]), .feature_threshold(feature_thresholds[1412]), .feature_above(feature_aboves[1412]), .feature_below(feature_belows[1412]), .scan_win_std_dev(scan_win_std_dev[1412]), .feature_accum(feature_accums[1412]));
  accum_calculator ac1413(.scan_win(scan_win1413), .rectangle1_x(rectangle1_xs[1413]), .rectangle1_y(rectangle1_ys[1413]), .rectangle1_width(rectangle1_widths[1413]), .rectangle1_height(rectangle1_heights[1413]), .rectangle1_weight(rectangle1_weights[1413]), .rectangle2_x(rectangle2_xs[1413]), .rectangle2_y(rectangle2_ys[1413]), .rectangle2_width(rectangle2_widths[1413]), .rectangle2_height(rectangle2_heights[1413]), .rectangle2_weight(rectangle2_weights[1413]), .rectangle3_x(rectangle3_xs[1413]), .rectangle3_y(rectangle3_ys[1413]), .rectangle3_width(rectangle3_widths[1413]), .rectangle3_height(rectangle3_heights[1413]), .rectangle3_weight(rectangle3_weights[1413]), .feature_threshold(feature_thresholds[1413]), .feature_above(feature_aboves[1413]), .feature_below(feature_belows[1413]), .scan_win_std_dev(scan_win_std_dev[1413]), .feature_accum(feature_accums[1413]));
  accum_calculator ac1414(.scan_win(scan_win1414), .rectangle1_x(rectangle1_xs[1414]), .rectangle1_y(rectangle1_ys[1414]), .rectangle1_width(rectangle1_widths[1414]), .rectangle1_height(rectangle1_heights[1414]), .rectangle1_weight(rectangle1_weights[1414]), .rectangle2_x(rectangle2_xs[1414]), .rectangle2_y(rectangle2_ys[1414]), .rectangle2_width(rectangle2_widths[1414]), .rectangle2_height(rectangle2_heights[1414]), .rectangle2_weight(rectangle2_weights[1414]), .rectangle3_x(rectangle3_xs[1414]), .rectangle3_y(rectangle3_ys[1414]), .rectangle3_width(rectangle3_widths[1414]), .rectangle3_height(rectangle3_heights[1414]), .rectangle3_weight(rectangle3_weights[1414]), .feature_threshold(feature_thresholds[1414]), .feature_above(feature_aboves[1414]), .feature_below(feature_belows[1414]), .scan_win_std_dev(scan_win_std_dev[1414]), .feature_accum(feature_accums[1414]));
  accum_calculator ac1415(.scan_win(scan_win1415), .rectangle1_x(rectangle1_xs[1415]), .rectangle1_y(rectangle1_ys[1415]), .rectangle1_width(rectangle1_widths[1415]), .rectangle1_height(rectangle1_heights[1415]), .rectangle1_weight(rectangle1_weights[1415]), .rectangle2_x(rectangle2_xs[1415]), .rectangle2_y(rectangle2_ys[1415]), .rectangle2_width(rectangle2_widths[1415]), .rectangle2_height(rectangle2_heights[1415]), .rectangle2_weight(rectangle2_weights[1415]), .rectangle3_x(rectangle3_xs[1415]), .rectangle3_y(rectangle3_ys[1415]), .rectangle3_width(rectangle3_widths[1415]), .rectangle3_height(rectangle3_heights[1415]), .rectangle3_weight(rectangle3_weights[1415]), .feature_threshold(feature_thresholds[1415]), .feature_above(feature_aboves[1415]), .feature_below(feature_belows[1415]), .scan_win_std_dev(scan_win_std_dev[1415]), .feature_accum(feature_accums[1415]));
  accum_calculator ac1416(.scan_win(scan_win1416), .rectangle1_x(rectangle1_xs[1416]), .rectangle1_y(rectangle1_ys[1416]), .rectangle1_width(rectangle1_widths[1416]), .rectangle1_height(rectangle1_heights[1416]), .rectangle1_weight(rectangle1_weights[1416]), .rectangle2_x(rectangle2_xs[1416]), .rectangle2_y(rectangle2_ys[1416]), .rectangle2_width(rectangle2_widths[1416]), .rectangle2_height(rectangle2_heights[1416]), .rectangle2_weight(rectangle2_weights[1416]), .rectangle3_x(rectangle3_xs[1416]), .rectangle3_y(rectangle3_ys[1416]), .rectangle3_width(rectangle3_widths[1416]), .rectangle3_height(rectangle3_heights[1416]), .rectangle3_weight(rectangle3_weights[1416]), .feature_threshold(feature_thresholds[1416]), .feature_above(feature_aboves[1416]), .feature_below(feature_belows[1416]), .scan_win_std_dev(scan_win_std_dev[1416]), .feature_accum(feature_accums[1416]));
  accum_calculator ac1417(.scan_win(scan_win1417), .rectangle1_x(rectangle1_xs[1417]), .rectangle1_y(rectangle1_ys[1417]), .rectangle1_width(rectangle1_widths[1417]), .rectangle1_height(rectangle1_heights[1417]), .rectangle1_weight(rectangle1_weights[1417]), .rectangle2_x(rectangle2_xs[1417]), .rectangle2_y(rectangle2_ys[1417]), .rectangle2_width(rectangle2_widths[1417]), .rectangle2_height(rectangle2_heights[1417]), .rectangle2_weight(rectangle2_weights[1417]), .rectangle3_x(rectangle3_xs[1417]), .rectangle3_y(rectangle3_ys[1417]), .rectangle3_width(rectangle3_widths[1417]), .rectangle3_height(rectangle3_heights[1417]), .rectangle3_weight(rectangle3_weights[1417]), .feature_threshold(feature_thresholds[1417]), .feature_above(feature_aboves[1417]), .feature_below(feature_belows[1417]), .scan_win_std_dev(scan_win_std_dev[1417]), .feature_accum(feature_accums[1417]));
  accum_calculator ac1418(.scan_win(scan_win1418), .rectangle1_x(rectangle1_xs[1418]), .rectangle1_y(rectangle1_ys[1418]), .rectangle1_width(rectangle1_widths[1418]), .rectangle1_height(rectangle1_heights[1418]), .rectangle1_weight(rectangle1_weights[1418]), .rectangle2_x(rectangle2_xs[1418]), .rectangle2_y(rectangle2_ys[1418]), .rectangle2_width(rectangle2_widths[1418]), .rectangle2_height(rectangle2_heights[1418]), .rectangle2_weight(rectangle2_weights[1418]), .rectangle3_x(rectangle3_xs[1418]), .rectangle3_y(rectangle3_ys[1418]), .rectangle3_width(rectangle3_widths[1418]), .rectangle3_height(rectangle3_heights[1418]), .rectangle3_weight(rectangle3_weights[1418]), .feature_threshold(feature_thresholds[1418]), .feature_above(feature_aboves[1418]), .feature_below(feature_belows[1418]), .scan_win_std_dev(scan_win_std_dev[1418]), .feature_accum(feature_accums[1418]));
  accum_calculator ac1419(.scan_win(scan_win1419), .rectangle1_x(rectangle1_xs[1419]), .rectangle1_y(rectangle1_ys[1419]), .rectangle1_width(rectangle1_widths[1419]), .rectangle1_height(rectangle1_heights[1419]), .rectangle1_weight(rectangle1_weights[1419]), .rectangle2_x(rectangle2_xs[1419]), .rectangle2_y(rectangle2_ys[1419]), .rectangle2_width(rectangle2_widths[1419]), .rectangle2_height(rectangle2_heights[1419]), .rectangle2_weight(rectangle2_weights[1419]), .rectangle3_x(rectangle3_xs[1419]), .rectangle3_y(rectangle3_ys[1419]), .rectangle3_width(rectangle3_widths[1419]), .rectangle3_height(rectangle3_heights[1419]), .rectangle3_weight(rectangle3_weights[1419]), .feature_threshold(feature_thresholds[1419]), .feature_above(feature_aboves[1419]), .feature_below(feature_belows[1419]), .scan_win_std_dev(scan_win_std_dev[1419]), .feature_accum(feature_accums[1419]));
  accum_calculator ac1420(.scan_win(scan_win1420), .rectangle1_x(rectangle1_xs[1420]), .rectangle1_y(rectangle1_ys[1420]), .rectangle1_width(rectangle1_widths[1420]), .rectangle1_height(rectangle1_heights[1420]), .rectangle1_weight(rectangle1_weights[1420]), .rectangle2_x(rectangle2_xs[1420]), .rectangle2_y(rectangle2_ys[1420]), .rectangle2_width(rectangle2_widths[1420]), .rectangle2_height(rectangle2_heights[1420]), .rectangle2_weight(rectangle2_weights[1420]), .rectangle3_x(rectangle3_xs[1420]), .rectangle3_y(rectangle3_ys[1420]), .rectangle3_width(rectangle3_widths[1420]), .rectangle3_height(rectangle3_heights[1420]), .rectangle3_weight(rectangle3_weights[1420]), .feature_threshold(feature_thresholds[1420]), .feature_above(feature_aboves[1420]), .feature_below(feature_belows[1420]), .scan_win_std_dev(scan_win_std_dev[1420]), .feature_accum(feature_accums[1420]));
  accum_calculator ac1421(.scan_win(scan_win1421), .rectangle1_x(rectangle1_xs[1421]), .rectangle1_y(rectangle1_ys[1421]), .rectangle1_width(rectangle1_widths[1421]), .rectangle1_height(rectangle1_heights[1421]), .rectangle1_weight(rectangle1_weights[1421]), .rectangle2_x(rectangle2_xs[1421]), .rectangle2_y(rectangle2_ys[1421]), .rectangle2_width(rectangle2_widths[1421]), .rectangle2_height(rectangle2_heights[1421]), .rectangle2_weight(rectangle2_weights[1421]), .rectangle3_x(rectangle3_xs[1421]), .rectangle3_y(rectangle3_ys[1421]), .rectangle3_width(rectangle3_widths[1421]), .rectangle3_height(rectangle3_heights[1421]), .rectangle3_weight(rectangle3_weights[1421]), .feature_threshold(feature_thresholds[1421]), .feature_above(feature_aboves[1421]), .feature_below(feature_belows[1421]), .scan_win_std_dev(scan_win_std_dev[1421]), .feature_accum(feature_accums[1421]));
  accum_calculator ac1422(.scan_win(scan_win1422), .rectangle1_x(rectangle1_xs[1422]), .rectangle1_y(rectangle1_ys[1422]), .rectangle1_width(rectangle1_widths[1422]), .rectangle1_height(rectangle1_heights[1422]), .rectangle1_weight(rectangle1_weights[1422]), .rectangle2_x(rectangle2_xs[1422]), .rectangle2_y(rectangle2_ys[1422]), .rectangle2_width(rectangle2_widths[1422]), .rectangle2_height(rectangle2_heights[1422]), .rectangle2_weight(rectangle2_weights[1422]), .rectangle3_x(rectangle3_xs[1422]), .rectangle3_y(rectangle3_ys[1422]), .rectangle3_width(rectangle3_widths[1422]), .rectangle3_height(rectangle3_heights[1422]), .rectangle3_weight(rectangle3_weights[1422]), .feature_threshold(feature_thresholds[1422]), .feature_above(feature_aboves[1422]), .feature_below(feature_belows[1422]), .scan_win_std_dev(scan_win_std_dev[1422]), .feature_accum(feature_accums[1422]));
  accum_calculator ac1423(.scan_win(scan_win1423), .rectangle1_x(rectangle1_xs[1423]), .rectangle1_y(rectangle1_ys[1423]), .rectangle1_width(rectangle1_widths[1423]), .rectangle1_height(rectangle1_heights[1423]), .rectangle1_weight(rectangle1_weights[1423]), .rectangle2_x(rectangle2_xs[1423]), .rectangle2_y(rectangle2_ys[1423]), .rectangle2_width(rectangle2_widths[1423]), .rectangle2_height(rectangle2_heights[1423]), .rectangle2_weight(rectangle2_weights[1423]), .rectangle3_x(rectangle3_xs[1423]), .rectangle3_y(rectangle3_ys[1423]), .rectangle3_width(rectangle3_widths[1423]), .rectangle3_height(rectangle3_heights[1423]), .rectangle3_weight(rectangle3_weights[1423]), .feature_threshold(feature_thresholds[1423]), .feature_above(feature_aboves[1423]), .feature_below(feature_belows[1423]), .scan_win_std_dev(scan_win_std_dev[1423]), .feature_accum(feature_accums[1423]));
  accum_calculator ac1424(.scan_win(scan_win1424), .rectangle1_x(rectangle1_xs[1424]), .rectangle1_y(rectangle1_ys[1424]), .rectangle1_width(rectangle1_widths[1424]), .rectangle1_height(rectangle1_heights[1424]), .rectangle1_weight(rectangle1_weights[1424]), .rectangle2_x(rectangle2_xs[1424]), .rectangle2_y(rectangle2_ys[1424]), .rectangle2_width(rectangle2_widths[1424]), .rectangle2_height(rectangle2_heights[1424]), .rectangle2_weight(rectangle2_weights[1424]), .rectangle3_x(rectangle3_xs[1424]), .rectangle3_y(rectangle3_ys[1424]), .rectangle3_width(rectangle3_widths[1424]), .rectangle3_height(rectangle3_heights[1424]), .rectangle3_weight(rectangle3_weights[1424]), .feature_threshold(feature_thresholds[1424]), .feature_above(feature_aboves[1424]), .feature_below(feature_belows[1424]), .scan_win_std_dev(scan_win_std_dev[1424]), .feature_accum(feature_accums[1424]));
  accum_calculator ac1425(.scan_win(scan_win1425), .rectangle1_x(rectangle1_xs[1425]), .rectangle1_y(rectangle1_ys[1425]), .rectangle1_width(rectangle1_widths[1425]), .rectangle1_height(rectangle1_heights[1425]), .rectangle1_weight(rectangle1_weights[1425]), .rectangle2_x(rectangle2_xs[1425]), .rectangle2_y(rectangle2_ys[1425]), .rectangle2_width(rectangle2_widths[1425]), .rectangle2_height(rectangle2_heights[1425]), .rectangle2_weight(rectangle2_weights[1425]), .rectangle3_x(rectangle3_xs[1425]), .rectangle3_y(rectangle3_ys[1425]), .rectangle3_width(rectangle3_widths[1425]), .rectangle3_height(rectangle3_heights[1425]), .rectangle3_weight(rectangle3_weights[1425]), .feature_threshold(feature_thresholds[1425]), .feature_above(feature_aboves[1425]), .feature_below(feature_belows[1425]), .scan_win_std_dev(scan_win_std_dev[1425]), .feature_accum(feature_accums[1425]));
  accum_calculator ac1426(.scan_win(scan_win1426), .rectangle1_x(rectangle1_xs[1426]), .rectangle1_y(rectangle1_ys[1426]), .rectangle1_width(rectangle1_widths[1426]), .rectangle1_height(rectangle1_heights[1426]), .rectangle1_weight(rectangle1_weights[1426]), .rectangle2_x(rectangle2_xs[1426]), .rectangle2_y(rectangle2_ys[1426]), .rectangle2_width(rectangle2_widths[1426]), .rectangle2_height(rectangle2_heights[1426]), .rectangle2_weight(rectangle2_weights[1426]), .rectangle3_x(rectangle3_xs[1426]), .rectangle3_y(rectangle3_ys[1426]), .rectangle3_width(rectangle3_widths[1426]), .rectangle3_height(rectangle3_heights[1426]), .rectangle3_weight(rectangle3_weights[1426]), .feature_threshold(feature_thresholds[1426]), .feature_above(feature_aboves[1426]), .feature_below(feature_belows[1426]), .scan_win_std_dev(scan_win_std_dev[1426]), .feature_accum(feature_accums[1426]));
  accum_calculator ac1427(.scan_win(scan_win1427), .rectangle1_x(rectangle1_xs[1427]), .rectangle1_y(rectangle1_ys[1427]), .rectangle1_width(rectangle1_widths[1427]), .rectangle1_height(rectangle1_heights[1427]), .rectangle1_weight(rectangle1_weights[1427]), .rectangle2_x(rectangle2_xs[1427]), .rectangle2_y(rectangle2_ys[1427]), .rectangle2_width(rectangle2_widths[1427]), .rectangle2_height(rectangle2_heights[1427]), .rectangle2_weight(rectangle2_weights[1427]), .rectangle3_x(rectangle3_xs[1427]), .rectangle3_y(rectangle3_ys[1427]), .rectangle3_width(rectangle3_widths[1427]), .rectangle3_height(rectangle3_heights[1427]), .rectangle3_weight(rectangle3_weights[1427]), .feature_threshold(feature_thresholds[1427]), .feature_above(feature_aboves[1427]), .feature_below(feature_belows[1427]), .scan_win_std_dev(scan_win_std_dev[1427]), .feature_accum(feature_accums[1427]));
  accum_calculator ac1428(.scan_win(scan_win1428), .rectangle1_x(rectangle1_xs[1428]), .rectangle1_y(rectangle1_ys[1428]), .rectangle1_width(rectangle1_widths[1428]), .rectangle1_height(rectangle1_heights[1428]), .rectangle1_weight(rectangle1_weights[1428]), .rectangle2_x(rectangle2_xs[1428]), .rectangle2_y(rectangle2_ys[1428]), .rectangle2_width(rectangle2_widths[1428]), .rectangle2_height(rectangle2_heights[1428]), .rectangle2_weight(rectangle2_weights[1428]), .rectangle3_x(rectangle3_xs[1428]), .rectangle3_y(rectangle3_ys[1428]), .rectangle3_width(rectangle3_widths[1428]), .rectangle3_height(rectangle3_heights[1428]), .rectangle3_weight(rectangle3_weights[1428]), .feature_threshold(feature_thresholds[1428]), .feature_above(feature_aboves[1428]), .feature_below(feature_belows[1428]), .scan_win_std_dev(scan_win_std_dev[1428]), .feature_accum(feature_accums[1428]));
  accum_calculator ac1429(.scan_win(scan_win1429), .rectangle1_x(rectangle1_xs[1429]), .rectangle1_y(rectangle1_ys[1429]), .rectangle1_width(rectangle1_widths[1429]), .rectangle1_height(rectangle1_heights[1429]), .rectangle1_weight(rectangle1_weights[1429]), .rectangle2_x(rectangle2_xs[1429]), .rectangle2_y(rectangle2_ys[1429]), .rectangle2_width(rectangle2_widths[1429]), .rectangle2_height(rectangle2_heights[1429]), .rectangle2_weight(rectangle2_weights[1429]), .rectangle3_x(rectangle3_xs[1429]), .rectangle3_y(rectangle3_ys[1429]), .rectangle3_width(rectangle3_widths[1429]), .rectangle3_height(rectangle3_heights[1429]), .rectangle3_weight(rectangle3_weights[1429]), .feature_threshold(feature_thresholds[1429]), .feature_above(feature_aboves[1429]), .feature_below(feature_belows[1429]), .scan_win_std_dev(scan_win_std_dev[1429]), .feature_accum(feature_accums[1429]));
  accum_calculator ac1430(.scan_win(scan_win1430), .rectangle1_x(rectangle1_xs[1430]), .rectangle1_y(rectangle1_ys[1430]), .rectangle1_width(rectangle1_widths[1430]), .rectangle1_height(rectangle1_heights[1430]), .rectangle1_weight(rectangle1_weights[1430]), .rectangle2_x(rectangle2_xs[1430]), .rectangle2_y(rectangle2_ys[1430]), .rectangle2_width(rectangle2_widths[1430]), .rectangle2_height(rectangle2_heights[1430]), .rectangle2_weight(rectangle2_weights[1430]), .rectangle3_x(rectangle3_xs[1430]), .rectangle3_y(rectangle3_ys[1430]), .rectangle3_width(rectangle3_widths[1430]), .rectangle3_height(rectangle3_heights[1430]), .rectangle3_weight(rectangle3_weights[1430]), .feature_threshold(feature_thresholds[1430]), .feature_above(feature_aboves[1430]), .feature_below(feature_belows[1430]), .scan_win_std_dev(scan_win_std_dev[1430]), .feature_accum(feature_accums[1430]));
  accum_calculator ac1431(.scan_win(scan_win1431), .rectangle1_x(rectangle1_xs[1431]), .rectangle1_y(rectangle1_ys[1431]), .rectangle1_width(rectangle1_widths[1431]), .rectangle1_height(rectangle1_heights[1431]), .rectangle1_weight(rectangle1_weights[1431]), .rectangle2_x(rectangle2_xs[1431]), .rectangle2_y(rectangle2_ys[1431]), .rectangle2_width(rectangle2_widths[1431]), .rectangle2_height(rectangle2_heights[1431]), .rectangle2_weight(rectangle2_weights[1431]), .rectangle3_x(rectangle3_xs[1431]), .rectangle3_y(rectangle3_ys[1431]), .rectangle3_width(rectangle3_widths[1431]), .rectangle3_height(rectangle3_heights[1431]), .rectangle3_weight(rectangle3_weights[1431]), .feature_threshold(feature_thresholds[1431]), .feature_above(feature_aboves[1431]), .feature_below(feature_belows[1431]), .scan_win_std_dev(scan_win_std_dev[1431]), .feature_accum(feature_accums[1431]));
  accum_calculator ac1432(.scan_win(scan_win1432), .rectangle1_x(rectangle1_xs[1432]), .rectangle1_y(rectangle1_ys[1432]), .rectangle1_width(rectangle1_widths[1432]), .rectangle1_height(rectangle1_heights[1432]), .rectangle1_weight(rectangle1_weights[1432]), .rectangle2_x(rectangle2_xs[1432]), .rectangle2_y(rectangle2_ys[1432]), .rectangle2_width(rectangle2_widths[1432]), .rectangle2_height(rectangle2_heights[1432]), .rectangle2_weight(rectangle2_weights[1432]), .rectangle3_x(rectangle3_xs[1432]), .rectangle3_y(rectangle3_ys[1432]), .rectangle3_width(rectangle3_widths[1432]), .rectangle3_height(rectangle3_heights[1432]), .rectangle3_weight(rectangle3_weights[1432]), .feature_threshold(feature_thresholds[1432]), .feature_above(feature_aboves[1432]), .feature_below(feature_belows[1432]), .scan_win_std_dev(scan_win_std_dev[1432]), .feature_accum(feature_accums[1432]));
  accum_calculator ac1433(.scan_win(scan_win1433), .rectangle1_x(rectangle1_xs[1433]), .rectangle1_y(rectangle1_ys[1433]), .rectangle1_width(rectangle1_widths[1433]), .rectangle1_height(rectangle1_heights[1433]), .rectangle1_weight(rectangle1_weights[1433]), .rectangle2_x(rectangle2_xs[1433]), .rectangle2_y(rectangle2_ys[1433]), .rectangle2_width(rectangle2_widths[1433]), .rectangle2_height(rectangle2_heights[1433]), .rectangle2_weight(rectangle2_weights[1433]), .rectangle3_x(rectangle3_xs[1433]), .rectangle3_y(rectangle3_ys[1433]), .rectangle3_width(rectangle3_widths[1433]), .rectangle3_height(rectangle3_heights[1433]), .rectangle3_weight(rectangle3_weights[1433]), .feature_threshold(feature_thresholds[1433]), .feature_above(feature_aboves[1433]), .feature_below(feature_belows[1433]), .scan_win_std_dev(scan_win_std_dev[1433]), .feature_accum(feature_accums[1433]));
  accum_calculator ac1434(.scan_win(scan_win1434), .rectangle1_x(rectangle1_xs[1434]), .rectangle1_y(rectangle1_ys[1434]), .rectangle1_width(rectangle1_widths[1434]), .rectangle1_height(rectangle1_heights[1434]), .rectangle1_weight(rectangle1_weights[1434]), .rectangle2_x(rectangle2_xs[1434]), .rectangle2_y(rectangle2_ys[1434]), .rectangle2_width(rectangle2_widths[1434]), .rectangle2_height(rectangle2_heights[1434]), .rectangle2_weight(rectangle2_weights[1434]), .rectangle3_x(rectangle3_xs[1434]), .rectangle3_y(rectangle3_ys[1434]), .rectangle3_width(rectangle3_widths[1434]), .rectangle3_height(rectangle3_heights[1434]), .rectangle3_weight(rectangle3_weights[1434]), .feature_threshold(feature_thresholds[1434]), .feature_above(feature_aboves[1434]), .feature_below(feature_belows[1434]), .scan_win_std_dev(scan_win_std_dev[1434]), .feature_accum(feature_accums[1434]));
  accum_calculator ac1435(.scan_win(scan_win1435), .rectangle1_x(rectangle1_xs[1435]), .rectangle1_y(rectangle1_ys[1435]), .rectangle1_width(rectangle1_widths[1435]), .rectangle1_height(rectangle1_heights[1435]), .rectangle1_weight(rectangle1_weights[1435]), .rectangle2_x(rectangle2_xs[1435]), .rectangle2_y(rectangle2_ys[1435]), .rectangle2_width(rectangle2_widths[1435]), .rectangle2_height(rectangle2_heights[1435]), .rectangle2_weight(rectangle2_weights[1435]), .rectangle3_x(rectangle3_xs[1435]), .rectangle3_y(rectangle3_ys[1435]), .rectangle3_width(rectangle3_widths[1435]), .rectangle3_height(rectangle3_heights[1435]), .rectangle3_weight(rectangle3_weights[1435]), .feature_threshold(feature_thresholds[1435]), .feature_above(feature_aboves[1435]), .feature_below(feature_belows[1435]), .scan_win_std_dev(scan_win_std_dev[1435]), .feature_accum(feature_accums[1435]));
  accum_calculator ac1436(.scan_win(scan_win1436), .rectangle1_x(rectangle1_xs[1436]), .rectangle1_y(rectangle1_ys[1436]), .rectangle1_width(rectangle1_widths[1436]), .rectangle1_height(rectangle1_heights[1436]), .rectangle1_weight(rectangle1_weights[1436]), .rectangle2_x(rectangle2_xs[1436]), .rectangle2_y(rectangle2_ys[1436]), .rectangle2_width(rectangle2_widths[1436]), .rectangle2_height(rectangle2_heights[1436]), .rectangle2_weight(rectangle2_weights[1436]), .rectangle3_x(rectangle3_xs[1436]), .rectangle3_y(rectangle3_ys[1436]), .rectangle3_width(rectangle3_widths[1436]), .rectangle3_height(rectangle3_heights[1436]), .rectangle3_weight(rectangle3_weights[1436]), .feature_threshold(feature_thresholds[1436]), .feature_above(feature_aboves[1436]), .feature_below(feature_belows[1436]), .scan_win_std_dev(scan_win_std_dev[1436]), .feature_accum(feature_accums[1436]));
  accum_calculator ac1437(.scan_win(scan_win1437), .rectangle1_x(rectangle1_xs[1437]), .rectangle1_y(rectangle1_ys[1437]), .rectangle1_width(rectangle1_widths[1437]), .rectangle1_height(rectangle1_heights[1437]), .rectangle1_weight(rectangle1_weights[1437]), .rectangle2_x(rectangle2_xs[1437]), .rectangle2_y(rectangle2_ys[1437]), .rectangle2_width(rectangle2_widths[1437]), .rectangle2_height(rectangle2_heights[1437]), .rectangle2_weight(rectangle2_weights[1437]), .rectangle3_x(rectangle3_xs[1437]), .rectangle3_y(rectangle3_ys[1437]), .rectangle3_width(rectangle3_widths[1437]), .rectangle3_height(rectangle3_heights[1437]), .rectangle3_weight(rectangle3_weights[1437]), .feature_threshold(feature_thresholds[1437]), .feature_above(feature_aboves[1437]), .feature_below(feature_belows[1437]), .scan_win_std_dev(scan_win_std_dev[1437]), .feature_accum(feature_accums[1437]));
  accum_calculator ac1438(.scan_win(scan_win1438), .rectangle1_x(rectangle1_xs[1438]), .rectangle1_y(rectangle1_ys[1438]), .rectangle1_width(rectangle1_widths[1438]), .rectangle1_height(rectangle1_heights[1438]), .rectangle1_weight(rectangle1_weights[1438]), .rectangle2_x(rectangle2_xs[1438]), .rectangle2_y(rectangle2_ys[1438]), .rectangle2_width(rectangle2_widths[1438]), .rectangle2_height(rectangle2_heights[1438]), .rectangle2_weight(rectangle2_weights[1438]), .rectangle3_x(rectangle3_xs[1438]), .rectangle3_y(rectangle3_ys[1438]), .rectangle3_width(rectangle3_widths[1438]), .rectangle3_height(rectangle3_heights[1438]), .rectangle3_weight(rectangle3_weights[1438]), .feature_threshold(feature_thresholds[1438]), .feature_above(feature_aboves[1438]), .feature_below(feature_belows[1438]), .scan_win_std_dev(scan_win_std_dev[1438]), .feature_accum(feature_accums[1438]));
  accum_calculator ac1439(.scan_win(scan_win1439), .rectangle1_x(rectangle1_xs[1439]), .rectangle1_y(rectangle1_ys[1439]), .rectangle1_width(rectangle1_widths[1439]), .rectangle1_height(rectangle1_heights[1439]), .rectangle1_weight(rectangle1_weights[1439]), .rectangle2_x(rectangle2_xs[1439]), .rectangle2_y(rectangle2_ys[1439]), .rectangle2_width(rectangle2_widths[1439]), .rectangle2_height(rectangle2_heights[1439]), .rectangle2_weight(rectangle2_weights[1439]), .rectangle3_x(rectangle3_xs[1439]), .rectangle3_y(rectangle3_ys[1439]), .rectangle3_width(rectangle3_widths[1439]), .rectangle3_height(rectangle3_heights[1439]), .rectangle3_weight(rectangle3_weights[1439]), .feature_threshold(feature_thresholds[1439]), .feature_above(feature_aboves[1439]), .feature_below(feature_belows[1439]), .scan_win_std_dev(scan_win_std_dev[1439]), .feature_accum(feature_accums[1439]));
  accum_calculator ac1440(.scan_win(scan_win1440), .rectangle1_x(rectangle1_xs[1440]), .rectangle1_y(rectangle1_ys[1440]), .rectangle1_width(rectangle1_widths[1440]), .rectangle1_height(rectangle1_heights[1440]), .rectangle1_weight(rectangle1_weights[1440]), .rectangle2_x(rectangle2_xs[1440]), .rectangle2_y(rectangle2_ys[1440]), .rectangle2_width(rectangle2_widths[1440]), .rectangle2_height(rectangle2_heights[1440]), .rectangle2_weight(rectangle2_weights[1440]), .rectangle3_x(rectangle3_xs[1440]), .rectangle3_y(rectangle3_ys[1440]), .rectangle3_width(rectangle3_widths[1440]), .rectangle3_height(rectangle3_heights[1440]), .rectangle3_weight(rectangle3_weights[1440]), .feature_threshold(feature_thresholds[1440]), .feature_above(feature_aboves[1440]), .feature_below(feature_belows[1440]), .scan_win_std_dev(scan_win_std_dev[1440]), .feature_accum(feature_accums[1440]));
  accum_calculator ac1441(.scan_win(scan_win1441), .rectangle1_x(rectangle1_xs[1441]), .rectangle1_y(rectangle1_ys[1441]), .rectangle1_width(rectangle1_widths[1441]), .rectangle1_height(rectangle1_heights[1441]), .rectangle1_weight(rectangle1_weights[1441]), .rectangle2_x(rectangle2_xs[1441]), .rectangle2_y(rectangle2_ys[1441]), .rectangle2_width(rectangle2_widths[1441]), .rectangle2_height(rectangle2_heights[1441]), .rectangle2_weight(rectangle2_weights[1441]), .rectangle3_x(rectangle3_xs[1441]), .rectangle3_y(rectangle3_ys[1441]), .rectangle3_width(rectangle3_widths[1441]), .rectangle3_height(rectangle3_heights[1441]), .rectangle3_weight(rectangle3_weights[1441]), .feature_threshold(feature_thresholds[1441]), .feature_above(feature_aboves[1441]), .feature_below(feature_belows[1441]), .scan_win_std_dev(scan_win_std_dev[1441]), .feature_accum(feature_accums[1441]));
  accum_calculator ac1442(.scan_win(scan_win1442), .rectangle1_x(rectangle1_xs[1442]), .rectangle1_y(rectangle1_ys[1442]), .rectangle1_width(rectangle1_widths[1442]), .rectangle1_height(rectangle1_heights[1442]), .rectangle1_weight(rectangle1_weights[1442]), .rectangle2_x(rectangle2_xs[1442]), .rectangle2_y(rectangle2_ys[1442]), .rectangle2_width(rectangle2_widths[1442]), .rectangle2_height(rectangle2_heights[1442]), .rectangle2_weight(rectangle2_weights[1442]), .rectangle3_x(rectangle3_xs[1442]), .rectangle3_y(rectangle3_ys[1442]), .rectangle3_width(rectangle3_widths[1442]), .rectangle3_height(rectangle3_heights[1442]), .rectangle3_weight(rectangle3_weights[1442]), .feature_threshold(feature_thresholds[1442]), .feature_above(feature_aboves[1442]), .feature_below(feature_belows[1442]), .scan_win_std_dev(scan_win_std_dev[1442]), .feature_accum(feature_accums[1442]));
  accum_calculator ac1443(.scan_win(scan_win1443), .rectangle1_x(rectangle1_xs[1443]), .rectangle1_y(rectangle1_ys[1443]), .rectangle1_width(rectangle1_widths[1443]), .rectangle1_height(rectangle1_heights[1443]), .rectangle1_weight(rectangle1_weights[1443]), .rectangle2_x(rectangle2_xs[1443]), .rectangle2_y(rectangle2_ys[1443]), .rectangle2_width(rectangle2_widths[1443]), .rectangle2_height(rectangle2_heights[1443]), .rectangle2_weight(rectangle2_weights[1443]), .rectangle3_x(rectangle3_xs[1443]), .rectangle3_y(rectangle3_ys[1443]), .rectangle3_width(rectangle3_widths[1443]), .rectangle3_height(rectangle3_heights[1443]), .rectangle3_weight(rectangle3_weights[1443]), .feature_threshold(feature_thresholds[1443]), .feature_above(feature_aboves[1443]), .feature_below(feature_belows[1443]), .scan_win_std_dev(scan_win_std_dev[1443]), .feature_accum(feature_accums[1443]));
  accum_calculator ac1444(.scan_win(scan_win1444), .rectangle1_x(rectangle1_xs[1444]), .rectangle1_y(rectangle1_ys[1444]), .rectangle1_width(rectangle1_widths[1444]), .rectangle1_height(rectangle1_heights[1444]), .rectangle1_weight(rectangle1_weights[1444]), .rectangle2_x(rectangle2_xs[1444]), .rectangle2_y(rectangle2_ys[1444]), .rectangle2_width(rectangle2_widths[1444]), .rectangle2_height(rectangle2_heights[1444]), .rectangle2_weight(rectangle2_weights[1444]), .rectangle3_x(rectangle3_xs[1444]), .rectangle3_y(rectangle3_ys[1444]), .rectangle3_width(rectangle3_widths[1444]), .rectangle3_height(rectangle3_heights[1444]), .rectangle3_weight(rectangle3_weights[1444]), .feature_threshold(feature_thresholds[1444]), .feature_above(feature_aboves[1444]), .feature_below(feature_belows[1444]), .scan_win_std_dev(scan_win_std_dev[1444]), .feature_accum(feature_accums[1444]));
  accum_calculator ac1445(.scan_win(scan_win1445), .rectangle1_x(rectangle1_xs[1445]), .rectangle1_y(rectangle1_ys[1445]), .rectangle1_width(rectangle1_widths[1445]), .rectangle1_height(rectangle1_heights[1445]), .rectangle1_weight(rectangle1_weights[1445]), .rectangle2_x(rectangle2_xs[1445]), .rectangle2_y(rectangle2_ys[1445]), .rectangle2_width(rectangle2_widths[1445]), .rectangle2_height(rectangle2_heights[1445]), .rectangle2_weight(rectangle2_weights[1445]), .rectangle3_x(rectangle3_xs[1445]), .rectangle3_y(rectangle3_ys[1445]), .rectangle3_width(rectangle3_widths[1445]), .rectangle3_height(rectangle3_heights[1445]), .rectangle3_weight(rectangle3_weights[1445]), .feature_threshold(feature_thresholds[1445]), .feature_above(feature_aboves[1445]), .feature_below(feature_belows[1445]), .scan_win_std_dev(scan_win_std_dev[1445]), .feature_accum(feature_accums[1445]));
  accum_calculator ac1446(.scan_win(scan_win1446), .rectangle1_x(rectangle1_xs[1446]), .rectangle1_y(rectangle1_ys[1446]), .rectangle1_width(rectangle1_widths[1446]), .rectangle1_height(rectangle1_heights[1446]), .rectangle1_weight(rectangle1_weights[1446]), .rectangle2_x(rectangle2_xs[1446]), .rectangle2_y(rectangle2_ys[1446]), .rectangle2_width(rectangle2_widths[1446]), .rectangle2_height(rectangle2_heights[1446]), .rectangle2_weight(rectangle2_weights[1446]), .rectangle3_x(rectangle3_xs[1446]), .rectangle3_y(rectangle3_ys[1446]), .rectangle3_width(rectangle3_widths[1446]), .rectangle3_height(rectangle3_heights[1446]), .rectangle3_weight(rectangle3_weights[1446]), .feature_threshold(feature_thresholds[1446]), .feature_above(feature_aboves[1446]), .feature_below(feature_belows[1446]), .scan_win_std_dev(scan_win_std_dev[1446]), .feature_accum(feature_accums[1446]));
  accum_calculator ac1447(.scan_win(scan_win1447), .rectangle1_x(rectangle1_xs[1447]), .rectangle1_y(rectangle1_ys[1447]), .rectangle1_width(rectangle1_widths[1447]), .rectangle1_height(rectangle1_heights[1447]), .rectangle1_weight(rectangle1_weights[1447]), .rectangle2_x(rectangle2_xs[1447]), .rectangle2_y(rectangle2_ys[1447]), .rectangle2_width(rectangle2_widths[1447]), .rectangle2_height(rectangle2_heights[1447]), .rectangle2_weight(rectangle2_weights[1447]), .rectangle3_x(rectangle3_xs[1447]), .rectangle3_y(rectangle3_ys[1447]), .rectangle3_width(rectangle3_widths[1447]), .rectangle3_height(rectangle3_heights[1447]), .rectangle3_weight(rectangle3_weights[1447]), .feature_threshold(feature_thresholds[1447]), .feature_above(feature_aboves[1447]), .feature_below(feature_belows[1447]), .scan_win_std_dev(scan_win_std_dev[1447]), .feature_accum(feature_accums[1447]));
  accum_calculator ac1448(.scan_win(scan_win1448), .rectangle1_x(rectangle1_xs[1448]), .rectangle1_y(rectangle1_ys[1448]), .rectangle1_width(rectangle1_widths[1448]), .rectangle1_height(rectangle1_heights[1448]), .rectangle1_weight(rectangle1_weights[1448]), .rectangle2_x(rectangle2_xs[1448]), .rectangle2_y(rectangle2_ys[1448]), .rectangle2_width(rectangle2_widths[1448]), .rectangle2_height(rectangle2_heights[1448]), .rectangle2_weight(rectangle2_weights[1448]), .rectangle3_x(rectangle3_xs[1448]), .rectangle3_y(rectangle3_ys[1448]), .rectangle3_width(rectangle3_widths[1448]), .rectangle3_height(rectangle3_heights[1448]), .rectangle3_weight(rectangle3_weights[1448]), .feature_threshold(feature_thresholds[1448]), .feature_above(feature_aboves[1448]), .feature_below(feature_belows[1448]), .scan_win_std_dev(scan_win_std_dev[1448]), .feature_accum(feature_accums[1448]));
  accum_calculator ac1449(.scan_win(scan_win1449), .rectangle1_x(rectangle1_xs[1449]), .rectangle1_y(rectangle1_ys[1449]), .rectangle1_width(rectangle1_widths[1449]), .rectangle1_height(rectangle1_heights[1449]), .rectangle1_weight(rectangle1_weights[1449]), .rectangle2_x(rectangle2_xs[1449]), .rectangle2_y(rectangle2_ys[1449]), .rectangle2_width(rectangle2_widths[1449]), .rectangle2_height(rectangle2_heights[1449]), .rectangle2_weight(rectangle2_weights[1449]), .rectangle3_x(rectangle3_xs[1449]), .rectangle3_y(rectangle3_ys[1449]), .rectangle3_width(rectangle3_widths[1449]), .rectangle3_height(rectangle3_heights[1449]), .rectangle3_weight(rectangle3_weights[1449]), .feature_threshold(feature_thresholds[1449]), .feature_above(feature_aboves[1449]), .feature_below(feature_belows[1449]), .scan_win_std_dev(scan_win_std_dev[1449]), .feature_accum(feature_accums[1449]));
  accum_calculator ac1450(.scan_win(scan_win1450), .rectangle1_x(rectangle1_xs[1450]), .rectangle1_y(rectangle1_ys[1450]), .rectangle1_width(rectangle1_widths[1450]), .rectangle1_height(rectangle1_heights[1450]), .rectangle1_weight(rectangle1_weights[1450]), .rectangle2_x(rectangle2_xs[1450]), .rectangle2_y(rectangle2_ys[1450]), .rectangle2_width(rectangle2_widths[1450]), .rectangle2_height(rectangle2_heights[1450]), .rectangle2_weight(rectangle2_weights[1450]), .rectangle3_x(rectangle3_xs[1450]), .rectangle3_y(rectangle3_ys[1450]), .rectangle3_width(rectangle3_widths[1450]), .rectangle3_height(rectangle3_heights[1450]), .rectangle3_weight(rectangle3_weights[1450]), .feature_threshold(feature_thresholds[1450]), .feature_above(feature_aboves[1450]), .feature_below(feature_belows[1450]), .scan_win_std_dev(scan_win_std_dev[1450]), .feature_accum(feature_accums[1450]));
  accum_calculator ac1451(.scan_win(scan_win1451), .rectangle1_x(rectangle1_xs[1451]), .rectangle1_y(rectangle1_ys[1451]), .rectangle1_width(rectangle1_widths[1451]), .rectangle1_height(rectangle1_heights[1451]), .rectangle1_weight(rectangle1_weights[1451]), .rectangle2_x(rectangle2_xs[1451]), .rectangle2_y(rectangle2_ys[1451]), .rectangle2_width(rectangle2_widths[1451]), .rectangle2_height(rectangle2_heights[1451]), .rectangle2_weight(rectangle2_weights[1451]), .rectangle3_x(rectangle3_xs[1451]), .rectangle3_y(rectangle3_ys[1451]), .rectangle3_width(rectangle3_widths[1451]), .rectangle3_height(rectangle3_heights[1451]), .rectangle3_weight(rectangle3_weights[1451]), .feature_threshold(feature_thresholds[1451]), .feature_above(feature_aboves[1451]), .feature_below(feature_belows[1451]), .scan_win_std_dev(scan_win_std_dev[1451]), .feature_accum(feature_accums[1451]));
  accum_calculator ac1452(.scan_win(scan_win1452), .rectangle1_x(rectangle1_xs[1452]), .rectangle1_y(rectangle1_ys[1452]), .rectangle1_width(rectangle1_widths[1452]), .rectangle1_height(rectangle1_heights[1452]), .rectangle1_weight(rectangle1_weights[1452]), .rectangle2_x(rectangle2_xs[1452]), .rectangle2_y(rectangle2_ys[1452]), .rectangle2_width(rectangle2_widths[1452]), .rectangle2_height(rectangle2_heights[1452]), .rectangle2_weight(rectangle2_weights[1452]), .rectangle3_x(rectangle3_xs[1452]), .rectangle3_y(rectangle3_ys[1452]), .rectangle3_width(rectangle3_widths[1452]), .rectangle3_height(rectangle3_heights[1452]), .rectangle3_weight(rectangle3_weights[1452]), .feature_threshold(feature_thresholds[1452]), .feature_above(feature_aboves[1452]), .feature_below(feature_belows[1452]), .scan_win_std_dev(scan_win_std_dev[1452]), .feature_accum(feature_accums[1452]));
  accum_calculator ac1453(.scan_win(scan_win1453), .rectangle1_x(rectangle1_xs[1453]), .rectangle1_y(rectangle1_ys[1453]), .rectangle1_width(rectangle1_widths[1453]), .rectangle1_height(rectangle1_heights[1453]), .rectangle1_weight(rectangle1_weights[1453]), .rectangle2_x(rectangle2_xs[1453]), .rectangle2_y(rectangle2_ys[1453]), .rectangle2_width(rectangle2_widths[1453]), .rectangle2_height(rectangle2_heights[1453]), .rectangle2_weight(rectangle2_weights[1453]), .rectangle3_x(rectangle3_xs[1453]), .rectangle3_y(rectangle3_ys[1453]), .rectangle3_width(rectangle3_widths[1453]), .rectangle3_height(rectangle3_heights[1453]), .rectangle3_weight(rectangle3_weights[1453]), .feature_threshold(feature_thresholds[1453]), .feature_above(feature_aboves[1453]), .feature_below(feature_belows[1453]), .scan_win_std_dev(scan_win_std_dev[1453]), .feature_accum(feature_accums[1453]));
  accum_calculator ac1454(.scan_win(scan_win1454), .rectangle1_x(rectangle1_xs[1454]), .rectangle1_y(rectangle1_ys[1454]), .rectangle1_width(rectangle1_widths[1454]), .rectangle1_height(rectangle1_heights[1454]), .rectangle1_weight(rectangle1_weights[1454]), .rectangle2_x(rectangle2_xs[1454]), .rectangle2_y(rectangle2_ys[1454]), .rectangle2_width(rectangle2_widths[1454]), .rectangle2_height(rectangle2_heights[1454]), .rectangle2_weight(rectangle2_weights[1454]), .rectangle3_x(rectangle3_xs[1454]), .rectangle3_y(rectangle3_ys[1454]), .rectangle3_width(rectangle3_widths[1454]), .rectangle3_height(rectangle3_heights[1454]), .rectangle3_weight(rectangle3_weights[1454]), .feature_threshold(feature_thresholds[1454]), .feature_above(feature_aboves[1454]), .feature_below(feature_belows[1454]), .scan_win_std_dev(scan_win_std_dev[1454]), .feature_accum(feature_accums[1454]));
  accum_calculator ac1455(.scan_win(scan_win1455), .rectangle1_x(rectangle1_xs[1455]), .rectangle1_y(rectangle1_ys[1455]), .rectangle1_width(rectangle1_widths[1455]), .rectangle1_height(rectangle1_heights[1455]), .rectangle1_weight(rectangle1_weights[1455]), .rectangle2_x(rectangle2_xs[1455]), .rectangle2_y(rectangle2_ys[1455]), .rectangle2_width(rectangle2_widths[1455]), .rectangle2_height(rectangle2_heights[1455]), .rectangle2_weight(rectangle2_weights[1455]), .rectangle3_x(rectangle3_xs[1455]), .rectangle3_y(rectangle3_ys[1455]), .rectangle3_width(rectangle3_widths[1455]), .rectangle3_height(rectangle3_heights[1455]), .rectangle3_weight(rectangle3_weights[1455]), .feature_threshold(feature_thresholds[1455]), .feature_above(feature_aboves[1455]), .feature_below(feature_belows[1455]), .scan_win_std_dev(scan_win_std_dev[1455]), .feature_accum(feature_accums[1455]));
  accum_calculator ac1456(.scan_win(scan_win1456), .rectangle1_x(rectangle1_xs[1456]), .rectangle1_y(rectangle1_ys[1456]), .rectangle1_width(rectangle1_widths[1456]), .rectangle1_height(rectangle1_heights[1456]), .rectangle1_weight(rectangle1_weights[1456]), .rectangle2_x(rectangle2_xs[1456]), .rectangle2_y(rectangle2_ys[1456]), .rectangle2_width(rectangle2_widths[1456]), .rectangle2_height(rectangle2_heights[1456]), .rectangle2_weight(rectangle2_weights[1456]), .rectangle3_x(rectangle3_xs[1456]), .rectangle3_y(rectangle3_ys[1456]), .rectangle3_width(rectangle3_widths[1456]), .rectangle3_height(rectangle3_heights[1456]), .rectangle3_weight(rectangle3_weights[1456]), .feature_threshold(feature_thresholds[1456]), .feature_above(feature_aboves[1456]), .feature_below(feature_belows[1456]), .scan_win_std_dev(scan_win_std_dev[1456]), .feature_accum(feature_accums[1456]));
  accum_calculator ac1457(.scan_win(scan_win1457), .rectangle1_x(rectangle1_xs[1457]), .rectangle1_y(rectangle1_ys[1457]), .rectangle1_width(rectangle1_widths[1457]), .rectangle1_height(rectangle1_heights[1457]), .rectangle1_weight(rectangle1_weights[1457]), .rectangle2_x(rectangle2_xs[1457]), .rectangle2_y(rectangle2_ys[1457]), .rectangle2_width(rectangle2_widths[1457]), .rectangle2_height(rectangle2_heights[1457]), .rectangle2_weight(rectangle2_weights[1457]), .rectangle3_x(rectangle3_xs[1457]), .rectangle3_y(rectangle3_ys[1457]), .rectangle3_width(rectangle3_widths[1457]), .rectangle3_height(rectangle3_heights[1457]), .rectangle3_weight(rectangle3_weights[1457]), .feature_threshold(feature_thresholds[1457]), .feature_above(feature_aboves[1457]), .feature_below(feature_belows[1457]), .scan_win_std_dev(scan_win_std_dev[1457]), .feature_accum(feature_accums[1457]));
  accum_calculator ac1458(.scan_win(scan_win1458), .rectangle1_x(rectangle1_xs[1458]), .rectangle1_y(rectangle1_ys[1458]), .rectangle1_width(rectangle1_widths[1458]), .rectangle1_height(rectangle1_heights[1458]), .rectangle1_weight(rectangle1_weights[1458]), .rectangle2_x(rectangle2_xs[1458]), .rectangle2_y(rectangle2_ys[1458]), .rectangle2_width(rectangle2_widths[1458]), .rectangle2_height(rectangle2_heights[1458]), .rectangle2_weight(rectangle2_weights[1458]), .rectangle3_x(rectangle3_xs[1458]), .rectangle3_y(rectangle3_ys[1458]), .rectangle3_width(rectangle3_widths[1458]), .rectangle3_height(rectangle3_heights[1458]), .rectangle3_weight(rectangle3_weights[1458]), .feature_threshold(feature_thresholds[1458]), .feature_above(feature_aboves[1458]), .feature_below(feature_belows[1458]), .scan_win_std_dev(scan_win_std_dev[1458]), .feature_accum(feature_accums[1458]));
  accum_calculator ac1459(.scan_win(scan_win1459), .rectangle1_x(rectangle1_xs[1459]), .rectangle1_y(rectangle1_ys[1459]), .rectangle1_width(rectangle1_widths[1459]), .rectangle1_height(rectangle1_heights[1459]), .rectangle1_weight(rectangle1_weights[1459]), .rectangle2_x(rectangle2_xs[1459]), .rectangle2_y(rectangle2_ys[1459]), .rectangle2_width(rectangle2_widths[1459]), .rectangle2_height(rectangle2_heights[1459]), .rectangle2_weight(rectangle2_weights[1459]), .rectangle3_x(rectangle3_xs[1459]), .rectangle3_y(rectangle3_ys[1459]), .rectangle3_width(rectangle3_widths[1459]), .rectangle3_height(rectangle3_heights[1459]), .rectangle3_weight(rectangle3_weights[1459]), .feature_threshold(feature_thresholds[1459]), .feature_above(feature_aboves[1459]), .feature_below(feature_belows[1459]), .scan_win_std_dev(scan_win_std_dev[1459]), .feature_accum(feature_accums[1459]));
  accum_calculator ac1460(.scan_win(scan_win1460), .rectangle1_x(rectangle1_xs[1460]), .rectangle1_y(rectangle1_ys[1460]), .rectangle1_width(rectangle1_widths[1460]), .rectangle1_height(rectangle1_heights[1460]), .rectangle1_weight(rectangle1_weights[1460]), .rectangle2_x(rectangle2_xs[1460]), .rectangle2_y(rectangle2_ys[1460]), .rectangle2_width(rectangle2_widths[1460]), .rectangle2_height(rectangle2_heights[1460]), .rectangle2_weight(rectangle2_weights[1460]), .rectangle3_x(rectangle3_xs[1460]), .rectangle3_y(rectangle3_ys[1460]), .rectangle3_width(rectangle3_widths[1460]), .rectangle3_height(rectangle3_heights[1460]), .rectangle3_weight(rectangle3_weights[1460]), .feature_threshold(feature_thresholds[1460]), .feature_above(feature_aboves[1460]), .feature_below(feature_belows[1460]), .scan_win_std_dev(scan_win_std_dev[1460]), .feature_accum(feature_accums[1460]));
  accum_calculator ac1461(.scan_win(scan_win1461), .rectangle1_x(rectangle1_xs[1461]), .rectangle1_y(rectangle1_ys[1461]), .rectangle1_width(rectangle1_widths[1461]), .rectangle1_height(rectangle1_heights[1461]), .rectangle1_weight(rectangle1_weights[1461]), .rectangle2_x(rectangle2_xs[1461]), .rectangle2_y(rectangle2_ys[1461]), .rectangle2_width(rectangle2_widths[1461]), .rectangle2_height(rectangle2_heights[1461]), .rectangle2_weight(rectangle2_weights[1461]), .rectangle3_x(rectangle3_xs[1461]), .rectangle3_y(rectangle3_ys[1461]), .rectangle3_width(rectangle3_widths[1461]), .rectangle3_height(rectangle3_heights[1461]), .rectangle3_weight(rectangle3_weights[1461]), .feature_threshold(feature_thresholds[1461]), .feature_above(feature_aboves[1461]), .feature_below(feature_belows[1461]), .scan_win_std_dev(scan_win_std_dev[1461]), .feature_accum(feature_accums[1461]));
  accum_calculator ac1462(.scan_win(scan_win1462), .rectangle1_x(rectangle1_xs[1462]), .rectangle1_y(rectangle1_ys[1462]), .rectangle1_width(rectangle1_widths[1462]), .rectangle1_height(rectangle1_heights[1462]), .rectangle1_weight(rectangle1_weights[1462]), .rectangle2_x(rectangle2_xs[1462]), .rectangle2_y(rectangle2_ys[1462]), .rectangle2_width(rectangle2_widths[1462]), .rectangle2_height(rectangle2_heights[1462]), .rectangle2_weight(rectangle2_weights[1462]), .rectangle3_x(rectangle3_xs[1462]), .rectangle3_y(rectangle3_ys[1462]), .rectangle3_width(rectangle3_widths[1462]), .rectangle3_height(rectangle3_heights[1462]), .rectangle3_weight(rectangle3_weights[1462]), .feature_threshold(feature_thresholds[1462]), .feature_above(feature_aboves[1462]), .feature_below(feature_belows[1462]), .scan_win_std_dev(scan_win_std_dev[1462]), .feature_accum(feature_accums[1462]));
  accum_calculator ac1463(.scan_win(scan_win1463), .rectangle1_x(rectangle1_xs[1463]), .rectangle1_y(rectangle1_ys[1463]), .rectangle1_width(rectangle1_widths[1463]), .rectangle1_height(rectangle1_heights[1463]), .rectangle1_weight(rectangle1_weights[1463]), .rectangle2_x(rectangle2_xs[1463]), .rectangle2_y(rectangle2_ys[1463]), .rectangle2_width(rectangle2_widths[1463]), .rectangle2_height(rectangle2_heights[1463]), .rectangle2_weight(rectangle2_weights[1463]), .rectangle3_x(rectangle3_xs[1463]), .rectangle3_y(rectangle3_ys[1463]), .rectangle3_width(rectangle3_widths[1463]), .rectangle3_height(rectangle3_heights[1463]), .rectangle3_weight(rectangle3_weights[1463]), .feature_threshold(feature_thresholds[1463]), .feature_above(feature_aboves[1463]), .feature_below(feature_belows[1463]), .scan_win_std_dev(scan_win_std_dev[1463]), .feature_accum(feature_accums[1463]));
  accum_calculator ac1464(.scan_win(scan_win1464), .rectangle1_x(rectangle1_xs[1464]), .rectangle1_y(rectangle1_ys[1464]), .rectangle1_width(rectangle1_widths[1464]), .rectangle1_height(rectangle1_heights[1464]), .rectangle1_weight(rectangle1_weights[1464]), .rectangle2_x(rectangle2_xs[1464]), .rectangle2_y(rectangle2_ys[1464]), .rectangle2_width(rectangle2_widths[1464]), .rectangle2_height(rectangle2_heights[1464]), .rectangle2_weight(rectangle2_weights[1464]), .rectangle3_x(rectangle3_xs[1464]), .rectangle3_y(rectangle3_ys[1464]), .rectangle3_width(rectangle3_widths[1464]), .rectangle3_height(rectangle3_heights[1464]), .rectangle3_weight(rectangle3_weights[1464]), .feature_threshold(feature_thresholds[1464]), .feature_above(feature_aboves[1464]), .feature_below(feature_belows[1464]), .scan_win_std_dev(scan_win_std_dev[1464]), .feature_accum(feature_accums[1464]));
  accum_calculator ac1465(.scan_win(scan_win1465), .rectangle1_x(rectangle1_xs[1465]), .rectangle1_y(rectangle1_ys[1465]), .rectangle1_width(rectangle1_widths[1465]), .rectangle1_height(rectangle1_heights[1465]), .rectangle1_weight(rectangle1_weights[1465]), .rectangle2_x(rectangle2_xs[1465]), .rectangle2_y(rectangle2_ys[1465]), .rectangle2_width(rectangle2_widths[1465]), .rectangle2_height(rectangle2_heights[1465]), .rectangle2_weight(rectangle2_weights[1465]), .rectangle3_x(rectangle3_xs[1465]), .rectangle3_y(rectangle3_ys[1465]), .rectangle3_width(rectangle3_widths[1465]), .rectangle3_height(rectangle3_heights[1465]), .rectangle3_weight(rectangle3_weights[1465]), .feature_threshold(feature_thresholds[1465]), .feature_above(feature_aboves[1465]), .feature_below(feature_belows[1465]), .scan_win_std_dev(scan_win_std_dev[1465]), .feature_accum(feature_accums[1465]));
  accum_calculator ac1466(.scan_win(scan_win1466), .rectangle1_x(rectangle1_xs[1466]), .rectangle1_y(rectangle1_ys[1466]), .rectangle1_width(rectangle1_widths[1466]), .rectangle1_height(rectangle1_heights[1466]), .rectangle1_weight(rectangle1_weights[1466]), .rectangle2_x(rectangle2_xs[1466]), .rectangle2_y(rectangle2_ys[1466]), .rectangle2_width(rectangle2_widths[1466]), .rectangle2_height(rectangle2_heights[1466]), .rectangle2_weight(rectangle2_weights[1466]), .rectangle3_x(rectangle3_xs[1466]), .rectangle3_y(rectangle3_ys[1466]), .rectangle3_width(rectangle3_widths[1466]), .rectangle3_height(rectangle3_heights[1466]), .rectangle3_weight(rectangle3_weights[1466]), .feature_threshold(feature_thresholds[1466]), .feature_above(feature_aboves[1466]), .feature_below(feature_belows[1466]), .scan_win_std_dev(scan_win_std_dev[1466]), .feature_accum(feature_accums[1466]));
  accum_calculator ac1467(.scan_win(scan_win1467), .rectangle1_x(rectangle1_xs[1467]), .rectangle1_y(rectangle1_ys[1467]), .rectangle1_width(rectangle1_widths[1467]), .rectangle1_height(rectangle1_heights[1467]), .rectangle1_weight(rectangle1_weights[1467]), .rectangle2_x(rectangle2_xs[1467]), .rectangle2_y(rectangle2_ys[1467]), .rectangle2_width(rectangle2_widths[1467]), .rectangle2_height(rectangle2_heights[1467]), .rectangle2_weight(rectangle2_weights[1467]), .rectangle3_x(rectangle3_xs[1467]), .rectangle3_y(rectangle3_ys[1467]), .rectangle3_width(rectangle3_widths[1467]), .rectangle3_height(rectangle3_heights[1467]), .rectangle3_weight(rectangle3_weights[1467]), .feature_threshold(feature_thresholds[1467]), .feature_above(feature_aboves[1467]), .feature_below(feature_belows[1467]), .scan_win_std_dev(scan_win_std_dev[1467]), .feature_accum(feature_accums[1467]));
  accum_calculator ac1468(.scan_win(scan_win1468), .rectangle1_x(rectangle1_xs[1468]), .rectangle1_y(rectangle1_ys[1468]), .rectangle1_width(rectangle1_widths[1468]), .rectangle1_height(rectangle1_heights[1468]), .rectangle1_weight(rectangle1_weights[1468]), .rectangle2_x(rectangle2_xs[1468]), .rectangle2_y(rectangle2_ys[1468]), .rectangle2_width(rectangle2_widths[1468]), .rectangle2_height(rectangle2_heights[1468]), .rectangle2_weight(rectangle2_weights[1468]), .rectangle3_x(rectangle3_xs[1468]), .rectangle3_y(rectangle3_ys[1468]), .rectangle3_width(rectangle3_widths[1468]), .rectangle3_height(rectangle3_heights[1468]), .rectangle3_weight(rectangle3_weights[1468]), .feature_threshold(feature_thresholds[1468]), .feature_above(feature_aboves[1468]), .feature_below(feature_belows[1468]), .scan_win_std_dev(scan_win_std_dev[1468]), .feature_accum(feature_accums[1468]));
  accum_calculator ac1469(.scan_win(scan_win1469), .rectangle1_x(rectangle1_xs[1469]), .rectangle1_y(rectangle1_ys[1469]), .rectangle1_width(rectangle1_widths[1469]), .rectangle1_height(rectangle1_heights[1469]), .rectangle1_weight(rectangle1_weights[1469]), .rectangle2_x(rectangle2_xs[1469]), .rectangle2_y(rectangle2_ys[1469]), .rectangle2_width(rectangle2_widths[1469]), .rectangle2_height(rectangle2_heights[1469]), .rectangle2_weight(rectangle2_weights[1469]), .rectangle3_x(rectangle3_xs[1469]), .rectangle3_y(rectangle3_ys[1469]), .rectangle3_width(rectangle3_widths[1469]), .rectangle3_height(rectangle3_heights[1469]), .rectangle3_weight(rectangle3_weights[1469]), .feature_threshold(feature_thresholds[1469]), .feature_above(feature_aboves[1469]), .feature_below(feature_belows[1469]), .scan_win_std_dev(scan_win_std_dev[1469]), .feature_accum(feature_accums[1469]));
  accum_calculator ac1470(.scan_win(scan_win1470), .rectangle1_x(rectangle1_xs[1470]), .rectangle1_y(rectangle1_ys[1470]), .rectangle1_width(rectangle1_widths[1470]), .rectangle1_height(rectangle1_heights[1470]), .rectangle1_weight(rectangle1_weights[1470]), .rectangle2_x(rectangle2_xs[1470]), .rectangle2_y(rectangle2_ys[1470]), .rectangle2_width(rectangle2_widths[1470]), .rectangle2_height(rectangle2_heights[1470]), .rectangle2_weight(rectangle2_weights[1470]), .rectangle3_x(rectangle3_xs[1470]), .rectangle3_y(rectangle3_ys[1470]), .rectangle3_width(rectangle3_widths[1470]), .rectangle3_height(rectangle3_heights[1470]), .rectangle3_weight(rectangle3_weights[1470]), .feature_threshold(feature_thresholds[1470]), .feature_above(feature_aboves[1470]), .feature_below(feature_belows[1470]), .scan_win_std_dev(scan_win_std_dev[1470]), .feature_accum(feature_accums[1470]));
  accum_calculator ac1471(.scan_win(scan_win1471), .rectangle1_x(rectangle1_xs[1471]), .rectangle1_y(rectangle1_ys[1471]), .rectangle1_width(rectangle1_widths[1471]), .rectangle1_height(rectangle1_heights[1471]), .rectangle1_weight(rectangle1_weights[1471]), .rectangle2_x(rectangle2_xs[1471]), .rectangle2_y(rectangle2_ys[1471]), .rectangle2_width(rectangle2_widths[1471]), .rectangle2_height(rectangle2_heights[1471]), .rectangle2_weight(rectangle2_weights[1471]), .rectangle3_x(rectangle3_xs[1471]), .rectangle3_y(rectangle3_ys[1471]), .rectangle3_width(rectangle3_widths[1471]), .rectangle3_height(rectangle3_heights[1471]), .rectangle3_weight(rectangle3_weights[1471]), .feature_threshold(feature_thresholds[1471]), .feature_above(feature_aboves[1471]), .feature_below(feature_belows[1471]), .scan_win_std_dev(scan_win_std_dev[1471]), .feature_accum(feature_accums[1471]));
  accum_calculator ac1472(.scan_win(scan_win1472), .rectangle1_x(rectangle1_xs[1472]), .rectangle1_y(rectangle1_ys[1472]), .rectangle1_width(rectangle1_widths[1472]), .rectangle1_height(rectangle1_heights[1472]), .rectangle1_weight(rectangle1_weights[1472]), .rectangle2_x(rectangle2_xs[1472]), .rectangle2_y(rectangle2_ys[1472]), .rectangle2_width(rectangle2_widths[1472]), .rectangle2_height(rectangle2_heights[1472]), .rectangle2_weight(rectangle2_weights[1472]), .rectangle3_x(rectangle3_xs[1472]), .rectangle3_y(rectangle3_ys[1472]), .rectangle3_width(rectangle3_widths[1472]), .rectangle3_height(rectangle3_heights[1472]), .rectangle3_weight(rectangle3_weights[1472]), .feature_threshold(feature_thresholds[1472]), .feature_above(feature_aboves[1472]), .feature_below(feature_belows[1472]), .scan_win_std_dev(scan_win_std_dev[1472]), .feature_accum(feature_accums[1472]));
  accum_calculator ac1473(.scan_win(scan_win1473), .rectangle1_x(rectangle1_xs[1473]), .rectangle1_y(rectangle1_ys[1473]), .rectangle1_width(rectangle1_widths[1473]), .rectangle1_height(rectangle1_heights[1473]), .rectangle1_weight(rectangle1_weights[1473]), .rectangle2_x(rectangle2_xs[1473]), .rectangle2_y(rectangle2_ys[1473]), .rectangle2_width(rectangle2_widths[1473]), .rectangle2_height(rectangle2_heights[1473]), .rectangle2_weight(rectangle2_weights[1473]), .rectangle3_x(rectangle3_xs[1473]), .rectangle3_y(rectangle3_ys[1473]), .rectangle3_width(rectangle3_widths[1473]), .rectangle3_height(rectangle3_heights[1473]), .rectangle3_weight(rectangle3_weights[1473]), .feature_threshold(feature_thresholds[1473]), .feature_above(feature_aboves[1473]), .feature_below(feature_belows[1473]), .scan_win_std_dev(scan_win_std_dev[1473]), .feature_accum(feature_accums[1473]));
  accum_calculator ac1474(.scan_win(scan_win1474), .rectangle1_x(rectangle1_xs[1474]), .rectangle1_y(rectangle1_ys[1474]), .rectangle1_width(rectangle1_widths[1474]), .rectangle1_height(rectangle1_heights[1474]), .rectangle1_weight(rectangle1_weights[1474]), .rectangle2_x(rectangle2_xs[1474]), .rectangle2_y(rectangle2_ys[1474]), .rectangle2_width(rectangle2_widths[1474]), .rectangle2_height(rectangle2_heights[1474]), .rectangle2_weight(rectangle2_weights[1474]), .rectangle3_x(rectangle3_xs[1474]), .rectangle3_y(rectangle3_ys[1474]), .rectangle3_width(rectangle3_widths[1474]), .rectangle3_height(rectangle3_heights[1474]), .rectangle3_weight(rectangle3_weights[1474]), .feature_threshold(feature_thresholds[1474]), .feature_above(feature_aboves[1474]), .feature_below(feature_belows[1474]), .scan_win_std_dev(scan_win_std_dev[1474]), .feature_accum(feature_accums[1474]));
  accum_calculator ac1475(.scan_win(scan_win1475), .rectangle1_x(rectangle1_xs[1475]), .rectangle1_y(rectangle1_ys[1475]), .rectangle1_width(rectangle1_widths[1475]), .rectangle1_height(rectangle1_heights[1475]), .rectangle1_weight(rectangle1_weights[1475]), .rectangle2_x(rectangle2_xs[1475]), .rectangle2_y(rectangle2_ys[1475]), .rectangle2_width(rectangle2_widths[1475]), .rectangle2_height(rectangle2_heights[1475]), .rectangle2_weight(rectangle2_weights[1475]), .rectangle3_x(rectangle3_xs[1475]), .rectangle3_y(rectangle3_ys[1475]), .rectangle3_width(rectangle3_widths[1475]), .rectangle3_height(rectangle3_heights[1475]), .rectangle3_weight(rectangle3_weights[1475]), .feature_threshold(feature_thresholds[1475]), .feature_above(feature_aboves[1475]), .feature_below(feature_belows[1475]), .scan_win_std_dev(scan_win_std_dev[1475]), .feature_accum(feature_accums[1475]));
  accum_calculator ac1476(.scan_win(scan_win1476), .rectangle1_x(rectangle1_xs[1476]), .rectangle1_y(rectangle1_ys[1476]), .rectangle1_width(rectangle1_widths[1476]), .rectangle1_height(rectangle1_heights[1476]), .rectangle1_weight(rectangle1_weights[1476]), .rectangle2_x(rectangle2_xs[1476]), .rectangle2_y(rectangle2_ys[1476]), .rectangle2_width(rectangle2_widths[1476]), .rectangle2_height(rectangle2_heights[1476]), .rectangle2_weight(rectangle2_weights[1476]), .rectangle3_x(rectangle3_xs[1476]), .rectangle3_y(rectangle3_ys[1476]), .rectangle3_width(rectangle3_widths[1476]), .rectangle3_height(rectangle3_heights[1476]), .rectangle3_weight(rectangle3_weights[1476]), .feature_threshold(feature_thresholds[1476]), .feature_above(feature_aboves[1476]), .feature_below(feature_belows[1476]), .scan_win_std_dev(scan_win_std_dev[1476]), .feature_accum(feature_accums[1476]));
  accum_calculator ac1477(.scan_win(scan_win1477), .rectangle1_x(rectangle1_xs[1477]), .rectangle1_y(rectangle1_ys[1477]), .rectangle1_width(rectangle1_widths[1477]), .rectangle1_height(rectangle1_heights[1477]), .rectangle1_weight(rectangle1_weights[1477]), .rectangle2_x(rectangle2_xs[1477]), .rectangle2_y(rectangle2_ys[1477]), .rectangle2_width(rectangle2_widths[1477]), .rectangle2_height(rectangle2_heights[1477]), .rectangle2_weight(rectangle2_weights[1477]), .rectangle3_x(rectangle3_xs[1477]), .rectangle3_y(rectangle3_ys[1477]), .rectangle3_width(rectangle3_widths[1477]), .rectangle3_height(rectangle3_heights[1477]), .rectangle3_weight(rectangle3_weights[1477]), .feature_threshold(feature_thresholds[1477]), .feature_above(feature_aboves[1477]), .feature_below(feature_belows[1477]), .scan_win_std_dev(scan_win_std_dev[1477]), .feature_accum(feature_accums[1477]));
  accum_calculator ac1478(.scan_win(scan_win1478), .rectangle1_x(rectangle1_xs[1478]), .rectangle1_y(rectangle1_ys[1478]), .rectangle1_width(rectangle1_widths[1478]), .rectangle1_height(rectangle1_heights[1478]), .rectangle1_weight(rectangle1_weights[1478]), .rectangle2_x(rectangle2_xs[1478]), .rectangle2_y(rectangle2_ys[1478]), .rectangle2_width(rectangle2_widths[1478]), .rectangle2_height(rectangle2_heights[1478]), .rectangle2_weight(rectangle2_weights[1478]), .rectangle3_x(rectangle3_xs[1478]), .rectangle3_y(rectangle3_ys[1478]), .rectangle3_width(rectangle3_widths[1478]), .rectangle3_height(rectangle3_heights[1478]), .rectangle3_weight(rectangle3_weights[1478]), .feature_threshold(feature_thresholds[1478]), .feature_above(feature_aboves[1478]), .feature_below(feature_belows[1478]), .scan_win_std_dev(scan_win_std_dev[1478]), .feature_accum(feature_accums[1478]));
  accum_calculator ac1479(.scan_win(scan_win1479), .rectangle1_x(rectangle1_xs[1479]), .rectangle1_y(rectangle1_ys[1479]), .rectangle1_width(rectangle1_widths[1479]), .rectangle1_height(rectangle1_heights[1479]), .rectangle1_weight(rectangle1_weights[1479]), .rectangle2_x(rectangle2_xs[1479]), .rectangle2_y(rectangle2_ys[1479]), .rectangle2_width(rectangle2_widths[1479]), .rectangle2_height(rectangle2_heights[1479]), .rectangle2_weight(rectangle2_weights[1479]), .rectangle3_x(rectangle3_xs[1479]), .rectangle3_y(rectangle3_ys[1479]), .rectangle3_width(rectangle3_widths[1479]), .rectangle3_height(rectangle3_heights[1479]), .rectangle3_weight(rectangle3_weights[1479]), .feature_threshold(feature_thresholds[1479]), .feature_above(feature_aboves[1479]), .feature_below(feature_belows[1479]), .scan_win_std_dev(scan_win_std_dev[1479]), .feature_accum(feature_accums[1479]));
  accum_calculator ac1480(.scan_win(scan_win1480), .rectangle1_x(rectangle1_xs[1480]), .rectangle1_y(rectangle1_ys[1480]), .rectangle1_width(rectangle1_widths[1480]), .rectangle1_height(rectangle1_heights[1480]), .rectangle1_weight(rectangle1_weights[1480]), .rectangle2_x(rectangle2_xs[1480]), .rectangle2_y(rectangle2_ys[1480]), .rectangle2_width(rectangle2_widths[1480]), .rectangle2_height(rectangle2_heights[1480]), .rectangle2_weight(rectangle2_weights[1480]), .rectangle3_x(rectangle3_xs[1480]), .rectangle3_y(rectangle3_ys[1480]), .rectangle3_width(rectangle3_widths[1480]), .rectangle3_height(rectangle3_heights[1480]), .rectangle3_weight(rectangle3_weights[1480]), .feature_threshold(feature_thresholds[1480]), .feature_above(feature_aboves[1480]), .feature_below(feature_belows[1480]), .scan_win_std_dev(scan_win_std_dev[1480]), .feature_accum(feature_accums[1480]));
  accum_calculator ac1481(.scan_win(scan_win1481), .rectangle1_x(rectangle1_xs[1481]), .rectangle1_y(rectangle1_ys[1481]), .rectangle1_width(rectangle1_widths[1481]), .rectangle1_height(rectangle1_heights[1481]), .rectangle1_weight(rectangle1_weights[1481]), .rectangle2_x(rectangle2_xs[1481]), .rectangle2_y(rectangle2_ys[1481]), .rectangle2_width(rectangle2_widths[1481]), .rectangle2_height(rectangle2_heights[1481]), .rectangle2_weight(rectangle2_weights[1481]), .rectangle3_x(rectangle3_xs[1481]), .rectangle3_y(rectangle3_ys[1481]), .rectangle3_width(rectangle3_widths[1481]), .rectangle3_height(rectangle3_heights[1481]), .rectangle3_weight(rectangle3_weights[1481]), .feature_threshold(feature_thresholds[1481]), .feature_above(feature_aboves[1481]), .feature_below(feature_belows[1481]), .scan_win_std_dev(scan_win_std_dev[1481]), .feature_accum(feature_accums[1481]));
  accum_calculator ac1482(.scan_win(scan_win1482), .rectangle1_x(rectangle1_xs[1482]), .rectangle1_y(rectangle1_ys[1482]), .rectangle1_width(rectangle1_widths[1482]), .rectangle1_height(rectangle1_heights[1482]), .rectangle1_weight(rectangle1_weights[1482]), .rectangle2_x(rectangle2_xs[1482]), .rectangle2_y(rectangle2_ys[1482]), .rectangle2_width(rectangle2_widths[1482]), .rectangle2_height(rectangle2_heights[1482]), .rectangle2_weight(rectangle2_weights[1482]), .rectangle3_x(rectangle3_xs[1482]), .rectangle3_y(rectangle3_ys[1482]), .rectangle3_width(rectangle3_widths[1482]), .rectangle3_height(rectangle3_heights[1482]), .rectangle3_weight(rectangle3_weights[1482]), .feature_threshold(feature_thresholds[1482]), .feature_above(feature_aboves[1482]), .feature_below(feature_belows[1482]), .scan_win_std_dev(scan_win_std_dev[1482]), .feature_accum(feature_accums[1482]));
  accum_calculator ac1483(.scan_win(scan_win1483), .rectangle1_x(rectangle1_xs[1483]), .rectangle1_y(rectangle1_ys[1483]), .rectangle1_width(rectangle1_widths[1483]), .rectangle1_height(rectangle1_heights[1483]), .rectangle1_weight(rectangle1_weights[1483]), .rectangle2_x(rectangle2_xs[1483]), .rectangle2_y(rectangle2_ys[1483]), .rectangle2_width(rectangle2_widths[1483]), .rectangle2_height(rectangle2_heights[1483]), .rectangle2_weight(rectangle2_weights[1483]), .rectangle3_x(rectangle3_xs[1483]), .rectangle3_y(rectangle3_ys[1483]), .rectangle3_width(rectangle3_widths[1483]), .rectangle3_height(rectangle3_heights[1483]), .rectangle3_weight(rectangle3_weights[1483]), .feature_threshold(feature_thresholds[1483]), .feature_above(feature_aboves[1483]), .feature_below(feature_belows[1483]), .scan_win_std_dev(scan_win_std_dev[1483]), .feature_accum(feature_accums[1483]));
  accum_calculator ac1484(.scan_win(scan_win1484), .rectangle1_x(rectangle1_xs[1484]), .rectangle1_y(rectangle1_ys[1484]), .rectangle1_width(rectangle1_widths[1484]), .rectangle1_height(rectangle1_heights[1484]), .rectangle1_weight(rectangle1_weights[1484]), .rectangle2_x(rectangle2_xs[1484]), .rectangle2_y(rectangle2_ys[1484]), .rectangle2_width(rectangle2_widths[1484]), .rectangle2_height(rectangle2_heights[1484]), .rectangle2_weight(rectangle2_weights[1484]), .rectangle3_x(rectangle3_xs[1484]), .rectangle3_y(rectangle3_ys[1484]), .rectangle3_width(rectangle3_widths[1484]), .rectangle3_height(rectangle3_heights[1484]), .rectangle3_weight(rectangle3_weights[1484]), .feature_threshold(feature_thresholds[1484]), .feature_above(feature_aboves[1484]), .feature_below(feature_belows[1484]), .scan_win_std_dev(scan_win_std_dev[1484]), .feature_accum(feature_accums[1484]));
  accum_calculator ac1485(.scan_win(scan_win1485), .rectangle1_x(rectangle1_xs[1485]), .rectangle1_y(rectangle1_ys[1485]), .rectangle1_width(rectangle1_widths[1485]), .rectangle1_height(rectangle1_heights[1485]), .rectangle1_weight(rectangle1_weights[1485]), .rectangle2_x(rectangle2_xs[1485]), .rectangle2_y(rectangle2_ys[1485]), .rectangle2_width(rectangle2_widths[1485]), .rectangle2_height(rectangle2_heights[1485]), .rectangle2_weight(rectangle2_weights[1485]), .rectangle3_x(rectangle3_xs[1485]), .rectangle3_y(rectangle3_ys[1485]), .rectangle3_width(rectangle3_widths[1485]), .rectangle3_height(rectangle3_heights[1485]), .rectangle3_weight(rectangle3_weights[1485]), .feature_threshold(feature_thresholds[1485]), .feature_above(feature_aboves[1485]), .feature_below(feature_belows[1485]), .scan_win_std_dev(scan_win_std_dev[1485]), .feature_accum(feature_accums[1485]));
  accum_calculator ac1486(.scan_win(scan_win1486), .rectangle1_x(rectangle1_xs[1486]), .rectangle1_y(rectangle1_ys[1486]), .rectangle1_width(rectangle1_widths[1486]), .rectangle1_height(rectangle1_heights[1486]), .rectangle1_weight(rectangle1_weights[1486]), .rectangle2_x(rectangle2_xs[1486]), .rectangle2_y(rectangle2_ys[1486]), .rectangle2_width(rectangle2_widths[1486]), .rectangle2_height(rectangle2_heights[1486]), .rectangle2_weight(rectangle2_weights[1486]), .rectangle3_x(rectangle3_xs[1486]), .rectangle3_y(rectangle3_ys[1486]), .rectangle3_width(rectangle3_widths[1486]), .rectangle3_height(rectangle3_heights[1486]), .rectangle3_weight(rectangle3_weights[1486]), .feature_threshold(feature_thresholds[1486]), .feature_above(feature_aboves[1486]), .feature_below(feature_belows[1486]), .scan_win_std_dev(scan_win_std_dev[1486]), .feature_accum(feature_accums[1486]));
  accum_calculator ac1487(.scan_win(scan_win1487), .rectangle1_x(rectangle1_xs[1487]), .rectangle1_y(rectangle1_ys[1487]), .rectangle1_width(rectangle1_widths[1487]), .rectangle1_height(rectangle1_heights[1487]), .rectangle1_weight(rectangle1_weights[1487]), .rectangle2_x(rectangle2_xs[1487]), .rectangle2_y(rectangle2_ys[1487]), .rectangle2_width(rectangle2_widths[1487]), .rectangle2_height(rectangle2_heights[1487]), .rectangle2_weight(rectangle2_weights[1487]), .rectangle3_x(rectangle3_xs[1487]), .rectangle3_y(rectangle3_ys[1487]), .rectangle3_width(rectangle3_widths[1487]), .rectangle3_height(rectangle3_heights[1487]), .rectangle3_weight(rectangle3_weights[1487]), .feature_threshold(feature_thresholds[1487]), .feature_above(feature_aboves[1487]), .feature_below(feature_belows[1487]), .scan_win_std_dev(scan_win_std_dev[1487]), .feature_accum(feature_accums[1487]));
  accum_calculator ac1488(.scan_win(scan_win1488), .rectangle1_x(rectangle1_xs[1488]), .rectangle1_y(rectangle1_ys[1488]), .rectangle1_width(rectangle1_widths[1488]), .rectangle1_height(rectangle1_heights[1488]), .rectangle1_weight(rectangle1_weights[1488]), .rectangle2_x(rectangle2_xs[1488]), .rectangle2_y(rectangle2_ys[1488]), .rectangle2_width(rectangle2_widths[1488]), .rectangle2_height(rectangle2_heights[1488]), .rectangle2_weight(rectangle2_weights[1488]), .rectangle3_x(rectangle3_xs[1488]), .rectangle3_y(rectangle3_ys[1488]), .rectangle3_width(rectangle3_widths[1488]), .rectangle3_height(rectangle3_heights[1488]), .rectangle3_weight(rectangle3_weights[1488]), .feature_threshold(feature_thresholds[1488]), .feature_above(feature_aboves[1488]), .feature_below(feature_belows[1488]), .scan_win_std_dev(scan_win_std_dev[1488]), .feature_accum(feature_accums[1488]));
  accum_calculator ac1489(.scan_win(scan_win1489), .rectangle1_x(rectangle1_xs[1489]), .rectangle1_y(rectangle1_ys[1489]), .rectangle1_width(rectangle1_widths[1489]), .rectangle1_height(rectangle1_heights[1489]), .rectangle1_weight(rectangle1_weights[1489]), .rectangle2_x(rectangle2_xs[1489]), .rectangle2_y(rectangle2_ys[1489]), .rectangle2_width(rectangle2_widths[1489]), .rectangle2_height(rectangle2_heights[1489]), .rectangle2_weight(rectangle2_weights[1489]), .rectangle3_x(rectangle3_xs[1489]), .rectangle3_y(rectangle3_ys[1489]), .rectangle3_width(rectangle3_widths[1489]), .rectangle3_height(rectangle3_heights[1489]), .rectangle3_weight(rectangle3_weights[1489]), .feature_threshold(feature_thresholds[1489]), .feature_above(feature_aboves[1489]), .feature_below(feature_belows[1489]), .scan_win_std_dev(scan_win_std_dev[1489]), .feature_accum(feature_accums[1489]));
  accum_calculator ac1490(.scan_win(scan_win1490), .rectangle1_x(rectangle1_xs[1490]), .rectangle1_y(rectangle1_ys[1490]), .rectangle1_width(rectangle1_widths[1490]), .rectangle1_height(rectangle1_heights[1490]), .rectangle1_weight(rectangle1_weights[1490]), .rectangle2_x(rectangle2_xs[1490]), .rectangle2_y(rectangle2_ys[1490]), .rectangle2_width(rectangle2_widths[1490]), .rectangle2_height(rectangle2_heights[1490]), .rectangle2_weight(rectangle2_weights[1490]), .rectangle3_x(rectangle3_xs[1490]), .rectangle3_y(rectangle3_ys[1490]), .rectangle3_width(rectangle3_widths[1490]), .rectangle3_height(rectangle3_heights[1490]), .rectangle3_weight(rectangle3_weights[1490]), .feature_threshold(feature_thresholds[1490]), .feature_above(feature_aboves[1490]), .feature_below(feature_belows[1490]), .scan_win_std_dev(scan_win_std_dev[1490]), .feature_accum(feature_accums[1490]));
  accum_calculator ac1491(.scan_win(scan_win1491), .rectangle1_x(rectangle1_xs[1491]), .rectangle1_y(rectangle1_ys[1491]), .rectangle1_width(rectangle1_widths[1491]), .rectangle1_height(rectangle1_heights[1491]), .rectangle1_weight(rectangle1_weights[1491]), .rectangle2_x(rectangle2_xs[1491]), .rectangle2_y(rectangle2_ys[1491]), .rectangle2_width(rectangle2_widths[1491]), .rectangle2_height(rectangle2_heights[1491]), .rectangle2_weight(rectangle2_weights[1491]), .rectangle3_x(rectangle3_xs[1491]), .rectangle3_y(rectangle3_ys[1491]), .rectangle3_width(rectangle3_widths[1491]), .rectangle3_height(rectangle3_heights[1491]), .rectangle3_weight(rectangle3_weights[1491]), .feature_threshold(feature_thresholds[1491]), .feature_above(feature_aboves[1491]), .feature_below(feature_belows[1491]), .scan_win_std_dev(scan_win_std_dev[1491]), .feature_accum(feature_accums[1491]));
  accum_calculator ac1492(.scan_win(scan_win1492), .rectangle1_x(rectangle1_xs[1492]), .rectangle1_y(rectangle1_ys[1492]), .rectangle1_width(rectangle1_widths[1492]), .rectangle1_height(rectangle1_heights[1492]), .rectangle1_weight(rectangle1_weights[1492]), .rectangle2_x(rectangle2_xs[1492]), .rectangle2_y(rectangle2_ys[1492]), .rectangle2_width(rectangle2_widths[1492]), .rectangle2_height(rectangle2_heights[1492]), .rectangle2_weight(rectangle2_weights[1492]), .rectangle3_x(rectangle3_xs[1492]), .rectangle3_y(rectangle3_ys[1492]), .rectangle3_width(rectangle3_widths[1492]), .rectangle3_height(rectangle3_heights[1492]), .rectangle3_weight(rectangle3_weights[1492]), .feature_threshold(feature_thresholds[1492]), .feature_above(feature_aboves[1492]), .feature_below(feature_belows[1492]), .scan_win_std_dev(scan_win_std_dev[1492]), .feature_accum(feature_accums[1492]));
  accum_calculator ac1493(.scan_win(scan_win1493), .rectangle1_x(rectangle1_xs[1493]), .rectangle1_y(rectangle1_ys[1493]), .rectangle1_width(rectangle1_widths[1493]), .rectangle1_height(rectangle1_heights[1493]), .rectangle1_weight(rectangle1_weights[1493]), .rectangle2_x(rectangle2_xs[1493]), .rectangle2_y(rectangle2_ys[1493]), .rectangle2_width(rectangle2_widths[1493]), .rectangle2_height(rectangle2_heights[1493]), .rectangle2_weight(rectangle2_weights[1493]), .rectangle3_x(rectangle3_xs[1493]), .rectangle3_y(rectangle3_ys[1493]), .rectangle3_width(rectangle3_widths[1493]), .rectangle3_height(rectangle3_heights[1493]), .rectangle3_weight(rectangle3_weights[1493]), .feature_threshold(feature_thresholds[1493]), .feature_above(feature_aboves[1493]), .feature_below(feature_belows[1493]), .scan_win_std_dev(scan_win_std_dev[1493]), .feature_accum(feature_accums[1493]));
  accum_calculator ac1494(.scan_win(scan_win1494), .rectangle1_x(rectangle1_xs[1494]), .rectangle1_y(rectangle1_ys[1494]), .rectangle1_width(rectangle1_widths[1494]), .rectangle1_height(rectangle1_heights[1494]), .rectangle1_weight(rectangle1_weights[1494]), .rectangle2_x(rectangle2_xs[1494]), .rectangle2_y(rectangle2_ys[1494]), .rectangle2_width(rectangle2_widths[1494]), .rectangle2_height(rectangle2_heights[1494]), .rectangle2_weight(rectangle2_weights[1494]), .rectangle3_x(rectangle3_xs[1494]), .rectangle3_y(rectangle3_ys[1494]), .rectangle3_width(rectangle3_widths[1494]), .rectangle3_height(rectangle3_heights[1494]), .rectangle3_weight(rectangle3_weights[1494]), .feature_threshold(feature_thresholds[1494]), .feature_above(feature_aboves[1494]), .feature_below(feature_belows[1494]), .scan_win_std_dev(scan_win_std_dev[1494]), .feature_accum(feature_accums[1494]));
  accum_calculator ac1495(.scan_win(scan_win1495), .rectangle1_x(rectangle1_xs[1495]), .rectangle1_y(rectangle1_ys[1495]), .rectangle1_width(rectangle1_widths[1495]), .rectangle1_height(rectangle1_heights[1495]), .rectangle1_weight(rectangle1_weights[1495]), .rectangle2_x(rectangle2_xs[1495]), .rectangle2_y(rectangle2_ys[1495]), .rectangle2_width(rectangle2_widths[1495]), .rectangle2_height(rectangle2_heights[1495]), .rectangle2_weight(rectangle2_weights[1495]), .rectangle3_x(rectangle3_xs[1495]), .rectangle3_y(rectangle3_ys[1495]), .rectangle3_width(rectangle3_widths[1495]), .rectangle3_height(rectangle3_heights[1495]), .rectangle3_weight(rectangle3_weights[1495]), .feature_threshold(feature_thresholds[1495]), .feature_above(feature_aboves[1495]), .feature_below(feature_belows[1495]), .scan_win_std_dev(scan_win_std_dev[1495]), .feature_accum(feature_accums[1495]));
  accum_calculator ac1496(.scan_win(scan_win1496), .rectangle1_x(rectangle1_xs[1496]), .rectangle1_y(rectangle1_ys[1496]), .rectangle1_width(rectangle1_widths[1496]), .rectangle1_height(rectangle1_heights[1496]), .rectangle1_weight(rectangle1_weights[1496]), .rectangle2_x(rectangle2_xs[1496]), .rectangle2_y(rectangle2_ys[1496]), .rectangle2_width(rectangle2_widths[1496]), .rectangle2_height(rectangle2_heights[1496]), .rectangle2_weight(rectangle2_weights[1496]), .rectangle3_x(rectangle3_xs[1496]), .rectangle3_y(rectangle3_ys[1496]), .rectangle3_width(rectangle3_widths[1496]), .rectangle3_height(rectangle3_heights[1496]), .rectangle3_weight(rectangle3_weights[1496]), .feature_threshold(feature_thresholds[1496]), .feature_above(feature_aboves[1496]), .feature_below(feature_belows[1496]), .scan_win_std_dev(scan_win_std_dev[1496]), .feature_accum(feature_accums[1496]));
  accum_calculator ac1497(.scan_win(scan_win1497), .rectangle1_x(rectangle1_xs[1497]), .rectangle1_y(rectangle1_ys[1497]), .rectangle1_width(rectangle1_widths[1497]), .rectangle1_height(rectangle1_heights[1497]), .rectangle1_weight(rectangle1_weights[1497]), .rectangle2_x(rectangle2_xs[1497]), .rectangle2_y(rectangle2_ys[1497]), .rectangle2_width(rectangle2_widths[1497]), .rectangle2_height(rectangle2_heights[1497]), .rectangle2_weight(rectangle2_weights[1497]), .rectangle3_x(rectangle3_xs[1497]), .rectangle3_y(rectangle3_ys[1497]), .rectangle3_width(rectangle3_widths[1497]), .rectangle3_height(rectangle3_heights[1497]), .rectangle3_weight(rectangle3_weights[1497]), .feature_threshold(feature_thresholds[1497]), .feature_above(feature_aboves[1497]), .feature_below(feature_belows[1497]), .scan_win_std_dev(scan_win_std_dev[1497]), .feature_accum(feature_accums[1497]));
  accum_calculator ac1498(.scan_win(scan_win1498), .rectangle1_x(rectangle1_xs[1498]), .rectangle1_y(rectangle1_ys[1498]), .rectangle1_width(rectangle1_widths[1498]), .rectangle1_height(rectangle1_heights[1498]), .rectangle1_weight(rectangle1_weights[1498]), .rectangle2_x(rectangle2_xs[1498]), .rectangle2_y(rectangle2_ys[1498]), .rectangle2_width(rectangle2_widths[1498]), .rectangle2_height(rectangle2_heights[1498]), .rectangle2_weight(rectangle2_weights[1498]), .rectangle3_x(rectangle3_xs[1498]), .rectangle3_y(rectangle3_ys[1498]), .rectangle3_width(rectangle3_widths[1498]), .rectangle3_height(rectangle3_heights[1498]), .rectangle3_weight(rectangle3_weights[1498]), .feature_threshold(feature_thresholds[1498]), .feature_above(feature_aboves[1498]), .feature_below(feature_belows[1498]), .scan_win_std_dev(scan_win_std_dev[1498]), .feature_accum(feature_accums[1498]));
  accum_calculator ac1499(.scan_win(scan_win1499), .rectangle1_x(rectangle1_xs[1499]), .rectangle1_y(rectangle1_ys[1499]), .rectangle1_width(rectangle1_widths[1499]), .rectangle1_height(rectangle1_heights[1499]), .rectangle1_weight(rectangle1_weights[1499]), .rectangle2_x(rectangle2_xs[1499]), .rectangle2_y(rectangle2_ys[1499]), .rectangle2_width(rectangle2_widths[1499]), .rectangle2_height(rectangle2_heights[1499]), .rectangle2_weight(rectangle2_weights[1499]), .rectangle3_x(rectangle3_xs[1499]), .rectangle3_y(rectangle3_ys[1499]), .rectangle3_width(rectangle3_widths[1499]), .rectangle3_height(rectangle3_heights[1499]), .rectangle3_weight(rectangle3_weights[1499]), .feature_threshold(feature_thresholds[1499]), .feature_above(feature_aboves[1499]), .feature_below(feature_belows[1499]), .scan_win_std_dev(scan_win_std_dev[1499]), .feature_accum(feature_accums[1499]));
  accum_calculator ac1500(.scan_win(scan_win1500), .rectangle1_x(rectangle1_xs[1500]), .rectangle1_y(rectangle1_ys[1500]), .rectangle1_width(rectangle1_widths[1500]), .rectangle1_height(rectangle1_heights[1500]), .rectangle1_weight(rectangle1_weights[1500]), .rectangle2_x(rectangle2_xs[1500]), .rectangle2_y(rectangle2_ys[1500]), .rectangle2_width(rectangle2_widths[1500]), .rectangle2_height(rectangle2_heights[1500]), .rectangle2_weight(rectangle2_weights[1500]), .rectangle3_x(rectangle3_xs[1500]), .rectangle3_y(rectangle3_ys[1500]), .rectangle3_width(rectangle3_widths[1500]), .rectangle3_height(rectangle3_heights[1500]), .rectangle3_weight(rectangle3_weights[1500]), .feature_threshold(feature_thresholds[1500]), .feature_above(feature_aboves[1500]), .feature_below(feature_belows[1500]), .scan_win_std_dev(scan_win_std_dev[1500]), .feature_accum(feature_accums[1500]));
  accum_calculator ac1501(.scan_win(scan_win1501), .rectangle1_x(rectangle1_xs[1501]), .rectangle1_y(rectangle1_ys[1501]), .rectangle1_width(rectangle1_widths[1501]), .rectangle1_height(rectangle1_heights[1501]), .rectangle1_weight(rectangle1_weights[1501]), .rectangle2_x(rectangle2_xs[1501]), .rectangle2_y(rectangle2_ys[1501]), .rectangle2_width(rectangle2_widths[1501]), .rectangle2_height(rectangle2_heights[1501]), .rectangle2_weight(rectangle2_weights[1501]), .rectangle3_x(rectangle3_xs[1501]), .rectangle3_y(rectangle3_ys[1501]), .rectangle3_width(rectangle3_widths[1501]), .rectangle3_height(rectangle3_heights[1501]), .rectangle3_weight(rectangle3_weights[1501]), .feature_threshold(feature_thresholds[1501]), .feature_above(feature_aboves[1501]), .feature_below(feature_belows[1501]), .scan_win_std_dev(scan_win_std_dev[1501]), .feature_accum(feature_accums[1501]));
  accum_calculator ac1502(.scan_win(scan_win1502), .rectangle1_x(rectangle1_xs[1502]), .rectangle1_y(rectangle1_ys[1502]), .rectangle1_width(rectangle1_widths[1502]), .rectangle1_height(rectangle1_heights[1502]), .rectangle1_weight(rectangle1_weights[1502]), .rectangle2_x(rectangle2_xs[1502]), .rectangle2_y(rectangle2_ys[1502]), .rectangle2_width(rectangle2_widths[1502]), .rectangle2_height(rectangle2_heights[1502]), .rectangle2_weight(rectangle2_weights[1502]), .rectangle3_x(rectangle3_xs[1502]), .rectangle3_y(rectangle3_ys[1502]), .rectangle3_width(rectangle3_widths[1502]), .rectangle3_height(rectangle3_heights[1502]), .rectangle3_weight(rectangle3_weights[1502]), .feature_threshold(feature_thresholds[1502]), .feature_above(feature_aboves[1502]), .feature_below(feature_belows[1502]), .scan_win_std_dev(scan_win_std_dev[1502]), .feature_accum(feature_accums[1502]));
  accum_calculator ac1503(.scan_win(scan_win1503), .rectangle1_x(rectangle1_xs[1503]), .rectangle1_y(rectangle1_ys[1503]), .rectangle1_width(rectangle1_widths[1503]), .rectangle1_height(rectangle1_heights[1503]), .rectangle1_weight(rectangle1_weights[1503]), .rectangle2_x(rectangle2_xs[1503]), .rectangle2_y(rectangle2_ys[1503]), .rectangle2_width(rectangle2_widths[1503]), .rectangle2_height(rectangle2_heights[1503]), .rectangle2_weight(rectangle2_weights[1503]), .rectangle3_x(rectangle3_xs[1503]), .rectangle3_y(rectangle3_ys[1503]), .rectangle3_width(rectangle3_widths[1503]), .rectangle3_height(rectangle3_heights[1503]), .rectangle3_weight(rectangle3_weights[1503]), .feature_threshold(feature_thresholds[1503]), .feature_above(feature_aboves[1503]), .feature_below(feature_belows[1503]), .scan_win_std_dev(scan_win_std_dev[1503]), .feature_accum(feature_accums[1503]));
  accum_calculator ac1504(.scan_win(scan_win1504), .rectangle1_x(rectangle1_xs[1504]), .rectangle1_y(rectangle1_ys[1504]), .rectangle1_width(rectangle1_widths[1504]), .rectangle1_height(rectangle1_heights[1504]), .rectangle1_weight(rectangle1_weights[1504]), .rectangle2_x(rectangle2_xs[1504]), .rectangle2_y(rectangle2_ys[1504]), .rectangle2_width(rectangle2_widths[1504]), .rectangle2_height(rectangle2_heights[1504]), .rectangle2_weight(rectangle2_weights[1504]), .rectangle3_x(rectangle3_xs[1504]), .rectangle3_y(rectangle3_ys[1504]), .rectangle3_width(rectangle3_widths[1504]), .rectangle3_height(rectangle3_heights[1504]), .rectangle3_weight(rectangle3_weights[1504]), .feature_threshold(feature_thresholds[1504]), .feature_above(feature_aboves[1504]), .feature_below(feature_belows[1504]), .scan_win_std_dev(scan_win_std_dev[1504]), .feature_accum(feature_accums[1504]));
  accum_calculator ac1505(.scan_win(scan_win1505), .rectangle1_x(rectangle1_xs[1505]), .rectangle1_y(rectangle1_ys[1505]), .rectangle1_width(rectangle1_widths[1505]), .rectangle1_height(rectangle1_heights[1505]), .rectangle1_weight(rectangle1_weights[1505]), .rectangle2_x(rectangle2_xs[1505]), .rectangle2_y(rectangle2_ys[1505]), .rectangle2_width(rectangle2_widths[1505]), .rectangle2_height(rectangle2_heights[1505]), .rectangle2_weight(rectangle2_weights[1505]), .rectangle3_x(rectangle3_xs[1505]), .rectangle3_y(rectangle3_ys[1505]), .rectangle3_width(rectangle3_widths[1505]), .rectangle3_height(rectangle3_heights[1505]), .rectangle3_weight(rectangle3_weights[1505]), .feature_threshold(feature_thresholds[1505]), .feature_above(feature_aboves[1505]), .feature_below(feature_belows[1505]), .scan_win_std_dev(scan_win_std_dev[1505]), .feature_accum(feature_accums[1505]));
  accum_calculator ac1506(.scan_win(scan_win1506), .rectangle1_x(rectangle1_xs[1506]), .rectangle1_y(rectangle1_ys[1506]), .rectangle1_width(rectangle1_widths[1506]), .rectangle1_height(rectangle1_heights[1506]), .rectangle1_weight(rectangle1_weights[1506]), .rectangle2_x(rectangle2_xs[1506]), .rectangle2_y(rectangle2_ys[1506]), .rectangle2_width(rectangle2_widths[1506]), .rectangle2_height(rectangle2_heights[1506]), .rectangle2_weight(rectangle2_weights[1506]), .rectangle3_x(rectangle3_xs[1506]), .rectangle3_y(rectangle3_ys[1506]), .rectangle3_width(rectangle3_widths[1506]), .rectangle3_height(rectangle3_heights[1506]), .rectangle3_weight(rectangle3_weights[1506]), .feature_threshold(feature_thresholds[1506]), .feature_above(feature_aboves[1506]), .feature_below(feature_belows[1506]), .scan_win_std_dev(scan_win_std_dev[1506]), .feature_accum(feature_accums[1506]));
  accum_calculator ac1507(.scan_win(scan_win1507), .rectangle1_x(rectangle1_xs[1507]), .rectangle1_y(rectangle1_ys[1507]), .rectangle1_width(rectangle1_widths[1507]), .rectangle1_height(rectangle1_heights[1507]), .rectangle1_weight(rectangle1_weights[1507]), .rectangle2_x(rectangle2_xs[1507]), .rectangle2_y(rectangle2_ys[1507]), .rectangle2_width(rectangle2_widths[1507]), .rectangle2_height(rectangle2_heights[1507]), .rectangle2_weight(rectangle2_weights[1507]), .rectangle3_x(rectangle3_xs[1507]), .rectangle3_y(rectangle3_ys[1507]), .rectangle3_width(rectangle3_widths[1507]), .rectangle3_height(rectangle3_heights[1507]), .rectangle3_weight(rectangle3_weights[1507]), .feature_threshold(feature_thresholds[1507]), .feature_above(feature_aboves[1507]), .feature_below(feature_belows[1507]), .scan_win_std_dev(scan_win_std_dev[1507]), .feature_accum(feature_accums[1507]));
  accum_calculator ac1508(.scan_win(scan_win1508), .rectangle1_x(rectangle1_xs[1508]), .rectangle1_y(rectangle1_ys[1508]), .rectangle1_width(rectangle1_widths[1508]), .rectangle1_height(rectangle1_heights[1508]), .rectangle1_weight(rectangle1_weights[1508]), .rectangle2_x(rectangle2_xs[1508]), .rectangle2_y(rectangle2_ys[1508]), .rectangle2_width(rectangle2_widths[1508]), .rectangle2_height(rectangle2_heights[1508]), .rectangle2_weight(rectangle2_weights[1508]), .rectangle3_x(rectangle3_xs[1508]), .rectangle3_y(rectangle3_ys[1508]), .rectangle3_width(rectangle3_widths[1508]), .rectangle3_height(rectangle3_heights[1508]), .rectangle3_weight(rectangle3_weights[1508]), .feature_threshold(feature_thresholds[1508]), .feature_above(feature_aboves[1508]), .feature_below(feature_belows[1508]), .scan_win_std_dev(scan_win_std_dev[1508]), .feature_accum(feature_accums[1508]));
  accum_calculator ac1509(.scan_win(scan_win1509), .rectangle1_x(rectangle1_xs[1509]), .rectangle1_y(rectangle1_ys[1509]), .rectangle1_width(rectangle1_widths[1509]), .rectangle1_height(rectangle1_heights[1509]), .rectangle1_weight(rectangle1_weights[1509]), .rectangle2_x(rectangle2_xs[1509]), .rectangle2_y(rectangle2_ys[1509]), .rectangle2_width(rectangle2_widths[1509]), .rectangle2_height(rectangle2_heights[1509]), .rectangle2_weight(rectangle2_weights[1509]), .rectangle3_x(rectangle3_xs[1509]), .rectangle3_y(rectangle3_ys[1509]), .rectangle3_width(rectangle3_widths[1509]), .rectangle3_height(rectangle3_heights[1509]), .rectangle3_weight(rectangle3_weights[1509]), .feature_threshold(feature_thresholds[1509]), .feature_above(feature_aboves[1509]), .feature_below(feature_belows[1509]), .scan_win_std_dev(scan_win_std_dev[1509]), .feature_accum(feature_accums[1509]));
  accum_calculator ac1510(.scan_win(scan_win1510), .rectangle1_x(rectangle1_xs[1510]), .rectangle1_y(rectangle1_ys[1510]), .rectangle1_width(rectangle1_widths[1510]), .rectangle1_height(rectangle1_heights[1510]), .rectangle1_weight(rectangle1_weights[1510]), .rectangle2_x(rectangle2_xs[1510]), .rectangle2_y(rectangle2_ys[1510]), .rectangle2_width(rectangle2_widths[1510]), .rectangle2_height(rectangle2_heights[1510]), .rectangle2_weight(rectangle2_weights[1510]), .rectangle3_x(rectangle3_xs[1510]), .rectangle3_y(rectangle3_ys[1510]), .rectangle3_width(rectangle3_widths[1510]), .rectangle3_height(rectangle3_heights[1510]), .rectangle3_weight(rectangle3_weights[1510]), .feature_threshold(feature_thresholds[1510]), .feature_above(feature_aboves[1510]), .feature_below(feature_belows[1510]), .scan_win_std_dev(scan_win_std_dev[1510]), .feature_accum(feature_accums[1510]));
  accum_calculator ac1511(.scan_win(scan_win1511), .rectangle1_x(rectangle1_xs[1511]), .rectangle1_y(rectangle1_ys[1511]), .rectangle1_width(rectangle1_widths[1511]), .rectangle1_height(rectangle1_heights[1511]), .rectangle1_weight(rectangle1_weights[1511]), .rectangle2_x(rectangle2_xs[1511]), .rectangle2_y(rectangle2_ys[1511]), .rectangle2_width(rectangle2_widths[1511]), .rectangle2_height(rectangle2_heights[1511]), .rectangle2_weight(rectangle2_weights[1511]), .rectangle3_x(rectangle3_xs[1511]), .rectangle3_y(rectangle3_ys[1511]), .rectangle3_width(rectangle3_widths[1511]), .rectangle3_height(rectangle3_heights[1511]), .rectangle3_weight(rectangle3_weights[1511]), .feature_threshold(feature_thresholds[1511]), .feature_above(feature_aboves[1511]), .feature_below(feature_belows[1511]), .scan_win_std_dev(scan_win_std_dev[1511]), .feature_accum(feature_accums[1511]));
  accum_calculator ac1512(.scan_win(scan_win1512), .rectangle1_x(rectangle1_xs[1512]), .rectangle1_y(rectangle1_ys[1512]), .rectangle1_width(rectangle1_widths[1512]), .rectangle1_height(rectangle1_heights[1512]), .rectangle1_weight(rectangle1_weights[1512]), .rectangle2_x(rectangle2_xs[1512]), .rectangle2_y(rectangle2_ys[1512]), .rectangle2_width(rectangle2_widths[1512]), .rectangle2_height(rectangle2_heights[1512]), .rectangle2_weight(rectangle2_weights[1512]), .rectangle3_x(rectangle3_xs[1512]), .rectangle3_y(rectangle3_ys[1512]), .rectangle3_width(rectangle3_widths[1512]), .rectangle3_height(rectangle3_heights[1512]), .rectangle3_weight(rectangle3_weights[1512]), .feature_threshold(feature_thresholds[1512]), .feature_above(feature_aboves[1512]), .feature_below(feature_belows[1512]), .scan_win_std_dev(scan_win_std_dev[1512]), .feature_accum(feature_accums[1512]));
  accum_calculator ac1513(.scan_win(scan_win1513), .rectangle1_x(rectangle1_xs[1513]), .rectangle1_y(rectangle1_ys[1513]), .rectangle1_width(rectangle1_widths[1513]), .rectangle1_height(rectangle1_heights[1513]), .rectangle1_weight(rectangle1_weights[1513]), .rectangle2_x(rectangle2_xs[1513]), .rectangle2_y(rectangle2_ys[1513]), .rectangle2_width(rectangle2_widths[1513]), .rectangle2_height(rectangle2_heights[1513]), .rectangle2_weight(rectangle2_weights[1513]), .rectangle3_x(rectangle3_xs[1513]), .rectangle3_y(rectangle3_ys[1513]), .rectangle3_width(rectangle3_widths[1513]), .rectangle3_height(rectangle3_heights[1513]), .rectangle3_weight(rectangle3_weights[1513]), .feature_threshold(feature_thresholds[1513]), .feature_above(feature_aboves[1513]), .feature_below(feature_belows[1513]), .scan_win_std_dev(scan_win_std_dev[1513]), .feature_accum(feature_accums[1513]));
  accum_calculator ac1514(.scan_win(scan_win1514), .rectangle1_x(rectangle1_xs[1514]), .rectangle1_y(rectangle1_ys[1514]), .rectangle1_width(rectangle1_widths[1514]), .rectangle1_height(rectangle1_heights[1514]), .rectangle1_weight(rectangle1_weights[1514]), .rectangle2_x(rectangle2_xs[1514]), .rectangle2_y(rectangle2_ys[1514]), .rectangle2_width(rectangle2_widths[1514]), .rectangle2_height(rectangle2_heights[1514]), .rectangle2_weight(rectangle2_weights[1514]), .rectangle3_x(rectangle3_xs[1514]), .rectangle3_y(rectangle3_ys[1514]), .rectangle3_width(rectangle3_widths[1514]), .rectangle3_height(rectangle3_heights[1514]), .rectangle3_weight(rectangle3_weights[1514]), .feature_threshold(feature_thresholds[1514]), .feature_above(feature_aboves[1514]), .feature_below(feature_belows[1514]), .scan_win_std_dev(scan_win_std_dev[1514]), .feature_accum(feature_accums[1514]));
  accum_calculator ac1515(.scan_win(scan_win1515), .rectangle1_x(rectangle1_xs[1515]), .rectangle1_y(rectangle1_ys[1515]), .rectangle1_width(rectangle1_widths[1515]), .rectangle1_height(rectangle1_heights[1515]), .rectangle1_weight(rectangle1_weights[1515]), .rectangle2_x(rectangle2_xs[1515]), .rectangle2_y(rectangle2_ys[1515]), .rectangle2_width(rectangle2_widths[1515]), .rectangle2_height(rectangle2_heights[1515]), .rectangle2_weight(rectangle2_weights[1515]), .rectangle3_x(rectangle3_xs[1515]), .rectangle3_y(rectangle3_ys[1515]), .rectangle3_width(rectangle3_widths[1515]), .rectangle3_height(rectangle3_heights[1515]), .rectangle3_weight(rectangle3_weights[1515]), .feature_threshold(feature_thresholds[1515]), .feature_above(feature_aboves[1515]), .feature_below(feature_belows[1515]), .scan_win_std_dev(scan_win_std_dev[1515]), .feature_accum(feature_accums[1515]));
  accum_calculator ac1516(.scan_win(scan_win1516), .rectangle1_x(rectangle1_xs[1516]), .rectangle1_y(rectangle1_ys[1516]), .rectangle1_width(rectangle1_widths[1516]), .rectangle1_height(rectangle1_heights[1516]), .rectangle1_weight(rectangle1_weights[1516]), .rectangle2_x(rectangle2_xs[1516]), .rectangle2_y(rectangle2_ys[1516]), .rectangle2_width(rectangle2_widths[1516]), .rectangle2_height(rectangle2_heights[1516]), .rectangle2_weight(rectangle2_weights[1516]), .rectangle3_x(rectangle3_xs[1516]), .rectangle3_y(rectangle3_ys[1516]), .rectangle3_width(rectangle3_widths[1516]), .rectangle3_height(rectangle3_heights[1516]), .rectangle3_weight(rectangle3_weights[1516]), .feature_threshold(feature_thresholds[1516]), .feature_above(feature_aboves[1516]), .feature_below(feature_belows[1516]), .scan_win_std_dev(scan_win_std_dev[1516]), .feature_accum(feature_accums[1516]));
  accum_calculator ac1517(.scan_win(scan_win1517), .rectangle1_x(rectangle1_xs[1517]), .rectangle1_y(rectangle1_ys[1517]), .rectangle1_width(rectangle1_widths[1517]), .rectangle1_height(rectangle1_heights[1517]), .rectangle1_weight(rectangle1_weights[1517]), .rectangle2_x(rectangle2_xs[1517]), .rectangle2_y(rectangle2_ys[1517]), .rectangle2_width(rectangle2_widths[1517]), .rectangle2_height(rectangle2_heights[1517]), .rectangle2_weight(rectangle2_weights[1517]), .rectangle3_x(rectangle3_xs[1517]), .rectangle3_y(rectangle3_ys[1517]), .rectangle3_width(rectangle3_widths[1517]), .rectangle3_height(rectangle3_heights[1517]), .rectangle3_weight(rectangle3_weights[1517]), .feature_threshold(feature_thresholds[1517]), .feature_above(feature_aboves[1517]), .feature_below(feature_belows[1517]), .scan_win_std_dev(scan_win_std_dev[1517]), .feature_accum(feature_accums[1517]));
  accum_calculator ac1518(.scan_win(scan_win1518), .rectangle1_x(rectangle1_xs[1518]), .rectangle1_y(rectangle1_ys[1518]), .rectangle1_width(rectangle1_widths[1518]), .rectangle1_height(rectangle1_heights[1518]), .rectangle1_weight(rectangle1_weights[1518]), .rectangle2_x(rectangle2_xs[1518]), .rectangle2_y(rectangle2_ys[1518]), .rectangle2_width(rectangle2_widths[1518]), .rectangle2_height(rectangle2_heights[1518]), .rectangle2_weight(rectangle2_weights[1518]), .rectangle3_x(rectangle3_xs[1518]), .rectangle3_y(rectangle3_ys[1518]), .rectangle3_width(rectangle3_widths[1518]), .rectangle3_height(rectangle3_heights[1518]), .rectangle3_weight(rectangle3_weights[1518]), .feature_threshold(feature_thresholds[1518]), .feature_above(feature_aboves[1518]), .feature_below(feature_belows[1518]), .scan_win_std_dev(scan_win_std_dev[1518]), .feature_accum(feature_accums[1518]));
  accum_calculator ac1519(.scan_win(scan_win1519), .rectangle1_x(rectangle1_xs[1519]), .rectangle1_y(rectangle1_ys[1519]), .rectangle1_width(rectangle1_widths[1519]), .rectangle1_height(rectangle1_heights[1519]), .rectangle1_weight(rectangle1_weights[1519]), .rectangle2_x(rectangle2_xs[1519]), .rectangle2_y(rectangle2_ys[1519]), .rectangle2_width(rectangle2_widths[1519]), .rectangle2_height(rectangle2_heights[1519]), .rectangle2_weight(rectangle2_weights[1519]), .rectangle3_x(rectangle3_xs[1519]), .rectangle3_y(rectangle3_ys[1519]), .rectangle3_width(rectangle3_widths[1519]), .rectangle3_height(rectangle3_heights[1519]), .rectangle3_weight(rectangle3_weights[1519]), .feature_threshold(feature_thresholds[1519]), .feature_above(feature_aboves[1519]), .feature_below(feature_belows[1519]), .scan_win_std_dev(scan_win_std_dev[1519]), .feature_accum(feature_accums[1519]));
  accum_calculator ac1520(.scan_win(scan_win1520), .rectangle1_x(rectangle1_xs[1520]), .rectangle1_y(rectangle1_ys[1520]), .rectangle1_width(rectangle1_widths[1520]), .rectangle1_height(rectangle1_heights[1520]), .rectangle1_weight(rectangle1_weights[1520]), .rectangle2_x(rectangle2_xs[1520]), .rectangle2_y(rectangle2_ys[1520]), .rectangle2_width(rectangle2_widths[1520]), .rectangle2_height(rectangle2_heights[1520]), .rectangle2_weight(rectangle2_weights[1520]), .rectangle3_x(rectangle3_xs[1520]), .rectangle3_y(rectangle3_ys[1520]), .rectangle3_width(rectangle3_widths[1520]), .rectangle3_height(rectangle3_heights[1520]), .rectangle3_weight(rectangle3_weights[1520]), .feature_threshold(feature_thresholds[1520]), .feature_above(feature_aboves[1520]), .feature_below(feature_belows[1520]), .scan_win_std_dev(scan_win_std_dev[1520]), .feature_accum(feature_accums[1520]));
  accum_calculator ac1521(.scan_win(scan_win1521), .rectangle1_x(rectangle1_xs[1521]), .rectangle1_y(rectangle1_ys[1521]), .rectangle1_width(rectangle1_widths[1521]), .rectangle1_height(rectangle1_heights[1521]), .rectangle1_weight(rectangle1_weights[1521]), .rectangle2_x(rectangle2_xs[1521]), .rectangle2_y(rectangle2_ys[1521]), .rectangle2_width(rectangle2_widths[1521]), .rectangle2_height(rectangle2_heights[1521]), .rectangle2_weight(rectangle2_weights[1521]), .rectangle3_x(rectangle3_xs[1521]), .rectangle3_y(rectangle3_ys[1521]), .rectangle3_width(rectangle3_widths[1521]), .rectangle3_height(rectangle3_heights[1521]), .rectangle3_weight(rectangle3_weights[1521]), .feature_threshold(feature_thresholds[1521]), .feature_above(feature_aboves[1521]), .feature_below(feature_belows[1521]), .scan_win_std_dev(scan_win_std_dev[1521]), .feature_accum(feature_accums[1521]));
  accum_calculator ac1522(.scan_win(scan_win1522), .rectangle1_x(rectangle1_xs[1522]), .rectangle1_y(rectangle1_ys[1522]), .rectangle1_width(rectangle1_widths[1522]), .rectangle1_height(rectangle1_heights[1522]), .rectangle1_weight(rectangle1_weights[1522]), .rectangle2_x(rectangle2_xs[1522]), .rectangle2_y(rectangle2_ys[1522]), .rectangle2_width(rectangle2_widths[1522]), .rectangle2_height(rectangle2_heights[1522]), .rectangle2_weight(rectangle2_weights[1522]), .rectangle3_x(rectangle3_xs[1522]), .rectangle3_y(rectangle3_ys[1522]), .rectangle3_width(rectangle3_widths[1522]), .rectangle3_height(rectangle3_heights[1522]), .rectangle3_weight(rectangle3_weights[1522]), .feature_threshold(feature_thresholds[1522]), .feature_above(feature_aboves[1522]), .feature_below(feature_belows[1522]), .scan_win_std_dev(scan_win_std_dev[1522]), .feature_accum(feature_accums[1522]));
  accum_calculator ac1523(.scan_win(scan_win1523), .rectangle1_x(rectangle1_xs[1523]), .rectangle1_y(rectangle1_ys[1523]), .rectangle1_width(rectangle1_widths[1523]), .rectangle1_height(rectangle1_heights[1523]), .rectangle1_weight(rectangle1_weights[1523]), .rectangle2_x(rectangle2_xs[1523]), .rectangle2_y(rectangle2_ys[1523]), .rectangle2_width(rectangle2_widths[1523]), .rectangle2_height(rectangle2_heights[1523]), .rectangle2_weight(rectangle2_weights[1523]), .rectangle3_x(rectangle3_xs[1523]), .rectangle3_y(rectangle3_ys[1523]), .rectangle3_width(rectangle3_widths[1523]), .rectangle3_height(rectangle3_heights[1523]), .rectangle3_weight(rectangle3_weights[1523]), .feature_threshold(feature_thresholds[1523]), .feature_above(feature_aboves[1523]), .feature_below(feature_belows[1523]), .scan_win_std_dev(scan_win_std_dev[1523]), .feature_accum(feature_accums[1523]));
  accum_calculator ac1524(.scan_win(scan_win1524), .rectangle1_x(rectangle1_xs[1524]), .rectangle1_y(rectangle1_ys[1524]), .rectangle1_width(rectangle1_widths[1524]), .rectangle1_height(rectangle1_heights[1524]), .rectangle1_weight(rectangle1_weights[1524]), .rectangle2_x(rectangle2_xs[1524]), .rectangle2_y(rectangle2_ys[1524]), .rectangle2_width(rectangle2_widths[1524]), .rectangle2_height(rectangle2_heights[1524]), .rectangle2_weight(rectangle2_weights[1524]), .rectangle3_x(rectangle3_xs[1524]), .rectangle3_y(rectangle3_ys[1524]), .rectangle3_width(rectangle3_widths[1524]), .rectangle3_height(rectangle3_heights[1524]), .rectangle3_weight(rectangle3_weights[1524]), .feature_threshold(feature_thresholds[1524]), .feature_above(feature_aboves[1524]), .feature_below(feature_belows[1524]), .scan_win_std_dev(scan_win_std_dev[1524]), .feature_accum(feature_accums[1524]));
  accum_calculator ac1525(.scan_win(scan_win1525), .rectangle1_x(rectangle1_xs[1525]), .rectangle1_y(rectangle1_ys[1525]), .rectangle1_width(rectangle1_widths[1525]), .rectangle1_height(rectangle1_heights[1525]), .rectangle1_weight(rectangle1_weights[1525]), .rectangle2_x(rectangle2_xs[1525]), .rectangle2_y(rectangle2_ys[1525]), .rectangle2_width(rectangle2_widths[1525]), .rectangle2_height(rectangle2_heights[1525]), .rectangle2_weight(rectangle2_weights[1525]), .rectangle3_x(rectangle3_xs[1525]), .rectangle3_y(rectangle3_ys[1525]), .rectangle3_width(rectangle3_widths[1525]), .rectangle3_height(rectangle3_heights[1525]), .rectangle3_weight(rectangle3_weights[1525]), .feature_threshold(feature_thresholds[1525]), .feature_above(feature_aboves[1525]), .feature_below(feature_belows[1525]), .scan_win_std_dev(scan_win_std_dev[1525]), .feature_accum(feature_accums[1525]));
  accum_calculator ac1526(.scan_win(scan_win1526), .rectangle1_x(rectangle1_xs[1526]), .rectangle1_y(rectangle1_ys[1526]), .rectangle1_width(rectangle1_widths[1526]), .rectangle1_height(rectangle1_heights[1526]), .rectangle1_weight(rectangle1_weights[1526]), .rectangle2_x(rectangle2_xs[1526]), .rectangle2_y(rectangle2_ys[1526]), .rectangle2_width(rectangle2_widths[1526]), .rectangle2_height(rectangle2_heights[1526]), .rectangle2_weight(rectangle2_weights[1526]), .rectangle3_x(rectangle3_xs[1526]), .rectangle3_y(rectangle3_ys[1526]), .rectangle3_width(rectangle3_widths[1526]), .rectangle3_height(rectangle3_heights[1526]), .rectangle3_weight(rectangle3_weights[1526]), .feature_threshold(feature_thresholds[1526]), .feature_above(feature_aboves[1526]), .feature_below(feature_belows[1526]), .scan_win_std_dev(scan_win_std_dev[1526]), .feature_accum(feature_accums[1526]));
  accum_calculator ac1527(.scan_win(scan_win1527), .rectangle1_x(rectangle1_xs[1527]), .rectangle1_y(rectangle1_ys[1527]), .rectangle1_width(rectangle1_widths[1527]), .rectangle1_height(rectangle1_heights[1527]), .rectangle1_weight(rectangle1_weights[1527]), .rectangle2_x(rectangle2_xs[1527]), .rectangle2_y(rectangle2_ys[1527]), .rectangle2_width(rectangle2_widths[1527]), .rectangle2_height(rectangle2_heights[1527]), .rectangle2_weight(rectangle2_weights[1527]), .rectangle3_x(rectangle3_xs[1527]), .rectangle3_y(rectangle3_ys[1527]), .rectangle3_width(rectangle3_widths[1527]), .rectangle3_height(rectangle3_heights[1527]), .rectangle3_weight(rectangle3_weights[1527]), .feature_threshold(feature_thresholds[1527]), .feature_above(feature_aboves[1527]), .feature_below(feature_belows[1527]), .scan_win_std_dev(scan_win_std_dev[1527]), .feature_accum(feature_accums[1527]));
  accum_calculator ac1528(.scan_win(scan_win1528), .rectangle1_x(rectangle1_xs[1528]), .rectangle1_y(rectangle1_ys[1528]), .rectangle1_width(rectangle1_widths[1528]), .rectangle1_height(rectangle1_heights[1528]), .rectangle1_weight(rectangle1_weights[1528]), .rectangle2_x(rectangle2_xs[1528]), .rectangle2_y(rectangle2_ys[1528]), .rectangle2_width(rectangle2_widths[1528]), .rectangle2_height(rectangle2_heights[1528]), .rectangle2_weight(rectangle2_weights[1528]), .rectangle3_x(rectangle3_xs[1528]), .rectangle3_y(rectangle3_ys[1528]), .rectangle3_width(rectangle3_widths[1528]), .rectangle3_height(rectangle3_heights[1528]), .rectangle3_weight(rectangle3_weights[1528]), .feature_threshold(feature_thresholds[1528]), .feature_above(feature_aboves[1528]), .feature_below(feature_belows[1528]), .scan_win_std_dev(scan_win_std_dev[1528]), .feature_accum(feature_accums[1528]));
  accum_calculator ac1529(.scan_win(scan_win1529), .rectangle1_x(rectangle1_xs[1529]), .rectangle1_y(rectangle1_ys[1529]), .rectangle1_width(rectangle1_widths[1529]), .rectangle1_height(rectangle1_heights[1529]), .rectangle1_weight(rectangle1_weights[1529]), .rectangle2_x(rectangle2_xs[1529]), .rectangle2_y(rectangle2_ys[1529]), .rectangle2_width(rectangle2_widths[1529]), .rectangle2_height(rectangle2_heights[1529]), .rectangle2_weight(rectangle2_weights[1529]), .rectangle3_x(rectangle3_xs[1529]), .rectangle3_y(rectangle3_ys[1529]), .rectangle3_width(rectangle3_widths[1529]), .rectangle3_height(rectangle3_heights[1529]), .rectangle3_weight(rectangle3_weights[1529]), .feature_threshold(feature_thresholds[1529]), .feature_above(feature_aboves[1529]), .feature_below(feature_belows[1529]), .scan_win_std_dev(scan_win_std_dev[1529]), .feature_accum(feature_accums[1529]));
  accum_calculator ac1530(.scan_win(scan_win1530), .rectangle1_x(rectangle1_xs[1530]), .rectangle1_y(rectangle1_ys[1530]), .rectangle1_width(rectangle1_widths[1530]), .rectangle1_height(rectangle1_heights[1530]), .rectangle1_weight(rectangle1_weights[1530]), .rectangle2_x(rectangle2_xs[1530]), .rectangle2_y(rectangle2_ys[1530]), .rectangle2_width(rectangle2_widths[1530]), .rectangle2_height(rectangle2_heights[1530]), .rectangle2_weight(rectangle2_weights[1530]), .rectangle3_x(rectangle3_xs[1530]), .rectangle3_y(rectangle3_ys[1530]), .rectangle3_width(rectangle3_widths[1530]), .rectangle3_height(rectangle3_heights[1530]), .rectangle3_weight(rectangle3_weights[1530]), .feature_threshold(feature_thresholds[1530]), .feature_above(feature_aboves[1530]), .feature_below(feature_belows[1530]), .scan_win_std_dev(scan_win_std_dev[1530]), .feature_accum(feature_accums[1530]));
  accum_calculator ac1531(.scan_win(scan_win1531), .rectangle1_x(rectangle1_xs[1531]), .rectangle1_y(rectangle1_ys[1531]), .rectangle1_width(rectangle1_widths[1531]), .rectangle1_height(rectangle1_heights[1531]), .rectangle1_weight(rectangle1_weights[1531]), .rectangle2_x(rectangle2_xs[1531]), .rectangle2_y(rectangle2_ys[1531]), .rectangle2_width(rectangle2_widths[1531]), .rectangle2_height(rectangle2_heights[1531]), .rectangle2_weight(rectangle2_weights[1531]), .rectangle3_x(rectangle3_xs[1531]), .rectangle3_y(rectangle3_ys[1531]), .rectangle3_width(rectangle3_widths[1531]), .rectangle3_height(rectangle3_heights[1531]), .rectangle3_weight(rectangle3_weights[1531]), .feature_threshold(feature_thresholds[1531]), .feature_above(feature_aboves[1531]), .feature_below(feature_belows[1531]), .scan_win_std_dev(scan_win_std_dev[1531]), .feature_accum(feature_accums[1531]));
  accum_calculator ac1532(.scan_win(scan_win1532), .rectangle1_x(rectangle1_xs[1532]), .rectangle1_y(rectangle1_ys[1532]), .rectangle1_width(rectangle1_widths[1532]), .rectangle1_height(rectangle1_heights[1532]), .rectangle1_weight(rectangle1_weights[1532]), .rectangle2_x(rectangle2_xs[1532]), .rectangle2_y(rectangle2_ys[1532]), .rectangle2_width(rectangle2_widths[1532]), .rectangle2_height(rectangle2_heights[1532]), .rectangle2_weight(rectangle2_weights[1532]), .rectangle3_x(rectangle3_xs[1532]), .rectangle3_y(rectangle3_ys[1532]), .rectangle3_width(rectangle3_widths[1532]), .rectangle3_height(rectangle3_heights[1532]), .rectangle3_weight(rectangle3_weights[1532]), .feature_threshold(feature_thresholds[1532]), .feature_above(feature_aboves[1532]), .feature_below(feature_belows[1532]), .scan_win_std_dev(scan_win_std_dev[1532]), .feature_accum(feature_accums[1532]));
  accum_calculator ac1533(.scan_win(scan_win1533), .rectangle1_x(rectangle1_xs[1533]), .rectangle1_y(rectangle1_ys[1533]), .rectangle1_width(rectangle1_widths[1533]), .rectangle1_height(rectangle1_heights[1533]), .rectangle1_weight(rectangle1_weights[1533]), .rectangle2_x(rectangle2_xs[1533]), .rectangle2_y(rectangle2_ys[1533]), .rectangle2_width(rectangle2_widths[1533]), .rectangle2_height(rectangle2_heights[1533]), .rectangle2_weight(rectangle2_weights[1533]), .rectangle3_x(rectangle3_xs[1533]), .rectangle3_y(rectangle3_ys[1533]), .rectangle3_width(rectangle3_widths[1533]), .rectangle3_height(rectangle3_heights[1533]), .rectangle3_weight(rectangle3_weights[1533]), .feature_threshold(feature_thresholds[1533]), .feature_above(feature_aboves[1533]), .feature_below(feature_belows[1533]), .scan_win_std_dev(scan_win_std_dev[1533]), .feature_accum(feature_accums[1533]));
  accum_calculator ac1534(.scan_win(scan_win1534), .rectangle1_x(rectangle1_xs[1534]), .rectangle1_y(rectangle1_ys[1534]), .rectangle1_width(rectangle1_widths[1534]), .rectangle1_height(rectangle1_heights[1534]), .rectangle1_weight(rectangle1_weights[1534]), .rectangle2_x(rectangle2_xs[1534]), .rectangle2_y(rectangle2_ys[1534]), .rectangle2_width(rectangle2_widths[1534]), .rectangle2_height(rectangle2_heights[1534]), .rectangle2_weight(rectangle2_weights[1534]), .rectangle3_x(rectangle3_xs[1534]), .rectangle3_y(rectangle3_ys[1534]), .rectangle3_width(rectangle3_widths[1534]), .rectangle3_height(rectangle3_heights[1534]), .rectangle3_weight(rectangle3_weights[1534]), .feature_threshold(feature_thresholds[1534]), .feature_above(feature_aboves[1534]), .feature_below(feature_belows[1534]), .scan_win_std_dev(scan_win_std_dev[1534]), .feature_accum(feature_accums[1534]));
  accum_calculator ac1535(.scan_win(scan_win1535), .rectangle1_x(rectangle1_xs[1535]), .rectangle1_y(rectangle1_ys[1535]), .rectangle1_width(rectangle1_widths[1535]), .rectangle1_height(rectangle1_heights[1535]), .rectangle1_weight(rectangle1_weights[1535]), .rectangle2_x(rectangle2_xs[1535]), .rectangle2_y(rectangle2_ys[1535]), .rectangle2_width(rectangle2_widths[1535]), .rectangle2_height(rectangle2_heights[1535]), .rectangle2_weight(rectangle2_weights[1535]), .rectangle3_x(rectangle3_xs[1535]), .rectangle3_y(rectangle3_ys[1535]), .rectangle3_width(rectangle3_widths[1535]), .rectangle3_height(rectangle3_heights[1535]), .rectangle3_weight(rectangle3_weights[1535]), .feature_threshold(feature_thresholds[1535]), .feature_above(feature_aboves[1535]), .feature_below(feature_belows[1535]), .scan_win_std_dev(scan_win_std_dev[1535]), .feature_accum(feature_accums[1535]));
  accum_calculator ac1536(.scan_win(scan_win1536), .rectangle1_x(rectangle1_xs[1536]), .rectangle1_y(rectangle1_ys[1536]), .rectangle1_width(rectangle1_widths[1536]), .rectangle1_height(rectangle1_heights[1536]), .rectangle1_weight(rectangle1_weights[1536]), .rectangle2_x(rectangle2_xs[1536]), .rectangle2_y(rectangle2_ys[1536]), .rectangle2_width(rectangle2_widths[1536]), .rectangle2_height(rectangle2_heights[1536]), .rectangle2_weight(rectangle2_weights[1536]), .rectangle3_x(rectangle3_xs[1536]), .rectangle3_y(rectangle3_ys[1536]), .rectangle3_width(rectangle3_widths[1536]), .rectangle3_height(rectangle3_heights[1536]), .rectangle3_weight(rectangle3_weights[1536]), .feature_threshold(feature_thresholds[1536]), .feature_above(feature_aboves[1536]), .feature_below(feature_belows[1536]), .scan_win_std_dev(scan_win_std_dev[1536]), .feature_accum(feature_accums[1536]));
  accum_calculator ac1537(.scan_win(scan_win1537), .rectangle1_x(rectangle1_xs[1537]), .rectangle1_y(rectangle1_ys[1537]), .rectangle1_width(rectangle1_widths[1537]), .rectangle1_height(rectangle1_heights[1537]), .rectangle1_weight(rectangle1_weights[1537]), .rectangle2_x(rectangle2_xs[1537]), .rectangle2_y(rectangle2_ys[1537]), .rectangle2_width(rectangle2_widths[1537]), .rectangle2_height(rectangle2_heights[1537]), .rectangle2_weight(rectangle2_weights[1537]), .rectangle3_x(rectangle3_xs[1537]), .rectangle3_y(rectangle3_ys[1537]), .rectangle3_width(rectangle3_widths[1537]), .rectangle3_height(rectangle3_heights[1537]), .rectangle3_weight(rectangle3_weights[1537]), .feature_threshold(feature_thresholds[1537]), .feature_above(feature_aboves[1537]), .feature_below(feature_belows[1537]), .scan_win_std_dev(scan_win_std_dev[1537]), .feature_accum(feature_accums[1537]));
  accum_calculator ac1538(.scan_win(scan_win1538), .rectangle1_x(rectangle1_xs[1538]), .rectangle1_y(rectangle1_ys[1538]), .rectangle1_width(rectangle1_widths[1538]), .rectangle1_height(rectangle1_heights[1538]), .rectangle1_weight(rectangle1_weights[1538]), .rectangle2_x(rectangle2_xs[1538]), .rectangle2_y(rectangle2_ys[1538]), .rectangle2_width(rectangle2_widths[1538]), .rectangle2_height(rectangle2_heights[1538]), .rectangle2_weight(rectangle2_weights[1538]), .rectangle3_x(rectangle3_xs[1538]), .rectangle3_y(rectangle3_ys[1538]), .rectangle3_width(rectangle3_widths[1538]), .rectangle3_height(rectangle3_heights[1538]), .rectangle3_weight(rectangle3_weights[1538]), .feature_threshold(feature_thresholds[1538]), .feature_above(feature_aboves[1538]), .feature_below(feature_belows[1538]), .scan_win_std_dev(scan_win_std_dev[1538]), .feature_accum(feature_accums[1538]));
  accum_calculator ac1539(.scan_win(scan_win1539), .rectangle1_x(rectangle1_xs[1539]), .rectangle1_y(rectangle1_ys[1539]), .rectangle1_width(rectangle1_widths[1539]), .rectangle1_height(rectangle1_heights[1539]), .rectangle1_weight(rectangle1_weights[1539]), .rectangle2_x(rectangle2_xs[1539]), .rectangle2_y(rectangle2_ys[1539]), .rectangle2_width(rectangle2_widths[1539]), .rectangle2_height(rectangle2_heights[1539]), .rectangle2_weight(rectangle2_weights[1539]), .rectangle3_x(rectangle3_xs[1539]), .rectangle3_y(rectangle3_ys[1539]), .rectangle3_width(rectangle3_widths[1539]), .rectangle3_height(rectangle3_heights[1539]), .rectangle3_weight(rectangle3_weights[1539]), .feature_threshold(feature_thresholds[1539]), .feature_above(feature_aboves[1539]), .feature_below(feature_belows[1539]), .scan_win_std_dev(scan_win_std_dev[1539]), .feature_accum(feature_accums[1539]));
  accum_calculator ac1540(.scan_win(scan_win1540), .rectangle1_x(rectangle1_xs[1540]), .rectangle1_y(rectangle1_ys[1540]), .rectangle1_width(rectangle1_widths[1540]), .rectangle1_height(rectangle1_heights[1540]), .rectangle1_weight(rectangle1_weights[1540]), .rectangle2_x(rectangle2_xs[1540]), .rectangle2_y(rectangle2_ys[1540]), .rectangle2_width(rectangle2_widths[1540]), .rectangle2_height(rectangle2_heights[1540]), .rectangle2_weight(rectangle2_weights[1540]), .rectangle3_x(rectangle3_xs[1540]), .rectangle3_y(rectangle3_ys[1540]), .rectangle3_width(rectangle3_widths[1540]), .rectangle3_height(rectangle3_heights[1540]), .rectangle3_weight(rectangle3_weights[1540]), .feature_threshold(feature_thresholds[1540]), .feature_above(feature_aboves[1540]), .feature_below(feature_belows[1540]), .scan_win_std_dev(scan_win_std_dev[1540]), .feature_accum(feature_accums[1540]));
  accum_calculator ac1541(.scan_win(scan_win1541), .rectangle1_x(rectangle1_xs[1541]), .rectangle1_y(rectangle1_ys[1541]), .rectangle1_width(rectangle1_widths[1541]), .rectangle1_height(rectangle1_heights[1541]), .rectangle1_weight(rectangle1_weights[1541]), .rectangle2_x(rectangle2_xs[1541]), .rectangle2_y(rectangle2_ys[1541]), .rectangle2_width(rectangle2_widths[1541]), .rectangle2_height(rectangle2_heights[1541]), .rectangle2_weight(rectangle2_weights[1541]), .rectangle3_x(rectangle3_xs[1541]), .rectangle3_y(rectangle3_ys[1541]), .rectangle3_width(rectangle3_widths[1541]), .rectangle3_height(rectangle3_heights[1541]), .rectangle3_weight(rectangle3_weights[1541]), .feature_threshold(feature_thresholds[1541]), .feature_above(feature_aboves[1541]), .feature_below(feature_belows[1541]), .scan_win_std_dev(scan_win_std_dev[1541]), .feature_accum(feature_accums[1541]));
  accum_calculator ac1542(.scan_win(scan_win1542), .rectangle1_x(rectangle1_xs[1542]), .rectangle1_y(rectangle1_ys[1542]), .rectangle1_width(rectangle1_widths[1542]), .rectangle1_height(rectangle1_heights[1542]), .rectangle1_weight(rectangle1_weights[1542]), .rectangle2_x(rectangle2_xs[1542]), .rectangle2_y(rectangle2_ys[1542]), .rectangle2_width(rectangle2_widths[1542]), .rectangle2_height(rectangle2_heights[1542]), .rectangle2_weight(rectangle2_weights[1542]), .rectangle3_x(rectangle3_xs[1542]), .rectangle3_y(rectangle3_ys[1542]), .rectangle3_width(rectangle3_widths[1542]), .rectangle3_height(rectangle3_heights[1542]), .rectangle3_weight(rectangle3_weights[1542]), .feature_threshold(feature_thresholds[1542]), .feature_above(feature_aboves[1542]), .feature_below(feature_belows[1542]), .scan_win_std_dev(scan_win_std_dev[1542]), .feature_accum(feature_accums[1542]));
  accum_calculator ac1543(.scan_win(scan_win1543), .rectangle1_x(rectangle1_xs[1543]), .rectangle1_y(rectangle1_ys[1543]), .rectangle1_width(rectangle1_widths[1543]), .rectangle1_height(rectangle1_heights[1543]), .rectangle1_weight(rectangle1_weights[1543]), .rectangle2_x(rectangle2_xs[1543]), .rectangle2_y(rectangle2_ys[1543]), .rectangle2_width(rectangle2_widths[1543]), .rectangle2_height(rectangle2_heights[1543]), .rectangle2_weight(rectangle2_weights[1543]), .rectangle3_x(rectangle3_xs[1543]), .rectangle3_y(rectangle3_ys[1543]), .rectangle3_width(rectangle3_widths[1543]), .rectangle3_height(rectangle3_heights[1543]), .rectangle3_weight(rectangle3_weights[1543]), .feature_threshold(feature_thresholds[1543]), .feature_above(feature_aboves[1543]), .feature_below(feature_belows[1543]), .scan_win_std_dev(scan_win_std_dev[1543]), .feature_accum(feature_accums[1543]));
  accum_calculator ac1544(.scan_win(scan_win1544), .rectangle1_x(rectangle1_xs[1544]), .rectangle1_y(rectangle1_ys[1544]), .rectangle1_width(rectangle1_widths[1544]), .rectangle1_height(rectangle1_heights[1544]), .rectangle1_weight(rectangle1_weights[1544]), .rectangle2_x(rectangle2_xs[1544]), .rectangle2_y(rectangle2_ys[1544]), .rectangle2_width(rectangle2_widths[1544]), .rectangle2_height(rectangle2_heights[1544]), .rectangle2_weight(rectangle2_weights[1544]), .rectangle3_x(rectangle3_xs[1544]), .rectangle3_y(rectangle3_ys[1544]), .rectangle3_width(rectangle3_widths[1544]), .rectangle3_height(rectangle3_heights[1544]), .rectangle3_weight(rectangle3_weights[1544]), .feature_threshold(feature_thresholds[1544]), .feature_above(feature_aboves[1544]), .feature_below(feature_belows[1544]), .scan_win_std_dev(scan_win_std_dev[1544]), .feature_accum(feature_accums[1544]));
  accum_calculator ac1545(.scan_win(scan_win1545), .rectangle1_x(rectangle1_xs[1545]), .rectangle1_y(rectangle1_ys[1545]), .rectangle1_width(rectangle1_widths[1545]), .rectangle1_height(rectangle1_heights[1545]), .rectangle1_weight(rectangle1_weights[1545]), .rectangle2_x(rectangle2_xs[1545]), .rectangle2_y(rectangle2_ys[1545]), .rectangle2_width(rectangle2_widths[1545]), .rectangle2_height(rectangle2_heights[1545]), .rectangle2_weight(rectangle2_weights[1545]), .rectangle3_x(rectangle3_xs[1545]), .rectangle3_y(rectangle3_ys[1545]), .rectangle3_width(rectangle3_widths[1545]), .rectangle3_height(rectangle3_heights[1545]), .rectangle3_weight(rectangle3_weights[1545]), .feature_threshold(feature_thresholds[1545]), .feature_above(feature_aboves[1545]), .feature_below(feature_belows[1545]), .scan_win_std_dev(scan_win_std_dev[1545]), .feature_accum(feature_accums[1545]));
  accum_calculator ac1546(.scan_win(scan_win1546), .rectangle1_x(rectangle1_xs[1546]), .rectangle1_y(rectangle1_ys[1546]), .rectangle1_width(rectangle1_widths[1546]), .rectangle1_height(rectangle1_heights[1546]), .rectangle1_weight(rectangle1_weights[1546]), .rectangle2_x(rectangle2_xs[1546]), .rectangle2_y(rectangle2_ys[1546]), .rectangle2_width(rectangle2_widths[1546]), .rectangle2_height(rectangle2_heights[1546]), .rectangle2_weight(rectangle2_weights[1546]), .rectangle3_x(rectangle3_xs[1546]), .rectangle3_y(rectangle3_ys[1546]), .rectangle3_width(rectangle3_widths[1546]), .rectangle3_height(rectangle3_heights[1546]), .rectangle3_weight(rectangle3_weights[1546]), .feature_threshold(feature_thresholds[1546]), .feature_above(feature_aboves[1546]), .feature_below(feature_belows[1546]), .scan_win_std_dev(scan_win_std_dev[1546]), .feature_accum(feature_accums[1546]));
  accum_calculator ac1547(.scan_win(scan_win1547), .rectangle1_x(rectangle1_xs[1547]), .rectangle1_y(rectangle1_ys[1547]), .rectangle1_width(rectangle1_widths[1547]), .rectangle1_height(rectangle1_heights[1547]), .rectangle1_weight(rectangle1_weights[1547]), .rectangle2_x(rectangle2_xs[1547]), .rectangle2_y(rectangle2_ys[1547]), .rectangle2_width(rectangle2_widths[1547]), .rectangle2_height(rectangle2_heights[1547]), .rectangle2_weight(rectangle2_weights[1547]), .rectangle3_x(rectangle3_xs[1547]), .rectangle3_y(rectangle3_ys[1547]), .rectangle3_width(rectangle3_widths[1547]), .rectangle3_height(rectangle3_heights[1547]), .rectangle3_weight(rectangle3_weights[1547]), .feature_threshold(feature_thresholds[1547]), .feature_above(feature_aboves[1547]), .feature_below(feature_belows[1547]), .scan_win_std_dev(scan_win_std_dev[1547]), .feature_accum(feature_accums[1547]));
  accum_calculator ac1548(.scan_win(scan_win1548), .rectangle1_x(rectangle1_xs[1548]), .rectangle1_y(rectangle1_ys[1548]), .rectangle1_width(rectangle1_widths[1548]), .rectangle1_height(rectangle1_heights[1548]), .rectangle1_weight(rectangle1_weights[1548]), .rectangle2_x(rectangle2_xs[1548]), .rectangle2_y(rectangle2_ys[1548]), .rectangle2_width(rectangle2_widths[1548]), .rectangle2_height(rectangle2_heights[1548]), .rectangle2_weight(rectangle2_weights[1548]), .rectangle3_x(rectangle3_xs[1548]), .rectangle3_y(rectangle3_ys[1548]), .rectangle3_width(rectangle3_widths[1548]), .rectangle3_height(rectangle3_heights[1548]), .rectangle3_weight(rectangle3_weights[1548]), .feature_threshold(feature_thresholds[1548]), .feature_above(feature_aboves[1548]), .feature_below(feature_belows[1548]), .scan_win_std_dev(scan_win_std_dev[1548]), .feature_accum(feature_accums[1548]));
  accum_calculator ac1549(.scan_win(scan_win1549), .rectangle1_x(rectangle1_xs[1549]), .rectangle1_y(rectangle1_ys[1549]), .rectangle1_width(rectangle1_widths[1549]), .rectangle1_height(rectangle1_heights[1549]), .rectangle1_weight(rectangle1_weights[1549]), .rectangle2_x(rectangle2_xs[1549]), .rectangle2_y(rectangle2_ys[1549]), .rectangle2_width(rectangle2_widths[1549]), .rectangle2_height(rectangle2_heights[1549]), .rectangle2_weight(rectangle2_weights[1549]), .rectangle3_x(rectangle3_xs[1549]), .rectangle3_y(rectangle3_ys[1549]), .rectangle3_width(rectangle3_widths[1549]), .rectangle3_height(rectangle3_heights[1549]), .rectangle3_weight(rectangle3_weights[1549]), .feature_threshold(feature_thresholds[1549]), .feature_above(feature_aboves[1549]), .feature_below(feature_belows[1549]), .scan_win_std_dev(scan_win_std_dev[1549]), .feature_accum(feature_accums[1549]));
  accum_calculator ac1550(.scan_win(scan_win1550), .rectangle1_x(rectangle1_xs[1550]), .rectangle1_y(rectangle1_ys[1550]), .rectangle1_width(rectangle1_widths[1550]), .rectangle1_height(rectangle1_heights[1550]), .rectangle1_weight(rectangle1_weights[1550]), .rectangle2_x(rectangle2_xs[1550]), .rectangle2_y(rectangle2_ys[1550]), .rectangle2_width(rectangle2_widths[1550]), .rectangle2_height(rectangle2_heights[1550]), .rectangle2_weight(rectangle2_weights[1550]), .rectangle3_x(rectangle3_xs[1550]), .rectangle3_y(rectangle3_ys[1550]), .rectangle3_width(rectangle3_widths[1550]), .rectangle3_height(rectangle3_heights[1550]), .rectangle3_weight(rectangle3_weights[1550]), .feature_threshold(feature_thresholds[1550]), .feature_above(feature_aboves[1550]), .feature_below(feature_belows[1550]), .scan_win_std_dev(scan_win_std_dev[1550]), .feature_accum(feature_accums[1550]));
  accum_calculator ac1551(.scan_win(scan_win1551), .rectangle1_x(rectangle1_xs[1551]), .rectangle1_y(rectangle1_ys[1551]), .rectangle1_width(rectangle1_widths[1551]), .rectangle1_height(rectangle1_heights[1551]), .rectangle1_weight(rectangle1_weights[1551]), .rectangle2_x(rectangle2_xs[1551]), .rectangle2_y(rectangle2_ys[1551]), .rectangle2_width(rectangle2_widths[1551]), .rectangle2_height(rectangle2_heights[1551]), .rectangle2_weight(rectangle2_weights[1551]), .rectangle3_x(rectangle3_xs[1551]), .rectangle3_y(rectangle3_ys[1551]), .rectangle3_width(rectangle3_widths[1551]), .rectangle3_height(rectangle3_heights[1551]), .rectangle3_weight(rectangle3_weights[1551]), .feature_threshold(feature_thresholds[1551]), .feature_above(feature_aboves[1551]), .feature_below(feature_belows[1551]), .scan_win_std_dev(scan_win_std_dev[1551]), .feature_accum(feature_accums[1551]));
  accum_calculator ac1552(.scan_win(scan_win1552), .rectangle1_x(rectangle1_xs[1552]), .rectangle1_y(rectangle1_ys[1552]), .rectangle1_width(rectangle1_widths[1552]), .rectangle1_height(rectangle1_heights[1552]), .rectangle1_weight(rectangle1_weights[1552]), .rectangle2_x(rectangle2_xs[1552]), .rectangle2_y(rectangle2_ys[1552]), .rectangle2_width(rectangle2_widths[1552]), .rectangle2_height(rectangle2_heights[1552]), .rectangle2_weight(rectangle2_weights[1552]), .rectangle3_x(rectangle3_xs[1552]), .rectangle3_y(rectangle3_ys[1552]), .rectangle3_width(rectangle3_widths[1552]), .rectangle3_height(rectangle3_heights[1552]), .rectangle3_weight(rectangle3_weights[1552]), .feature_threshold(feature_thresholds[1552]), .feature_above(feature_aboves[1552]), .feature_below(feature_belows[1552]), .scan_win_std_dev(scan_win_std_dev[1552]), .feature_accum(feature_accums[1552]));
  accum_calculator ac1553(.scan_win(scan_win1553), .rectangle1_x(rectangle1_xs[1553]), .rectangle1_y(rectangle1_ys[1553]), .rectangle1_width(rectangle1_widths[1553]), .rectangle1_height(rectangle1_heights[1553]), .rectangle1_weight(rectangle1_weights[1553]), .rectangle2_x(rectangle2_xs[1553]), .rectangle2_y(rectangle2_ys[1553]), .rectangle2_width(rectangle2_widths[1553]), .rectangle2_height(rectangle2_heights[1553]), .rectangle2_weight(rectangle2_weights[1553]), .rectangle3_x(rectangle3_xs[1553]), .rectangle3_y(rectangle3_ys[1553]), .rectangle3_width(rectangle3_widths[1553]), .rectangle3_height(rectangle3_heights[1553]), .rectangle3_weight(rectangle3_weights[1553]), .feature_threshold(feature_thresholds[1553]), .feature_above(feature_aboves[1553]), .feature_below(feature_belows[1553]), .scan_win_std_dev(scan_win_std_dev[1553]), .feature_accum(feature_accums[1553]));
  accum_calculator ac1554(.scan_win(scan_win1554), .rectangle1_x(rectangle1_xs[1554]), .rectangle1_y(rectangle1_ys[1554]), .rectangle1_width(rectangle1_widths[1554]), .rectangle1_height(rectangle1_heights[1554]), .rectangle1_weight(rectangle1_weights[1554]), .rectangle2_x(rectangle2_xs[1554]), .rectangle2_y(rectangle2_ys[1554]), .rectangle2_width(rectangle2_widths[1554]), .rectangle2_height(rectangle2_heights[1554]), .rectangle2_weight(rectangle2_weights[1554]), .rectangle3_x(rectangle3_xs[1554]), .rectangle3_y(rectangle3_ys[1554]), .rectangle3_width(rectangle3_widths[1554]), .rectangle3_height(rectangle3_heights[1554]), .rectangle3_weight(rectangle3_weights[1554]), .feature_threshold(feature_thresholds[1554]), .feature_above(feature_aboves[1554]), .feature_below(feature_belows[1554]), .scan_win_std_dev(scan_win_std_dev[1554]), .feature_accum(feature_accums[1554]));
  accum_calculator ac1555(.scan_win(scan_win1555), .rectangle1_x(rectangle1_xs[1555]), .rectangle1_y(rectangle1_ys[1555]), .rectangle1_width(rectangle1_widths[1555]), .rectangle1_height(rectangle1_heights[1555]), .rectangle1_weight(rectangle1_weights[1555]), .rectangle2_x(rectangle2_xs[1555]), .rectangle2_y(rectangle2_ys[1555]), .rectangle2_width(rectangle2_widths[1555]), .rectangle2_height(rectangle2_heights[1555]), .rectangle2_weight(rectangle2_weights[1555]), .rectangle3_x(rectangle3_xs[1555]), .rectangle3_y(rectangle3_ys[1555]), .rectangle3_width(rectangle3_widths[1555]), .rectangle3_height(rectangle3_heights[1555]), .rectangle3_weight(rectangle3_weights[1555]), .feature_threshold(feature_thresholds[1555]), .feature_above(feature_aboves[1555]), .feature_below(feature_belows[1555]), .scan_win_std_dev(scan_win_std_dev[1555]), .feature_accum(feature_accums[1555]));
  accum_calculator ac1556(.scan_win(scan_win1556), .rectangle1_x(rectangle1_xs[1556]), .rectangle1_y(rectangle1_ys[1556]), .rectangle1_width(rectangle1_widths[1556]), .rectangle1_height(rectangle1_heights[1556]), .rectangle1_weight(rectangle1_weights[1556]), .rectangle2_x(rectangle2_xs[1556]), .rectangle2_y(rectangle2_ys[1556]), .rectangle2_width(rectangle2_widths[1556]), .rectangle2_height(rectangle2_heights[1556]), .rectangle2_weight(rectangle2_weights[1556]), .rectangle3_x(rectangle3_xs[1556]), .rectangle3_y(rectangle3_ys[1556]), .rectangle3_width(rectangle3_widths[1556]), .rectangle3_height(rectangle3_heights[1556]), .rectangle3_weight(rectangle3_weights[1556]), .feature_threshold(feature_thresholds[1556]), .feature_above(feature_aboves[1556]), .feature_below(feature_belows[1556]), .scan_win_std_dev(scan_win_std_dev[1556]), .feature_accum(feature_accums[1556]));
  accum_calculator ac1557(.scan_win(scan_win1557), .rectangle1_x(rectangle1_xs[1557]), .rectangle1_y(rectangle1_ys[1557]), .rectangle1_width(rectangle1_widths[1557]), .rectangle1_height(rectangle1_heights[1557]), .rectangle1_weight(rectangle1_weights[1557]), .rectangle2_x(rectangle2_xs[1557]), .rectangle2_y(rectangle2_ys[1557]), .rectangle2_width(rectangle2_widths[1557]), .rectangle2_height(rectangle2_heights[1557]), .rectangle2_weight(rectangle2_weights[1557]), .rectangle3_x(rectangle3_xs[1557]), .rectangle3_y(rectangle3_ys[1557]), .rectangle3_width(rectangle3_widths[1557]), .rectangle3_height(rectangle3_heights[1557]), .rectangle3_weight(rectangle3_weights[1557]), .feature_threshold(feature_thresholds[1557]), .feature_above(feature_aboves[1557]), .feature_below(feature_belows[1557]), .scan_win_std_dev(scan_win_std_dev[1557]), .feature_accum(feature_accums[1557]));
  accum_calculator ac1558(.scan_win(scan_win1558), .rectangle1_x(rectangle1_xs[1558]), .rectangle1_y(rectangle1_ys[1558]), .rectangle1_width(rectangle1_widths[1558]), .rectangle1_height(rectangle1_heights[1558]), .rectangle1_weight(rectangle1_weights[1558]), .rectangle2_x(rectangle2_xs[1558]), .rectangle2_y(rectangle2_ys[1558]), .rectangle2_width(rectangle2_widths[1558]), .rectangle2_height(rectangle2_heights[1558]), .rectangle2_weight(rectangle2_weights[1558]), .rectangle3_x(rectangle3_xs[1558]), .rectangle3_y(rectangle3_ys[1558]), .rectangle3_width(rectangle3_widths[1558]), .rectangle3_height(rectangle3_heights[1558]), .rectangle3_weight(rectangle3_weights[1558]), .feature_threshold(feature_thresholds[1558]), .feature_above(feature_aboves[1558]), .feature_below(feature_belows[1558]), .scan_win_std_dev(scan_win_std_dev[1558]), .feature_accum(feature_accums[1558]));
  accum_calculator ac1559(.scan_win(scan_win1559), .rectangle1_x(rectangle1_xs[1559]), .rectangle1_y(rectangle1_ys[1559]), .rectangle1_width(rectangle1_widths[1559]), .rectangle1_height(rectangle1_heights[1559]), .rectangle1_weight(rectangle1_weights[1559]), .rectangle2_x(rectangle2_xs[1559]), .rectangle2_y(rectangle2_ys[1559]), .rectangle2_width(rectangle2_widths[1559]), .rectangle2_height(rectangle2_heights[1559]), .rectangle2_weight(rectangle2_weights[1559]), .rectangle3_x(rectangle3_xs[1559]), .rectangle3_y(rectangle3_ys[1559]), .rectangle3_width(rectangle3_widths[1559]), .rectangle3_height(rectangle3_heights[1559]), .rectangle3_weight(rectangle3_weights[1559]), .feature_threshold(feature_thresholds[1559]), .feature_above(feature_aboves[1559]), .feature_below(feature_belows[1559]), .scan_win_std_dev(scan_win_std_dev[1559]), .feature_accum(feature_accums[1559]));
  accum_calculator ac1560(.scan_win(scan_win1560), .rectangle1_x(rectangle1_xs[1560]), .rectangle1_y(rectangle1_ys[1560]), .rectangle1_width(rectangle1_widths[1560]), .rectangle1_height(rectangle1_heights[1560]), .rectangle1_weight(rectangle1_weights[1560]), .rectangle2_x(rectangle2_xs[1560]), .rectangle2_y(rectangle2_ys[1560]), .rectangle2_width(rectangle2_widths[1560]), .rectangle2_height(rectangle2_heights[1560]), .rectangle2_weight(rectangle2_weights[1560]), .rectangle3_x(rectangle3_xs[1560]), .rectangle3_y(rectangle3_ys[1560]), .rectangle3_width(rectangle3_widths[1560]), .rectangle3_height(rectangle3_heights[1560]), .rectangle3_weight(rectangle3_weights[1560]), .feature_threshold(feature_thresholds[1560]), .feature_above(feature_aboves[1560]), .feature_below(feature_belows[1560]), .scan_win_std_dev(scan_win_std_dev[1560]), .feature_accum(feature_accums[1560]));
  accum_calculator ac1561(.scan_win(scan_win1561), .rectangle1_x(rectangle1_xs[1561]), .rectangle1_y(rectangle1_ys[1561]), .rectangle1_width(rectangle1_widths[1561]), .rectangle1_height(rectangle1_heights[1561]), .rectangle1_weight(rectangle1_weights[1561]), .rectangle2_x(rectangle2_xs[1561]), .rectangle2_y(rectangle2_ys[1561]), .rectangle2_width(rectangle2_widths[1561]), .rectangle2_height(rectangle2_heights[1561]), .rectangle2_weight(rectangle2_weights[1561]), .rectangle3_x(rectangle3_xs[1561]), .rectangle3_y(rectangle3_ys[1561]), .rectangle3_width(rectangle3_widths[1561]), .rectangle3_height(rectangle3_heights[1561]), .rectangle3_weight(rectangle3_weights[1561]), .feature_threshold(feature_thresholds[1561]), .feature_above(feature_aboves[1561]), .feature_below(feature_belows[1561]), .scan_win_std_dev(scan_win_std_dev[1561]), .feature_accum(feature_accums[1561]));
  accum_calculator ac1562(.scan_win(scan_win1562), .rectangle1_x(rectangle1_xs[1562]), .rectangle1_y(rectangle1_ys[1562]), .rectangle1_width(rectangle1_widths[1562]), .rectangle1_height(rectangle1_heights[1562]), .rectangle1_weight(rectangle1_weights[1562]), .rectangle2_x(rectangle2_xs[1562]), .rectangle2_y(rectangle2_ys[1562]), .rectangle2_width(rectangle2_widths[1562]), .rectangle2_height(rectangle2_heights[1562]), .rectangle2_weight(rectangle2_weights[1562]), .rectangle3_x(rectangle3_xs[1562]), .rectangle3_y(rectangle3_ys[1562]), .rectangle3_width(rectangle3_widths[1562]), .rectangle3_height(rectangle3_heights[1562]), .rectangle3_weight(rectangle3_weights[1562]), .feature_threshold(feature_thresholds[1562]), .feature_above(feature_aboves[1562]), .feature_below(feature_belows[1562]), .scan_win_std_dev(scan_win_std_dev[1562]), .feature_accum(feature_accums[1562]));
  accum_calculator ac1563(.scan_win(scan_win1563), .rectangle1_x(rectangle1_xs[1563]), .rectangle1_y(rectangle1_ys[1563]), .rectangle1_width(rectangle1_widths[1563]), .rectangle1_height(rectangle1_heights[1563]), .rectangle1_weight(rectangle1_weights[1563]), .rectangle2_x(rectangle2_xs[1563]), .rectangle2_y(rectangle2_ys[1563]), .rectangle2_width(rectangle2_widths[1563]), .rectangle2_height(rectangle2_heights[1563]), .rectangle2_weight(rectangle2_weights[1563]), .rectangle3_x(rectangle3_xs[1563]), .rectangle3_y(rectangle3_ys[1563]), .rectangle3_width(rectangle3_widths[1563]), .rectangle3_height(rectangle3_heights[1563]), .rectangle3_weight(rectangle3_weights[1563]), .feature_threshold(feature_thresholds[1563]), .feature_above(feature_aboves[1563]), .feature_below(feature_belows[1563]), .scan_win_std_dev(scan_win_std_dev[1563]), .feature_accum(feature_accums[1563]));
  accum_calculator ac1564(.scan_win(scan_win1564), .rectangle1_x(rectangle1_xs[1564]), .rectangle1_y(rectangle1_ys[1564]), .rectangle1_width(rectangle1_widths[1564]), .rectangle1_height(rectangle1_heights[1564]), .rectangle1_weight(rectangle1_weights[1564]), .rectangle2_x(rectangle2_xs[1564]), .rectangle2_y(rectangle2_ys[1564]), .rectangle2_width(rectangle2_widths[1564]), .rectangle2_height(rectangle2_heights[1564]), .rectangle2_weight(rectangle2_weights[1564]), .rectangle3_x(rectangle3_xs[1564]), .rectangle3_y(rectangle3_ys[1564]), .rectangle3_width(rectangle3_widths[1564]), .rectangle3_height(rectangle3_heights[1564]), .rectangle3_weight(rectangle3_weights[1564]), .feature_threshold(feature_thresholds[1564]), .feature_above(feature_aboves[1564]), .feature_below(feature_belows[1564]), .scan_win_std_dev(scan_win_std_dev[1564]), .feature_accum(feature_accums[1564]));
  accum_calculator ac1565(.scan_win(scan_win1565), .rectangle1_x(rectangle1_xs[1565]), .rectangle1_y(rectangle1_ys[1565]), .rectangle1_width(rectangle1_widths[1565]), .rectangle1_height(rectangle1_heights[1565]), .rectangle1_weight(rectangle1_weights[1565]), .rectangle2_x(rectangle2_xs[1565]), .rectangle2_y(rectangle2_ys[1565]), .rectangle2_width(rectangle2_widths[1565]), .rectangle2_height(rectangle2_heights[1565]), .rectangle2_weight(rectangle2_weights[1565]), .rectangle3_x(rectangle3_xs[1565]), .rectangle3_y(rectangle3_ys[1565]), .rectangle3_width(rectangle3_widths[1565]), .rectangle3_height(rectangle3_heights[1565]), .rectangle3_weight(rectangle3_weights[1565]), .feature_threshold(feature_thresholds[1565]), .feature_above(feature_aboves[1565]), .feature_below(feature_belows[1565]), .scan_win_std_dev(scan_win_std_dev[1565]), .feature_accum(feature_accums[1565]));
  accum_calculator ac1566(.scan_win(scan_win1566), .rectangle1_x(rectangle1_xs[1566]), .rectangle1_y(rectangle1_ys[1566]), .rectangle1_width(rectangle1_widths[1566]), .rectangle1_height(rectangle1_heights[1566]), .rectangle1_weight(rectangle1_weights[1566]), .rectangle2_x(rectangle2_xs[1566]), .rectangle2_y(rectangle2_ys[1566]), .rectangle2_width(rectangle2_widths[1566]), .rectangle2_height(rectangle2_heights[1566]), .rectangle2_weight(rectangle2_weights[1566]), .rectangle3_x(rectangle3_xs[1566]), .rectangle3_y(rectangle3_ys[1566]), .rectangle3_width(rectangle3_widths[1566]), .rectangle3_height(rectangle3_heights[1566]), .rectangle3_weight(rectangle3_weights[1566]), .feature_threshold(feature_thresholds[1566]), .feature_above(feature_aboves[1566]), .feature_below(feature_belows[1566]), .scan_win_std_dev(scan_win_std_dev[1566]), .feature_accum(feature_accums[1566]));
  accum_calculator ac1567(.scan_win(scan_win1567), .rectangle1_x(rectangle1_xs[1567]), .rectangle1_y(rectangle1_ys[1567]), .rectangle1_width(rectangle1_widths[1567]), .rectangle1_height(rectangle1_heights[1567]), .rectangle1_weight(rectangle1_weights[1567]), .rectangle2_x(rectangle2_xs[1567]), .rectangle2_y(rectangle2_ys[1567]), .rectangle2_width(rectangle2_widths[1567]), .rectangle2_height(rectangle2_heights[1567]), .rectangle2_weight(rectangle2_weights[1567]), .rectangle3_x(rectangle3_xs[1567]), .rectangle3_y(rectangle3_ys[1567]), .rectangle3_width(rectangle3_widths[1567]), .rectangle3_height(rectangle3_heights[1567]), .rectangle3_weight(rectangle3_weights[1567]), .feature_threshold(feature_thresholds[1567]), .feature_above(feature_aboves[1567]), .feature_below(feature_belows[1567]), .scan_win_std_dev(scan_win_std_dev[1567]), .feature_accum(feature_accums[1567]));
  accum_calculator ac1568(.scan_win(scan_win1568), .rectangle1_x(rectangle1_xs[1568]), .rectangle1_y(rectangle1_ys[1568]), .rectangle1_width(rectangle1_widths[1568]), .rectangle1_height(rectangle1_heights[1568]), .rectangle1_weight(rectangle1_weights[1568]), .rectangle2_x(rectangle2_xs[1568]), .rectangle2_y(rectangle2_ys[1568]), .rectangle2_width(rectangle2_widths[1568]), .rectangle2_height(rectangle2_heights[1568]), .rectangle2_weight(rectangle2_weights[1568]), .rectangle3_x(rectangle3_xs[1568]), .rectangle3_y(rectangle3_ys[1568]), .rectangle3_width(rectangle3_widths[1568]), .rectangle3_height(rectangle3_heights[1568]), .rectangle3_weight(rectangle3_weights[1568]), .feature_threshold(feature_thresholds[1568]), .feature_above(feature_aboves[1568]), .feature_below(feature_belows[1568]), .scan_win_std_dev(scan_win_std_dev[1568]), .feature_accum(feature_accums[1568]));
  accum_calculator ac1569(.scan_win(scan_win1569), .rectangle1_x(rectangle1_xs[1569]), .rectangle1_y(rectangle1_ys[1569]), .rectangle1_width(rectangle1_widths[1569]), .rectangle1_height(rectangle1_heights[1569]), .rectangle1_weight(rectangle1_weights[1569]), .rectangle2_x(rectangle2_xs[1569]), .rectangle2_y(rectangle2_ys[1569]), .rectangle2_width(rectangle2_widths[1569]), .rectangle2_height(rectangle2_heights[1569]), .rectangle2_weight(rectangle2_weights[1569]), .rectangle3_x(rectangle3_xs[1569]), .rectangle3_y(rectangle3_ys[1569]), .rectangle3_width(rectangle3_widths[1569]), .rectangle3_height(rectangle3_heights[1569]), .rectangle3_weight(rectangle3_weights[1569]), .feature_threshold(feature_thresholds[1569]), .feature_above(feature_aboves[1569]), .feature_below(feature_belows[1569]), .scan_win_std_dev(scan_win_std_dev[1569]), .feature_accum(feature_accums[1569]));
  accum_calculator ac1570(.scan_win(scan_win1570), .rectangle1_x(rectangle1_xs[1570]), .rectangle1_y(rectangle1_ys[1570]), .rectangle1_width(rectangle1_widths[1570]), .rectangle1_height(rectangle1_heights[1570]), .rectangle1_weight(rectangle1_weights[1570]), .rectangle2_x(rectangle2_xs[1570]), .rectangle2_y(rectangle2_ys[1570]), .rectangle2_width(rectangle2_widths[1570]), .rectangle2_height(rectangle2_heights[1570]), .rectangle2_weight(rectangle2_weights[1570]), .rectangle3_x(rectangle3_xs[1570]), .rectangle3_y(rectangle3_ys[1570]), .rectangle3_width(rectangle3_widths[1570]), .rectangle3_height(rectangle3_heights[1570]), .rectangle3_weight(rectangle3_weights[1570]), .feature_threshold(feature_thresholds[1570]), .feature_above(feature_aboves[1570]), .feature_below(feature_belows[1570]), .scan_win_std_dev(scan_win_std_dev[1570]), .feature_accum(feature_accums[1570]));
  accum_calculator ac1571(.scan_win(scan_win1571), .rectangle1_x(rectangle1_xs[1571]), .rectangle1_y(rectangle1_ys[1571]), .rectangle1_width(rectangle1_widths[1571]), .rectangle1_height(rectangle1_heights[1571]), .rectangle1_weight(rectangle1_weights[1571]), .rectangle2_x(rectangle2_xs[1571]), .rectangle2_y(rectangle2_ys[1571]), .rectangle2_width(rectangle2_widths[1571]), .rectangle2_height(rectangle2_heights[1571]), .rectangle2_weight(rectangle2_weights[1571]), .rectangle3_x(rectangle3_xs[1571]), .rectangle3_y(rectangle3_ys[1571]), .rectangle3_width(rectangle3_widths[1571]), .rectangle3_height(rectangle3_heights[1571]), .rectangle3_weight(rectangle3_weights[1571]), .feature_threshold(feature_thresholds[1571]), .feature_above(feature_aboves[1571]), .feature_below(feature_belows[1571]), .scan_win_std_dev(scan_win_std_dev[1571]), .feature_accum(feature_accums[1571]));
  accum_calculator ac1572(.scan_win(scan_win1572), .rectangle1_x(rectangle1_xs[1572]), .rectangle1_y(rectangle1_ys[1572]), .rectangle1_width(rectangle1_widths[1572]), .rectangle1_height(rectangle1_heights[1572]), .rectangle1_weight(rectangle1_weights[1572]), .rectangle2_x(rectangle2_xs[1572]), .rectangle2_y(rectangle2_ys[1572]), .rectangle2_width(rectangle2_widths[1572]), .rectangle2_height(rectangle2_heights[1572]), .rectangle2_weight(rectangle2_weights[1572]), .rectangle3_x(rectangle3_xs[1572]), .rectangle3_y(rectangle3_ys[1572]), .rectangle3_width(rectangle3_widths[1572]), .rectangle3_height(rectangle3_heights[1572]), .rectangle3_weight(rectangle3_weights[1572]), .feature_threshold(feature_thresholds[1572]), .feature_above(feature_aboves[1572]), .feature_below(feature_belows[1572]), .scan_win_std_dev(scan_win_std_dev[1572]), .feature_accum(feature_accums[1572]));
  accum_calculator ac1573(.scan_win(scan_win1573), .rectangle1_x(rectangle1_xs[1573]), .rectangle1_y(rectangle1_ys[1573]), .rectangle1_width(rectangle1_widths[1573]), .rectangle1_height(rectangle1_heights[1573]), .rectangle1_weight(rectangle1_weights[1573]), .rectangle2_x(rectangle2_xs[1573]), .rectangle2_y(rectangle2_ys[1573]), .rectangle2_width(rectangle2_widths[1573]), .rectangle2_height(rectangle2_heights[1573]), .rectangle2_weight(rectangle2_weights[1573]), .rectangle3_x(rectangle3_xs[1573]), .rectangle3_y(rectangle3_ys[1573]), .rectangle3_width(rectangle3_widths[1573]), .rectangle3_height(rectangle3_heights[1573]), .rectangle3_weight(rectangle3_weights[1573]), .feature_threshold(feature_thresholds[1573]), .feature_above(feature_aboves[1573]), .feature_below(feature_belows[1573]), .scan_win_std_dev(scan_win_std_dev[1573]), .feature_accum(feature_accums[1573]));
  accum_calculator ac1574(.scan_win(scan_win1574), .rectangle1_x(rectangle1_xs[1574]), .rectangle1_y(rectangle1_ys[1574]), .rectangle1_width(rectangle1_widths[1574]), .rectangle1_height(rectangle1_heights[1574]), .rectangle1_weight(rectangle1_weights[1574]), .rectangle2_x(rectangle2_xs[1574]), .rectangle2_y(rectangle2_ys[1574]), .rectangle2_width(rectangle2_widths[1574]), .rectangle2_height(rectangle2_heights[1574]), .rectangle2_weight(rectangle2_weights[1574]), .rectangle3_x(rectangle3_xs[1574]), .rectangle3_y(rectangle3_ys[1574]), .rectangle3_width(rectangle3_widths[1574]), .rectangle3_height(rectangle3_heights[1574]), .rectangle3_weight(rectangle3_weights[1574]), .feature_threshold(feature_thresholds[1574]), .feature_above(feature_aboves[1574]), .feature_below(feature_belows[1574]), .scan_win_std_dev(scan_win_std_dev[1574]), .feature_accum(feature_accums[1574]));
  accum_calculator ac1575(.scan_win(scan_win1575), .rectangle1_x(rectangle1_xs[1575]), .rectangle1_y(rectangle1_ys[1575]), .rectangle1_width(rectangle1_widths[1575]), .rectangle1_height(rectangle1_heights[1575]), .rectangle1_weight(rectangle1_weights[1575]), .rectangle2_x(rectangle2_xs[1575]), .rectangle2_y(rectangle2_ys[1575]), .rectangle2_width(rectangle2_widths[1575]), .rectangle2_height(rectangle2_heights[1575]), .rectangle2_weight(rectangle2_weights[1575]), .rectangle3_x(rectangle3_xs[1575]), .rectangle3_y(rectangle3_ys[1575]), .rectangle3_width(rectangle3_widths[1575]), .rectangle3_height(rectangle3_heights[1575]), .rectangle3_weight(rectangle3_weights[1575]), .feature_threshold(feature_thresholds[1575]), .feature_above(feature_aboves[1575]), .feature_below(feature_belows[1575]), .scan_win_std_dev(scan_win_std_dev[1575]), .feature_accum(feature_accums[1575]));
  accum_calculator ac1576(.scan_win(scan_win1576), .rectangle1_x(rectangle1_xs[1576]), .rectangle1_y(rectangle1_ys[1576]), .rectangle1_width(rectangle1_widths[1576]), .rectangle1_height(rectangle1_heights[1576]), .rectangle1_weight(rectangle1_weights[1576]), .rectangle2_x(rectangle2_xs[1576]), .rectangle2_y(rectangle2_ys[1576]), .rectangle2_width(rectangle2_widths[1576]), .rectangle2_height(rectangle2_heights[1576]), .rectangle2_weight(rectangle2_weights[1576]), .rectangle3_x(rectangle3_xs[1576]), .rectangle3_y(rectangle3_ys[1576]), .rectangle3_width(rectangle3_widths[1576]), .rectangle3_height(rectangle3_heights[1576]), .rectangle3_weight(rectangle3_weights[1576]), .feature_threshold(feature_thresholds[1576]), .feature_above(feature_aboves[1576]), .feature_below(feature_belows[1576]), .scan_win_std_dev(scan_win_std_dev[1576]), .feature_accum(feature_accums[1576]));
  accum_calculator ac1577(.scan_win(scan_win1577), .rectangle1_x(rectangle1_xs[1577]), .rectangle1_y(rectangle1_ys[1577]), .rectangle1_width(rectangle1_widths[1577]), .rectangle1_height(rectangle1_heights[1577]), .rectangle1_weight(rectangle1_weights[1577]), .rectangle2_x(rectangle2_xs[1577]), .rectangle2_y(rectangle2_ys[1577]), .rectangle2_width(rectangle2_widths[1577]), .rectangle2_height(rectangle2_heights[1577]), .rectangle2_weight(rectangle2_weights[1577]), .rectangle3_x(rectangle3_xs[1577]), .rectangle3_y(rectangle3_ys[1577]), .rectangle3_width(rectangle3_widths[1577]), .rectangle3_height(rectangle3_heights[1577]), .rectangle3_weight(rectangle3_weights[1577]), .feature_threshold(feature_thresholds[1577]), .feature_above(feature_aboves[1577]), .feature_below(feature_belows[1577]), .scan_win_std_dev(scan_win_std_dev[1577]), .feature_accum(feature_accums[1577]));
  accum_calculator ac1578(.scan_win(scan_win1578), .rectangle1_x(rectangle1_xs[1578]), .rectangle1_y(rectangle1_ys[1578]), .rectangle1_width(rectangle1_widths[1578]), .rectangle1_height(rectangle1_heights[1578]), .rectangle1_weight(rectangle1_weights[1578]), .rectangle2_x(rectangle2_xs[1578]), .rectangle2_y(rectangle2_ys[1578]), .rectangle2_width(rectangle2_widths[1578]), .rectangle2_height(rectangle2_heights[1578]), .rectangle2_weight(rectangle2_weights[1578]), .rectangle3_x(rectangle3_xs[1578]), .rectangle3_y(rectangle3_ys[1578]), .rectangle3_width(rectangle3_widths[1578]), .rectangle3_height(rectangle3_heights[1578]), .rectangle3_weight(rectangle3_weights[1578]), .feature_threshold(feature_thresholds[1578]), .feature_above(feature_aboves[1578]), .feature_below(feature_belows[1578]), .scan_win_std_dev(scan_win_std_dev[1578]), .feature_accum(feature_accums[1578]));
  accum_calculator ac1579(.scan_win(scan_win1579), .rectangle1_x(rectangle1_xs[1579]), .rectangle1_y(rectangle1_ys[1579]), .rectangle1_width(rectangle1_widths[1579]), .rectangle1_height(rectangle1_heights[1579]), .rectangle1_weight(rectangle1_weights[1579]), .rectangle2_x(rectangle2_xs[1579]), .rectangle2_y(rectangle2_ys[1579]), .rectangle2_width(rectangle2_widths[1579]), .rectangle2_height(rectangle2_heights[1579]), .rectangle2_weight(rectangle2_weights[1579]), .rectangle3_x(rectangle3_xs[1579]), .rectangle3_y(rectangle3_ys[1579]), .rectangle3_width(rectangle3_widths[1579]), .rectangle3_height(rectangle3_heights[1579]), .rectangle3_weight(rectangle3_weights[1579]), .feature_threshold(feature_thresholds[1579]), .feature_above(feature_aboves[1579]), .feature_below(feature_belows[1579]), .scan_win_std_dev(scan_win_std_dev[1579]), .feature_accum(feature_accums[1579]));
  accum_calculator ac1580(.scan_win(scan_win1580), .rectangle1_x(rectangle1_xs[1580]), .rectangle1_y(rectangle1_ys[1580]), .rectangle1_width(rectangle1_widths[1580]), .rectangle1_height(rectangle1_heights[1580]), .rectangle1_weight(rectangle1_weights[1580]), .rectangle2_x(rectangle2_xs[1580]), .rectangle2_y(rectangle2_ys[1580]), .rectangle2_width(rectangle2_widths[1580]), .rectangle2_height(rectangle2_heights[1580]), .rectangle2_weight(rectangle2_weights[1580]), .rectangle3_x(rectangle3_xs[1580]), .rectangle3_y(rectangle3_ys[1580]), .rectangle3_width(rectangle3_widths[1580]), .rectangle3_height(rectangle3_heights[1580]), .rectangle3_weight(rectangle3_weights[1580]), .feature_threshold(feature_thresholds[1580]), .feature_above(feature_aboves[1580]), .feature_below(feature_belows[1580]), .scan_win_std_dev(scan_win_std_dev[1580]), .feature_accum(feature_accums[1580]));
  accum_calculator ac1581(.scan_win(scan_win1581), .rectangle1_x(rectangle1_xs[1581]), .rectangle1_y(rectangle1_ys[1581]), .rectangle1_width(rectangle1_widths[1581]), .rectangle1_height(rectangle1_heights[1581]), .rectangle1_weight(rectangle1_weights[1581]), .rectangle2_x(rectangle2_xs[1581]), .rectangle2_y(rectangle2_ys[1581]), .rectangle2_width(rectangle2_widths[1581]), .rectangle2_height(rectangle2_heights[1581]), .rectangle2_weight(rectangle2_weights[1581]), .rectangle3_x(rectangle3_xs[1581]), .rectangle3_y(rectangle3_ys[1581]), .rectangle3_width(rectangle3_widths[1581]), .rectangle3_height(rectangle3_heights[1581]), .rectangle3_weight(rectangle3_weights[1581]), .feature_threshold(feature_thresholds[1581]), .feature_above(feature_aboves[1581]), .feature_below(feature_belows[1581]), .scan_win_std_dev(scan_win_std_dev[1581]), .feature_accum(feature_accums[1581]));
  accum_calculator ac1582(.scan_win(scan_win1582), .rectangle1_x(rectangle1_xs[1582]), .rectangle1_y(rectangle1_ys[1582]), .rectangle1_width(rectangle1_widths[1582]), .rectangle1_height(rectangle1_heights[1582]), .rectangle1_weight(rectangle1_weights[1582]), .rectangle2_x(rectangle2_xs[1582]), .rectangle2_y(rectangle2_ys[1582]), .rectangle2_width(rectangle2_widths[1582]), .rectangle2_height(rectangle2_heights[1582]), .rectangle2_weight(rectangle2_weights[1582]), .rectangle3_x(rectangle3_xs[1582]), .rectangle3_y(rectangle3_ys[1582]), .rectangle3_width(rectangle3_widths[1582]), .rectangle3_height(rectangle3_heights[1582]), .rectangle3_weight(rectangle3_weights[1582]), .feature_threshold(feature_thresholds[1582]), .feature_above(feature_aboves[1582]), .feature_below(feature_belows[1582]), .scan_win_std_dev(scan_win_std_dev[1582]), .feature_accum(feature_accums[1582]));
  accum_calculator ac1583(.scan_win(scan_win1583), .rectangle1_x(rectangle1_xs[1583]), .rectangle1_y(rectangle1_ys[1583]), .rectangle1_width(rectangle1_widths[1583]), .rectangle1_height(rectangle1_heights[1583]), .rectangle1_weight(rectangle1_weights[1583]), .rectangle2_x(rectangle2_xs[1583]), .rectangle2_y(rectangle2_ys[1583]), .rectangle2_width(rectangle2_widths[1583]), .rectangle2_height(rectangle2_heights[1583]), .rectangle2_weight(rectangle2_weights[1583]), .rectangle3_x(rectangle3_xs[1583]), .rectangle3_y(rectangle3_ys[1583]), .rectangle3_width(rectangle3_widths[1583]), .rectangle3_height(rectangle3_heights[1583]), .rectangle3_weight(rectangle3_weights[1583]), .feature_threshold(feature_thresholds[1583]), .feature_above(feature_aboves[1583]), .feature_below(feature_belows[1583]), .scan_win_std_dev(scan_win_std_dev[1583]), .feature_accum(feature_accums[1583]));
  accum_calculator ac1584(.scan_win(scan_win1584), .rectangle1_x(rectangle1_xs[1584]), .rectangle1_y(rectangle1_ys[1584]), .rectangle1_width(rectangle1_widths[1584]), .rectangle1_height(rectangle1_heights[1584]), .rectangle1_weight(rectangle1_weights[1584]), .rectangle2_x(rectangle2_xs[1584]), .rectangle2_y(rectangle2_ys[1584]), .rectangle2_width(rectangle2_widths[1584]), .rectangle2_height(rectangle2_heights[1584]), .rectangle2_weight(rectangle2_weights[1584]), .rectangle3_x(rectangle3_xs[1584]), .rectangle3_y(rectangle3_ys[1584]), .rectangle3_width(rectangle3_widths[1584]), .rectangle3_height(rectangle3_heights[1584]), .rectangle3_weight(rectangle3_weights[1584]), .feature_threshold(feature_thresholds[1584]), .feature_above(feature_aboves[1584]), .feature_below(feature_belows[1584]), .scan_win_std_dev(scan_win_std_dev[1584]), .feature_accum(feature_accums[1584]));
  accum_calculator ac1585(.scan_win(scan_win1585), .rectangle1_x(rectangle1_xs[1585]), .rectangle1_y(rectangle1_ys[1585]), .rectangle1_width(rectangle1_widths[1585]), .rectangle1_height(rectangle1_heights[1585]), .rectangle1_weight(rectangle1_weights[1585]), .rectangle2_x(rectangle2_xs[1585]), .rectangle2_y(rectangle2_ys[1585]), .rectangle2_width(rectangle2_widths[1585]), .rectangle2_height(rectangle2_heights[1585]), .rectangle2_weight(rectangle2_weights[1585]), .rectangle3_x(rectangle3_xs[1585]), .rectangle3_y(rectangle3_ys[1585]), .rectangle3_width(rectangle3_widths[1585]), .rectangle3_height(rectangle3_heights[1585]), .rectangle3_weight(rectangle3_weights[1585]), .feature_threshold(feature_thresholds[1585]), .feature_above(feature_aboves[1585]), .feature_below(feature_belows[1585]), .scan_win_std_dev(scan_win_std_dev[1585]), .feature_accum(feature_accums[1585]));
  accum_calculator ac1586(.scan_win(scan_win1586), .rectangle1_x(rectangle1_xs[1586]), .rectangle1_y(rectangle1_ys[1586]), .rectangle1_width(rectangle1_widths[1586]), .rectangle1_height(rectangle1_heights[1586]), .rectangle1_weight(rectangle1_weights[1586]), .rectangle2_x(rectangle2_xs[1586]), .rectangle2_y(rectangle2_ys[1586]), .rectangle2_width(rectangle2_widths[1586]), .rectangle2_height(rectangle2_heights[1586]), .rectangle2_weight(rectangle2_weights[1586]), .rectangle3_x(rectangle3_xs[1586]), .rectangle3_y(rectangle3_ys[1586]), .rectangle3_width(rectangle3_widths[1586]), .rectangle3_height(rectangle3_heights[1586]), .rectangle3_weight(rectangle3_weights[1586]), .feature_threshold(feature_thresholds[1586]), .feature_above(feature_aboves[1586]), .feature_below(feature_belows[1586]), .scan_win_std_dev(scan_win_std_dev[1586]), .feature_accum(feature_accums[1586]));
  accum_calculator ac1587(.scan_win(scan_win1587), .rectangle1_x(rectangle1_xs[1587]), .rectangle1_y(rectangle1_ys[1587]), .rectangle1_width(rectangle1_widths[1587]), .rectangle1_height(rectangle1_heights[1587]), .rectangle1_weight(rectangle1_weights[1587]), .rectangle2_x(rectangle2_xs[1587]), .rectangle2_y(rectangle2_ys[1587]), .rectangle2_width(rectangle2_widths[1587]), .rectangle2_height(rectangle2_heights[1587]), .rectangle2_weight(rectangle2_weights[1587]), .rectangle3_x(rectangle3_xs[1587]), .rectangle3_y(rectangle3_ys[1587]), .rectangle3_width(rectangle3_widths[1587]), .rectangle3_height(rectangle3_heights[1587]), .rectangle3_weight(rectangle3_weights[1587]), .feature_threshold(feature_thresholds[1587]), .feature_above(feature_aboves[1587]), .feature_below(feature_belows[1587]), .scan_win_std_dev(scan_win_std_dev[1587]), .feature_accum(feature_accums[1587]));
  accum_calculator ac1588(.scan_win(scan_win1588), .rectangle1_x(rectangle1_xs[1588]), .rectangle1_y(rectangle1_ys[1588]), .rectangle1_width(rectangle1_widths[1588]), .rectangle1_height(rectangle1_heights[1588]), .rectangle1_weight(rectangle1_weights[1588]), .rectangle2_x(rectangle2_xs[1588]), .rectangle2_y(rectangle2_ys[1588]), .rectangle2_width(rectangle2_widths[1588]), .rectangle2_height(rectangle2_heights[1588]), .rectangle2_weight(rectangle2_weights[1588]), .rectangle3_x(rectangle3_xs[1588]), .rectangle3_y(rectangle3_ys[1588]), .rectangle3_width(rectangle3_widths[1588]), .rectangle3_height(rectangle3_heights[1588]), .rectangle3_weight(rectangle3_weights[1588]), .feature_threshold(feature_thresholds[1588]), .feature_above(feature_aboves[1588]), .feature_below(feature_belows[1588]), .scan_win_std_dev(scan_win_std_dev[1588]), .feature_accum(feature_accums[1588]));
  accum_calculator ac1589(.scan_win(scan_win1589), .rectangle1_x(rectangle1_xs[1589]), .rectangle1_y(rectangle1_ys[1589]), .rectangle1_width(rectangle1_widths[1589]), .rectangle1_height(rectangle1_heights[1589]), .rectangle1_weight(rectangle1_weights[1589]), .rectangle2_x(rectangle2_xs[1589]), .rectangle2_y(rectangle2_ys[1589]), .rectangle2_width(rectangle2_widths[1589]), .rectangle2_height(rectangle2_heights[1589]), .rectangle2_weight(rectangle2_weights[1589]), .rectangle3_x(rectangle3_xs[1589]), .rectangle3_y(rectangle3_ys[1589]), .rectangle3_width(rectangle3_widths[1589]), .rectangle3_height(rectangle3_heights[1589]), .rectangle3_weight(rectangle3_weights[1589]), .feature_threshold(feature_thresholds[1589]), .feature_above(feature_aboves[1589]), .feature_below(feature_belows[1589]), .scan_win_std_dev(scan_win_std_dev[1589]), .feature_accum(feature_accums[1589]));
  accum_calculator ac1590(.scan_win(scan_win1590), .rectangle1_x(rectangle1_xs[1590]), .rectangle1_y(rectangle1_ys[1590]), .rectangle1_width(rectangle1_widths[1590]), .rectangle1_height(rectangle1_heights[1590]), .rectangle1_weight(rectangle1_weights[1590]), .rectangle2_x(rectangle2_xs[1590]), .rectangle2_y(rectangle2_ys[1590]), .rectangle2_width(rectangle2_widths[1590]), .rectangle2_height(rectangle2_heights[1590]), .rectangle2_weight(rectangle2_weights[1590]), .rectangle3_x(rectangle3_xs[1590]), .rectangle3_y(rectangle3_ys[1590]), .rectangle3_width(rectangle3_widths[1590]), .rectangle3_height(rectangle3_heights[1590]), .rectangle3_weight(rectangle3_weights[1590]), .feature_threshold(feature_thresholds[1590]), .feature_above(feature_aboves[1590]), .feature_below(feature_belows[1590]), .scan_win_std_dev(scan_win_std_dev[1590]), .feature_accum(feature_accums[1590]));
  accum_calculator ac1591(.scan_win(scan_win1591), .rectangle1_x(rectangle1_xs[1591]), .rectangle1_y(rectangle1_ys[1591]), .rectangle1_width(rectangle1_widths[1591]), .rectangle1_height(rectangle1_heights[1591]), .rectangle1_weight(rectangle1_weights[1591]), .rectangle2_x(rectangle2_xs[1591]), .rectangle2_y(rectangle2_ys[1591]), .rectangle2_width(rectangle2_widths[1591]), .rectangle2_height(rectangle2_heights[1591]), .rectangle2_weight(rectangle2_weights[1591]), .rectangle3_x(rectangle3_xs[1591]), .rectangle3_y(rectangle3_ys[1591]), .rectangle3_width(rectangle3_widths[1591]), .rectangle3_height(rectangle3_heights[1591]), .rectangle3_weight(rectangle3_weights[1591]), .feature_threshold(feature_thresholds[1591]), .feature_above(feature_aboves[1591]), .feature_below(feature_belows[1591]), .scan_win_std_dev(scan_win_std_dev[1591]), .feature_accum(feature_accums[1591]));
  accum_calculator ac1592(.scan_win(scan_win1592), .rectangle1_x(rectangle1_xs[1592]), .rectangle1_y(rectangle1_ys[1592]), .rectangle1_width(rectangle1_widths[1592]), .rectangle1_height(rectangle1_heights[1592]), .rectangle1_weight(rectangle1_weights[1592]), .rectangle2_x(rectangle2_xs[1592]), .rectangle2_y(rectangle2_ys[1592]), .rectangle2_width(rectangle2_widths[1592]), .rectangle2_height(rectangle2_heights[1592]), .rectangle2_weight(rectangle2_weights[1592]), .rectangle3_x(rectangle3_xs[1592]), .rectangle3_y(rectangle3_ys[1592]), .rectangle3_width(rectangle3_widths[1592]), .rectangle3_height(rectangle3_heights[1592]), .rectangle3_weight(rectangle3_weights[1592]), .feature_threshold(feature_thresholds[1592]), .feature_above(feature_aboves[1592]), .feature_below(feature_belows[1592]), .scan_win_std_dev(scan_win_std_dev[1592]), .feature_accum(feature_accums[1592]));
  accum_calculator ac1593(.scan_win(scan_win1593), .rectangle1_x(rectangle1_xs[1593]), .rectangle1_y(rectangle1_ys[1593]), .rectangle1_width(rectangle1_widths[1593]), .rectangle1_height(rectangle1_heights[1593]), .rectangle1_weight(rectangle1_weights[1593]), .rectangle2_x(rectangle2_xs[1593]), .rectangle2_y(rectangle2_ys[1593]), .rectangle2_width(rectangle2_widths[1593]), .rectangle2_height(rectangle2_heights[1593]), .rectangle2_weight(rectangle2_weights[1593]), .rectangle3_x(rectangle3_xs[1593]), .rectangle3_y(rectangle3_ys[1593]), .rectangle3_width(rectangle3_widths[1593]), .rectangle3_height(rectangle3_heights[1593]), .rectangle3_weight(rectangle3_weights[1593]), .feature_threshold(feature_thresholds[1593]), .feature_above(feature_aboves[1593]), .feature_below(feature_belows[1593]), .scan_win_std_dev(scan_win_std_dev[1593]), .feature_accum(feature_accums[1593]));
  accum_calculator ac1594(.scan_win(scan_win1594), .rectangle1_x(rectangle1_xs[1594]), .rectangle1_y(rectangle1_ys[1594]), .rectangle1_width(rectangle1_widths[1594]), .rectangle1_height(rectangle1_heights[1594]), .rectangle1_weight(rectangle1_weights[1594]), .rectangle2_x(rectangle2_xs[1594]), .rectangle2_y(rectangle2_ys[1594]), .rectangle2_width(rectangle2_widths[1594]), .rectangle2_height(rectangle2_heights[1594]), .rectangle2_weight(rectangle2_weights[1594]), .rectangle3_x(rectangle3_xs[1594]), .rectangle3_y(rectangle3_ys[1594]), .rectangle3_width(rectangle3_widths[1594]), .rectangle3_height(rectangle3_heights[1594]), .rectangle3_weight(rectangle3_weights[1594]), .feature_threshold(feature_thresholds[1594]), .feature_above(feature_aboves[1594]), .feature_below(feature_belows[1594]), .scan_win_std_dev(scan_win_std_dev[1594]), .feature_accum(feature_accums[1594]));
  accum_calculator ac1595(.scan_win(scan_win1595), .rectangle1_x(rectangle1_xs[1595]), .rectangle1_y(rectangle1_ys[1595]), .rectangle1_width(rectangle1_widths[1595]), .rectangle1_height(rectangle1_heights[1595]), .rectangle1_weight(rectangle1_weights[1595]), .rectangle2_x(rectangle2_xs[1595]), .rectangle2_y(rectangle2_ys[1595]), .rectangle2_width(rectangle2_widths[1595]), .rectangle2_height(rectangle2_heights[1595]), .rectangle2_weight(rectangle2_weights[1595]), .rectangle3_x(rectangle3_xs[1595]), .rectangle3_y(rectangle3_ys[1595]), .rectangle3_width(rectangle3_widths[1595]), .rectangle3_height(rectangle3_heights[1595]), .rectangle3_weight(rectangle3_weights[1595]), .feature_threshold(feature_thresholds[1595]), .feature_above(feature_aboves[1595]), .feature_below(feature_belows[1595]), .scan_win_std_dev(scan_win_std_dev[1595]), .feature_accum(feature_accums[1595]));
  accum_calculator ac1596(.scan_win(scan_win1596), .rectangle1_x(rectangle1_xs[1596]), .rectangle1_y(rectangle1_ys[1596]), .rectangle1_width(rectangle1_widths[1596]), .rectangle1_height(rectangle1_heights[1596]), .rectangle1_weight(rectangle1_weights[1596]), .rectangle2_x(rectangle2_xs[1596]), .rectangle2_y(rectangle2_ys[1596]), .rectangle2_width(rectangle2_widths[1596]), .rectangle2_height(rectangle2_heights[1596]), .rectangle2_weight(rectangle2_weights[1596]), .rectangle3_x(rectangle3_xs[1596]), .rectangle3_y(rectangle3_ys[1596]), .rectangle3_width(rectangle3_widths[1596]), .rectangle3_height(rectangle3_heights[1596]), .rectangle3_weight(rectangle3_weights[1596]), .feature_threshold(feature_thresholds[1596]), .feature_above(feature_aboves[1596]), .feature_below(feature_belows[1596]), .scan_win_std_dev(scan_win_std_dev[1596]), .feature_accum(feature_accums[1596]));
  accum_calculator ac1597(.scan_win(scan_win1597), .rectangle1_x(rectangle1_xs[1597]), .rectangle1_y(rectangle1_ys[1597]), .rectangle1_width(rectangle1_widths[1597]), .rectangle1_height(rectangle1_heights[1597]), .rectangle1_weight(rectangle1_weights[1597]), .rectangle2_x(rectangle2_xs[1597]), .rectangle2_y(rectangle2_ys[1597]), .rectangle2_width(rectangle2_widths[1597]), .rectangle2_height(rectangle2_heights[1597]), .rectangle2_weight(rectangle2_weights[1597]), .rectangle3_x(rectangle3_xs[1597]), .rectangle3_y(rectangle3_ys[1597]), .rectangle3_width(rectangle3_widths[1597]), .rectangle3_height(rectangle3_heights[1597]), .rectangle3_weight(rectangle3_weights[1597]), .feature_threshold(feature_thresholds[1597]), .feature_above(feature_aboves[1597]), .feature_below(feature_belows[1597]), .scan_win_std_dev(scan_win_std_dev[1597]), .feature_accum(feature_accums[1597]));
  accum_calculator ac1598(.scan_win(scan_win1598), .rectangle1_x(rectangle1_xs[1598]), .rectangle1_y(rectangle1_ys[1598]), .rectangle1_width(rectangle1_widths[1598]), .rectangle1_height(rectangle1_heights[1598]), .rectangle1_weight(rectangle1_weights[1598]), .rectangle2_x(rectangle2_xs[1598]), .rectangle2_y(rectangle2_ys[1598]), .rectangle2_width(rectangle2_widths[1598]), .rectangle2_height(rectangle2_heights[1598]), .rectangle2_weight(rectangle2_weights[1598]), .rectangle3_x(rectangle3_xs[1598]), .rectangle3_y(rectangle3_ys[1598]), .rectangle3_width(rectangle3_widths[1598]), .rectangle3_height(rectangle3_heights[1598]), .rectangle3_weight(rectangle3_weights[1598]), .feature_threshold(feature_thresholds[1598]), .feature_above(feature_aboves[1598]), .feature_below(feature_belows[1598]), .scan_win_std_dev(scan_win_std_dev[1598]), .feature_accum(feature_accums[1598]));
  accum_calculator ac1599(.scan_win(scan_win1599), .rectangle1_x(rectangle1_xs[1599]), .rectangle1_y(rectangle1_ys[1599]), .rectangle1_width(rectangle1_widths[1599]), .rectangle1_height(rectangle1_heights[1599]), .rectangle1_weight(rectangle1_weights[1599]), .rectangle2_x(rectangle2_xs[1599]), .rectangle2_y(rectangle2_ys[1599]), .rectangle2_width(rectangle2_widths[1599]), .rectangle2_height(rectangle2_heights[1599]), .rectangle2_weight(rectangle2_weights[1599]), .rectangle3_x(rectangle3_xs[1599]), .rectangle3_y(rectangle3_ys[1599]), .rectangle3_width(rectangle3_widths[1599]), .rectangle3_height(rectangle3_heights[1599]), .rectangle3_weight(rectangle3_weights[1599]), .feature_threshold(feature_thresholds[1599]), .feature_above(feature_aboves[1599]), .feature_below(feature_belows[1599]), .scan_win_std_dev(scan_win_std_dev[1599]), .feature_accum(feature_accums[1599]));
  accum_calculator ac1600(.scan_win(scan_win1600), .rectangle1_x(rectangle1_xs[1600]), .rectangle1_y(rectangle1_ys[1600]), .rectangle1_width(rectangle1_widths[1600]), .rectangle1_height(rectangle1_heights[1600]), .rectangle1_weight(rectangle1_weights[1600]), .rectangle2_x(rectangle2_xs[1600]), .rectangle2_y(rectangle2_ys[1600]), .rectangle2_width(rectangle2_widths[1600]), .rectangle2_height(rectangle2_heights[1600]), .rectangle2_weight(rectangle2_weights[1600]), .rectangle3_x(rectangle3_xs[1600]), .rectangle3_y(rectangle3_ys[1600]), .rectangle3_width(rectangle3_widths[1600]), .rectangle3_height(rectangle3_heights[1600]), .rectangle3_weight(rectangle3_weights[1600]), .feature_threshold(feature_thresholds[1600]), .feature_above(feature_aboves[1600]), .feature_below(feature_belows[1600]), .scan_win_std_dev(scan_win_std_dev[1600]), .feature_accum(feature_accums[1600]));
  accum_calculator ac1601(.scan_win(scan_win1601), .rectangle1_x(rectangle1_xs[1601]), .rectangle1_y(rectangle1_ys[1601]), .rectangle1_width(rectangle1_widths[1601]), .rectangle1_height(rectangle1_heights[1601]), .rectangle1_weight(rectangle1_weights[1601]), .rectangle2_x(rectangle2_xs[1601]), .rectangle2_y(rectangle2_ys[1601]), .rectangle2_width(rectangle2_widths[1601]), .rectangle2_height(rectangle2_heights[1601]), .rectangle2_weight(rectangle2_weights[1601]), .rectangle3_x(rectangle3_xs[1601]), .rectangle3_y(rectangle3_ys[1601]), .rectangle3_width(rectangle3_widths[1601]), .rectangle3_height(rectangle3_heights[1601]), .rectangle3_weight(rectangle3_weights[1601]), .feature_threshold(feature_thresholds[1601]), .feature_above(feature_aboves[1601]), .feature_below(feature_belows[1601]), .scan_win_std_dev(scan_win_std_dev[1601]), .feature_accum(feature_accums[1601]));
  accum_calculator ac1602(.scan_win(scan_win1602), .rectangle1_x(rectangle1_xs[1602]), .rectangle1_y(rectangle1_ys[1602]), .rectangle1_width(rectangle1_widths[1602]), .rectangle1_height(rectangle1_heights[1602]), .rectangle1_weight(rectangle1_weights[1602]), .rectangle2_x(rectangle2_xs[1602]), .rectangle2_y(rectangle2_ys[1602]), .rectangle2_width(rectangle2_widths[1602]), .rectangle2_height(rectangle2_heights[1602]), .rectangle2_weight(rectangle2_weights[1602]), .rectangle3_x(rectangle3_xs[1602]), .rectangle3_y(rectangle3_ys[1602]), .rectangle3_width(rectangle3_widths[1602]), .rectangle3_height(rectangle3_heights[1602]), .rectangle3_weight(rectangle3_weights[1602]), .feature_threshold(feature_thresholds[1602]), .feature_above(feature_aboves[1602]), .feature_below(feature_belows[1602]), .scan_win_std_dev(scan_win_std_dev[1602]), .feature_accum(feature_accums[1602]));
  accum_calculator ac1603(.scan_win(scan_win1603), .rectangle1_x(rectangle1_xs[1603]), .rectangle1_y(rectangle1_ys[1603]), .rectangle1_width(rectangle1_widths[1603]), .rectangle1_height(rectangle1_heights[1603]), .rectangle1_weight(rectangle1_weights[1603]), .rectangle2_x(rectangle2_xs[1603]), .rectangle2_y(rectangle2_ys[1603]), .rectangle2_width(rectangle2_widths[1603]), .rectangle2_height(rectangle2_heights[1603]), .rectangle2_weight(rectangle2_weights[1603]), .rectangle3_x(rectangle3_xs[1603]), .rectangle3_y(rectangle3_ys[1603]), .rectangle3_width(rectangle3_widths[1603]), .rectangle3_height(rectangle3_heights[1603]), .rectangle3_weight(rectangle3_weights[1603]), .feature_threshold(feature_thresholds[1603]), .feature_above(feature_aboves[1603]), .feature_below(feature_belows[1603]), .scan_win_std_dev(scan_win_std_dev[1603]), .feature_accum(feature_accums[1603]));
  accum_calculator ac1604(.scan_win(scan_win1604), .rectangle1_x(rectangle1_xs[1604]), .rectangle1_y(rectangle1_ys[1604]), .rectangle1_width(rectangle1_widths[1604]), .rectangle1_height(rectangle1_heights[1604]), .rectangle1_weight(rectangle1_weights[1604]), .rectangle2_x(rectangle2_xs[1604]), .rectangle2_y(rectangle2_ys[1604]), .rectangle2_width(rectangle2_widths[1604]), .rectangle2_height(rectangle2_heights[1604]), .rectangle2_weight(rectangle2_weights[1604]), .rectangle3_x(rectangle3_xs[1604]), .rectangle3_y(rectangle3_ys[1604]), .rectangle3_width(rectangle3_widths[1604]), .rectangle3_height(rectangle3_heights[1604]), .rectangle3_weight(rectangle3_weights[1604]), .feature_threshold(feature_thresholds[1604]), .feature_above(feature_aboves[1604]), .feature_below(feature_belows[1604]), .scan_win_std_dev(scan_win_std_dev[1604]), .feature_accum(feature_accums[1604]));
  accum_calculator ac1605(.scan_win(scan_win1605), .rectangle1_x(rectangle1_xs[1605]), .rectangle1_y(rectangle1_ys[1605]), .rectangle1_width(rectangle1_widths[1605]), .rectangle1_height(rectangle1_heights[1605]), .rectangle1_weight(rectangle1_weights[1605]), .rectangle2_x(rectangle2_xs[1605]), .rectangle2_y(rectangle2_ys[1605]), .rectangle2_width(rectangle2_widths[1605]), .rectangle2_height(rectangle2_heights[1605]), .rectangle2_weight(rectangle2_weights[1605]), .rectangle3_x(rectangle3_xs[1605]), .rectangle3_y(rectangle3_ys[1605]), .rectangle3_width(rectangle3_widths[1605]), .rectangle3_height(rectangle3_heights[1605]), .rectangle3_weight(rectangle3_weights[1605]), .feature_threshold(feature_thresholds[1605]), .feature_above(feature_aboves[1605]), .feature_below(feature_belows[1605]), .scan_win_std_dev(scan_win_std_dev[1605]), .feature_accum(feature_accums[1605]));
  accum_calculator ac1606(.scan_win(scan_win1606), .rectangle1_x(rectangle1_xs[1606]), .rectangle1_y(rectangle1_ys[1606]), .rectangle1_width(rectangle1_widths[1606]), .rectangle1_height(rectangle1_heights[1606]), .rectangle1_weight(rectangle1_weights[1606]), .rectangle2_x(rectangle2_xs[1606]), .rectangle2_y(rectangle2_ys[1606]), .rectangle2_width(rectangle2_widths[1606]), .rectangle2_height(rectangle2_heights[1606]), .rectangle2_weight(rectangle2_weights[1606]), .rectangle3_x(rectangle3_xs[1606]), .rectangle3_y(rectangle3_ys[1606]), .rectangle3_width(rectangle3_widths[1606]), .rectangle3_height(rectangle3_heights[1606]), .rectangle3_weight(rectangle3_weights[1606]), .feature_threshold(feature_thresholds[1606]), .feature_above(feature_aboves[1606]), .feature_below(feature_belows[1606]), .scan_win_std_dev(scan_win_std_dev[1606]), .feature_accum(feature_accums[1606]));
  accum_calculator ac1607(.scan_win(scan_win1607), .rectangle1_x(rectangle1_xs[1607]), .rectangle1_y(rectangle1_ys[1607]), .rectangle1_width(rectangle1_widths[1607]), .rectangle1_height(rectangle1_heights[1607]), .rectangle1_weight(rectangle1_weights[1607]), .rectangle2_x(rectangle2_xs[1607]), .rectangle2_y(rectangle2_ys[1607]), .rectangle2_width(rectangle2_widths[1607]), .rectangle2_height(rectangle2_heights[1607]), .rectangle2_weight(rectangle2_weights[1607]), .rectangle3_x(rectangle3_xs[1607]), .rectangle3_y(rectangle3_ys[1607]), .rectangle3_width(rectangle3_widths[1607]), .rectangle3_height(rectangle3_heights[1607]), .rectangle3_weight(rectangle3_weights[1607]), .feature_threshold(feature_thresholds[1607]), .feature_above(feature_aboves[1607]), .feature_below(feature_belows[1607]), .scan_win_std_dev(scan_win_std_dev[1607]), .feature_accum(feature_accums[1607]));
  accum_calculator ac1608(.scan_win(scan_win1608), .rectangle1_x(rectangle1_xs[1608]), .rectangle1_y(rectangle1_ys[1608]), .rectangle1_width(rectangle1_widths[1608]), .rectangle1_height(rectangle1_heights[1608]), .rectangle1_weight(rectangle1_weights[1608]), .rectangle2_x(rectangle2_xs[1608]), .rectangle2_y(rectangle2_ys[1608]), .rectangle2_width(rectangle2_widths[1608]), .rectangle2_height(rectangle2_heights[1608]), .rectangle2_weight(rectangle2_weights[1608]), .rectangle3_x(rectangle3_xs[1608]), .rectangle3_y(rectangle3_ys[1608]), .rectangle3_width(rectangle3_widths[1608]), .rectangle3_height(rectangle3_heights[1608]), .rectangle3_weight(rectangle3_weights[1608]), .feature_threshold(feature_thresholds[1608]), .feature_above(feature_aboves[1608]), .feature_below(feature_belows[1608]), .scan_win_std_dev(scan_win_std_dev[1608]), .feature_accum(feature_accums[1608]));
  accum_calculator ac1609(.scan_win(scan_win1609), .rectangle1_x(rectangle1_xs[1609]), .rectangle1_y(rectangle1_ys[1609]), .rectangle1_width(rectangle1_widths[1609]), .rectangle1_height(rectangle1_heights[1609]), .rectangle1_weight(rectangle1_weights[1609]), .rectangle2_x(rectangle2_xs[1609]), .rectangle2_y(rectangle2_ys[1609]), .rectangle2_width(rectangle2_widths[1609]), .rectangle2_height(rectangle2_heights[1609]), .rectangle2_weight(rectangle2_weights[1609]), .rectangle3_x(rectangle3_xs[1609]), .rectangle3_y(rectangle3_ys[1609]), .rectangle3_width(rectangle3_widths[1609]), .rectangle3_height(rectangle3_heights[1609]), .rectangle3_weight(rectangle3_weights[1609]), .feature_threshold(feature_thresholds[1609]), .feature_above(feature_aboves[1609]), .feature_below(feature_belows[1609]), .scan_win_std_dev(scan_win_std_dev[1609]), .feature_accum(feature_accums[1609]));
  accum_calculator ac1610(.scan_win(scan_win1610), .rectangle1_x(rectangle1_xs[1610]), .rectangle1_y(rectangle1_ys[1610]), .rectangle1_width(rectangle1_widths[1610]), .rectangle1_height(rectangle1_heights[1610]), .rectangle1_weight(rectangle1_weights[1610]), .rectangle2_x(rectangle2_xs[1610]), .rectangle2_y(rectangle2_ys[1610]), .rectangle2_width(rectangle2_widths[1610]), .rectangle2_height(rectangle2_heights[1610]), .rectangle2_weight(rectangle2_weights[1610]), .rectangle3_x(rectangle3_xs[1610]), .rectangle3_y(rectangle3_ys[1610]), .rectangle3_width(rectangle3_widths[1610]), .rectangle3_height(rectangle3_heights[1610]), .rectangle3_weight(rectangle3_weights[1610]), .feature_threshold(feature_thresholds[1610]), .feature_above(feature_aboves[1610]), .feature_below(feature_belows[1610]), .scan_win_std_dev(scan_win_std_dev[1610]), .feature_accum(feature_accums[1610]));
  accum_calculator ac1611(.scan_win(scan_win1611), .rectangle1_x(rectangle1_xs[1611]), .rectangle1_y(rectangle1_ys[1611]), .rectangle1_width(rectangle1_widths[1611]), .rectangle1_height(rectangle1_heights[1611]), .rectangle1_weight(rectangle1_weights[1611]), .rectangle2_x(rectangle2_xs[1611]), .rectangle2_y(rectangle2_ys[1611]), .rectangle2_width(rectangle2_widths[1611]), .rectangle2_height(rectangle2_heights[1611]), .rectangle2_weight(rectangle2_weights[1611]), .rectangle3_x(rectangle3_xs[1611]), .rectangle3_y(rectangle3_ys[1611]), .rectangle3_width(rectangle3_widths[1611]), .rectangle3_height(rectangle3_heights[1611]), .rectangle3_weight(rectangle3_weights[1611]), .feature_threshold(feature_thresholds[1611]), .feature_above(feature_aboves[1611]), .feature_below(feature_belows[1611]), .scan_win_std_dev(scan_win_std_dev[1611]), .feature_accum(feature_accums[1611]));
  accum_calculator ac1612(.scan_win(scan_win1612), .rectangle1_x(rectangle1_xs[1612]), .rectangle1_y(rectangle1_ys[1612]), .rectangle1_width(rectangle1_widths[1612]), .rectangle1_height(rectangle1_heights[1612]), .rectangle1_weight(rectangle1_weights[1612]), .rectangle2_x(rectangle2_xs[1612]), .rectangle2_y(rectangle2_ys[1612]), .rectangle2_width(rectangle2_widths[1612]), .rectangle2_height(rectangle2_heights[1612]), .rectangle2_weight(rectangle2_weights[1612]), .rectangle3_x(rectangle3_xs[1612]), .rectangle3_y(rectangle3_ys[1612]), .rectangle3_width(rectangle3_widths[1612]), .rectangle3_height(rectangle3_heights[1612]), .rectangle3_weight(rectangle3_weights[1612]), .feature_threshold(feature_thresholds[1612]), .feature_above(feature_aboves[1612]), .feature_below(feature_belows[1612]), .scan_win_std_dev(scan_win_std_dev[1612]), .feature_accum(feature_accums[1612]));
  accum_calculator ac1613(.scan_win(scan_win1613), .rectangle1_x(rectangle1_xs[1613]), .rectangle1_y(rectangle1_ys[1613]), .rectangle1_width(rectangle1_widths[1613]), .rectangle1_height(rectangle1_heights[1613]), .rectangle1_weight(rectangle1_weights[1613]), .rectangle2_x(rectangle2_xs[1613]), .rectangle2_y(rectangle2_ys[1613]), .rectangle2_width(rectangle2_widths[1613]), .rectangle2_height(rectangle2_heights[1613]), .rectangle2_weight(rectangle2_weights[1613]), .rectangle3_x(rectangle3_xs[1613]), .rectangle3_y(rectangle3_ys[1613]), .rectangle3_width(rectangle3_widths[1613]), .rectangle3_height(rectangle3_heights[1613]), .rectangle3_weight(rectangle3_weights[1613]), .feature_threshold(feature_thresholds[1613]), .feature_above(feature_aboves[1613]), .feature_below(feature_belows[1613]), .scan_win_std_dev(scan_win_std_dev[1613]), .feature_accum(feature_accums[1613]));
  accum_calculator ac1614(.scan_win(scan_win1614), .rectangle1_x(rectangle1_xs[1614]), .rectangle1_y(rectangle1_ys[1614]), .rectangle1_width(rectangle1_widths[1614]), .rectangle1_height(rectangle1_heights[1614]), .rectangle1_weight(rectangle1_weights[1614]), .rectangle2_x(rectangle2_xs[1614]), .rectangle2_y(rectangle2_ys[1614]), .rectangle2_width(rectangle2_widths[1614]), .rectangle2_height(rectangle2_heights[1614]), .rectangle2_weight(rectangle2_weights[1614]), .rectangle3_x(rectangle3_xs[1614]), .rectangle3_y(rectangle3_ys[1614]), .rectangle3_width(rectangle3_widths[1614]), .rectangle3_height(rectangle3_heights[1614]), .rectangle3_weight(rectangle3_weights[1614]), .feature_threshold(feature_thresholds[1614]), .feature_above(feature_aboves[1614]), .feature_below(feature_belows[1614]), .scan_win_std_dev(scan_win_std_dev[1614]), .feature_accum(feature_accums[1614]));
  accum_calculator ac1615(.scan_win(scan_win1615), .rectangle1_x(rectangle1_xs[1615]), .rectangle1_y(rectangle1_ys[1615]), .rectangle1_width(rectangle1_widths[1615]), .rectangle1_height(rectangle1_heights[1615]), .rectangle1_weight(rectangle1_weights[1615]), .rectangle2_x(rectangle2_xs[1615]), .rectangle2_y(rectangle2_ys[1615]), .rectangle2_width(rectangle2_widths[1615]), .rectangle2_height(rectangle2_heights[1615]), .rectangle2_weight(rectangle2_weights[1615]), .rectangle3_x(rectangle3_xs[1615]), .rectangle3_y(rectangle3_ys[1615]), .rectangle3_width(rectangle3_widths[1615]), .rectangle3_height(rectangle3_heights[1615]), .rectangle3_weight(rectangle3_weights[1615]), .feature_threshold(feature_thresholds[1615]), .feature_above(feature_aboves[1615]), .feature_below(feature_belows[1615]), .scan_win_std_dev(scan_win_std_dev[1615]), .feature_accum(feature_accums[1615]));
  accum_calculator ac1616(.scan_win(scan_win1616), .rectangle1_x(rectangle1_xs[1616]), .rectangle1_y(rectangle1_ys[1616]), .rectangle1_width(rectangle1_widths[1616]), .rectangle1_height(rectangle1_heights[1616]), .rectangle1_weight(rectangle1_weights[1616]), .rectangle2_x(rectangle2_xs[1616]), .rectangle2_y(rectangle2_ys[1616]), .rectangle2_width(rectangle2_widths[1616]), .rectangle2_height(rectangle2_heights[1616]), .rectangle2_weight(rectangle2_weights[1616]), .rectangle3_x(rectangle3_xs[1616]), .rectangle3_y(rectangle3_ys[1616]), .rectangle3_width(rectangle3_widths[1616]), .rectangle3_height(rectangle3_heights[1616]), .rectangle3_weight(rectangle3_weights[1616]), .feature_threshold(feature_thresholds[1616]), .feature_above(feature_aboves[1616]), .feature_below(feature_belows[1616]), .scan_win_std_dev(scan_win_std_dev[1616]), .feature_accum(feature_accums[1616]));
  accum_calculator ac1617(.scan_win(scan_win1617), .rectangle1_x(rectangle1_xs[1617]), .rectangle1_y(rectangle1_ys[1617]), .rectangle1_width(rectangle1_widths[1617]), .rectangle1_height(rectangle1_heights[1617]), .rectangle1_weight(rectangle1_weights[1617]), .rectangle2_x(rectangle2_xs[1617]), .rectangle2_y(rectangle2_ys[1617]), .rectangle2_width(rectangle2_widths[1617]), .rectangle2_height(rectangle2_heights[1617]), .rectangle2_weight(rectangle2_weights[1617]), .rectangle3_x(rectangle3_xs[1617]), .rectangle3_y(rectangle3_ys[1617]), .rectangle3_width(rectangle3_widths[1617]), .rectangle3_height(rectangle3_heights[1617]), .rectangle3_weight(rectangle3_weights[1617]), .feature_threshold(feature_thresholds[1617]), .feature_above(feature_aboves[1617]), .feature_below(feature_belows[1617]), .scan_win_std_dev(scan_win_std_dev[1617]), .feature_accum(feature_accums[1617]));
  accum_calculator ac1618(.scan_win(scan_win1618), .rectangle1_x(rectangle1_xs[1618]), .rectangle1_y(rectangle1_ys[1618]), .rectangle1_width(rectangle1_widths[1618]), .rectangle1_height(rectangle1_heights[1618]), .rectangle1_weight(rectangle1_weights[1618]), .rectangle2_x(rectangle2_xs[1618]), .rectangle2_y(rectangle2_ys[1618]), .rectangle2_width(rectangle2_widths[1618]), .rectangle2_height(rectangle2_heights[1618]), .rectangle2_weight(rectangle2_weights[1618]), .rectangle3_x(rectangle3_xs[1618]), .rectangle3_y(rectangle3_ys[1618]), .rectangle3_width(rectangle3_widths[1618]), .rectangle3_height(rectangle3_heights[1618]), .rectangle3_weight(rectangle3_weights[1618]), .feature_threshold(feature_thresholds[1618]), .feature_above(feature_aboves[1618]), .feature_below(feature_belows[1618]), .scan_win_std_dev(scan_win_std_dev[1618]), .feature_accum(feature_accums[1618]));
  accum_calculator ac1619(.scan_win(scan_win1619), .rectangle1_x(rectangle1_xs[1619]), .rectangle1_y(rectangle1_ys[1619]), .rectangle1_width(rectangle1_widths[1619]), .rectangle1_height(rectangle1_heights[1619]), .rectangle1_weight(rectangle1_weights[1619]), .rectangle2_x(rectangle2_xs[1619]), .rectangle2_y(rectangle2_ys[1619]), .rectangle2_width(rectangle2_widths[1619]), .rectangle2_height(rectangle2_heights[1619]), .rectangle2_weight(rectangle2_weights[1619]), .rectangle3_x(rectangle3_xs[1619]), .rectangle3_y(rectangle3_ys[1619]), .rectangle3_width(rectangle3_widths[1619]), .rectangle3_height(rectangle3_heights[1619]), .rectangle3_weight(rectangle3_weights[1619]), .feature_threshold(feature_thresholds[1619]), .feature_above(feature_aboves[1619]), .feature_below(feature_belows[1619]), .scan_win_std_dev(scan_win_std_dev[1619]), .feature_accum(feature_accums[1619]));
  accum_calculator ac1620(.scan_win(scan_win1620), .rectangle1_x(rectangle1_xs[1620]), .rectangle1_y(rectangle1_ys[1620]), .rectangle1_width(rectangle1_widths[1620]), .rectangle1_height(rectangle1_heights[1620]), .rectangle1_weight(rectangle1_weights[1620]), .rectangle2_x(rectangle2_xs[1620]), .rectangle2_y(rectangle2_ys[1620]), .rectangle2_width(rectangle2_widths[1620]), .rectangle2_height(rectangle2_heights[1620]), .rectangle2_weight(rectangle2_weights[1620]), .rectangle3_x(rectangle3_xs[1620]), .rectangle3_y(rectangle3_ys[1620]), .rectangle3_width(rectangle3_widths[1620]), .rectangle3_height(rectangle3_heights[1620]), .rectangle3_weight(rectangle3_weights[1620]), .feature_threshold(feature_thresholds[1620]), .feature_above(feature_aboves[1620]), .feature_below(feature_belows[1620]), .scan_win_std_dev(scan_win_std_dev[1620]), .feature_accum(feature_accums[1620]));
  accum_calculator ac1621(.scan_win(scan_win1621), .rectangle1_x(rectangle1_xs[1621]), .rectangle1_y(rectangle1_ys[1621]), .rectangle1_width(rectangle1_widths[1621]), .rectangle1_height(rectangle1_heights[1621]), .rectangle1_weight(rectangle1_weights[1621]), .rectangle2_x(rectangle2_xs[1621]), .rectangle2_y(rectangle2_ys[1621]), .rectangle2_width(rectangle2_widths[1621]), .rectangle2_height(rectangle2_heights[1621]), .rectangle2_weight(rectangle2_weights[1621]), .rectangle3_x(rectangle3_xs[1621]), .rectangle3_y(rectangle3_ys[1621]), .rectangle3_width(rectangle3_widths[1621]), .rectangle3_height(rectangle3_heights[1621]), .rectangle3_weight(rectangle3_weights[1621]), .feature_threshold(feature_thresholds[1621]), .feature_above(feature_aboves[1621]), .feature_below(feature_belows[1621]), .scan_win_std_dev(scan_win_std_dev[1621]), .feature_accum(feature_accums[1621]));
  accum_calculator ac1622(.scan_win(scan_win1622), .rectangle1_x(rectangle1_xs[1622]), .rectangle1_y(rectangle1_ys[1622]), .rectangle1_width(rectangle1_widths[1622]), .rectangle1_height(rectangle1_heights[1622]), .rectangle1_weight(rectangle1_weights[1622]), .rectangle2_x(rectangle2_xs[1622]), .rectangle2_y(rectangle2_ys[1622]), .rectangle2_width(rectangle2_widths[1622]), .rectangle2_height(rectangle2_heights[1622]), .rectangle2_weight(rectangle2_weights[1622]), .rectangle3_x(rectangle3_xs[1622]), .rectangle3_y(rectangle3_ys[1622]), .rectangle3_width(rectangle3_widths[1622]), .rectangle3_height(rectangle3_heights[1622]), .rectangle3_weight(rectangle3_weights[1622]), .feature_threshold(feature_thresholds[1622]), .feature_above(feature_aboves[1622]), .feature_below(feature_belows[1622]), .scan_win_std_dev(scan_win_std_dev[1622]), .feature_accum(feature_accums[1622]));
  accum_calculator ac1623(.scan_win(scan_win1623), .rectangle1_x(rectangle1_xs[1623]), .rectangle1_y(rectangle1_ys[1623]), .rectangle1_width(rectangle1_widths[1623]), .rectangle1_height(rectangle1_heights[1623]), .rectangle1_weight(rectangle1_weights[1623]), .rectangle2_x(rectangle2_xs[1623]), .rectangle2_y(rectangle2_ys[1623]), .rectangle2_width(rectangle2_widths[1623]), .rectangle2_height(rectangle2_heights[1623]), .rectangle2_weight(rectangle2_weights[1623]), .rectangle3_x(rectangle3_xs[1623]), .rectangle3_y(rectangle3_ys[1623]), .rectangle3_width(rectangle3_widths[1623]), .rectangle3_height(rectangle3_heights[1623]), .rectangle3_weight(rectangle3_weights[1623]), .feature_threshold(feature_thresholds[1623]), .feature_above(feature_aboves[1623]), .feature_below(feature_belows[1623]), .scan_win_std_dev(scan_win_std_dev[1623]), .feature_accum(feature_accums[1623]));
  accum_calculator ac1624(.scan_win(scan_win1624), .rectangle1_x(rectangle1_xs[1624]), .rectangle1_y(rectangle1_ys[1624]), .rectangle1_width(rectangle1_widths[1624]), .rectangle1_height(rectangle1_heights[1624]), .rectangle1_weight(rectangle1_weights[1624]), .rectangle2_x(rectangle2_xs[1624]), .rectangle2_y(rectangle2_ys[1624]), .rectangle2_width(rectangle2_widths[1624]), .rectangle2_height(rectangle2_heights[1624]), .rectangle2_weight(rectangle2_weights[1624]), .rectangle3_x(rectangle3_xs[1624]), .rectangle3_y(rectangle3_ys[1624]), .rectangle3_width(rectangle3_widths[1624]), .rectangle3_height(rectangle3_heights[1624]), .rectangle3_weight(rectangle3_weights[1624]), .feature_threshold(feature_thresholds[1624]), .feature_above(feature_aboves[1624]), .feature_below(feature_belows[1624]), .scan_win_std_dev(scan_win_std_dev[1624]), .feature_accum(feature_accums[1624]));
  accum_calculator ac1625(.scan_win(scan_win1625), .rectangle1_x(rectangle1_xs[1625]), .rectangle1_y(rectangle1_ys[1625]), .rectangle1_width(rectangle1_widths[1625]), .rectangle1_height(rectangle1_heights[1625]), .rectangle1_weight(rectangle1_weights[1625]), .rectangle2_x(rectangle2_xs[1625]), .rectangle2_y(rectangle2_ys[1625]), .rectangle2_width(rectangle2_widths[1625]), .rectangle2_height(rectangle2_heights[1625]), .rectangle2_weight(rectangle2_weights[1625]), .rectangle3_x(rectangle3_xs[1625]), .rectangle3_y(rectangle3_ys[1625]), .rectangle3_width(rectangle3_widths[1625]), .rectangle3_height(rectangle3_heights[1625]), .rectangle3_weight(rectangle3_weights[1625]), .feature_threshold(feature_thresholds[1625]), .feature_above(feature_aboves[1625]), .feature_below(feature_belows[1625]), .scan_win_std_dev(scan_win_std_dev[1625]), .feature_accum(feature_accums[1625]));
  accum_calculator ac1626(.scan_win(scan_win1626), .rectangle1_x(rectangle1_xs[1626]), .rectangle1_y(rectangle1_ys[1626]), .rectangle1_width(rectangle1_widths[1626]), .rectangle1_height(rectangle1_heights[1626]), .rectangle1_weight(rectangle1_weights[1626]), .rectangle2_x(rectangle2_xs[1626]), .rectangle2_y(rectangle2_ys[1626]), .rectangle2_width(rectangle2_widths[1626]), .rectangle2_height(rectangle2_heights[1626]), .rectangle2_weight(rectangle2_weights[1626]), .rectangle3_x(rectangle3_xs[1626]), .rectangle3_y(rectangle3_ys[1626]), .rectangle3_width(rectangle3_widths[1626]), .rectangle3_height(rectangle3_heights[1626]), .rectangle3_weight(rectangle3_weights[1626]), .feature_threshold(feature_thresholds[1626]), .feature_above(feature_aboves[1626]), .feature_below(feature_belows[1626]), .scan_win_std_dev(scan_win_std_dev[1626]), .feature_accum(feature_accums[1626]));
  accum_calculator ac1627(.scan_win(scan_win1627), .rectangle1_x(rectangle1_xs[1627]), .rectangle1_y(rectangle1_ys[1627]), .rectangle1_width(rectangle1_widths[1627]), .rectangle1_height(rectangle1_heights[1627]), .rectangle1_weight(rectangle1_weights[1627]), .rectangle2_x(rectangle2_xs[1627]), .rectangle2_y(rectangle2_ys[1627]), .rectangle2_width(rectangle2_widths[1627]), .rectangle2_height(rectangle2_heights[1627]), .rectangle2_weight(rectangle2_weights[1627]), .rectangle3_x(rectangle3_xs[1627]), .rectangle3_y(rectangle3_ys[1627]), .rectangle3_width(rectangle3_widths[1627]), .rectangle3_height(rectangle3_heights[1627]), .rectangle3_weight(rectangle3_weights[1627]), .feature_threshold(feature_thresholds[1627]), .feature_above(feature_aboves[1627]), .feature_below(feature_belows[1627]), .scan_win_std_dev(scan_win_std_dev[1627]), .feature_accum(feature_accums[1627]));
  accum_calculator ac1628(.scan_win(scan_win1628), .rectangle1_x(rectangle1_xs[1628]), .rectangle1_y(rectangle1_ys[1628]), .rectangle1_width(rectangle1_widths[1628]), .rectangle1_height(rectangle1_heights[1628]), .rectangle1_weight(rectangle1_weights[1628]), .rectangle2_x(rectangle2_xs[1628]), .rectangle2_y(rectangle2_ys[1628]), .rectangle2_width(rectangle2_widths[1628]), .rectangle2_height(rectangle2_heights[1628]), .rectangle2_weight(rectangle2_weights[1628]), .rectangle3_x(rectangle3_xs[1628]), .rectangle3_y(rectangle3_ys[1628]), .rectangle3_width(rectangle3_widths[1628]), .rectangle3_height(rectangle3_heights[1628]), .rectangle3_weight(rectangle3_weights[1628]), .feature_threshold(feature_thresholds[1628]), .feature_above(feature_aboves[1628]), .feature_below(feature_belows[1628]), .scan_win_std_dev(scan_win_std_dev[1628]), .feature_accum(feature_accums[1628]));
  accum_calculator ac1629(.scan_win(scan_win1629), .rectangle1_x(rectangle1_xs[1629]), .rectangle1_y(rectangle1_ys[1629]), .rectangle1_width(rectangle1_widths[1629]), .rectangle1_height(rectangle1_heights[1629]), .rectangle1_weight(rectangle1_weights[1629]), .rectangle2_x(rectangle2_xs[1629]), .rectangle2_y(rectangle2_ys[1629]), .rectangle2_width(rectangle2_widths[1629]), .rectangle2_height(rectangle2_heights[1629]), .rectangle2_weight(rectangle2_weights[1629]), .rectangle3_x(rectangle3_xs[1629]), .rectangle3_y(rectangle3_ys[1629]), .rectangle3_width(rectangle3_widths[1629]), .rectangle3_height(rectangle3_heights[1629]), .rectangle3_weight(rectangle3_weights[1629]), .feature_threshold(feature_thresholds[1629]), .feature_above(feature_aboves[1629]), .feature_below(feature_belows[1629]), .scan_win_std_dev(scan_win_std_dev[1629]), .feature_accum(feature_accums[1629]));
  accum_calculator ac1630(.scan_win(scan_win1630), .rectangle1_x(rectangle1_xs[1630]), .rectangle1_y(rectangle1_ys[1630]), .rectangle1_width(rectangle1_widths[1630]), .rectangle1_height(rectangle1_heights[1630]), .rectangle1_weight(rectangle1_weights[1630]), .rectangle2_x(rectangle2_xs[1630]), .rectangle2_y(rectangle2_ys[1630]), .rectangle2_width(rectangle2_widths[1630]), .rectangle2_height(rectangle2_heights[1630]), .rectangle2_weight(rectangle2_weights[1630]), .rectangle3_x(rectangle3_xs[1630]), .rectangle3_y(rectangle3_ys[1630]), .rectangle3_width(rectangle3_widths[1630]), .rectangle3_height(rectangle3_heights[1630]), .rectangle3_weight(rectangle3_weights[1630]), .feature_threshold(feature_thresholds[1630]), .feature_above(feature_aboves[1630]), .feature_below(feature_belows[1630]), .scan_win_std_dev(scan_win_std_dev[1630]), .feature_accum(feature_accums[1630]));
  accum_calculator ac1631(.scan_win(scan_win1631), .rectangle1_x(rectangle1_xs[1631]), .rectangle1_y(rectangle1_ys[1631]), .rectangle1_width(rectangle1_widths[1631]), .rectangle1_height(rectangle1_heights[1631]), .rectangle1_weight(rectangle1_weights[1631]), .rectangle2_x(rectangle2_xs[1631]), .rectangle2_y(rectangle2_ys[1631]), .rectangle2_width(rectangle2_widths[1631]), .rectangle2_height(rectangle2_heights[1631]), .rectangle2_weight(rectangle2_weights[1631]), .rectangle3_x(rectangle3_xs[1631]), .rectangle3_y(rectangle3_ys[1631]), .rectangle3_width(rectangle3_widths[1631]), .rectangle3_height(rectangle3_heights[1631]), .rectangle3_weight(rectangle3_weights[1631]), .feature_threshold(feature_thresholds[1631]), .feature_above(feature_aboves[1631]), .feature_below(feature_belows[1631]), .scan_win_std_dev(scan_win_std_dev[1631]), .feature_accum(feature_accums[1631]));
  accum_calculator ac1632(.scan_win(scan_win1632), .rectangle1_x(rectangle1_xs[1632]), .rectangle1_y(rectangle1_ys[1632]), .rectangle1_width(rectangle1_widths[1632]), .rectangle1_height(rectangle1_heights[1632]), .rectangle1_weight(rectangle1_weights[1632]), .rectangle2_x(rectangle2_xs[1632]), .rectangle2_y(rectangle2_ys[1632]), .rectangle2_width(rectangle2_widths[1632]), .rectangle2_height(rectangle2_heights[1632]), .rectangle2_weight(rectangle2_weights[1632]), .rectangle3_x(rectangle3_xs[1632]), .rectangle3_y(rectangle3_ys[1632]), .rectangle3_width(rectangle3_widths[1632]), .rectangle3_height(rectangle3_heights[1632]), .rectangle3_weight(rectangle3_weights[1632]), .feature_threshold(feature_thresholds[1632]), .feature_above(feature_aboves[1632]), .feature_below(feature_belows[1632]), .scan_win_std_dev(scan_win_std_dev[1632]), .feature_accum(feature_accums[1632]));
  accum_calculator ac1633(.scan_win(scan_win1633), .rectangle1_x(rectangle1_xs[1633]), .rectangle1_y(rectangle1_ys[1633]), .rectangle1_width(rectangle1_widths[1633]), .rectangle1_height(rectangle1_heights[1633]), .rectangle1_weight(rectangle1_weights[1633]), .rectangle2_x(rectangle2_xs[1633]), .rectangle2_y(rectangle2_ys[1633]), .rectangle2_width(rectangle2_widths[1633]), .rectangle2_height(rectangle2_heights[1633]), .rectangle2_weight(rectangle2_weights[1633]), .rectangle3_x(rectangle3_xs[1633]), .rectangle3_y(rectangle3_ys[1633]), .rectangle3_width(rectangle3_widths[1633]), .rectangle3_height(rectangle3_heights[1633]), .rectangle3_weight(rectangle3_weights[1633]), .feature_threshold(feature_thresholds[1633]), .feature_above(feature_aboves[1633]), .feature_below(feature_belows[1633]), .scan_win_std_dev(scan_win_std_dev[1633]), .feature_accum(feature_accums[1633]));
  accum_calculator ac1634(.scan_win(scan_win1634), .rectangle1_x(rectangle1_xs[1634]), .rectangle1_y(rectangle1_ys[1634]), .rectangle1_width(rectangle1_widths[1634]), .rectangle1_height(rectangle1_heights[1634]), .rectangle1_weight(rectangle1_weights[1634]), .rectangle2_x(rectangle2_xs[1634]), .rectangle2_y(rectangle2_ys[1634]), .rectangle2_width(rectangle2_widths[1634]), .rectangle2_height(rectangle2_heights[1634]), .rectangle2_weight(rectangle2_weights[1634]), .rectangle3_x(rectangle3_xs[1634]), .rectangle3_y(rectangle3_ys[1634]), .rectangle3_width(rectangle3_widths[1634]), .rectangle3_height(rectangle3_heights[1634]), .rectangle3_weight(rectangle3_weights[1634]), .feature_threshold(feature_thresholds[1634]), .feature_above(feature_aboves[1634]), .feature_below(feature_belows[1634]), .scan_win_std_dev(scan_win_std_dev[1634]), .feature_accum(feature_accums[1634]));
  accum_calculator ac1635(.scan_win(scan_win1635), .rectangle1_x(rectangle1_xs[1635]), .rectangle1_y(rectangle1_ys[1635]), .rectangle1_width(rectangle1_widths[1635]), .rectangle1_height(rectangle1_heights[1635]), .rectangle1_weight(rectangle1_weights[1635]), .rectangle2_x(rectangle2_xs[1635]), .rectangle2_y(rectangle2_ys[1635]), .rectangle2_width(rectangle2_widths[1635]), .rectangle2_height(rectangle2_heights[1635]), .rectangle2_weight(rectangle2_weights[1635]), .rectangle3_x(rectangle3_xs[1635]), .rectangle3_y(rectangle3_ys[1635]), .rectangle3_width(rectangle3_widths[1635]), .rectangle3_height(rectangle3_heights[1635]), .rectangle3_weight(rectangle3_weights[1635]), .feature_threshold(feature_thresholds[1635]), .feature_above(feature_aboves[1635]), .feature_below(feature_belows[1635]), .scan_win_std_dev(scan_win_std_dev[1635]), .feature_accum(feature_accums[1635]));
  accum_calculator ac1636(.scan_win(scan_win1636), .rectangle1_x(rectangle1_xs[1636]), .rectangle1_y(rectangle1_ys[1636]), .rectangle1_width(rectangle1_widths[1636]), .rectangle1_height(rectangle1_heights[1636]), .rectangle1_weight(rectangle1_weights[1636]), .rectangle2_x(rectangle2_xs[1636]), .rectangle2_y(rectangle2_ys[1636]), .rectangle2_width(rectangle2_widths[1636]), .rectangle2_height(rectangle2_heights[1636]), .rectangle2_weight(rectangle2_weights[1636]), .rectangle3_x(rectangle3_xs[1636]), .rectangle3_y(rectangle3_ys[1636]), .rectangle3_width(rectangle3_widths[1636]), .rectangle3_height(rectangle3_heights[1636]), .rectangle3_weight(rectangle3_weights[1636]), .feature_threshold(feature_thresholds[1636]), .feature_above(feature_aboves[1636]), .feature_below(feature_belows[1636]), .scan_win_std_dev(scan_win_std_dev[1636]), .feature_accum(feature_accums[1636]));
  accum_calculator ac1637(.scan_win(scan_win1637), .rectangle1_x(rectangle1_xs[1637]), .rectangle1_y(rectangle1_ys[1637]), .rectangle1_width(rectangle1_widths[1637]), .rectangle1_height(rectangle1_heights[1637]), .rectangle1_weight(rectangle1_weights[1637]), .rectangle2_x(rectangle2_xs[1637]), .rectangle2_y(rectangle2_ys[1637]), .rectangle2_width(rectangle2_widths[1637]), .rectangle2_height(rectangle2_heights[1637]), .rectangle2_weight(rectangle2_weights[1637]), .rectangle3_x(rectangle3_xs[1637]), .rectangle3_y(rectangle3_ys[1637]), .rectangle3_width(rectangle3_widths[1637]), .rectangle3_height(rectangle3_heights[1637]), .rectangle3_weight(rectangle3_weights[1637]), .feature_threshold(feature_thresholds[1637]), .feature_above(feature_aboves[1637]), .feature_below(feature_belows[1637]), .scan_win_std_dev(scan_win_std_dev[1637]), .feature_accum(feature_accums[1637]));
  accum_calculator ac1638(.scan_win(scan_win1638), .rectangle1_x(rectangle1_xs[1638]), .rectangle1_y(rectangle1_ys[1638]), .rectangle1_width(rectangle1_widths[1638]), .rectangle1_height(rectangle1_heights[1638]), .rectangle1_weight(rectangle1_weights[1638]), .rectangle2_x(rectangle2_xs[1638]), .rectangle2_y(rectangle2_ys[1638]), .rectangle2_width(rectangle2_widths[1638]), .rectangle2_height(rectangle2_heights[1638]), .rectangle2_weight(rectangle2_weights[1638]), .rectangle3_x(rectangle3_xs[1638]), .rectangle3_y(rectangle3_ys[1638]), .rectangle3_width(rectangle3_widths[1638]), .rectangle3_height(rectangle3_heights[1638]), .rectangle3_weight(rectangle3_weights[1638]), .feature_threshold(feature_thresholds[1638]), .feature_above(feature_aboves[1638]), .feature_below(feature_belows[1638]), .scan_win_std_dev(scan_win_std_dev[1638]), .feature_accum(feature_accums[1638]));
  accum_calculator ac1639(.scan_win(scan_win1639), .rectangle1_x(rectangle1_xs[1639]), .rectangle1_y(rectangle1_ys[1639]), .rectangle1_width(rectangle1_widths[1639]), .rectangle1_height(rectangle1_heights[1639]), .rectangle1_weight(rectangle1_weights[1639]), .rectangle2_x(rectangle2_xs[1639]), .rectangle2_y(rectangle2_ys[1639]), .rectangle2_width(rectangle2_widths[1639]), .rectangle2_height(rectangle2_heights[1639]), .rectangle2_weight(rectangle2_weights[1639]), .rectangle3_x(rectangle3_xs[1639]), .rectangle3_y(rectangle3_ys[1639]), .rectangle3_width(rectangle3_widths[1639]), .rectangle3_height(rectangle3_heights[1639]), .rectangle3_weight(rectangle3_weights[1639]), .feature_threshold(feature_thresholds[1639]), .feature_above(feature_aboves[1639]), .feature_below(feature_belows[1639]), .scan_win_std_dev(scan_win_std_dev[1639]), .feature_accum(feature_accums[1639]));
  accum_calculator ac1640(.scan_win(scan_win1640), .rectangle1_x(rectangle1_xs[1640]), .rectangle1_y(rectangle1_ys[1640]), .rectangle1_width(rectangle1_widths[1640]), .rectangle1_height(rectangle1_heights[1640]), .rectangle1_weight(rectangle1_weights[1640]), .rectangle2_x(rectangle2_xs[1640]), .rectangle2_y(rectangle2_ys[1640]), .rectangle2_width(rectangle2_widths[1640]), .rectangle2_height(rectangle2_heights[1640]), .rectangle2_weight(rectangle2_weights[1640]), .rectangle3_x(rectangle3_xs[1640]), .rectangle3_y(rectangle3_ys[1640]), .rectangle3_width(rectangle3_widths[1640]), .rectangle3_height(rectangle3_heights[1640]), .rectangle3_weight(rectangle3_weights[1640]), .feature_threshold(feature_thresholds[1640]), .feature_above(feature_aboves[1640]), .feature_below(feature_belows[1640]), .scan_win_std_dev(scan_win_std_dev[1640]), .feature_accum(feature_accums[1640]));
  accum_calculator ac1641(.scan_win(scan_win1641), .rectangle1_x(rectangle1_xs[1641]), .rectangle1_y(rectangle1_ys[1641]), .rectangle1_width(rectangle1_widths[1641]), .rectangle1_height(rectangle1_heights[1641]), .rectangle1_weight(rectangle1_weights[1641]), .rectangle2_x(rectangle2_xs[1641]), .rectangle2_y(rectangle2_ys[1641]), .rectangle2_width(rectangle2_widths[1641]), .rectangle2_height(rectangle2_heights[1641]), .rectangle2_weight(rectangle2_weights[1641]), .rectangle3_x(rectangle3_xs[1641]), .rectangle3_y(rectangle3_ys[1641]), .rectangle3_width(rectangle3_widths[1641]), .rectangle3_height(rectangle3_heights[1641]), .rectangle3_weight(rectangle3_weights[1641]), .feature_threshold(feature_thresholds[1641]), .feature_above(feature_aboves[1641]), .feature_below(feature_belows[1641]), .scan_win_std_dev(scan_win_std_dev[1641]), .feature_accum(feature_accums[1641]));
  accum_calculator ac1642(.scan_win(scan_win1642), .rectangle1_x(rectangle1_xs[1642]), .rectangle1_y(rectangle1_ys[1642]), .rectangle1_width(rectangle1_widths[1642]), .rectangle1_height(rectangle1_heights[1642]), .rectangle1_weight(rectangle1_weights[1642]), .rectangle2_x(rectangle2_xs[1642]), .rectangle2_y(rectangle2_ys[1642]), .rectangle2_width(rectangle2_widths[1642]), .rectangle2_height(rectangle2_heights[1642]), .rectangle2_weight(rectangle2_weights[1642]), .rectangle3_x(rectangle3_xs[1642]), .rectangle3_y(rectangle3_ys[1642]), .rectangle3_width(rectangle3_widths[1642]), .rectangle3_height(rectangle3_heights[1642]), .rectangle3_weight(rectangle3_weights[1642]), .feature_threshold(feature_thresholds[1642]), .feature_above(feature_aboves[1642]), .feature_below(feature_belows[1642]), .scan_win_std_dev(scan_win_std_dev[1642]), .feature_accum(feature_accums[1642]));
  accum_calculator ac1643(.scan_win(scan_win1643), .rectangle1_x(rectangle1_xs[1643]), .rectangle1_y(rectangle1_ys[1643]), .rectangle1_width(rectangle1_widths[1643]), .rectangle1_height(rectangle1_heights[1643]), .rectangle1_weight(rectangle1_weights[1643]), .rectangle2_x(rectangle2_xs[1643]), .rectangle2_y(rectangle2_ys[1643]), .rectangle2_width(rectangle2_widths[1643]), .rectangle2_height(rectangle2_heights[1643]), .rectangle2_weight(rectangle2_weights[1643]), .rectangle3_x(rectangle3_xs[1643]), .rectangle3_y(rectangle3_ys[1643]), .rectangle3_width(rectangle3_widths[1643]), .rectangle3_height(rectangle3_heights[1643]), .rectangle3_weight(rectangle3_weights[1643]), .feature_threshold(feature_thresholds[1643]), .feature_above(feature_aboves[1643]), .feature_below(feature_belows[1643]), .scan_win_std_dev(scan_win_std_dev[1643]), .feature_accum(feature_accums[1643]));
  accum_calculator ac1644(.scan_win(scan_win1644), .rectangle1_x(rectangle1_xs[1644]), .rectangle1_y(rectangle1_ys[1644]), .rectangle1_width(rectangle1_widths[1644]), .rectangle1_height(rectangle1_heights[1644]), .rectangle1_weight(rectangle1_weights[1644]), .rectangle2_x(rectangle2_xs[1644]), .rectangle2_y(rectangle2_ys[1644]), .rectangle2_width(rectangle2_widths[1644]), .rectangle2_height(rectangle2_heights[1644]), .rectangle2_weight(rectangle2_weights[1644]), .rectangle3_x(rectangle3_xs[1644]), .rectangle3_y(rectangle3_ys[1644]), .rectangle3_width(rectangle3_widths[1644]), .rectangle3_height(rectangle3_heights[1644]), .rectangle3_weight(rectangle3_weights[1644]), .feature_threshold(feature_thresholds[1644]), .feature_above(feature_aboves[1644]), .feature_below(feature_belows[1644]), .scan_win_std_dev(scan_win_std_dev[1644]), .feature_accum(feature_accums[1644]));
  accum_calculator ac1645(.scan_win(scan_win1645), .rectangle1_x(rectangle1_xs[1645]), .rectangle1_y(rectangle1_ys[1645]), .rectangle1_width(rectangle1_widths[1645]), .rectangle1_height(rectangle1_heights[1645]), .rectangle1_weight(rectangle1_weights[1645]), .rectangle2_x(rectangle2_xs[1645]), .rectangle2_y(rectangle2_ys[1645]), .rectangle2_width(rectangle2_widths[1645]), .rectangle2_height(rectangle2_heights[1645]), .rectangle2_weight(rectangle2_weights[1645]), .rectangle3_x(rectangle3_xs[1645]), .rectangle3_y(rectangle3_ys[1645]), .rectangle3_width(rectangle3_widths[1645]), .rectangle3_height(rectangle3_heights[1645]), .rectangle3_weight(rectangle3_weights[1645]), .feature_threshold(feature_thresholds[1645]), .feature_above(feature_aboves[1645]), .feature_below(feature_belows[1645]), .scan_win_std_dev(scan_win_std_dev[1645]), .feature_accum(feature_accums[1645]));
  accum_calculator ac1646(.scan_win(scan_win1646), .rectangle1_x(rectangle1_xs[1646]), .rectangle1_y(rectangle1_ys[1646]), .rectangle1_width(rectangle1_widths[1646]), .rectangle1_height(rectangle1_heights[1646]), .rectangle1_weight(rectangle1_weights[1646]), .rectangle2_x(rectangle2_xs[1646]), .rectangle2_y(rectangle2_ys[1646]), .rectangle2_width(rectangle2_widths[1646]), .rectangle2_height(rectangle2_heights[1646]), .rectangle2_weight(rectangle2_weights[1646]), .rectangle3_x(rectangle3_xs[1646]), .rectangle3_y(rectangle3_ys[1646]), .rectangle3_width(rectangle3_widths[1646]), .rectangle3_height(rectangle3_heights[1646]), .rectangle3_weight(rectangle3_weights[1646]), .feature_threshold(feature_thresholds[1646]), .feature_above(feature_aboves[1646]), .feature_below(feature_belows[1646]), .scan_win_std_dev(scan_win_std_dev[1646]), .feature_accum(feature_accums[1646]));
  accum_calculator ac1647(.scan_win(scan_win1647), .rectangle1_x(rectangle1_xs[1647]), .rectangle1_y(rectangle1_ys[1647]), .rectangle1_width(rectangle1_widths[1647]), .rectangle1_height(rectangle1_heights[1647]), .rectangle1_weight(rectangle1_weights[1647]), .rectangle2_x(rectangle2_xs[1647]), .rectangle2_y(rectangle2_ys[1647]), .rectangle2_width(rectangle2_widths[1647]), .rectangle2_height(rectangle2_heights[1647]), .rectangle2_weight(rectangle2_weights[1647]), .rectangle3_x(rectangle3_xs[1647]), .rectangle3_y(rectangle3_ys[1647]), .rectangle3_width(rectangle3_widths[1647]), .rectangle3_height(rectangle3_heights[1647]), .rectangle3_weight(rectangle3_weights[1647]), .feature_threshold(feature_thresholds[1647]), .feature_above(feature_aboves[1647]), .feature_below(feature_belows[1647]), .scan_win_std_dev(scan_win_std_dev[1647]), .feature_accum(feature_accums[1647]));
  accum_calculator ac1648(.scan_win(scan_win1648), .rectangle1_x(rectangle1_xs[1648]), .rectangle1_y(rectangle1_ys[1648]), .rectangle1_width(rectangle1_widths[1648]), .rectangle1_height(rectangle1_heights[1648]), .rectangle1_weight(rectangle1_weights[1648]), .rectangle2_x(rectangle2_xs[1648]), .rectangle2_y(rectangle2_ys[1648]), .rectangle2_width(rectangle2_widths[1648]), .rectangle2_height(rectangle2_heights[1648]), .rectangle2_weight(rectangle2_weights[1648]), .rectangle3_x(rectangle3_xs[1648]), .rectangle3_y(rectangle3_ys[1648]), .rectangle3_width(rectangle3_widths[1648]), .rectangle3_height(rectangle3_heights[1648]), .rectangle3_weight(rectangle3_weights[1648]), .feature_threshold(feature_thresholds[1648]), .feature_above(feature_aboves[1648]), .feature_below(feature_belows[1648]), .scan_win_std_dev(scan_win_std_dev[1648]), .feature_accum(feature_accums[1648]));
  accum_calculator ac1649(.scan_win(scan_win1649), .rectangle1_x(rectangle1_xs[1649]), .rectangle1_y(rectangle1_ys[1649]), .rectangle1_width(rectangle1_widths[1649]), .rectangle1_height(rectangle1_heights[1649]), .rectangle1_weight(rectangle1_weights[1649]), .rectangle2_x(rectangle2_xs[1649]), .rectangle2_y(rectangle2_ys[1649]), .rectangle2_width(rectangle2_widths[1649]), .rectangle2_height(rectangle2_heights[1649]), .rectangle2_weight(rectangle2_weights[1649]), .rectangle3_x(rectangle3_xs[1649]), .rectangle3_y(rectangle3_ys[1649]), .rectangle3_width(rectangle3_widths[1649]), .rectangle3_height(rectangle3_heights[1649]), .rectangle3_weight(rectangle3_weights[1649]), .feature_threshold(feature_thresholds[1649]), .feature_above(feature_aboves[1649]), .feature_below(feature_belows[1649]), .scan_win_std_dev(scan_win_std_dev[1649]), .feature_accum(feature_accums[1649]));
  accum_calculator ac1650(.scan_win(scan_win1650), .rectangle1_x(rectangle1_xs[1650]), .rectangle1_y(rectangle1_ys[1650]), .rectangle1_width(rectangle1_widths[1650]), .rectangle1_height(rectangle1_heights[1650]), .rectangle1_weight(rectangle1_weights[1650]), .rectangle2_x(rectangle2_xs[1650]), .rectangle2_y(rectangle2_ys[1650]), .rectangle2_width(rectangle2_widths[1650]), .rectangle2_height(rectangle2_heights[1650]), .rectangle2_weight(rectangle2_weights[1650]), .rectangle3_x(rectangle3_xs[1650]), .rectangle3_y(rectangle3_ys[1650]), .rectangle3_width(rectangle3_widths[1650]), .rectangle3_height(rectangle3_heights[1650]), .rectangle3_weight(rectangle3_weights[1650]), .feature_threshold(feature_thresholds[1650]), .feature_above(feature_aboves[1650]), .feature_below(feature_belows[1650]), .scan_win_std_dev(scan_win_std_dev[1650]), .feature_accum(feature_accums[1650]));
  accum_calculator ac1651(.scan_win(scan_win1651), .rectangle1_x(rectangle1_xs[1651]), .rectangle1_y(rectangle1_ys[1651]), .rectangle1_width(rectangle1_widths[1651]), .rectangle1_height(rectangle1_heights[1651]), .rectangle1_weight(rectangle1_weights[1651]), .rectangle2_x(rectangle2_xs[1651]), .rectangle2_y(rectangle2_ys[1651]), .rectangle2_width(rectangle2_widths[1651]), .rectangle2_height(rectangle2_heights[1651]), .rectangle2_weight(rectangle2_weights[1651]), .rectangle3_x(rectangle3_xs[1651]), .rectangle3_y(rectangle3_ys[1651]), .rectangle3_width(rectangle3_widths[1651]), .rectangle3_height(rectangle3_heights[1651]), .rectangle3_weight(rectangle3_weights[1651]), .feature_threshold(feature_thresholds[1651]), .feature_above(feature_aboves[1651]), .feature_below(feature_belows[1651]), .scan_win_std_dev(scan_win_std_dev[1651]), .feature_accum(feature_accums[1651]));
  accum_calculator ac1652(.scan_win(scan_win1652), .rectangle1_x(rectangle1_xs[1652]), .rectangle1_y(rectangle1_ys[1652]), .rectangle1_width(rectangle1_widths[1652]), .rectangle1_height(rectangle1_heights[1652]), .rectangle1_weight(rectangle1_weights[1652]), .rectangle2_x(rectangle2_xs[1652]), .rectangle2_y(rectangle2_ys[1652]), .rectangle2_width(rectangle2_widths[1652]), .rectangle2_height(rectangle2_heights[1652]), .rectangle2_weight(rectangle2_weights[1652]), .rectangle3_x(rectangle3_xs[1652]), .rectangle3_y(rectangle3_ys[1652]), .rectangle3_width(rectangle3_widths[1652]), .rectangle3_height(rectangle3_heights[1652]), .rectangle3_weight(rectangle3_weights[1652]), .feature_threshold(feature_thresholds[1652]), .feature_above(feature_aboves[1652]), .feature_below(feature_belows[1652]), .scan_win_std_dev(scan_win_std_dev[1652]), .feature_accum(feature_accums[1652]));
  accum_calculator ac1653(.scan_win(scan_win1653), .rectangle1_x(rectangle1_xs[1653]), .rectangle1_y(rectangle1_ys[1653]), .rectangle1_width(rectangle1_widths[1653]), .rectangle1_height(rectangle1_heights[1653]), .rectangle1_weight(rectangle1_weights[1653]), .rectangle2_x(rectangle2_xs[1653]), .rectangle2_y(rectangle2_ys[1653]), .rectangle2_width(rectangle2_widths[1653]), .rectangle2_height(rectangle2_heights[1653]), .rectangle2_weight(rectangle2_weights[1653]), .rectangle3_x(rectangle3_xs[1653]), .rectangle3_y(rectangle3_ys[1653]), .rectangle3_width(rectangle3_widths[1653]), .rectangle3_height(rectangle3_heights[1653]), .rectangle3_weight(rectangle3_weights[1653]), .feature_threshold(feature_thresholds[1653]), .feature_above(feature_aboves[1653]), .feature_below(feature_belows[1653]), .scan_win_std_dev(scan_win_std_dev[1653]), .feature_accum(feature_accums[1653]));
  accum_calculator ac1654(.scan_win(scan_win1654), .rectangle1_x(rectangle1_xs[1654]), .rectangle1_y(rectangle1_ys[1654]), .rectangle1_width(rectangle1_widths[1654]), .rectangle1_height(rectangle1_heights[1654]), .rectangle1_weight(rectangle1_weights[1654]), .rectangle2_x(rectangle2_xs[1654]), .rectangle2_y(rectangle2_ys[1654]), .rectangle2_width(rectangle2_widths[1654]), .rectangle2_height(rectangle2_heights[1654]), .rectangle2_weight(rectangle2_weights[1654]), .rectangle3_x(rectangle3_xs[1654]), .rectangle3_y(rectangle3_ys[1654]), .rectangle3_width(rectangle3_widths[1654]), .rectangle3_height(rectangle3_heights[1654]), .rectangle3_weight(rectangle3_weights[1654]), .feature_threshold(feature_thresholds[1654]), .feature_above(feature_aboves[1654]), .feature_below(feature_belows[1654]), .scan_win_std_dev(scan_win_std_dev[1654]), .feature_accum(feature_accums[1654]));
  accum_calculator ac1655(.scan_win(scan_win1655), .rectangle1_x(rectangle1_xs[1655]), .rectangle1_y(rectangle1_ys[1655]), .rectangle1_width(rectangle1_widths[1655]), .rectangle1_height(rectangle1_heights[1655]), .rectangle1_weight(rectangle1_weights[1655]), .rectangle2_x(rectangle2_xs[1655]), .rectangle2_y(rectangle2_ys[1655]), .rectangle2_width(rectangle2_widths[1655]), .rectangle2_height(rectangle2_heights[1655]), .rectangle2_weight(rectangle2_weights[1655]), .rectangle3_x(rectangle3_xs[1655]), .rectangle3_y(rectangle3_ys[1655]), .rectangle3_width(rectangle3_widths[1655]), .rectangle3_height(rectangle3_heights[1655]), .rectangle3_weight(rectangle3_weights[1655]), .feature_threshold(feature_thresholds[1655]), .feature_above(feature_aboves[1655]), .feature_below(feature_belows[1655]), .scan_win_std_dev(scan_win_std_dev[1655]), .feature_accum(feature_accums[1655]));
  accum_calculator ac1656(.scan_win(scan_win1656), .rectangle1_x(rectangle1_xs[1656]), .rectangle1_y(rectangle1_ys[1656]), .rectangle1_width(rectangle1_widths[1656]), .rectangle1_height(rectangle1_heights[1656]), .rectangle1_weight(rectangle1_weights[1656]), .rectangle2_x(rectangle2_xs[1656]), .rectangle2_y(rectangle2_ys[1656]), .rectangle2_width(rectangle2_widths[1656]), .rectangle2_height(rectangle2_heights[1656]), .rectangle2_weight(rectangle2_weights[1656]), .rectangle3_x(rectangle3_xs[1656]), .rectangle3_y(rectangle3_ys[1656]), .rectangle3_width(rectangle3_widths[1656]), .rectangle3_height(rectangle3_heights[1656]), .rectangle3_weight(rectangle3_weights[1656]), .feature_threshold(feature_thresholds[1656]), .feature_above(feature_aboves[1656]), .feature_below(feature_belows[1656]), .scan_win_std_dev(scan_win_std_dev[1656]), .feature_accum(feature_accums[1656]));
  accum_calculator ac1657(.scan_win(scan_win1657), .rectangle1_x(rectangle1_xs[1657]), .rectangle1_y(rectangle1_ys[1657]), .rectangle1_width(rectangle1_widths[1657]), .rectangle1_height(rectangle1_heights[1657]), .rectangle1_weight(rectangle1_weights[1657]), .rectangle2_x(rectangle2_xs[1657]), .rectangle2_y(rectangle2_ys[1657]), .rectangle2_width(rectangle2_widths[1657]), .rectangle2_height(rectangle2_heights[1657]), .rectangle2_weight(rectangle2_weights[1657]), .rectangle3_x(rectangle3_xs[1657]), .rectangle3_y(rectangle3_ys[1657]), .rectangle3_width(rectangle3_widths[1657]), .rectangle3_height(rectangle3_heights[1657]), .rectangle3_weight(rectangle3_weights[1657]), .feature_threshold(feature_thresholds[1657]), .feature_above(feature_aboves[1657]), .feature_below(feature_belows[1657]), .scan_win_std_dev(scan_win_std_dev[1657]), .feature_accum(feature_accums[1657]));
  accum_calculator ac1658(.scan_win(scan_win1658), .rectangle1_x(rectangle1_xs[1658]), .rectangle1_y(rectangle1_ys[1658]), .rectangle1_width(rectangle1_widths[1658]), .rectangle1_height(rectangle1_heights[1658]), .rectangle1_weight(rectangle1_weights[1658]), .rectangle2_x(rectangle2_xs[1658]), .rectangle2_y(rectangle2_ys[1658]), .rectangle2_width(rectangle2_widths[1658]), .rectangle2_height(rectangle2_heights[1658]), .rectangle2_weight(rectangle2_weights[1658]), .rectangle3_x(rectangle3_xs[1658]), .rectangle3_y(rectangle3_ys[1658]), .rectangle3_width(rectangle3_widths[1658]), .rectangle3_height(rectangle3_heights[1658]), .rectangle3_weight(rectangle3_weights[1658]), .feature_threshold(feature_thresholds[1658]), .feature_above(feature_aboves[1658]), .feature_below(feature_belows[1658]), .scan_win_std_dev(scan_win_std_dev[1658]), .feature_accum(feature_accums[1658]));
  accum_calculator ac1659(.scan_win(scan_win1659), .rectangle1_x(rectangle1_xs[1659]), .rectangle1_y(rectangle1_ys[1659]), .rectangle1_width(rectangle1_widths[1659]), .rectangle1_height(rectangle1_heights[1659]), .rectangle1_weight(rectangle1_weights[1659]), .rectangle2_x(rectangle2_xs[1659]), .rectangle2_y(rectangle2_ys[1659]), .rectangle2_width(rectangle2_widths[1659]), .rectangle2_height(rectangle2_heights[1659]), .rectangle2_weight(rectangle2_weights[1659]), .rectangle3_x(rectangle3_xs[1659]), .rectangle3_y(rectangle3_ys[1659]), .rectangle3_width(rectangle3_widths[1659]), .rectangle3_height(rectangle3_heights[1659]), .rectangle3_weight(rectangle3_weights[1659]), .feature_threshold(feature_thresholds[1659]), .feature_above(feature_aboves[1659]), .feature_below(feature_belows[1659]), .scan_win_std_dev(scan_win_std_dev[1659]), .feature_accum(feature_accums[1659]));
  accum_calculator ac1660(.scan_win(scan_win1660), .rectangle1_x(rectangle1_xs[1660]), .rectangle1_y(rectangle1_ys[1660]), .rectangle1_width(rectangle1_widths[1660]), .rectangle1_height(rectangle1_heights[1660]), .rectangle1_weight(rectangle1_weights[1660]), .rectangle2_x(rectangle2_xs[1660]), .rectangle2_y(rectangle2_ys[1660]), .rectangle2_width(rectangle2_widths[1660]), .rectangle2_height(rectangle2_heights[1660]), .rectangle2_weight(rectangle2_weights[1660]), .rectangle3_x(rectangle3_xs[1660]), .rectangle3_y(rectangle3_ys[1660]), .rectangle3_width(rectangle3_widths[1660]), .rectangle3_height(rectangle3_heights[1660]), .rectangle3_weight(rectangle3_weights[1660]), .feature_threshold(feature_thresholds[1660]), .feature_above(feature_aboves[1660]), .feature_below(feature_belows[1660]), .scan_win_std_dev(scan_win_std_dev[1660]), .feature_accum(feature_accums[1660]));
  accum_calculator ac1661(.scan_win(scan_win1661), .rectangle1_x(rectangle1_xs[1661]), .rectangle1_y(rectangle1_ys[1661]), .rectangle1_width(rectangle1_widths[1661]), .rectangle1_height(rectangle1_heights[1661]), .rectangle1_weight(rectangle1_weights[1661]), .rectangle2_x(rectangle2_xs[1661]), .rectangle2_y(rectangle2_ys[1661]), .rectangle2_width(rectangle2_widths[1661]), .rectangle2_height(rectangle2_heights[1661]), .rectangle2_weight(rectangle2_weights[1661]), .rectangle3_x(rectangle3_xs[1661]), .rectangle3_y(rectangle3_ys[1661]), .rectangle3_width(rectangle3_widths[1661]), .rectangle3_height(rectangle3_heights[1661]), .rectangle3_weight(rectangle3_weights[1661]), .feature_threshold(feature_thresholds[1661]), .feature_above(feature_aboves[1661]), .feature_below(feature_belows[1661]), .scan_win_std_dev(scan_win_std_dev[1661]), .feature_accum(feature_accums[1661]));
  accum_calculator ac1662(.scan_win(scan_win1662), .rectangle1_x(rectangle1_xs[1662]), .rectangle1_y(rectangle1_ys[1662]), .rectangle1_width(rectangle1_widths[1662]), .rectangle1_height(rectangle1_heights[1662]), .rectangle1_weight(rectangle1_weights[1662]), .rectangle2_x(rectangle2_xs[1662]), .rectangle2_y(rectangle2_ys[1662]), .rectangle2_width(rectangle2_widths[1662]), .rectangle2_height(rectangle2_heights[1662]), .rectangle2_weight(rectangle2_weights[1662]), .rectangle3_x(rectangle3_xs[1662]), .rectangle3_y(rectangle3_ys[1662]), .rectangle3_width(rectangle3_widths[1662]), .rectangle3_height(rectangle3_heights[1662]), .rectangle3_weight(rectangle3_weights[1662]), .feature_threshold(feature_thresholds[1662]), .feature_above(feature_aboves[1662]), .feature_below(feature_belows[1662]), .scan_win_std_dev(scan_win_std_dev[1662]), .feature_accum(feature_accums[1662]));
  accum_calculator ac1663(.scan_win(scan_win1663), .rectangle1_x(rectangle1_xs[1663]), .rectangle1_y(rectangle1_ys[1663]), .rectangle1_width(rectangle1_widths[1663]), .rectangle1_height(rectangle1_heights[1663]), .rectangle1_weight(rectangle1_weights[1663]), .rectangle2_x(rectangle2_xs[1663]), .rectangle2_y(rectangle2_ys[1663]), .rectangle2_width(rectangle2_widths[1663]), .rectangle2_height(rectangle2_heights[1663]), .rectangle2_weight(rectangle2_weights[1663]), .rectangle3_x(rectangle3_xs[1663]), .rectangle3_y(rectangle3_ys[1663]), .rectangle3_width(rectangle3_widths[1663]), .rectangle3_height(rectangle3_heights[1663]), .rectangle3_weight(rectangle3_weights[1663]), .feature_threshold(feature_thresholds[1663]), .feature_above(feature_aboves[1663]), .feature_below(feature_belows[1663]), .scan_win_std_dev(scan_win_std_dev[1663]), .feature_accum(feature_accums[1663]));
  accum_calculator ac1664(.scan_win(scan_win1664), .rectangle1_x(rectangle1_xs[1664]), .rectangle1_y(rectangle1_ys[1664]), .rectangle1_width(rectangle1_widths[1664]), .rectangle1_height(rectangle1_heights[1664]), .rectangle1_weight(rectangle1_weights[1664]), .rectangle2_x(rectangle2_xs[1664]), .rectangle2_y(rectangle2_ys[1664]), .rectangle2_width(rectangle2_widths[1664]), .rectangle2_height(rectangle2_heights[1664]), .rectangle2_weight(rectangle2_weights[1664]), .rectangle3_x(rectangle3_xs[1664]), .rectangle3_y(rectangle3_ys[1664]), .rectangle3_width(rectangle3_widths[1664]), .rectangle3_height(rectangle3_heights[1664]), .rectangle3_weight(rectangle3_weights[1664]), .feature_threshold(feature_thresholds[1664]), .feature_above(feature_aboves[1664]), .feature_below(feature_belows[1664]), .scan_win_std_dev(scan_win_std_dev[1664]), .feature_accum(feature_accums[1664]));
  accum_calculator ac1665(.scan_win(scan_win1665), .rectangle1_x(rectangle1_xs[1665]), .rectangle1_y(rectangle1_ys[1665]), .rectangle1_width(rectangle1_widths[1665]), .rectangle1_height(rectangle1_heights[1665]), .rectangle1_weight(rectangle1_weights[1665]), .rectangle2_x(rectangle2_xs[1665]), .rectangle2_y(rectangle2_ys[1665]), .rectangle2_width(rectangle2_widths[1665]), .rectangle2_height(rectangle2_heights[1665]), .rectangle2_weight(rectangle2_weights[1665]), .rectangle3_x(rectangle3_xs[1665]), .rectangle3_y(rectangle3_ys[1665]), .rectangle3_width(rectangle3_widths[1665]), .rectangle3_height(rectangle3_heights[1665]), .rectangle3_weight(rectangle3_weights[1665]), .feature_threshold(feature_thresholds[1665]), .feature_above(feature_aboves[1665]), .feature_below(feature_belows[1665]), .scan_win_std_dev(scan_win_std_dev[1665]), .feature_accum(feature_accums[1665]));
  accum_calculator ac1666(.scan_win(scan_win1666), .rectangle1_x(rectangle1_xs[1666]), .rectangle1_y(rectangle1_ys[1666]), .rectangle1_width(rectangle1_widths[1666]), .rectangle1_height(rectangle1_heights[1666]), .rectangle1_weight(rectangle1_weights[1666]), .rectangle2_x(rectangle2_xs[1666]), .rectangle2_y(rectangle2_ys[1666]), .rectangle2_width(rectangle2_widths[1666]), .rectangle2_height(rectangle2_heights[1666]), .rectangle2_weight(rectangle2_weights[1666]), .rectangle3_x(rectangle3_xs[1666]), .rectangle3_y(rectangle3_ys[1666]), .rectangle3_width(rectangle3_widths[1666]), .rectangle3_height(rectangle3_heights[1666]), .rectangle3_weight(rectangle3_weights[1666]), .feature_threshold(feature_thresholds[1666]), .feature_above(feature_aboves[1666]), .feature_below(feature_belows[1666]), .scan_win_std_dev(scan_win_std_dev[1666]), .feature_accum(feature_accums[1666]));
  accum_calculator ac1667(.scan_win(scan_win1667), .rectangle1_x(rectangle1_xs[1667]), .rectangle1_y(rectangle1_ys[1667]), .rectangle1_width(rectangle1_widths[1667]), .rectangle1_height(rectangle1_heights[1667]), .rectangle1_weight(rectangle1_weights[1667]), .rectangle2_x(rectangle2_xs[1667]), .rectangle2_y(rectangle2_ys[1667]), .rectangle2_width(rectangle2_widths[1667]), .rectangle2_height(rectangle2_heights[1667]), .rectangle2_weight(rectangle2_weights[1667]), .rectangle3_x(rectangle3_xs[1667]), .rectangle3_y(rectangle3_ys[1667]), .rectangle3_width(rectangle3_widths[1667]), .rectangle3_height(rectangle3_heights[1667]), .rectangle3_weight(rectangle3_weights[1667]), .feature_threshold(feature_thresholds[1667]), .feature_above(feature_aboves[1667]), .feature_below(feature_belows[1667]), .scan_win_std_dev(scan_win_std_dev[1667]), .feature_accum(feature_accums[1667]));
  accum_calculator ac1668(.scan_win(scan_win1668), .rectangle1_x(rectangle1_xs[1668]), .rectangle1_y(rectangle1_ys[1668]), .rectangle1_width(rectangle1_widths[1668]), .rectangle1_height(rectangle1_heights[1668]), .rectangle1_weight(rectangle1_weights[1668]), .rectangle2_x(rectangle2_xs[1668]), .rectangle2_y(rectangle2_ys[1668]), .rectangle2_width(rectangle2_widths[1668]), .rectangle2_height(rectangle2_heights[1668]), .rectangle2_weight(rectangle2_weights[1668]), .rectangle3_x(rectangle3_xs[1668]), .rectangle3_y(rectangle3_ys[1668]), .rectangle3_width(rectangle3_widths[1668]), .rectangle3_height(rectangle3_heights[1668]), .rectangle3_weight(rectangle3_weights[1668]), .feature_threshold(feature_thresholds[1668]), .feature_above(feature_aboves[1668]), .feature_below(feature_belows[1668]), .scan_win_std_dev(scan_win_std_dev[1668]), .feature_accum(feature_accums[1668]));
  accum_calculator ac1669(.scan_win(scan_win1669), .rectangle1_x(rectangle1_xs[1669]), .rectangle1_y(rectangle1_ys[1669]), .rectangle1_width(rectangle1_widths[1669]), .rectangle1_height(rectangle1_heights[1669]), .rectangle1_weight(rectangle1_weights[1669]), .rectangle2_x(rectangle2_xs[1669]), .rectangle2_y(rectangle2_ys[1669]), .rectangle2_width(rectangle2_widths[1669]), .rectangle2_height(rectangle2_heights[1669]), .rectangle2_weight(rectangle2_weights[1669]), .rectangle3_x(rectangle3_xs[1669]), .rectangle3_y(rectangle3_ys[1669]), .rectangle3_width(rectangle3_widths[1669]), .rectangle3_height(rectangle3_heights[1669]), .rectangle3_weight(rectangle3_weights[1669]), .feature_threshold(feature_thresholds[1669]), .feature_above(feature_aboves[1669]), .feature_below(feature_belows[1669]), .scan_win_std_dev(scan_win_std_dev[1669]), .feature_accum(feature_accums[1669]));
  accum_calculator ac1670(.scan_win(scan_win1670), .rectangle1_x(rectangle1_xs[1670]), .rectangle1_y(rectangle1_ys[1670]), .rectangle1_width(rectangle1_widths[1670]), .rectangle1_height(rectangle1_heights[1670]), .rectangle1_weight(rectangle1_weights[1670]), .rectangle2_x(rectangle2_xs[1670]), .rectangle2_y(rectangle2_ys[1670]), .rectangle2_width(rectangle2_widths[1670]), .rectangle2_height(rectangle2_heights[1670]), .rectangle2_weight(rectangle2_weights[1670]), .rectangle3_x(rectangle3_xs[1670]), .rectangle3_y(rectangle3_ys[1670]), .rectangle3_width(rectangle3_widths[1670]), .rectangle3_height(rectangle3_heights[1670]), .rectangle3_weight(rectangle3_weights[1670]), .feature_threshold(feature_thresholds[1670]), .feature_above(feature_aboves[1670]), .feature_below(feature_belows[1670]), .scan_win_std_dev(scan_win_std_dev[1670]), .feature_accum(feature_accums[1670]));
  accum_calculator ac1671(.scan_win(scan_win1671), .rectangle1_x(rectangle1_xs[1671]), .rectangle1_y(rectangle1_ys[1671]), .rectangle1_width(rectangle1_widths[1671]), .rectangle1_height(rectangle1_heights[1671]), .rectangle1_weight(rectangle1_weights[1671]), .rectangle2_x(rectangle2_xs[1671]), .rectangle2_y(rectangle2_ys[1671]), .rectangle2_width(rectangle2_widths[1671]), .rectangle2_height(rectangle2_heights[1671]), .rectangle2_weight(rectangle2_weights[1671]), .rectangle3_x(rectangle3_xs[1671]), .rectangle3_y(rectangle3_ys[1671]), .rectangle3_width(rectangle3_widths[1671]), .rectangle3_height(rectangle3_heights[1671]), .rectangle3_weight(rectangle3_weights[1671]), .feature_threshold(feature_thresholds[1671]), .feature_above(feature_aboves[1671]), .feature_below(feature_belows[1671]), .scan_win_std_dev(scan_win_std_dev[1671]), .feature_accum(feature_accums[1671]));
  accum_calculator ac1672(.scan_win(scan_win1672), .rectangle1_x(rectangle1_xs[1672]), .rectangle1_y(rectangle1_ys[1672]), .rectangle1_width(rectangle1_widths[1672]), .rectangle1_height(rectangle1_heights[1672]), .rectangle1_weight(rectangle1_weights[1672]), .rectangle2_x(rectangle2_xs[1672]), .rectangle2_y(rectangle2_ys[1672]), .rectangle2_width(rectangle2_widths[1672]), .rectangle2_height(rectangle2_heights[1672]), .rectangle2_weight(rectangle2_weights[1672]), .rectangle3_x(rectangle3_xs[1672]), .rectangle3_y(rectangle3_ys[1672]), .rectangle3_width(rectangle3_widths[1672]), .rectangle3_height(rectangle3_heights[1672]), .rectangle3_weight(rectangle3_weights[1672]), .feature_threshold(feature_thresholds[1672]), .feature_above(feature_aboves[1672]), .feature_below(feature_belows[1672]), .scan_win_std_dev(scan_win_std_dev[1672]), .feature_accum(feature_accums[1672]));
  accum_calculator ac1673(.scan_win(scan_win1673), .rectangle1_x(rectangle1_xs[1673]), .rectangle1_y(rectangle1_ys[1673]), .rectangle1_width(rectangle1_widths[1673]), .rectangle1_height(rectangle1_heights[1673]), .rectangle1_weight(rectangle1_weights[1673]), .rectangle2_x(rectangle2_xs[1673]), .rectangle2_y(rectangle2_ys[1673]), .rectangle2_width(rectangle2_widths[1673]), .rectangle2_height(rectangle2_heights[1673]), .rectangle2_weight(rectangle2_weights[1673]), .rectangle3_x(rectangle3_xs[1673]), .rectangle3_y(rectangle3_ys[1673]), .rectangle3_width(rectangle3_widths[1673]), .rectangle3_height(rectangle3_heights[1673]), .rectangle3_weight(rectangle3_weights[1673]), .feature_threshold(feature_thresholds[1673]), .feature_above(feature_aboves[1673]), .feature_below(feature_belows[1673]), .scan_win_std_dev(scan_win_std_dev[1673]), .feature_accum(feature_accums[1673]));
  accum_calculator ac1674(.scan_win(scan_win1674), .rectangle1_x(rectangle1_xs[1674]), .rectangle1_y(rectangle1_ys[1674]), .rectangle1_width(rectangle1_widths[1674]), .rectangle1_height(rectangle1_heights[1674]), .rectangle1_weight(rectangle1_weights[1674]), .rectangle2_x(rectangle2_xs[1674]), .rectangle2_y(rectangle2_ys[1674]), .rectangle2_width(rectangle2_widths[1674]), .rectangle2_height(rectangle2_heights[1674]), .rectangle2_weight(rectangle2_weights[1674]), .rectangle3_x(rectangle3_xs[1674]), .rectangle3_y(rectangle3_ys[1674]), .rectangle3_width(rectangle3_widths[1674]), .rectangle3_height(rectangle3_heights[1674]), .rectangle3_weight(rectangle3_weights[1674]), .feature_threshold(feature_thresholds[1674]), .feature_above(feature_aboves[1674]), .feature_below(feature_belows[1674]), .scan_win_std_dev(scan_win_std_dev[1674]), .feature_accum(feature_accums[1674]));
  accum_calculator ac1675(.scan_win(scan_win1675), .rectangle1_x(rectangle1_xs[1675]), .rectangle1_y(rectangle1_ys[1675]), .rectangle1_width(rectangle1_widths[1675]), .rectangle1_height(rectangle1_heights[1675]), .rectangle1_weight(rectangle1_weights[1675]), .rectangle2_x(rectangle2_xs[1675]), .rectangle2_y(rectangle2_ys[1675]), .rectangle2_width(rectangle2_widths[1675]), .rectangle2_height(rectangle2_heights[1675]), .rectangle2_weight(rectangle2_weights[1675]), .rectangle3_x(rectangle3_xs[1675]), .rectangle3_y(rectangle3_ys[1675]), .rectangle3_width(rectangle3_widths[1675]), .rectangle3_height(rectangle3_heights[1675]), .rectangle3_weight(rectangle3_weights[1675]), .feature_threshold(feature_thresholds[1675]), .feature_above(feature_aboves[1675]), .feature_below(feature_belows[1675]), .scan_win_std_dev(scan_win_std_dev[1675]), .feature_accum(feature_accums[1675]));
  accum_calculator ac1676(.scan_win(scan_win1676), .rectangle1_x(rectangle1_xs[1676]), .rectangle1_y(rectangle1_ys[1676]), .rectangle1_width(rectangle1_widths[1676]), .rectangle1_height(rectangle1_heights[1676]), .rectangle1_weight(rectangle1_weights[1676]), .rectangle2_x(rectangle2_xs[1676]), .rectangle2_y(rectangle2_ys[1676]), .rectangle2_width(rectangle2_widths[1676]), .rectangle2_height(rectangle2_heights[1676]), .rectangle2_weight(rectangle2_weights[1676]), .rectangle3_x(rectangle3_xs[1676]), .rectangle3_y(rectangle3_ys[1676]), .rectangle3_width(rectangle3_widths[1676]), .rectangle3_height(rectangle3_heights[1676]), .rectangle3_weight(rectangle3_weights[1676]), .feature_threshold(feature_thresholds[1676]), .feature_above(feature_aboves[1676]), .feature_below(feature_belows[1676]), .scan_win_std_dev(scan_win_std_dev[1676]), .feature_accum(feature_accums[1676]));
  accum_calculator ac1677(.scan_win(scan_win1677), .rectangle1_x(rectangle1_xs[1677]), .rectangle1_y(rectangle1_ys[1677]), .rectangle1_width(rectangle1_widths[1677]), .rectangle1_height(rectangle1_heights[1677]), .rectangle1_weight(rectangle1_weights[1677]), .rectangle2_x(rectangle2_xs[1677]), .rectangle2_y(rectangle2_ys[1677]), .rectangle2_width(rectangle2_widths[1677]), .rectangle2_height(rectangle2_heights[1677]), .rectangle2_weight(rectangle2_weights[1677]), .rectangle3_x(rectangle3_xs[1677]), .rectangle3_y(rectangle3_ys[1677]), .rectangle3_width(rectangle3_widths[1677]), .rectangle3_height(rectangle3_heights[1677]), .rectangle3_weight(rectangle3_weights[1677]), .feature_threshold(feature_thresholds[1677]), .feature_above(feature_aboves[1677]), .feature_below(feature_belows[1677]), .scan_win_std_dev(scan_win_std_dev[1677]), .feature_accum(feature_accums[1677]));
  accum_calculator ac1678(.scan_win(scan_win1678), .rectangle1_x(rectangle1_xs[1678]), .rectangle1_y(rectangle1_ys[1678]), .rectangle1_width(rectangle1_widths[1678]), .rectangle1_height(rectangle1_heights[1678]), .rectangle1_weight(rectangle1_weights[1678]), .rectangle2_x(rectangle2_xs[1678]), .rectangle2_y(rectangle2_ys[1678]), .rectangle2_width(rectangle2_widths[1678]), .rectangle2_height(rectangle2_heights[1678]), .rectangle2_weight(rectangle2_weights[1678]), .rectangle3_x(rectangle3_xs[1678]), .rectangle3_y(rectangle3_ys[1678]), .rectangle3_width(rectangle3_widths[1678]), .rectangle3_height(rectangle3_heights[1678]), .rectangle3_weight(rectangle3_weights[1678]), .feature_threshold(feature_thresholds[1678]), .feature_above(feature_aboves[1678]), .feature_below(feature_belows[1678]), .scan_win_std_dev(scan_win_std_dev[1678]), .feature_accum(feature_accums[1678]));
  accum_calculator ac1679(.scan_win(scan_win1679), .rectangle1_x(rectangle1_xs[1679]), .rectangle1_y(rectangle1_ys[1679]), .rectangle1_width(rectangle1_widths[1679]), .rectangle1_height(rectangle1_heights[1679]), .rectangle1_weight(rectangle1_weights[1679]), .rectangle2_x(rectangle2_xs[1679]), .rectangle2_y(rectangle2_ys[1679]), .rectangle2_width(rectangle2_widths[1679]), .rectangle2_height(rectangle2_heights[1679]), .rectangle2_weight(rectangle2_weights[1679]), .rectangle3_x(rectangle3_xs[1679]), .rectangle3_y(rectangle3_ys[1679]), .rectangle3_width(rectangle3_widths[1679]), .rectangle3_height(rectangle3_heights[1679]), .rectangle3_weight(rectangle3_weights[1679]), .feature_threshold(feature_thresholds[1679]), .feature_above(feature_aboves[1679]), .feature_below(feature_belows[1679]), .scan_win_std_dev(scan_win_std_dev[1679]), .feature_accum(feature_accums[1679]));
  accum_calculator ac1680(.scan_win(scan_win1680), .rectangle1_x(rectangle1_xs[1680]), .rectangle1_y(rectangle1_ys[1680]), .rectangle1_width(rectangle1_widths[1680]), .rectangle1_height(rectangle1_heights[1680]), .rectangle1_weight(rectangle1_weights[1680]), .rectangle2_x(rectangle2_xs[1680]), .rectangle2_y(rectangle2_ys[1680]), .rectangle2_width(rectangle2_widths[1680]), .rectangle2_height(rectangle2_heights[1680]), .rectangle2_weight(rectangle2_weights[1680]), .rectangle3_x(rectangle3_xs[1680]), .rectangle3_y(rectangle3_ys[1680]), .rectangle3_width(rectangle3_widths[1680]), .rectangle3_height(rectangle3_heights[1680]), .rectangle3_weight(rectangle3_weights[1680]), .feature_threshold(feature_thresholds[1680]), .feature_above(feature_aboves[1680]), .feature_below(feature_belows[1680]), .scan_win_std_dev(scan_win_std_dev[1680]), .feature_accum(feature_accums[1680]));
  accum_calculator ac1681(.scan_win(scan_win1681), .rectangle1_x(rectangle1_xs[1681]), .rectangle1_y(rectangle1_ys[1681]), .rectangle1_width(rectangle1_widths[1681]), .rectangle1_height(rectangle1_heights[1681]), .rectangle1_weight(rectangle1_weights[1681]), .rectangle2_x(rectangle2_xs[1681]), .rectangle2_y(rectangle2_ys[1681]), .rectangle2_width(rectangle2_widths[1681]), .rectangle2_height(rectangle2_heights[1681]), .rectangle2_weight(rectangle2_weights[1681]), .rectangle3_x(rectangle3_xs[1681]), .rectangle3_y(rectangle3_ys[1681]), .rectangle3_width(rectangle3_widths[1681]), .rectangle3_height(rectangle3_heights[1681]), .rectangle3_weight(rectangle3_weights[1681]), .feature_threshold(feature_thresholds[1681]), .feature_above(feature_aboves[1681]), .feature_below(feature_belows[1681]), .scan_win_std_dev(scan_win_std_dev[1681]), .feature_accum(feature_accums[1681]));
  accum_calculator ac1682(.scan_win(scan_win1682), .rectangle1_x(rectangle1_xs[1682]), .rectangle1_y(rectangle1_ys[1682]), .rectangle1_width(rectangle1_widths[1682]), .rectangle1_height(rectangle1_heights[1682]), .rectangle1_weight(rectangle1_weights[1682]), .rectangle2_x(rectangle2_xs[1682]), .rectangle2_y(rectangle2_ys[1682]), .rectangle2_width(rectangle2_widths[1682]), .rectangle2_height(rectangle2_heights[1682]), .rectangle2_weight(rectangle2_weights[1682]), .rectangle3_x(rectangle3_xs[1682]), .rectangle3_y(rectangle3_ys[1682]), .rectangle3_width(rectangle3_widths[1682]), .rectangle3_height(rectangle3_heights[1682]), .rectangle3_weight(rectangle3_weights[1682]), .feature_threshold(feature_thresholds[1682]), .feature_above(feature_aboves[1682]), .feature_below(feature_belows[1682]), .scan_win_std_dev(scan_win_std_dev[1682]), .feature_accum(feature_accums[1682]));
  accum_calculator ac1683(.scan_win(scan_win1683), .rectangle1_x(rectangle1_xs[1683]), .rectangle1_y(rectangle1_ys[1683]), .rectangle1_width(rectangle1_widths[1683]), .rectangle1_height(rectangle1_heights[1683]), .rectangle1_weight(rectangle1_weights[1683]), .rectangle2_x(rectangle2_xs[1683]), .rectangle2_y(rectangle2_ys[1683]), .rectangle2_width(rectangle2_widths[1683]), .rectangle2_height(rectangle2_heights[1683]), .rectangle2_weight(rectangle2_weights[1683]), .rectangle3_x(rectangle3_xs[1683]), .rectangle3_y(rectangle3_ys[1683]), .rectangle3_width(rectangle3_widths[1683]), .rectangle3_height(rectangle3_heights[1683]), .rectangle3_weight(rectangle3_weights[1683]), .feature_threshold(feature_thresholds[1683]), .feature_above(feature_aboves[1683]), .feature_below(feature_belows[1683]), .scan_win_std_dev(scan_win_std_dev[1683]), .feature_accum(feature_accums[1683]));
  accum_calculator ac1684(.scan_win(scan_win1684), .rectangle1_x(rectangle1_xs[1684]), .rectangle1_y(rectangle1_ys[1684]), .rectangle1_width(rectangle1_widths[1684]), .rectangle1_height(rectangle1_heights[1684]), .rectangle1_weight(rectangle1_weights[1684]), .rectangle2_x(rectangle2_xs[1684]), .rectangle2_y(rectangle2_ys[1684]), .rectangle2_width(rectangle2_widths[1684]), .rectangle2_height(rectangle2_heights[1684]), .rectangle2_weight(rectangle2_weights[1684]), .rectangle3_x(rectangle3_xs[1684]), .rectangle3_y(rectangle3_ys[1684]), .rectangle3_width(rectangle3_widths[1684]), .rectangle3_height(rectangle3_heights[1684]), .rectangle3_weight(rectangle3_weights[1684]), .feature_threshold(feature_thresholds[1684]), .feature_above(feature_aboves[1684]), .feature_below(feature_belows[1684]), .scan_win_std_dev(scan_win_std_dev[1684]), .feature_accum(feature_accums[1684]));
  accum_calculator ac1685(.scan_win(scan_win1685), .rectangle1_x(rectangle1_xs[1685]), .rectangle1_y(rectangle1_ys[1685]), .rectangle1_width(rectangle1_widths[1685]), .rectangle1_height(rectangle1_heights[1685]), .rectangle1_weight(rectangle1_weights[1685]), .rectangle2_x(rectangle2_xs[1685]), .rectangle2_y(rectangle2_ys[1685]), .rectangle2_width(rectangle2_widths[1685]), .rectangle2_height(rectangle2_heights[1685]), .rectangle2_weight(rectangle2_weights[1685]), .rectangle3_x(rectangle3_xs[1685]), .rectangle3_y(rectangle3_ys[1685]), .rectangle3_width(rectangle3_widths[1685]), .rectangle3_height(rectangle3_heights[1685]), .rectangle3_weight(rectangle3_weights[1685]), .feature_threshold(feature_thresholds[1685]), .feature_above(feature_aboves[1685]), .feature_below(feature_belows[1685]), .scan_win_std_dev(scan_win_std_dev[1685]), .feature_accum(feature_accums[1685]));
  accum_calculator ac1686(.scan_win(scan_win1686), .rectangle1_x(rectangle1_xs[1686]), .rectangle1_y(rectangle1_ys[1686]), .rectangle1_width(rectangle1_widths[1686]), .rectangle1_height(rectangle1_heights[1686]), .rectangle1_weight(rectangle1_weights[1686]), .rectangle2_x(rectangle2_xs[1686]), .rectangle2_y(rectangle2_ys[1686]), .rectangle2_width(rectangle2_widths[1686]), .rectangle2_height(rectangle2_heights[1686]), .rectangle2_weight(rectangle2_weights[1686]), .rectangle3_x(rectangle3_xs[1686]), .rectangle3_y(rectangle3_ys[1686]), .rectangle3_width(rectangle3_widths[1686]), .rectangle3_height(rectangle3_heights[1686]), .rectangle3_weight(rectangle3_weights[1686]), .feature_threshold(feature_thresholds[1686]), .feature_above(feature_aboves[1686]), .feature_below(feature_belows[1686]), .scan_win_std_dev(scan_win_std_dev[1686]), .feature_accum(feature_accums[1686]));
  accum_calculator ac1687(.scan_win(scan_win1687), .rectangle1_x(rectangle1_xs[1687]), .rectangle1_y(rectangle1_ys[1687]), .rectangle1_width(rectangle1_widths[1687]), .rectangle1_height(rectangle1_heights[1687]), .rectangle1_weight(rectangle1_weights[1687]), .rectangle2_x(rectangle2_xs[1687]), .rectangle2_y(rectangle2_ys[1687]), .rectangle2_width(rectangle2_widths[1687]), .rectangle2_height(rectangle2_heights[1687]), .rectangle2_weight(rectangle2_weights[1687]), .rectangle3_x(rectangle3_xs[1687]), .rectangle3_y(rectangle3_ys[1687]), .rectangle3_width(rectangle3_widths[1687]), .rectangle3_height(rectangle3_heights[1687]), .rectangle3_weight(rectangle3_weights[1687]), .feature_threshold(feature_thresholds[1687]), .feature_above(feature_aboves[1687]), .feature_below(feature_belows[1687]), .scan_win_std_dev(scan_win_std_dev[1687]), .feature_accum(feature_accums[1687]));
  accum_calculator ac1688(.scan_win(scan_win1688), .rectangle1_x(rectangle1_xs[1688]), .rectangle1_y(rectangle1_ys[1688]), .rectangle1_width(rectangle1_widths[1688]), .rectangle1_height(rectangle1_heights[1688]), .rectangle1_weight(rectangle1_weights[1688]), .rectangle2_x(rectangle2_xs[1688]), .rectangle2_y(rectangle2_ys[1688]), .rectangle2_width(rectangle2_widths[1688]), .rectangle2_height(rectangle2_heights[1688]), .rectangle2_weight(rectangle2_weights[1688]), .rectangle3_x(rectangle3_xs[1688]), .rectangle3_y(rectangle3_ys[1688]), .rectangle3_width(rectangle3_widths[1688]), .rectangle3_height(rectangle3_heights[1688]), .rectangle3_weight(rectangle3_weights[1688]), .feature_threshold(feature_thresholds[1688]), .feature_above(feature_aboves[1688]), .feature_below(feature_belows[1688]), .scan_win_std_dev(scan_win_std_dev[1688]), .feature_accum(feature_accums[1688]));
  accum_calculator ac1689(.scan_win(scan_win1689), .rectangle1_x(rectangle1_xs[1689]), .rectangle1_y(rectangle1_ys[1689]), .rectangle1_width(rectangle1_widths[1689]), .rectangle1_height(rectangle1_heights[1689]), .rectangle1_weight(rectangle1_weights[1689]), .rectangle2_x(rectangle2_xs[1689]), .rectangle2_y(rectangle2_ys[1689]), .rectangle2_width(rectangle2_widths[1689]), .rectangle2_height(rectangle2_heights[1689]), .rectangle2_weight(rectangle2_weights[1689]), .rectangle3_x(rectangle3_xs[1689]), .rectangle3_y(rectangle3_ys[1689]), .rectangle3_width(rectangle3_widths[1689]), .rectangle3_height(rectangle3_heights[1689]), .rectangle3_weight(rectangle3_weights[1689]), .feature_threshold(feature_thresholds[1689]), .feature_above(feature_aboves[1689]), .feature_below(feature_belows[1689]), .scan_win_std_dev(scan_win_std_dev[1689]), .feature_accum(feature_accums[1689]));
  accum_calculator ac1690(.scan_win(scan_win1690), .rectangle1_x(rectangle1_xs[1690]), .rectangle1_y(rectangle1_ys[1690]), .rectangle1_width(rectangle1_widths[1690]), .rectangle1_height(rectangle1_heights[1690]), .rectangle1_weight(rectangle1_weights[1690]), .rectangle2_x(rectangle2_xs[1690]), .rectangle2_y(rectangle2_ys[1690]), .rectangle2_width(rectangle2_widths[1690]), .rectangle2_height(rectangle2_heights[1690]), .rectangle2_weight(rectangle2_weights[1690]), .rectangle3_x(rectangle3_xs[1690]), .rectangle3_y(rectangle3_ys[1690]), .rectangle3_width(rectangle3_widths[1690]), .rectangle3_height(rectangle3_heights[1690]), .rectangle3_weight(rectangle3_weights[1690]), .feature_threshold(feature_thresholds[1690]), .feature_above(feature_aboves[1690]), .feature_below(feature_belows[1690]), .scan_win_std_dev(scan_win_std_dev[1690]), .feature_accum(feature_accums[1690]));
  accum_calculator ac1691(.scan_win(scan_win1691), .rectangle1_x(rectangle1_xs[1691]), .rectangle1_y(rectangle1_ys[1691]), .rectangle1_width(rectangle1_widths[1691]), .rectangle1_height(rectangle1_heights[1691]), .rectangle1_weight(rectangle1_weights[1691]), .rectangle2_x(rectangle2_xs[1691]), .rectangle2_y(rectangle2_ys[1691]), .rectangle2_width(rectangle2_widths[1691]), .rectangle2_height(rectangle2_heights[1691]), .rectangle2_weight(rectangle2_weights[1691]), .rectangle3_x(rectangle3_xs[1691]), .rectangle3_y(rectangle3_ys[1691]), .rectangle3_width(rectangle3_widths[1691]), .rectangle3_height(rectangle3_heights[1691]), .rectangle3_weight(rectangle3_weights[1691]), .feature_threshold(feature_thresholds[1691]), .feature_above(feature_aboves[1691]), .feature_below(feature_belows[1691]), .scan_win_std_dev(scan_win_std_dev[1691]), .feature_accum(feature_accums[1691]));
  accum_calculator ac1692(.scan_win(scan_win1692), .rectangle1_x(rectangle1_xs[1692]), .rectangle1_y(rectangle1_ys[1692]), .rectangle1_width(rectangle1_widths[1692]), .rectangle1_height(rectangle1_heights[1692]), .rectangle1_weight(rectangle1_weights[1692]), .rectangle2_x(rectangle2_xs[1692]), .rectangle2_y(rectangle2_ys[1692]), .rectangle2_width(rectangle2_widths[1692]), .rectangle2_height(rectangle2_heights[1692]), .rectangle2_weight(rectangle2_weights[1692]), .rectangle3_x(rectangle3_xs[1692]), .rectangle3_y(rectangle3_ys[1692]), .rectangle3_width(rectangle3_widths[1692]), .rectangle3_height(rectangle3_heights[1692]), .rectangle3_weight(rectangle3_weights[1692]), .feature_threshold(feature_thresholds[1692]), .feature_above(feature_aboves[1692]), .feature_below(feature_belows[1692]), .scan_win_std_dev(scan_win_std_dev[1692]), .feature_accum(feature_accums[1692]));
  accum_calculator ac1693(.scan_win(scan_win1693), .rectangle1_x(rectangle1_xs[1693]), .rectangle1_y(rectangle1_ys[1693]), .rectangle1_width(rectangle1_widths[1693]), .rectangle1_height(rectangle1_heights[1693]), .rectangle1_weight(rectangle1_weights[1693]), .rectangle2_x(rectangle2_xs[1693]), .rectangle2_y(rectangle2_ys[1693]), .rectangle2_width(rectangle2_widths[1693]), .rectangle2_height(rectangle2_heights[1693]), .rectangle2_weight(rectangle2_weights[1693]), .rectangle3_x(rectangle3_xs[1693]), .rectangle3_y(rectangle3_ys[1693]), .rectangle3_width(rectangle3_widths[1693]), .rectangle3_height(rectangle3_heights[1693]), .rectangle3_weight(rectangle3_weights[1693]), .feature_threshold(feature_thresholds[1693]), .feature_above(feature_aboves[1693]), .feature_below(feature_belows[1693]), .scan_win_std_dev(scan_win_std_dev[1693]), .feature_accum(feature_accums[1693]));
  accum_calculator ac1694(.scan_win(scan_win1694), .rectangle1_x(rectangle1_xs[1694]), .rectangle1_y(rectangle1_ys[1694]), .rectangle1_width(rectangle1_widths[1694]), .rectangle1_height(rectangle1_heights[1694]), .rectangle1_weight(rectangle1_weights[1694]), .rectangle2_x(rectangle2_xs[1694]), .rectangle2_y(rectangle2_ys[1694]), .rectangle2_width(rectangle2_widths[1694]), .rectangle2_height(rectangle2_heights[1694]), .rectangle2_weight(rectangle2_weights[1694]), .rectangle3_x(rectangle3_xs[1694]), .rectangle3_y(rectangle3_ys[1694]), .rectangle3_width(rectangle3_widths[1694]), .rectangle3_height(rectangle3_heights[1694]), .rectangle3_weight(rectangle3_weights[1694]), .feature_threshold(feature_thresholds[1694]), .feature_above(feature_aboves[1694]), .feature_below(feature_belows[1694]), .scan_win_std_dev(scan_win_std_dev[1694]), .feature_accum(feature_accums[1694]));
  accum_calculator ac1695(.scan_win(scan_win1695), .rectangle1_x(rectangle1_xs[1695]), .rectangle1_y(rectangle1_ys[1695]), .rectangle1_width(rectangle1_widths[1695]), .rectangle1_height(rectangle1_heights[1695]), .rectangle1_weight(rectangle1_weights[1695]), .rectangle2_x(rectangle2_xs[1695]), .rectangle2_y(rectangle2_ys[1695]), .rectangle2_width(rectangle2_widths[1695]), .rectangle2_height(rectangle2_heights[1695]), .rectangle2_weight(rectangle2_weights[1695]), .rectangle3_x(rectangle3_xs[1695]), .rectangle3_y(rectangle3_ys[1695]), .rectangle3_width(rectangle3_widths[1695]), .rectangle3_height(rectangle3_heights[1695]), .rectangle3_weight(rectangle3_weights[1695]), .feature_threshold(feature_thresholds[1695]), .feature_above(feature_aboves[1695]), .feature_below(feature_belows[1695]), .scan_win_std_dev(scan_win_std_dev[1695]), .feature_accum(feature_accums[1695]));
  accum_calculator ac1696(.scan_win(scan_win1696), .rectangle1_x(rectangle1_xs[1696]), .rectangle1_y(rectangle1_ys[1696]), .rectangle1_width(rectangle1_widths[1696]), .rectangle1_height(rectangle1_heights[1696]), .rectangle1_weight(rectangle1_weights[1696]), .rectangle2_x(rectangle2_xs[1696]), .rectangle2_y(rectangle2_ys[1696]), .rectangle2_width(rectangle2_widths[1696]), .rectangle2_height(rectangle2_heights[1696]), .rectangle2_weight(rectangle2_weights[1696]), .rectangle3_x(rectangle3_xs[1696]), .rectangle3_y(rectangle3_ys[1696]), .rectangle3_width(rectangle3_widths[1696]), .rectangle3_height(rectangle3_heights[1696]), .rectangle3_weight(rectangle3_weights[1696]), .feature_threshold(feature_thresholds[1696]), .feature_above(feature_aboves[1696]), .feature_below(feature_belows[1696]), .scan_win_std_dev(scan_win_std_dev[1696]), .feature_accum(feature_accums[1696]));
  accum_calculator ac1697(.scan_win(scan_win1697), .rectangle1_x(rectangle1_xs[1697]), .rectangle1_y(rectangle1_ys[1697]), .rectangle1_width(rectangle1_widths[1697]), .rectangle1_height(rectangle1_heights[1697]), .rectangle1_weight(rectangle1_weights[1697]), .rectangle2_x(rectangle2_xs[1697]), .rectangle2_y(rectangle2_ys[1697]), .rectangle2_width(rectangle2_widths[1697]), .rectangle2_height(rectangle2_heights[1697]), .rectangle2_weight(rectangle2_weights[1697]), .rectangle3_x(rectangle3_xs[1697]), .rectangle3_y(rectangle3_ys[1697]), .rectangle3_width(rectangle3_widths[1697]), .rectangle3_height(rectangle3_heights[1697]), .rectangle3_weight(rectangle3_weights[1697]), .feature_threshold(feature_thresholds[1697]), .feature_above(feature_aboves[1697]), .feature_below(feature_belows[1697]), .scan_win_std_dev(scan_win_std_dev[1697]), .feature_accum(feature_accums[1697]));
  accum_calculator ac1698(.scan_win(scan_win1698), .rectangle1_x(rectangle1_xs[1698]), .rectangle1_y(rectangle1_ys[1698]), .rectangle1_width(rectangle1_widths[1698]), .rectangle1_height(rectangle1_heights[1698]), .rectangle1_weight(rectangle1_weights[1698]), .rectangle2_x(rectangle2_xs[1698]), .rectangle2_y(rectangle2_ys[1698]), .rectangle2_width(rectangle2_widths[1698]), .rectangle2_height(rectangle2_heights[1698]), .rectangle2_weight(rectangle2_weights[1698]), .rectangle3_x(rectangle3_xs[1698]), .rectangle3_y(rectangle3_ys[1698]), .rectangle3_width(rectangle3_widths[1698]), .rectangle3_height(rectangle3_heights[1698]), .rectangle3_weight(rectangle3_weights[1698]), .feature_threshold(feature_thresholds[1698]), .feature_above(feature_aboves[1698]), .feature_below(feature_belows[1698]), .scan_win_std_dev(scan_win_std_dev[1698]), .feature_accum(feature_accums[1698]));
  accum_calculator ac1699(.scan_win(scan_win1699), .rectangle1_x(rectangle1_xs[1699]), .rectangle1_y(rectangle1_ys[1699]), .rectangle1_width(rectangle1_widths[1699]), .rectangle1_height(rectangle1_heights[1699]), .rectangle1_weight(rectangle1_weights[1699]), .rectangle2_x(rectangle2_xs[1699]), .rectangle2_y(rectangle2_ys[1699]), .rectangle2_width(rectangle2_widths[1699]), .rectangle2_height(rectangle2_heights[1699]), .rectangle2_weight(rectangle2_weights[1699]), .rectangle3_x(rectangle3_xs[1699]), .rectangle3_y(rectangle3_ys[1699]), .rectangle3_width(rectangle3_widths[1699]), .rectangle3_height(rectangle3_heights[1699]), .rectangle3_weight(rectangle3_weights[1699]), .feature_threshold(feature_thresholds[1699]), .feature_above(feature_aboves[1699]), .feature_below(feature_belows[1699]), .scan_win_std_dev(scan_win_std_dev[1699]), .feature_accum(feature_accums[1699]));
  accum_calculator ac1700(.scan_win(scan_win1700), .rectangle1_x(rectangle1_xs[1700]), .rectangle1_y(rectangle1_ys[1700]), .rectangle1_width(rectangle1_widths[1700]), .rectangle1_height(rectangle1_heights[1700]), .rectangle1_weight(rectangle1_weights[1700]), .rectangle2_x(rectangle2_xs[1700]), .rectangle2_y(rectangle2_ys[1700]), .rectangle2_width(rectangle2_widths[1700]), .rectangle2_height(rectangle2_heights[1700]), .rectangle2_weight(rectangle2_weights[1700]), .rectangle3_x(rectangle3_xs[1700]), .rectangle3_y(rectangle3_ys[1700]), .rectangle3_width(rectangle3_widths[1700]), .rectangle3_height(rectangle3_heights[1700]), .rectangle3_weight(rectangle3_weights[1700]), .feature_threshold(feature_thresholds[1700]), .feature_above(feature_aboves[1700]), .feature_below(feature_belows[1700]), .scan_win_std_dev(scan_win_std_dev[1700]), .feature_accum(feature_accums[1700]));
  accum_calculator ac1701(.scan_win(scan_win1701), .rectangle1_x(rectangle1_xs[1701]), .rectangle1_y(rectangle1_ys[1701]), .rectangle1_width(rectangle1_widths[1701]), .rectangle1_height(rectangle1_heights[1701]), .rectangle1_weight(rectangle1_weights[1701]), .rectangle2_x(rectangle2_xs[1701]), .rectangle2_y(rectangle2_ys[1701]), .rectangle2_width(rectangle2_widths[1701]), .rectangle2_height(rectangle2_heights[1701]), .rectangle2_weight(rectangle2_weights[1701]), .rectangle3_x(rectangle3_xs[1701]), .rectangle3_y(rectangle3_ys[1701]), .rectangle3_width(rectangle3_widths[1701]), .rectangle3_height(rectangle3_heights[1701]), .rectangle3_weight(rectangle3_weights[1701]), .feature_threshold(feature_thresholds[1701]), .feature_above(feature_aboves[1701]), .feature_below(feature_belows[1701]), .scan_win_std_dev(scan_win_std_dev[1701]), .feature_accum(feature_accums[1701]));
  accum_calculator ac1702(.scan_win(scan_win1702), .rectangle1_x(rectangle1_xs[1702]), .rectangle1_y(rectangle1_ys[1702]), .rectangle1_width(rectangle1_widths[1702]), .rectangle1_height(rectangle1_heights[1702]), .rectangle1_weight(rectangle1_weights[1702]), .rectangle2_x(rectangle2_xs[1702]), .rectangle2_y(rectangle2_ys[1702]), .rectangle2_width(rectangle2_widths[1702]), .rectangle2_height(rectangle2_heights[1702]), .rectangle2_weight(rectangle2_weights[1702]), .rectangle3_x(rectangle3_xs[1702]), .rectangle3_y(rectangle3_ys[1702]), .rectangle3_width(rectangle3_widths[1702]), .rectangle3_height(rectangle3_heights[1702]), .rectangle3_weight(rectangle3_weights[1702]), .feature_threshold(feature_thresholds[1702]), .feature_above(feature_aboves[1702]), .feature_below(feature_belows[1702]), .scan_win_std_dev(scan_win_std_dev[1702]), .feature_accum(feature_accums[1702]));
  accum_calculator ac1703(.scan_win(scan_win1703), .rectangle1_x(rectangle1_xs[1703]), .rectangle1_y(rectangle1_ys[1703]), .rectangle1_width(rectangle1_widths[1703]), .rectangle1_height(rectangle1_heights[1703]), .rectangle1_weight(rectangle1_weights[1703]), .rectangle2_x(rectangle2_xs[1703]), .rectangle2_y(rectangle2_ys[1703]), .rectangle2_width(rectangle2_widths[1703]), .rectangle2_height(rectangle2_heights[1703]), .rectangle2_weight(rectangle2_weights[1703]), .rectangle3_x(rectangle3_xs[1703]), .rectangle3_y(rectangle3_ys[1703]), .rectangle3_width(rectangle3_widths[1703]), .rectangle3_height(rectangle3_heights[1703]), .rectangle3_weight(rectangle3_weights[1703]), .feature_threshold(feature_thresholds[1703]), .feature_above(feature_aboves[1703]), .feature_below(feature_belows[1703]), .scan_win_std_dev(scan_win_std_dev[1703]), .feature_accum(feature_accums[1703]));
  accum_calculator ac1704(.scan_win(scan_win1704), .rectangle1_x(rectangle1_xs[1704]), .rectangle1_y(rectangle1_ys[1704]), .rectangle1_width(rectangle1_widths[1704]), .rectangle1_height(rectangle1_heights[1704]), .rectangle1_weight(rectangle1_weights[1704]), .rectangle2_x(rectangle2_xs[1704]), .rectangle2_y(rectangle2_ys[1704]), .rectangle2_width(rectangle2_widths[1704]), .rectangle2_height(rectangle2_heights[1704]), .rectangle2_weight(rectangle2_weights[1704]), .rectangle3_x(rectangle3_xs[1704]), .rectangle3_y(rectangle3_ys[1704]), .rectangle3_width(rectangle3_widths[1704]), .rectangle3_height(rectangle3_heights[1704]), .rectangle3_weight(rectangle3_weights[1704]), .feature_threshold(feature_thresholds[1704]), .feature_above(feature_aboves[1704]), .feature_below(feature_belows[1704]), .scan_win_std_dev(scan_win_std_dev[1704]), .feature_accum(feature_accums[1704]));
  accum_calculator ac1705(.scan_win(scan_win1705), .rectangle1_x(rectangle1_xs[1705]), .rectangle1_y(rectangle1_ys[1705]), .rectangle1_width(rectangle1_widths[1705]), .rectangle1_height(rectangle1_heights[1705]), .rectangle1_weight(rectangle1_weights[1705]), .rectangle2_x(rectangle2_xs[1705]), .rectangle2_y(rectangle2_ys[1705]), .rectangle2_width(rectangle2_widths[1705]), .rectangle2_height(rectangle2_heights[1705]), .rectangle2_weight(rectangle2_weights[1705]), .rectangle3_x(rectangle3_xs[1705]), .rectangle3_y(rectangle3_ys[1705]), .rectangle3_width(rectangle3_widths[1705]), .rectangle3_height(rectangle3_heights[1705]), .rectangle3_weight(rectangle3_weights[1705]), .feature_threshold(feature_thresholds[1705]), .feature_above(feature_aboves[1705]), .feature_below(feature_belows[1705]), .scan_win_std_dev(scan_win_std_dev[1705]), .feature_accum(feature_accums[1705]));
  accum_calculator ac1706(.scan_win(scan_win1706), .rectangle1_x(rectangle1_xs[1706]), .rectangle1_y(rectangle1_ys[1706]), .rectangle1_width(rectangle1_widths[1706]), .rectangle1_height(rectangle1_heights[1706]), .rectangle1_weight(rectangle1_weights[1706]), .rectangle2_x(rectangle2_xs[1706]), .rectangle2_y(rectangle2_ys[1706]), .rectangle2_width(rectangle2_widths[1706]), .rectangle2_height(rectangle2_heights[1706]), .rectangle2_weight(rectangle2_weights[1706]), .rectangle3_x(rectangle3_xs[1706]), .rectangle3_y(rectangle3_ys[1706]), .rectangle3_width(rectangle3_widths[1706]), .rectangle3_height(rectangle3_heights[1706]), .rectangle3_weight(rectangle3_weights[1706]), .feature_threshold(feature_thresholds[1706]), .feature_above(feature_aboves[1706]), .feature_below(feature_belows[1706]), .scan_win_std_dev(scan_win_std_dev[1706]), .feature_accum(feature_accums[1706]));
  accum_calculator ac1707(.scan_win(scan_win1707), .rectangle1_x(rectangle1_xs[1707]), .rectangle1_y(rectangle1_ys[1707]), .rectangle1_width(rectangle1_widths[1707]), .rectangle1_height(rectangle1_heights[1707]), .rectangle1_weight(rectangle1_weights[1707]), .rectangle2_x(rectangle2_xs[1707]), .rectangle2_y(rectangle2_ys[1707]), .rectangle2_width(rectangle2_widths[1707]), .rectangle2_height(rectangle2_heights[1707]), .rectangle2_weight(rectangle2_weights[1707]), .rectangle3_x(rectangle3_xs[1707]), .rectangle3_y(rectangle3_ys[1707]), .rectangle3_width(rectangle3_widths[1707]), .rectangle3_height(rectangle3_heights[1707]), .rectangle3_weight(rectangle3_weights[1707]), .feature_threshold(feature_thresholds[1707]), .feature_above(feature_aboves[1707]), .feature_below(feature_belows[1707]), .scan_win_std_dev(scan_win_std_dev[1707]), .feature_accum(feature_accums[1707]));
  accum_calculator ac1708(.scan_win(scan_win1708), .rectangle1_x(rectangle1_xs[1708]), .rectangle1_y(rectangle1_ys[1708]), .rectangle1_width(rectangle1_widths[1708]), .rectangle1_height(rectangle1_heights[1708]), .rectangle1_weight(rectangle1_weights[1708]), .rectangle2_x(rectangle2_xs[1708]), .rectangle2_y(rectangle2_ys[1708]), .rectangle2_width(rectangle2_widths[1708]), .rectangle2_height(rectangle2_heights[1708]), .rectangle2_weight(rectangle2_weights[1708]), .rectangle3_x(rectangle3_xs[1708]), .rectangle3_y(rectangle3_ys[1708]), .rectangle3_width(rectangle3_widths[1708]), .rectangle3_height(rectangle3_heights[1708]), .rectangle3_weight(rectangle3_weights[1708]), .feature_threshold(feature_thresholds[1708]), .feature_above(feature_aboves[1708]), .feature_below(feature_belows[1708]), .scan_win_std_dev(scan_win_std_dev[1708]), .feature_accum(feature_accums[1708]));
  accum_calculator ac1709(.scan_win(scan_win1709), .rectangle1_x(rectangle1_xs[1709]), .rectangle1_y(rectangle1_ys[1709]), .rectangle1_width(rectangle1_widths[1709]), .rectangle1_height(rectangle1_heights[1709]), .rectangle1_weight(rectangle1_weights[1709]), .rectangle2_x(rectangle2_xs[1709]), .rectangle2_y(rectangle2_ys[1709]), .rectangle2_width(rectangle2_widths[1709]), .rectangle2_height(rectangle2_heights[1709]), .rectangle2_weight(rectangle2_weights[1709]), .rectangle3_x(rectangle3_xs[1709]), .rectangle3_y(rectangle3_ys[1709]), .rectangle3_width(rectangle3_widths[1709]), .rectangle3_height(rectangle3_heights[1709]), .rectangle3_weight(rectangle3_weights[1709]), .feature_threshold(feature_thresholds[1709]), .feature_above(feature_aboves[1709]), .feature_below(feature_belows[1709]), .scan_win_std_dev(scan_win_std_dev[1709]), .feature_accum(feature_accums[1709]));
  accum_calculator ac1710(.scan_win(scan_win1710), .rectangle1_x(rectangle1_xs[1710]), .rectangle1_y(rectangle1_ys[1710]), .rectangle1_width(rectangle1_widths[1710]), .rectangle1_height(rectangle1_heights[1710]), .rectangle1_weight(rectangle1_weights[1710]), .rectangle2_x(rectangle2_xs[1710]), .rectangle2_y(rectangle2_ys[1710]), .rectangle2_width(rectangle2_widths[1710]), .rectangle2_height(rectangle2_heights[1710]), .rectangle2_weight(rectangle2_weights[1710]), .rectangle3_x(rectangle3_xs[1710]), .rectangle3_y(rectangle3_ys[1710]), .rectangle3_width(rectangle3_widths[1710]), .rectangle3_height(rectangle3_heights[1710]), .rectangle3_weight(rectangle3_weights[1710]), .feature_threshold(feature_thresholds[1710]), .feature_above(feature_aboves[1710]), .feature_below(feature_belows[1710]), .scan_win_std_dev(scan_win_std_dev[1710]), .feature_accum(feature_accums[1710]));
  accum_calculator ac1711(.scan_win(scan_win1711), .rectangle1_x(rectangle1_xs[1711]), .rectangle1_y(rectangle1_ys[1711]), .rectangle1_width(rectangle1_widths[1711]), .rectangle1_height(rectangle1_heights[1711]), .rectangle1_weight(rectangle1_weights[1711]), .rectangle2_x(rectangle2_xs[1711]), .rectangle2_y(rectangle2_ys[1711]), .rectangle2_width(rectangle2_widths[1711]), .rectangle2_height(rectangle2_heights[1711]), .rectangle2_weight(rectangle2_weights[1711]), .rectangle3_x(rectangle3_xs[1711]), .rectangle3_y(rectangle3_ys[1711]), .rectangle3_width(rectangle3_widths[1711]), .rectangle3_height(rectangle3_heights[1711]), .rectangle3_weight(rectangle3_weights[1711]), .feature_threshold(feature_thresholds[1711]), .feature_above(feature_aboves[1711]), .feature_below(feature_belows[1711]), .scan_win_std_dev(scan_win_std_dev[1711]), .feature_accum(feature_accums[1711]));
  accum_calculator ac1712(.scan_win(scan_win1712), .rectangle1_x(rectangle1_xs[1712]), .rectangle1_y(rectangle1_ys[1712]), .rectangle1_width(rectangle1_widths[1712]), .rectangle1_height(rectangle1_heights[1712]), .rectangle1_weight(rectangle1_weights[1712]), .rectangle2_x(rectangle2_xs[1712]), .rectangle2_y(rectangle2_ys[1712]), .rectangle2_width(rectangle2_widths[1712]), .rectangle2_height(rectangle2_heights[1712]), .rectangle2_weight(rectangle2_weights[1712]), .rectangle3_x(rectangle3_xs[1712]), .rectangle3_y(rectangle3_ys[1712]), .rectangle3_width(rectangle3_widths[1712]), .rectangle3_height(rectangle3_heights[1712]), .rectangle3_weight(rectangle3_weights[1712]), .feature_threshold(feature_thresholds[1712]), .feature_above(feature_aboves[1712]), .feature_below(feature_belows[1712]), .scan_win_std_dev(scan_win_std_dev[1712]), .feature_accum(feature_accums[1712]));
  accum_calculator ac1713(.scan_win(scan_win1713), .rectangle1_x(rectangle1_xs[1713]), .rectangle1_y(rectangle1_ys[1713]), .rectangle1_width(rectangle1_widths[1713]), .rectangle1_height(rectangle1_heights[1713]), .rectangle1_weight(rectangle1_weights[1713]), .rectangle2_x(rectangle2_xs[1713]), .rectangle2_y(rectangle2_ys[1713]), .rectangle2_width(rectangle2_widths[1713]), .rectangle2_height(rectangle2_heights[1713]), .rectangle2_weight(rectangle2_weights[1713]), .rectangle3_x(rectangle3_xs[1713]), .rectangle3_y(rectangle3_ys[1713]), .rectangle3_width(rectangle3_widths[1713]), .rectangle3_height(rectangle3_heights[1713]), .rectangle3_weight(rectangle3_weights[1713]), .feature_threshold(feature_thresholds[1713]), .feature_above(feature_aboves[1713]), .feature_below(feature_belows[1713]), .scan_win_std_dev(scan_win_std_dev[1713]), .feature_accum(feature_accums[1713]));
  accum_calculator ac1714(.scan_win(scan_win1714), .rectangle1_x(rectangle1_xs[1714]), .rectangle1_y(rectangle1_ys[1714]), .rectangle1_width(rectangle1_widths[1714]), .rectangle1_height(rectangle1_heights[1714]), .rectangle1_weight(rectangle1_weights[1714]), .rectangle2_x(rectangle2_xs[1714]), .rectangle2_y(rectangle2_ys[1714]), .rectangle2_width(rectangle2_widths[1714]), .rectangle2_height(rectangle2_heights[1714]), .rectangle2_weight(rectangle2_weights[1714]), .rectangle3_x(rectangle3_xs[1714]), .rectangle3_y(rectangle3_ys[1714]), .rectangle3_width(rectangle3_widths[1714]), .rectangle3_height(rectangle3_heights[1714]), .rectangle3_weight(rectangle3_weights[1714]), .feature_threshold(feature_thresholds[1714]), .feature_above(feature_aboves[1714]), .feature_below(feature_belows[1714]), .scan_win_std_dev(scan_win_std_dev[1714]), .feature_accum(feature_accums[1714]));
  accum_calculator ac1715(.scan_win(scan_win1715), .rectangle1_x(rectangle1_xs[1715]), .rectangle1_y(rectangle1_ys[1715]), .rectangle1_width(rectangle1_widths[1715]), .rectangle1_height(rectangle1_heights[1715]), .rectangle1_weight(rectangle1_weights[1715]), .rectangle2_x(rectangle2_xs[1715]), .rectangle2_y(rectangle2_ys[1715]), .rectangle2_width(rectangle2_widths[1715]), .rectangle2_height(rectangle2_heights[1715]), .rectangle2_weight(rectangle2_weights[1715]), .rectangle3_x(rectangle3_xs[1715]), .rectangle3_y(rectangle3_ys[1715]), .rectangle3_width(rectangle3_widths[1715]), .rectangle3_height(rectangle3_heights[1715]), .rectangle3_weight(rectangle3_weights[1715]), .feature_threshold(feature_thresholds[1715]), .feature_above(feature_aboves[1715]), .feature_below(feature_belows[1715]), .scan_win_std_dev(scan_win_std_dev[1715]), .feature_accum(feature_accums[1715]));
  accum_calculator ac1716(.scan_win(scan_win1716), .rectangle1_x(rectangle1_xs[1716]), .rectangle1_y(rectangle1_ys[1716]), .rectangle1_width(rectangle1_widths[1716]), .rectangle1_height(rectangle1_heights[1716]), .rectangle1_weight(rectangle1_weights[1716]), .rectangle2_x(rectangle2_xs[1716]), .rectangle2_y(rectangle2_ys[1716]), .rectangle2_width(rectangle2_widths[1716]), .rectangle2_height(rectangle2_heights[1716]), .rectangle2_weight(rectangle2_weights[1716]), .rectangle3_x(rectangle3_xs[1716]), .rectangle3_y(rectangle3_ys[1716]), .rectangle3_width(rectangle3_widths[1716]), .rectangle3_height(rectangle3_heights[1716]), .rectangle3_weight(rectangle3_weights[1716]), .feature_threshold(feature_thresholds[1716]), .feature_above(feature_aboves[1716]), .feature_below(feature_belows[1716]), .scan_win_std_dev(scan_win_std_dev[1716]), .feature_accum(feature_accums[1716]));
  accum_calculator ac1717(.scan_win(scan_win1717), .rectangle1_x(rectangle1_xs[1717]), .rectangle1_y(rectangle1_ys[1717]), .rectangle1_width(rectangle1_widths[1717]), .rectangle1_height(rectangle1_heights[1717]), .rectangle1_weight(rectangle1_weights[1717]), .rectangle2_x(rectangle2_xs[1717]), .rectangle2_y(rectangle2_ys[1717]), .rectangle2_width(rectangle2_widths[1717]), .rectangle2_height(rectangle2_heights[1717]), .rectangle2_weight(rectangle2_weights[1717]), .rectangle3_x(rectangle3_xs[1717]), .rectangle3_y(rectangle3_ys[1717]), .rectangle3_width(rectangle3_widths[1717]), .rectangle3_height(rectangle3_heights[1717]), .rectangle3_weight(rectangle3_weights[1717]), .feature_threshold(feature_thresholds[1717]), .feature_above(feature_aboves[1717]), .feature_below(feature_belows[1717]), .scan_win_std_dev(scan_win_std_dev[1717]), .feature_accum(feature_accums[1717]));
  accum_calculator ac1718(.scan_win(scan_win1718), .rectangle1_x(rectangle1_xs[1718]), .rectangle1_y(rectangle1_ys[1718]), .rectangle1_width(rectangle1_widths[1718]), .rectangle1_height(rectangle1_heights[1718]), .rectangle1_weight(rectangle1_weights[1718]), .rectangle2_x(rectangle2_xs[1718]), .rectangle2_y(rectangle2_ys[1718]), .rectangle2_width(rectangle2_widths[1718]), .rectangle2_height(rectangle2_heights[1718]), .rectangle2_weight(rectangle2_weights[1718]), .rectangle3_x(rectangle3_xs[1718]), .rectangle3_y(rectangle3_ys[1718]), .rectangle3_width(rectangle3_widths[1718]), .rectangle3_height(rectangle3_heights[1718]), .rectangle3_weight(rectangle3_weights[1718]), .feature_threshold(feature_thresholds[1718]), .feature_above(feature_aboves[1718]), .feature_below(feature_belows[1718]), .scan_win_std_dev(scan_win_std_dev[1718]), .feature_accum(feature_accums[1718]));
  accum_calculator ac1719(.scan_win(scan_win1719), .rectangle1_x(rectangle1_xs[1719]), .rectangle1_y(rectangle1_ys[1719]), .rectangle1_width(rectangle1_widths[1719]), .rectangle1_height(rectangle1_heights[1719]), .rectangle1_weight(rectangle1_weights[1719]), .rectangle2_x(rectangle2_xs[1719]), .rectangle2_y(rectangle2_ys[1719]), .rectangle2_width(rectangle2_widths[1719]), .rectangle2_height(rectangle2_heights[1719]), .rectangle2_weight(rectangle2_weights[1719]), .rectangle3_x(rectangle3_xs[1719]), .rectangle3_y(rectangle3_ys[1719]), .rectangle3_width(rectangle3_widths[1719]), .rectangle3_height(rectangle3_heights[1719]), .rectangle3_weight(rectangle3_weights[1719]), .feature_threshold(feature_thresholds[1719]), .feature_above(feature_aboves[1719]), .feature_below(feature_belows[1719]), .scan_win_std_dev(scan_win_std_dev[1719]), .feature_accum(feature_accums[1719]));
  accum_calculator ac1720(.scan_win(scan_win1720), .rectangle1_x(rectangle1_xs[1720]), .rectangle1_y(rectangle1_ys[1720]), .rectangle1_width(rectangle1_widths[1720]), .rectangle1_height(rectangle1_heights[1720]), .rectangle1_weight(rectangle1_weights[1720]), .rectangle2_x(rectangle2_xs[1720]), .rectangle2_y(rectangle2_ys[1720]), .rectangle2_width(rectangle2_widths[1720]), .rectangle2_height(rectangle2_heights[1720]), .rectangle2_weight(rectangle2_weights[1720]), .rectangle3_x(rectangle3_xs[1720]), .rectangle3_y(rectangle3_ys[1720]), .rectangle3_width(rectangle3_widths[1720]), .rectangle3_height(rectangle3_heights[1720]), .rectangle3_weight(rectangle3_weights[1720]), .feature_threshold(feature_thresholds[1720]), .feature_above(feature_aboves[1720]), .feature_below(feature_belows[1720]), .scan_win_std_dev(scan_win_std_dev[1720]), .feature_accum(feature_accums[1720]));
  accum_calculator ac1721(.scan_win(scan_win1721), .rectangle1_x(rectangle1_xs[1721]), .rectangle1_y(rectangle1_ys[1721]), .rectangle1_width(rectangle1_widths[1721]), .rectangle1_height(rectangle1_heights[1721]), .rectangle1_weight(rectangle1_weights[1721]), .rectangle2_x(rectangle2_xs[1721]), .rectangle2_y(rectangle2_ys[1721]), .rectangle2_width(rectangle2_widths[1721]), .rectangle2_height(rectangle2_heights[1721]), .rectangle2_weight(rectangle2_weights[1721]), .rectangle3_x(rectangle3_xs[1721]), .rectangle3_y(rectangle3_ys[1721]), .rectangle3_width(rectangle3_widths[1721]), .rectangle3_height(rectangle3_heights[1721]), .rectangle3_weight(rectangle3_weights[1721]), .feature_threshold(feature_thresholds[1721]), .feature_above(feature_aboves[1721]), .feature_below(feature_belows[1721]), .scan_win_std_dev(scan_win_std_dev[1721]), .feature_accum(feature_accums[1721]));
  accum_calculator ac1722(.scan_win(scan_win1722), .rectangle1_x(rectangle1_xs[1722]), .rectangle1_y(rectangle1_ys[1722]), .rectangle1_width(rectangle1_widths[1722]), .rectangle1_height(rectangle1_heights[1722]), .rectangle1_weight(rectangle1_weights[1722]), .rectangle2_x(rectangle2_xs[1722]), .rectangle2_y(rectangle2_ys[1722]), .rectangle2_width(rectangle2_widths[1722]), .rectangle2_height(rectangle2_heights[1722]), .rectangle2_weight(rectangle2_weights[1722]), .rectangle3_x(rectangle3_xs[1722]), .rectangle3_y(rectangle3_ys[1722]), .rectangle3_width(rectangle3_widths[1722]), .rectangle3_height(rectangle3_heights[1722]), .rectangle3_weight(rectangle3_weights[1722]), .feature_threshold(feature_thresholds[1722]), .feature_above(feature_aboves[1722]), .feature_below(feature_belows[1722]), .scan_win_std_dev(scan_win_std_dev[1722]), .feature_accum(feature_accums[1722]));
  accum_calculator ac1723(.scan_win(scan_win1723), .rectangle1_x(rectangle1_xs[1723]), .rectangle1_y(rectangle1_ys[1723]), .rectangle1_width(rectangle1_widths[1723]), .rectangle1_height(rectangle1_heights[1723]), .rectangle1_weight(rectangle1_weights[1723]), .rectangle2_x(rectangle2_xs[1723]), .rectangle2_y(rectangle2_ys[1723]), .rectangle2_width(rectangle2_widths[1723]), .rectangle2_height(rectangle2_heights[1723]), .rectangle2_weight(rectangle2_weights[1723]), .rectangle3_x(rectangle3_xs[1723]), .rectangle3_y(rectangle3_ys[1723]), .rectangle3_width(rectangle3_widths[1723]), .rectangle3_height(rectangle3_heights[1723]), .rectangle3_weight(rectangle3_weights[1723]), .feature_threshold(feature_thresholds[1723]), .feature_above(feature_aboves[1723]), .feature_below(feature_belows[1723]), .scan_win_std_dev(scan_win_std_dev[1723]), .feature_accum(feature_accums[1723]));
  accum_calculator ac1724(.scan_win(scan_win1724), .rectangle1_x(rectangle1_xs[1724]), .rectangle1_y(rectangle1_ys[1724]), .rectangle1_width(rectangle1_widths[1724]), .rectangle1_height(rectangle1_heights[1724]), .rectangle1_weight(rectangle1_weights[1724]), .rectangle2_x(rectangle2_xs[1724]), .rectangle2_y(rectangle2_ys[1724]), .rectangle2_width(rectangle2_widths[1724]), .rectangle2_height(rectangle2_heights[1724]), .rectangle2_weight(rectangle2_weights[1724]), .rectangle3_x(rectangle3_xs[1724]), .rectangle3_y(rectangle3_ys[1724]), .rectangle3_width(rectangle3_widths[1724]), .rectangle3_height(rectangle3_heights[1724]), .rectangle3_weight(rectangle3_weights[1724]), .feature_threshold(feature_thresholds[1724]), .feature_above(feature_aboves[1724]), .feature_below(feature_belows[1724]), .scan_win_std_dev(scan_win_std_dev[1724]), .feature_accum(feature_accums[1724]));
  accum_calculator ac1725(.scan_win(scan_win1725), .rectangle1_x(rectangle1_xs[1725]), .rectangle1_y(rectangle1_ys[1725]), .rectangle1_width(rectangle1_widths[1725]), .rectangle1_height(rectangle1_heights[1725]), .rectangle1_weight(rectangle1_weights[1725]), .rectangle2_x(rectangle2_xs[1725]), .rectangle2_y(rectangle2_ys[1725]), .rectangle2_width(rectangle2_widths[1725]), .rectangle2_height(rectangle2_heights[1725]), .rectangle2_weight(rectangle2_weights[1725]), .rectangle3_x(rectangle3_xs[1725]), .rectangle3_y(rectangle3_ys[1725]), .rectangle3_width(rectangle3_widths[1725]), .rectangle3_height(rectangle3_heights[1725]), .rectangle3_weight(rectangle3_weights[1725]), .feature_threshold(feature_thresholds[1725]), .feature_above(feature_aboves[1725]), .feature_below(feature_belows[1725]), .scan_win_std_dev(scan_win_std_dev[1725]), .feature_accum(feature_accums[1725]));
  accum_calculator ac1726(.scan_win(scan_win1726), .rectangle1_x(rectangle1_xs[1726]), .rectangle1_y(rectangle1_ys[1726]), .rectangle1_width(rectangle1_widths[1726]), .rectangle1_height(rectangle1_heights[1726]), .rectangle1_weight(rectangle1_weights[1726]), .rectangle2_x(rectangle2_xs[1726]), .rectangle2_y(rectangle2_ys[1726]), .rectangle2_width(rectangle2_widths[1726]), .rectangle2_height(rectangle2_heights[1726]), .rectangle2_weight(rectangle2_weights[1726]), .rectangle3_x(rectangle3_xs[1726]), .rectangle3_y(rectangle3_ys[1726]), .rectangle3_width(rectangle3_widths[1726]), .rectangle3_height(rectangle3_heights[1726]), .rectangle3_weight(rectangle3_weights[1726]), .feature_threshold(feature_thresholds[1726]), .feature_above(feature_aboves[1726]), .feature_below(feature_belows[1726]), .scan_win_std_dev(scan_win_std_dev[1726]), .feature_accum(feature_accums[1726]));
  accum_calculator ac1727(.scan_win(scan_win1727), .rectangle1_x(rectangle1_xs[1727]), .rectangle1_y(rectangle1_ys[1727]), .rectangle1_width(rectangle1_widths[1727]), .rectangle1_height(rectangle1_heights[1727]), .rectangle1_weight(rectangle1_weights[1727]), .rectangle2_x(rectangle2_xs[1727]), .rectangle2_y(rectangle2_ys[1727]), .rectangle2_width(rectangle2_widths[1727]), .rectangle2_height(rectangle2_heights[1727]), .rectangle2_weight(rectangle2_weights[1727]), .rectangle3_x(rectangle3_xs[1727]), .rectangle3_y(rectangle3_ys[1727]), .rectangle3_width(rectangle3_widths[1727]), .rectangle3_height(rectangle3_heights[1727]), .rectangle3_weight(rectangle3_weights[1727]), .feature_threshold(feature_thresholds[1727]), .feature_above(feature_aboves[1727]), .feature_below(feature_belows[1727]), .scan_win_std_dev(scan_win_std_dev[1727]), .feature_accum(feature_accums[1727]));
  accum_calculator ac1728(.scan_win(scan_win1728), .rectangle1_x(rectangle1_xs[1728]), .rectangle1_y(rectangle1_ys[1728]), .rectangle1_width(rectangle1_widths[1728]), .rectangle1_height(rectangle1_heights[1728]), .rectangle1_weight(rectangle1_weights[1728]), .rectangle2_x(rectangle2_xs[1728]), .rectangle2_y(rectangle2_ys[1728]), .rectangle2_width(rectangle2_widths[1728]), .rectangle2_height(rectangle2_heights[1728]), .rectangle2_weight(rectangle2_weights[1728]), .rectangle3_x(rectangle3_xs[1728]), .rectangle3_y(rectangle3_ys[1728]), .rectangle3_width(rectangle3_widths[1728]), .rectangle3_height(rectangle3_heights[1728]), .rectangle3_weight(rectangle3_weights[1728]), .feature_threshold(feature_thresholds[1728]), .feature_above(feature_aboves[1728]), .feature_below(feature_belows[1728]), .scan_win_std_dev(scan_win_std_dev[1728]), .feature_accum(feature_accums[1728]));
  accum_calculator ac1729(.scan_win(scan_win1729), .rectangle1_x(rectangle1_xs[1729]), .rectangle1_y(rectangle1_ys[1729]), .rectangle1_width(rectangle1_widths[1729]), .rectangle1_height(rectangle1_heights[1729]), .rectangle1_weight(rectangle1_weights[1729]), .rectangle2_x(rectangle2_xs[1729]), .rectangle2_y(rectangle2_ys[1729]), .rectangle2_width(rectangle2_widths[1729]), .rectangle2_height(rectangle2_heights[1729]), .rectangle2_weight(rectangle2_weights[1729]), .rectangle3_x(rectangle3_xs[1729]), .rectangle3_y(rectangle3_ys[1729]), .rectangle3_width(rectangle3_widths[1729]), .rectangle3_height(rectangle3_heights[1729]), .rectangle3_weight(rectangle3_weights[1729]), .feature_threshold(feature_thresholds[1729]), .feature_above(feature_aboves[1729]), .feature_below(feature_belows[1729]), .scan_win_std_dev(scan_win_std_dev[1729]), .feature_accum(feature_accums[1729]));
  accum_calculator ac1730(.scan_win(scan_win1730), .rectangle1_x(rectangle1_xs[1730]), .rectangle1_y(rectangle1_ys[1730]), .rectangle1_width(rectangle1_widths[1730]), .rectangle1_height(rectangle1_heights[1730]), .rectangle1_weight(rectangle1_weights[1730]), .rectangle2_x(rectangle2_xs[1730]), .rectangle2_y(rectangle2_ys[1730]), .rectangle2_width(rectangle2_widths[1730]), .rectangle2_height(rectangle2_heights[1730]), .rectangle2_weight(rectangle2_weights[1730]), .rectangle3_x(rectangle3_xs[1730]), .rectangle3_y(rectangle3_ys[1730]), .rectangle3_width(rectangle3_widths[1730]), .rectangle3_height(rectangle3_heights[1730]), .rectangle3_weight(rectangle3_weights[1730]), .feature_threshold(feature_thresholds[1730]), .feature_above(feature_aboves[1730]), .feature_below(feature_belows[1730]), .scan_win_std_dev(scan_win_std_dev[1730]), .feature_accum(feature_accums[1730]));
  accum_calculator ac1731(.scan_win(scan_win1731), .rectangle1_x(rectangle1_xs[1731]), .rectangle1_y(rectangle1_ys[1731]), .rectangle1_width(rectangle1_widths[1731]), .rectangle1_height(rectangle1_heights[1731]), .rectangle1_weight(rectangle1_weights[1731]), .rectangle2_x(rectangle2_xs[1731]), .rectangle2_y(rectangle2_ys[1731]), .rectangle2_width(rectangle2_widths[1731]), .rectangle2_height(rectangle2_heights[1731]), .rectangle2_weight(rectangle2_weights[1731]), .rectangle3_x(rectangle3_xs[1731]), .rectangle3_y(rectangle3_ys[1731]), .rectangle3_width(rectangle3_widths[1731]), .rectangle3_height(rectangle3_heights[1731]), .rectangle3_weight(rectangle3_weights[1731]), .feature_threshold(feature_thresholds[1731]), .feature_above(feature_aboves[1731]), .feature_below(feature_belows[1731]), .scan_win_std_dev(scan_win_std_dev[1731]), .feature_accum(feature_accums[1731]));
  accum_calculator ac1732(.scan_win(scan_win1732), .rectangle1_x(rectangle1_xs[1732]), .rectangle1_y(rectangle1_ys[1732]), .rectangle1_width(rectangle1_widths[1732]), .rectangle1_height(rectangle1_heights[1732]), .rectangle1_weight(rectangle1_weights[1732]), .rectangle2_x(rectangle2_xs[1732]), .rectangle2_y(rectangle2_ys[1732]), .rectangle2_width(rectangle2_widths[1732]), .rectangle2_height(rectangle2_heights[1732]), .rectangle2_weight(rectangle2_weights[1732]), .rectangle3_x(rectangle3_xs[1732]), .rectangle3_y(rectangle3_ys[1732]), .rectangle3_width(rectangle3_widths[1732]), .rectangle3_height(rectangle3_heights[1732]), .rectangle3_weight(rectangle3_weights[1732]), .feature_threshold(feature_thresholds[1732]), .feature_above(feature_aboves[1732]), .feature_below(feature_belows[1732]), .scan_win_std_dev(scan_win_std_dev[1732]), .feature_accum(feature_accums[1732]));
  accum_calculator ac1733(.scan_win(scan_win1733), .rectangle1_x(rectangle1_xs[1733]), .rectangle1_y(rectangle1_ys[1733]), .rectangle1_width(rectangle1_widths[1733]), .rectangle1_height(rectangle1_heights[1733]), .rectangle1_weight(rectangle1_weights[1733]), .rectangle2_x(rectangle2_xs[1733]), .rectangle2_y(rectangle2_ys[1733]), .rectangle2_width(rectangle2_widths[1733]), .rectangle2_height(rectangle2_heights[1733]), .rectangle2_weight(rectangle2_weights[1733]), .rectangle3_x(rectangle3_xs[1733]), .rectangle3_y(rectangle3_ys[1733]), .rectangle3_width(rectangle3_widths[1733]), .rectangle3_height(rectangle3_heights[1733]), .rectangle3_weight(rectangle3_weights[1733]), .feature_threshold(feature_thresholds[1733]), .feature_above(feature_aboves[1733]), .feature_below(feature_belows[1733]), .scan_win_std_dev(scan_win_std_dev[1733]), .feature_accum(feature_accums[1733]));
  accum_calculator ac1734(.scan_win(scan_win1734), .rectangle1_x(rectangle1_xs[1734]), .rectangle1_y(rectangle1_ys[1734]), .rectangle1_width(rectangle1_widths[1734]), .rectangle1_height(rectangle1_heights[1734]), .rectangle1_weight(rectangle1_weights[1734]), .rectangle2_x(rectangle2_xs[1734]), .rectangle2_y(rectangle2_ys[1734]), .rectangle2_width(rectangle2_widths[1734]), .rectangle2_height(rectangle2_heights[1734]), .rectangle2_weight(rectangle2_weights[1734]), .rectangle3_x(rectangle3_xs[1734]), .rectangle3_y(rectangle3_ys[1734]), .rectangle3_width(rectangle3_widths[1734]), .rectangle3_height(rectangle3_heights[1734]), .rectangle3_weight(rectangle3_weights[1734]), .feature_threshold(feature_thresholds[1734]), .feature_above(feature_aboves[1734]), .feature_below(feature_belows[1734]), .scan_win_std_dev(scan_win_std_dev[1734]), .feature_accum(feature_accums[1734]));
  accum_calculator ac1735(.scan_win(scan_win1735), .rectangle1_x(rectangle1_xs[1735]), .rectangle1_y(rectangle1_ys[1735]), .rectangle1_width(rectangle1_widths[1735]), .rectangle1_height(rectangle1_heights[1735]), .rectangle1_weight(rectangle1_weights[1735]), .rectangle2_x(rectangle2_xs[1735]), .rectangle2_y(rectangle2_ys[1735]), .rectangle2_width(rectangle2_widths[1735]), .rectangle2_height(rectangle2_heights[1735]), .rectangle2_weight(rectangle2_weights[1735]), .rectangle3_x(rectangle3_xs[1735]), .rectangle3_y(rectangle3_ys[1735]), .rectangle3_width(rectangle3_widths[1735]), .rectangle3_height(rectangle3_heights[1735]), .rectangle3_weight(rectangle3_weights[1735]), .feature_threshold(feature_thresholds[1735]), .feature_above(feature_aboves[1735]), .feature_below(feature_belows[1735]), .scan_win_std_dev(scan_win_std_dev[1735]), .feature_accum(feature_accums[1735]));
  accum_calculator ac1736(.scan_win(scan_win1736), .rectangle1_x(rectangle1_xs[1736]), .rectangle1_y(rectangle1_ys[1736]), .rectangle1_width(rectangle1_widths[1736]), .rectangle1_height(rectangle1_heights[1736]), .rectangle1_weight(rectangle1_weights[1736]), .rectangle2_x(rectangle2_xs[1736]), .rectangle2_y(rectangle2_ys[1736]), .rectangle2_width(rectangle2_widths[1736]), .rectangle2_height(rectangle2_heights[1736]), .rectangle2_weight(rectangle2_weights[1736]), .rectangle3_x(rectangle3_xs[1736]), .rectangle3_y(rectangle3_ys[1736]), .rectangle3_width(rectangle3_widths[1736]), .rectangle3_height(rectangle3_heights[1736]), .rectangle3_weight(rectangle3_weights[1736]), .feature_threshold(feature_thresholds[1736]), .feature_above(feature_aboves[1736]), .feature_below(feature_belows[1736]), .scan_win_std_dev(scan_win_std_dev[1736]), .feature_accum(feature_accums[1736]));
  accum_calculator ac1737(.scan_win(scan_win1737), .rectangle1_x(rectangle1_xs[1737]), .rectangle1_y(rectangle1_ys[1737]), .rectangle1_width(rectangle1_widths[1737]), .rectangle1_height(rectangle1_heights[1737]), .rectangle1_weight(rectangle1_weights[1737]), .rectangle2_x(rectangle2_xs[1737]), .rectangle2_y(rectangle2_ys[1737]), .rectangle2_width(rectangle2_widths[1737]), .rectangle2_height(rectangle2_heights[1737]), .rectangle2_weight(rectangle2_weights[1737]), .rectangle3_x(rectangle3_xs[1737]), .rectangle3_y(rectangle3_ys[1737]), .rectangle3_width(rectangle3_widths[1737]), .rectangle3_height(rectangle3_heights[1737]), .rectangle3_weight(rectangle3_weights[1737]), .feature_threshold(feature_thresholds[1737]), .feature_above(feature_aboves[1737]), .feature_below(feature_belows[1737]), .scan_win_std_dev(scan_win_std_dev[1737]), .feature_accum(feature_accums[1737]));
  accum_calculator ac1738(.scan_win(scan_win1738), .rectangle1_x(rectangle1_xs[1738]), .rectangle1_y(rectangle1_ys[1738]), .rectangle1_width(rectangle1_widths[1738]), .rectangle1_height(rectangle1_heights[1738]), .rectangle1_weight(rectangle1_weights[1738]), .rectangle2_x(rectangle2_xs[1738]), .rectangle2_y(rectangle2_ys[1738]), .rectangle2_width(rectangle2_widths[1738]), .rectangle2_height(rectangle2_heights[1738]), .rectangle2_weight(rectangle2_weights[1738]), .rectangle3_x(rectangle3_xs[1738]), .rectangle3_y(rectangle3_ys[1738]), .rectangle3_width(rectangle3_widths[1738]), .rectangle3_height(rectangle3_heights[1738]), .rectangle3_weight(rectangle3_weights[1738]), .feature_threshold(feature_thresholds[1738]), .feature_above(feature_aboves[1738]), .feature_below(feature_belows[1738]), .scan_win_std_dev(scan_win_std_dev[1738]), .feature_accum(feature_accums[1738]));
  accum_calculator ac1739(.scan_win(scan_win1739), .rectangle1_x(rectangle1_xs[1739]), .rectangle1_y(rectangle1_ys[1739]), .rectangle1_width(rectangle1_widths[1739]), .rectangle1_height(rectangle1_heights[1739]), .rectangle1_weight(rectangle1_weights[1739]), .rectangle2_x(rectangle2_xs[1739]), .rectangle2_y(rectangle2_ys[1739]), .rectangle2_width(rectangle2_widths[1739]), .rectangle2_height(rectangle2_heights[1739]), .rectangle2_weight(rectangle2_weights[1739]), .rectangle3_x(rectangle3_xs[1739]), .rectangle3_y(rectangle3_ys[1739]), .rectangle3_width(rectangle3_widths[1739]), .rectangle3_height(rectangle3_heights[1739]), .rectangle3_weight(rectangle3_weights[1739]), .feature_threshold(feature_thresholds[1739]), .feature_above(feature_aboves[1739]), .feature_below(feature_belows[1739]), .scan_win_std_dev(scan_win_std_dev[1739]), .feature_accum(feature_accums[1739]));
  accum_calculator ac1740(.scan_win(scan_win1740), .rectangle1_x(rectangle1_xs[1740]), .rectangle1_y(rectangle1_ys[1740]), .rectangle1_width(rectangle1_widths[1740]), .rectangle1_height(rectangle1_heights[1740]), .rectangle1_weight(rectangle1_weights[1740]), .rectangle2_x(rectangle2_xs[1740]), .rectangle2_y(rectangle2_ys[1740]), .rectangle2_width(rectangle2_widths[1740]), .rectangle2_height(rectangle2_heights[1740]), .rectangle2_weight(rectangle2_weights[1740]), .rectangle3_x(rectangle3_xs[1740]), .rectangle3_y(rectangle3_ys[1740]), .rectangle3_width(rectangle3_widths[1740]), .rectangle3_height(rectangle3_heights[1740]), .rectangle3_weight(rectangle3_weights[1740]), .feature_threshold(feature_thresholds[1740]), .feature_above(feature_aboves[1740]), .feature_below(feature_belows[1740]), .scan_win_std_dev(scan_win_std_dev[1740]), .feature_accum(feature_accums[1740]));
  accum_calculator ac1741(.scan_win(scan_win1741), .rectangle1_x(rectangle1_xs[1741]), .rectangle1_y(rectangle1_ys[1741]), .rectangle1_width(rectangle1_widths[1741]), .rectangle1_height(rectangle1_heights[1741]), .rectangle1_weight(rectangle1_weights[1741]), .rectangle2_x(rectangle2_xs[1741]), .rectangle2_y(rectangle2_ys[1741]), .rectangle2_width(rectangle2_widths[1741]), .rectangle2_height(rectangle2_heights[1741]), .rectangle2_weight(rectangle2_weights[1741]), .rectangle3_x(rectangle3_xs[1741]), .rectangle3_y(rectangle3_ys[1741]), .rectangle3_width(rectangle3_widths[1741]), .rectangle3_height(rectangle3_heights[1741]), .rectangle3_weight(rectangle3_weights[1741]), .feature_threshold(feature_thresholds[1741]), .feature_above(feature_aboves[1741]), .feature_below(feature_belows[1741]), .scan_win_std_dev(scan_win_std_dev[1741]), .feature_accum(feature_accums[1741]));
  accum_calculator ac1742(.scan_win(scan_win1742), .rectangle1_x(rectangle1_xs[1742]), .rectangle1_y(rectangle1_ys[1742]), .rectangle1_width(rectangle1_widths[1742]), .rectangle1_height(rectangle1_heights[1742]), .rectangle1_weight(rectangle1_weights[1742]), .rectangle2_x(rectangle2_xs[1742]), .rectangle2_y(rectangle2_ys[1742]), .rectangle2_width(rectangle2_widths[1742]), .rectangle2_height(rectangle2_heights[1742]), .rectangle2_weight(rectangle2_weights[1742]), .rectangle3_x(rectangle3_xs[1742]), .rectangle3_y(rectangle3_ys[1742]), .rectangle3_width(rectangle3_widths[1742]), .rectangle3_height(rectangle3_heights[1742]), .rectangle3_weight(rectangle3_weights[1742]), .feature_threshold(feature_thresholds[1742]), .feature_above(feature_aboves[1742]), .feature_below(feature_belows[1742]), .scan_win_std_dev(scan_win_std_dev[1742]), .feature_accum(feature_accums[1742]));
  accum_calculator ac1743(.scan_win(scan_win1743), .rectangle1_x(rectangle1_xs[1743]), .rectangle1_y(rectangle1_ys[1743]), .rectangle1_width(rectangle1_widths[1743]), .rectangle1_height(rectangle1_heights[1743]), .rectangle1_weight(rectangle1_weights[1743]), .rectangle2_x(rectangle2_xs[1743]), .rectangle2_y(rectangle2_ys[1743]), .rectangle2_width(rectangle2_widths[1743]), .rectangle2_height(rectangle2_heights[1743]), .rectangle2_weight(rectangle2_weights[1743]), .rectangle3_x(rectangle3_xs[1743]), .rectangle3_y(rectangle3_ys[1743]), .rectangle3_width(rectangle3_widths[1743]), .rectangle3_height(rectangle3_heights[1743]), .rectangle3_weight(rectangle3_weights[1743]), .feature_threshold(feature_thresholds[1743]), .feature_above(feature_aboves[1743]), .feature_below(feature_belows[1743]), .scan_win_std_dev(scan_win_std_dev[1743]), .feature_accum(feature_accums[1743]));
  accum_calculator ac1744(.scan_win(scan_win1744), .rectangle1_x(rectangle1_xs[1744]), .rectangle1_y(rectangle1_ys[1744]), .rectangle1_width(rectangle1_widths[1744]), .rectangle1_height(rectangle1_heights[1744]), .rectangle1_weight(rectangle1_weights[1744]), .rectangle2_x(rectangle2_xs[1744]), .rectangle2_y(rectangle2_ys[1744]), .rectangle2_width(rectangle2_widths[1744]), .rectangle2_height(rectangle2_heights[1744]), .rectangle2_weight(rectangle2_weights[1744]), .rectangle3_x(rectangle3_xs[1744]), .rectangle3_y(rectangle3_ys[1744]), .rectangle3_width(rectangle3_widths[1744]), .rectangle3_height(rectangle3_heights[1744]), .rectangle3_weight(rectangle3_weights[1744]), .feature_threshold(feature_thresholds[1744]), .feature_above(feature_aboves[1744]), .feature_below(feature_belows[1744]), .scan_win_std_dev(scan_win_std_dev[1744]), .feature_accum(feature_accums[1744]));
  accum_calculator ac1745(.scan_win(scan_win1745), .rectangle1_x(rectangle1_xs[1745]), .rectangle1_y(rectangle1_ys[1745]), .rectangle1_width(rectangle1_widths[1745]), .rectangle1_height(rectangle1_heights[1745]), .rectangle1_weight(rectangle1_weights[1745]), .rectangle2_x(rectangle2_xs[1745]), .rectangle2_y(rectangle2_ys[1745]), .rectangle2_width(rectangle2_widths[1745]), .rectangle2_height(rectangle2_heights[1745]), .rectangle2_weight(rectangle2_weights[1745]), .rectangle3_x(rectangle3_xs[1745]), .rectangle3_y(rectangle3_ys[1745]), .rectangle3_width(rectangle3_widths[1745]), .rectangle3_height(rectangle3_heights[1745]), .rectangle3_weight(rectangle3_weights[1745]), .feature_threshold(feature_thresholds[1745]), .feature_above(feature_aboves[1745]), .feature_below(feature_belows[1745]), .scan_win_std_dev(scan_win_std_dev[1745]), .feature_accum(feature_accums[1745]));
  accum_calculator ac1746(.scan_win(scan_win1746), .rectangle1_x(rectangle1_xs[1746]), .rectangle1_y(rectangle1_ys[1746]), .rectangle1_width(rectangle1_widths[1746]), .rectangle1_height(rectangle1_heights[1746]), .rectangle1_weight(rectangle1_weights[1746]), .rectangle2_x(rectangle2_xs[1746]), .rectangle2_y(rectangle2_ys[1746]), .rectangle2_width(rectangle2_widths[1746]), .rectangle2_height(rectangle2_heights[1746]), .rectangle2_weight(rectangle2_weights[1746]), .rectangle3_x(rectangle3_xs[1746]), .rectangle3_y(rectangle3_ys[1746]), .rectangle3_width(rectangle3_widths[1746]), .rectangle3_height(rectangle3_heights[1746]), .rectangle3_weight(rectangle3_weights[1746]), .feature_threshold(feature_thresholds[1746]), .feature_above(feature_aboves[1746]), .feature_below(feature_belows[1746]), .scan_win_std_dev(scan_win_std_dev[1746]), .feature_accum(feature_accums[1746]));
  accum_calculator ac1747(.scan_win(scan_win1747), .rectangle1_x(rectangle1_xs[1747]), .rectangle1_y(rectangle1_ys[1747]), .rectangle1_width(rectangle1_widths[1747]), .rectangle1_height(rectangle1_heights[1747]), .rectangle1_weight(rectangle1_weights[1747]), .rectangle2_x(rectangle2_xs[1747]), .rectangle2_y(rectangle2_ys[1747]), .rectangle2_width(rectangle2_widths[1747]), .rectangle2_height(rectangle2_heights[1747]), .rectangle2_weight(rectangle2_weights[1747]), .rectangle3_x(rectangle3_xs[1747]), .rectangle3_y(rectangle3_ys[1747]), .rectangle3_width(rectangle3_widths[1747]), .rectangle3_height(rectangle3_heights[1747]), .rectangle3_weight(rectangle3_weights[1747]), .feature_threshold(feature_thresholds[1747]), .feature_above(feature_aboves[1747]), .feature_below(feature_belows[1747]), .scan_win_std_dev(scan_win_std_dev[1747]), .feature_accum(feature_accums[1747]));
  accum_calculator ac1748(.scan_win(scan_win1748), .rectangle1_x(rectangle1_xs[1748]), .rectangle1_y(rectangle1_ys[1748]), .rectangle1_width(rectangle1_widths[1748]), .rectangle1_height(rectangle1_heights[1748]), .rectangle1_weight(rectangle1_weights[1748]), .rectangle2_x(rectangle2_xs[1748]), .rectangle2_y(rectangle2_ys[1748]), .rectangle2_width(rectangle2_widths[1748]), .rectangle2_height(rectangle2_heights[1748]), .rectangle2_weight(rectangle2_weights[1748]), .rectangle3_x(rectangle3_xs[1748]), .rectangle3_y(rectangle3_ys[1748]), .rectangle3_width(rectangle3_widths[1748]), .rectangle3_height(rectangle3_heights[1748]), .rectangle3_weight(rectangle3_weights[1748]), .feature_threshold(feature_thresholds[1748]), .feature_above(feature_aboves[1748]), .feature_below(feature_belows[1748]), .scan_win_std_dev(scan_win_std_dev[1748]), .feature_accum(feature_accums[1748]));
  accum_calculator ac1749(.scan_win(scan_win1749), .rectangle1_x(rectangle1_xs[1749]), .rectangle1_y(rectangle1_ys[1749]), .rectangle1_width(rectangle1_widths[1749]), .rectangle1_height(rectangle1_heights[1749]), .rectangle1_weight(rectangle1_weights[1749]), .rectangle2_x(rectangle2_xs[1749]), .rectangle2_y(rectangle2_ys[1749]), .rectangle2_width(rectangle2_widths[1749]), .rectangle2_height(rectangle2_heights[1749]), .rectangle2_weight(rectangle2_weights[1749]), .rectangle3_x(rectangle3_xs[1749]), .rectangle3_y(rectangle3_ys[1749]), .rectangle3_width(rectangle3_widths[1749]), .rectangle3_height(rectangle3_heights[1749]), .rectangle3_weight(rectangle3_weights[1749]), .feature_threshold(feature_thresholds[1749]), .feature_above(feature_aboves[1749]), .feature_below(feature_belows[1749]), .scan_win_std_dev(scan_win_std_dev[1749]), .feature_accum(feature_accums[1749]));
  accum_calculator ac1750(.scan_win(scan_win1750), .rectangle1_x(rectangle1_xs[1750]), .rectangle1_y(rectangle1_ys[1750]), .rectangle1_width(rectangle1_widths[1750]), .rectangle1_height(rectangle1_heights[1750]), .rectangle1_weight(rectangle1_weights[1750]), .rectangle2_x(rectangle2_xs[1750]), .rectangle2_y(rectangle2_ys[1750]), .rectangle2_width(rectangle2_widths[1750]), .rectangle2_height(rectangle2_heights[1750]), .rectangle2_weight(rectangle2_weights[1750]), .rectangle3_x(rectangle3_xs[1750]), .rectangle3_y(rectangle3_ys[1750]), .rectangle3_width(rectangle3_widths[1750]), .rectangle3_height(rectangle3_heights[1750]), .rectangle3_weight(rectangle3_weights[1750]), .feature_threshold(feature_thresholds[1750]), .feature_above(feature_aboves[1750]), .feature_below(feature_belows[1750]), .scan_win_std_dev(scan_win_std_dev[1750]), .feature_accum(feature_accums[1750]));
  accum_calculator ac1751(.scan_win(scan_win1751), .rectangle1_x(rectangle1_xs[1751]), .rectangle1_y(rectangle1_ys[1751]), .rectangle1_width(rectangle1_widths[1751]), .rectangle1_height(rectangle1_heights[1751]), .rectangle1_weight(rectangle1_weights[1751]), .rectangle2_x(rectangle2_xs[1751]), .rectangle2_y(rectangle2_ys[1751]), .rectangle2_width(rectangle2_widths[1751]), .rectangle2_height(rectangle2_heights[1751]), .rectangle2_weight(rectangle2_weights[1751]), .rectangle3_x(rectangle3_xs[1751]), .rectangle3_y(rectangle3_ys[1751]), .rectangle3_width(rectangle3_widths[1751]), .rectangle3_height(rectangle3_heights[1751]), .rectangle3_weight(rectangle3_weights[1751]), .feature_threshold(feature_thresholds[1751]), .feature_above(feature_aboves[1751]), .feature_below(feature_belows[1751]), .scan_win_std_dev(scan_win_std_dev[1751]), .feature_accum(feature_accums[1751]));
  accum_calculator ac1752(.scan_win(scan_win1752), .rectangle1_x(rectangle1_xs[1752]), .rectangle1_y(rectangle1_ys[1752]), .rectangle1_width(rectangle1_widths[1752]), .rectangle1_height(rectangle1_heights[1752]), .rectangle1_weight(rectangle1_weights[1752]), .rectangle2_x(rectangle2_xs[1752]), .rectangle2_y(rectangle2_ys[1752]), .rectangle2_width(rectangle2_widths[1752]), .rectangle2_height(rectangle2_heights[1752]), .rectangle2_weight(rectangle2_weights[1752]), .rectangle3_x(rectangle3_xs[1752]), .rectangle3_y(rectangle3_ys[1752]), .rectangle3_width(rectangle3_widths[1752]), .rectangle3_height(rectangle3_heights[1752]), .rectangle3_weight(rectangle3_weights[1752]), .feature_threshold(feature_thresholds[1752]), .feature_above(feature_aboves[1752]), .feature_below(feature_belows[1752]), .scan_win_std_dev(scan_win_std_dev[1752]), .feature_accum(feature_accums[1752]));
  accum_calculator ac1753(.scan_win(scan_win1753), .rectangle1_x(rectangle1_xs[1753]), .rectangle1_y(rectangle1_ys[1753]), .rectangle1_width(rectangle1_widths[1753]), .rectangle1_height(rectangle1_heights[1753]), .rectangle1_weight(rectangle1_weights[1753]), .rectangle2_x(rectangle2_xs[1753]), .rectangle2_y(rectangle2_ys[1753]), .rectangle2_width(rectangle2_widths[1753]), .rectangle2_height(rectangle2_heights[1753]), .rectangle2_weight(rectangle2_weights[1753]), .rectangle3_x(rectangle3_xs[1753]), .rectangle3_y(rectangle3_ys[1753]), .rectangle3_width(rectangle3_widths[1753]), .rectangle3_height(rectangle3_heights[1753]), .rectangle3_weight(rectangle3_weights[1753]), .feature_threshold(feature_thresholds[1753]), .feature_above(feature_aboves[1753]), .feature_below(feature_belows[1753]), .scan_win_std_dev(scan_win_std_dev[1753]), .feature_accum(feature_accums[1753]));
  accum_calculator ac1754(.scan_win(scan_win1754), .rectangle1_x(rectangle1_xs[1754]), .rectangle1_y(rectangle1_ys[1754]), .rectangle1_width(rectangle1_widths[1754]), .rectangle1_height(rectangle1_heights[1754]), .rectangle1_weight(rectangle1_weights[1754]), .rectangle2_x(rectangle2_xs[1754]), .rectangle2_y(rectangle2_ys[1754]), .rectangle2_width(rectangle2_widths[1754]), .rectangle2_height(rectangle2_heights[1754]), .rectangle2_weight(rectangle2_weights[1754]), .rectangle3_x(rectangle3_xs[1754]), .rectangle3_y(rectangle3_ys[1754]), .rectangle3_width(rectangle3_widths[1754]), .rectangle3_height(rectangle3_heights[1754]), .rectangle3_weight(rectangle3_weights[1754]), .feature_threshold(feature_thresholds[1754]), .feature_above(feature_aboves[1754]), .feature_below(feature_belows[1754]), .scan_win_std_dev(scan_win_std_dev[1754]), .feature_accum(feature_accums[1754]));
  accum_calculator ac1755(.scan_win(scan_win1755), .rectangle1_x(rectangle1_xs[1755]), .rectangle1_y(rectangle1_ys[1755]), .rectangle1_width(rectangle1_widths[1755]), .rectangle1_height(rectangle1_heights[1755]), .rectangle1_weight(rectangle1_weights[1755]), .rectangle2_x(rectangle2_xs[1755]), .rectangle2_y(rectangle2_ys[1755]), .rectangle2_width(rectangle2_widths[1755]), .rectangle2_height(rectangle2_heights[1755]), .rectangle2_weight(rectangle2_weights[1755]), .rectangle3_x(rectangle3_xs[1755]), .rectangle3_y(rectangle3_ys[1755]), .rectangle3_width(rectangle3_widths[1755]), .rectangle3_height(rectangle3_heights[1755]), .rectangle3_weight(rectangle3_weights[1755]), .feature_threshold(feature_thresholds[1755]), .feature_above(feature_aboves[1755]), .feature_below(feature_belows[1755]), .scan_win_std_dev(scan_win_std_dev[1755]), .feature_accum(feature_accums[1755]));
  accum_calculator ac1756(.scan_win(scan_win1756), .rectangle1_x(rectangle1_xs[1756]), .rectangle1_y(rectangle1_ys[1756]), .rectangle1_width(rectangle1_widths[1756]), .rectangle1_height(rectangle1_heights[1756]), .rectangle1_weight(rectangle1_weights[1756]), .rectangle2_x(rectangle2_xs[1756]), .rectangle2_y(rectangle2_ys[1756]), .rectangle2_width(rectangle2_widths[1756]), .rectangle2_height(rectangle2_heights[1756]), .rectangle2_weight(rectangle2_weights[1756]), .rectangle3_x(rectangle3_xs[1756]), .rectangle3_y(rectangle3_ys[1756]), .rectangle3_width(rectangle3_widths[1756]), .rectangle3_height(rectangle3_heights[1756]), .rectangle3_weight(rectangle3_weights[1756]), .feature_threshold(feature_thresholds[1756]), .feature_above(feature_aboves[1756]), .feature_below(feature_belows[1756]), .scan_win_std_dev(scan_win_std_dev[1756]), .feature_accum(feature_accums[1756]));
  accum_calculator ac1757(.scan_win(scan_win1757), .rectangle1_x(rectangle1_xs[1757]), .rectangle1_y(rectangle1_ys[1757]), .rectangle1_width(rectangle1_widths[1757]), .rectangle1_height(rectangle1_heights[1757]), .rectangle1_weight(rectangle1_weights[1757]), .rectangle2_x(rectangle2_xs[1757]), .rectangle2_y(rectangle2_ys[1757]), .rectangle2_width(rectangle2_widths[1757]), .rectangle2_height(rectangle2_heights[1757]), .rectangle2_weight(rectangle2_weights[1757]), .rectangle3_x(rectangle3_xs[1757]), .rectangle3_y(rectangle3_ys[1757]), .rectangle3_width(rectangle3_widths[1757]), .rectangle3_height(rectangle3_heights[1757]), .rectangle3_weight(rectangle3_weights[1757]), .feature_threshold(feature_thresholds[1757]), .feature_above(feature_aboves[1757]), .feature_below(feature_belows[1757]), .scan_win_std_dev(scan_win_std_dev[1757]), .feature_accum(feature_accums[1757]));
  accum_calculator ac1758(.scan_win(scan_win1758), .rectangle1_x(rectangle1_xs[1758]), .rectangle1_y(rectangle1_ys[1758]), .rectangle1_width(rectangle1_widths[1758]), .rectangle1_height(rectangle1_heights[1758]), .rectangle1_weight(rectangle1_weights[1758]), .rectangle2_x(rectangle2_xs[1758]), .rectangle2_y(rectangle2_ys[1758]), .rectangle2_width(rectangle2_widths[1758]), .rectangle2_height(rectangle2_heights[1758]), .rectangle2_weight(rectangle2_weights[1758]), .rectangle3_x(rectangle3_xs[1758]), .rectangle3_y(rectangle3_ys[1758]), .rectangle3_width(rectangle3_widths[1758]), .rectangle3_height(rectangle3_heights[1758]), .rectangle3_weight(rectangle3_weights[1758]), .feature_threshold(feature_thresholds[1758]), .feature_above(feature_aboves[1758]), .feature_below(feature_belows[1758]), .scan_win_std_dev(scan_win_std_dev[1758]), .feature_accum(feature_accums[1758]));
  accum_calculator ac1759(.scan_win(scan_win1759), .rectangle1_x(rectangle1_xs[1759]), .rectangle1_y(rectangle1_ys[1759]), .rectangle1_width(rectangle1_widths[1759]), .rectangle1_height(rectangle1_heights[1759]), .rectangle1_weight(rectangle1_weights[1759]), .rectangle2_x(rectangle2_xs[1759]), .rectangle2_y(rectangle2_ys[1759]), .rectangle2_width(rectangle2_widths[1759]), .rectangle2_height(rectangle2_heights[1759]), .rectangle2_weight(rectangle2_weights[1759]), .rectangle3_x(rectangle3_xs[1759]), .rectangle3_y(rectangle3_ys[1759]), .rectangle3_width(rectangle3_widths[1759]), .rectangle3_height(rectangle3_heights[1759]), .rectangle3_weight(rectangle3_weights[1759]), .feature_threshold(feature_thresholds[1759]), .feature_above(feature_aboves[1759]), .feature_below(feature_belows[1759]), .scan_win_std_dev(scan_win_std_dev[1759]), .feature_accum(feature_accums[1759]));
  accum_calculator ac1760(.scan_win(scan_win1760), .rectangle1_x(rectangle1_xs[1760]), .rectangle1_y(rectangle1_ys[1760]), .rectangle1_width(rectangle1_widths[1760]), .rectangle1_height(rectangle1_heights[1760]), .rectangle1_weight(rectangle1_weights[1760]), .rectangle2_x(rectangle2_xs[1760]), .rectangle2_y(rectangle2_ys[1760]), .rectangle2_width(rectangle2_widths[1760]), .rectangle2_height(rectangle2_heights[1760]), .rectangle2_weight(rectangle2_weights[1760]), .rectangle3_x(rectangle3_xs[1760]), .rectangle3_y(rectangle3_ys[1760]), .rectangle3_width(rectangle3_widths[1760]), .rectangle3_height(rectangle3_heights[1760]), .rectangle3_weight(rectangle3_weights[1760]), .feature_threshold(feature_thresholds[1760]), .feature_above(feature_aboves[1760]), .feature_below(feature_belows[1760]), .scan_win_std_dev(scan_win_std_dev[1760]), .feature_accum(feature_accums[1760]));
  accum_calculator ac1761(.scan_win(scan_win1761), .rectangle1_x(rectangle1_xs[1761]), .rectangle1_y(rectangle1_ys[1761]), .rectangle1_width(rectangle1_widths[1761]), .rectangle1_height(rectangle1_heights[1761]), .rectangle1_weight(rectangle1_weights[1761]), .rectangle2_x(rectangle2_xs[1761]), .rectangle2_y(rectangle2_ys[1761]), .rectangle2_width(rectangle2_widths[1761]), .rectangle2_height(rectangle2_heights[1761]), .rectangle2_weight(rectangle2_weights[1761]), .rectangle3_x(rectangle3_xs[1761]), .rectangle3_y(rectangle3_ys[1761]), .rectangle3_width(rectangle3_widths[1761]), .rectangle3_height(rectangle3_heights[1761]), .rectangle3_weight(rectangle3_weights[1761]), .feature_threshold(feature_thresholds[1761]), .feature_above(feature_aboves[1761]), .feature_below(feature_belows[1761]), .scan_win_std_dev(scan_win_std_dev[1761]), .feature_accum(feature_accums[1761]));
  accum_calculator ac1762(.scan_win(scan_win1762), .rectangle1_x(rectangle1_xs[1762]), .rectangle1_y(rectangle1_ys[1762]), .rectangle1_width(rectangle1_widths[1762]), .rectangle1_height(rectangle1_heights[1762]), .rectangle1_weight(rectangle1_weights[1762]), .rectangle2_x(rectangle2_xs[1762]), .rectangle2_y(rectangle2_ys[1762]), .rectangle2_width(rectangle2_widths[1762]), .rectangle2_height(rectangle2_heights[1762]), .rectangle2_weight(rectangle2_weights[1762]), .rectangle3_x(rectangle3_xs[1762]), .rectangle3_y(rectangle3_ys[1762]), .rectangle3_width(rectangle3_widths[1762]), .rectangle3_height(rectangle3_heights[1762]), .rectangle3_weight(rectangle3_weights[1762]), .feature_threshold(feature_thresholds[1762]), .feature_above(feature_aboves[1762]), .feature_below(feature_belows[1762]), .scan_win_std_dev(scan_win_std_dev[1762]), .feature_accum(feature_accums[1762]));
  accum_calculator ac1763(.scan_win(scan_win1763), .rectangle1_x(rectangle1_xs[1763]), .rectangle1_y(rectangle1_ys[1763]), .rectangle1_width(rectangle1_widths[1763]), .rectangle1_height(rectangle1_heights[1763]), .rectangle1_weight(rectangle1_weights[1763]), .rectangle2_x(rectangle2_xs[1763]), .rectangle2_y(rectangle2_ys[1763]), .rectangle2_width(rectangle2_widths[1763]), .rectangle2_height(rectangle2_heights[1763]), .rectangle2_weight(rectangle2_weights[1763]), .rectangle3_x(rectangle3_xs[1763]), .rectangle3_y(rectangle3_ys[1763]), .rectangle3_width(rectangle3_widths[1763]), .rectangle3_height(rectangle3_heights[1763]), .rectangle3_weight(rectangle3_weights[1763]), .feature_threshold(feature_thresholds[1763]), .feature_above(feature_aboves[1763]), .feature_below(feature_belows[1763]), .scan_win_std_dev(scan_win_std_dev[1763]), .feature_accum(feature_accums[1763]));
  accum_calculator ac1764(.scan_win(scan_win1764), .rectangle1_x(rectangle1_xs[1764]), .rectangle1_y(rectangle1_ys[1764]), .rectangle1_width(rectangle1_widths[1764]), .rectangle1_height(rectangle1_heights[1764]), .rectangle1_weight(rectangle1_weights[1764]), .rectangle2_x(rectangle2_xs[1764]), .rectangle2_y(rectangle2_ys[1764]), .rectangle2_width(rectangle2_widths[1764]), .rectangle2_height(rectangle2_heights[1764]), .rectangle2_weight(rectangle2_weights[1764]), .rectangle3_x(rectangle3_xs[1764]), .rectangle3_y(rectangle3_ys[1764]), .rectangle3_width(rectangle3_widths[1764]), .rectangle3_height(rectangle3_heights[1764]), .rectangle3_weight(rectangle3_weights[1764]), .feature_threshold(feature_thresholds[1764]), .feature_above(feature_aboves[1764]), .feature_below(feature_belows[1764]), .scan_win_std_dev(scan_win_std_dev[1764]), .feature_accum(feature_accums[1764]));
  accum_calculator ac1765(.scan_win(scan_win1765), .rectangle1_x(rectangle1_xs[1765]), .rectangle1_y(rectangle1_ys[1765]), .rectangle1_width(rectangle1_widths[1765]), .rectangle1_height(rectangle1_heights[1765]), .rectangle1_weight(rectangle1_weights[1765]), .rectangle2_x(rectangle2_xs[1765]), .rectangle2_y(rectangle2_ys[1765]), .rectangle2_width(rectangle2_widths[1765]), .rectangle2_height(rectangle2_heights[1765]), .rectangle2_weight(rectangle2_weights[1765]), .rectangle3_x(rectangle3_xs[1765]), .rectangle3_y(rectangle3_ys[1765]), .rectangle3_width(rectangle3_widths[1765]), .rectangle3_height(rectangle3_heights[1765]), .rectangle3_weight(rectangle3_weights[1765]), .feature_threshold(feature_thresholds[1765]), .feature_above(feature_aboves[1765]), .feature_below(feature_belows[1765]), .scan_win_std_dev(scan_win_std_dev[1765]), .feature_accum(feature_accums[1765]));
  accum_calculator ac1766(.scan_win(scan_win1766), .rectangle1_x(rectangle1_xs[1766]), .rectangle1_y(rectangle1_ys[1766]), .rectangle1_width(rectangle1_widths[1766]), .rectangle1_height(rectangle1_heights[1766]), .rectangle1_weight(rectangle1_weights[1766]), .rectangle2_x(rectangle2_xs[1766]), .rectangle2_y(rectangle2_ys[1766]), .rectangle2_width(rectangle2_widths[1766]), .rectangle2_height(rectangle2_heights[1766]), .rectangle2_weight(rectangle2_weights[1766]), .rectangle3_x(rectangle3_xs[1766]), .rectangle3_y(rectangle3_ys[1766]), .rectangle3_width(rectangle3_widths[1766]), .rectangle3_height(rectangle3_heights[1766]), .rectangle3_weight(rectangle3_weights[1766]), .feature_threshold(feature_thresholds[1766]), .feature_above(feature_aboves[1766]), .feature_below(feature_belows[1766]), .scan_win_std_dev(scan_win_std_dev[1766]), .feature_accum(feature_accums[1766]));
  accum_calculator ac1767(.scan_win(scan_win1767), .rectangle1_x(rectangle1_xs[1767]), .rectangle1_y(rectangle1_ys[1767]), .rectangle1_width(rectangle1_widths[1767]), .rectangle1_height(rectangle1_heights[1767]), .rectangle1_weight(rectangle1_weights[1767]), .rectangle2_x(rectangle2_xs[1767]), .rectangle2_y(rectangle2_ys[1767]), .rectangle2_width(rectangle2_widths[1767]), .rectangle2_height(rectangle2_heights[1767]), .rectangle2_weight(rectangle2_weights[1767]), .rectangle3_x(rectangle3_xs[1767]), .rectangle3_y(rectangle3_ys[1767]), .rectangle3_width(rectangle3_widths[1767]), .rectangle3_height(rectangle3_heights[1767]), .rectangle3_weight(rectangle3_weights[1767]), .feature_threshold(feature_thresholds[1767]), .feature_above(feature_aboves[1767]), .feature_below(feature_belows[1767]), .scan_win_std_dev(scan_win_std_dev[1767]), .feature_accum(feature_accums[1767]));
  accum_calculator ac1768(.scan_win(scan_win1768), .rectangle1_x(rectangle1_xs[1768]), .rectangle1_y(rectangle1_ys[1768]), .rectangle1_width(rectangle1_widths[1768]), .rectangle1_height(rectangle1_heights[1768]), .rectangle1_weight(rectangle1_weights[1768]), .rectangle2_x(rectangle2_xs[1768]), .rectangle2_y(rectangle2_ys[1768]), .rectangle2_width(rectangle2_widths[1768]), .rectangle2_height(rectangle2_heights[1768]), .rectangle2_weight(rectangle2_weights[1768]), .rectangle3_x(rectangle3_xs[1768]), .rectangle3_y(rectangle3_ys[1768]), .rectangle3_width(rectangle3_widths[1768]), .rectangle3_height(rectangle3_heights[1768]), .rectangle3_weight(rectangle3_weights[1768]), .feature_threshold(feature_thresholds[1768]), .feature_above(feature_aboves[1768]), .feature_below(feature_belows[1768]), .scan_win_std_dev(scan_win_std_dev[1768]), .feature_accum(feature_accums[1768]));
  accum_calculator ac1769(.scan_win(scan_win1769), .rectangle1_x(rectangle1_xs[1769]), .rectangle1_y(rectangle1_ys[1769]), .rectangle1_width(rectangle1_widths[1769]), .rectangle1_height(rectangle1_heights[1769]), .rectangle1_weight(rectangle1_weights[1769]), .rectangle2_x(rectangle2_xs[1769]), .rectangle2_y(rectangle2_ys[1769]), .rectangle2_width(rectangle2_widths[1769]), .rectangle2_height(rectangle2_heights[1769]), .rectangle2_weight(rectangle2_weights[1769]), .rectangle3_x(rectangle3_xs[1769]), .rectangle3_y(rectangle3_ys[1769]), .rectangle3_width(rectangle3_widths[1769]), .rectangle3_height(rectangle3_heights[1769]), .rectangle3_weight(rectangle3_weights[1769]), .feature_threshold(feature_thresholds[1769]), .feature_above(feature_aboves[1769]), .feature_below(feature_belows[1769]), .scan_win_std_dev(scan_win_std_dev[1769]), .feature_accum(feature_accums[1769]));
  accum_calculator ac1770(.scan_win(scan_win1770), .rectangle1_x(rectangle1_xs[1770]), .rectangle1_y(rectangle1_ys[1770]), .rectangle1_width(rectangle1_widths[1770]), .rectangle1_height(rectangle1_heights[1770]), .rectangle1_weight(rectangle1_weights[1770]), .rectangle2_x(rectangle2_xs[1770]), .rectangle2_y(rectangle2_ys[1770]), .rectangle2_width(rectangle2_widths[1770]), .rectangle2_height(rectangle2_heights[1770]), .rectangle2_weight(rectangle2_weights[1770]), .rectangle3_x(rectangle3_xs[1770]), .rectangle3_y(rectangle3_ys[1770]), .rectangle3_width(rectangle3_widths[1770]), .rectangle3_height(rectangle3_heights[1770]), .rectangle3_weight(rectangle3_weights[1770]), .feature_threshold(feature_thresholds[1770]), .feature_above(feature_aboves[1770]), .feature_below(feature_belows[1770]), .scan_win_std_dev(scan_win_std_dev[1770]), .feature_accum(feature_accums[1770]));
  accum_calculator ac1771(.scan_win(scan_win1771), .rectangle1_x(rectangle1_xs[1771]), .rectangle1_y(rectangle1_ys[1771]), .rectangle1_width(rectangle1_widths[1771]), .rectangle1_height(rectangle1_heights[1771]), .rectangle1_weight(rectangle1_weights[1771]), .rectangle2_x(rectangle2_xs[1771]), .rectangle2_y(rectangle2_ys[1771]), .rectangle2_width(rectangle2_widths[1771]), .rectangle2_height(rectangle2_heights[1771]), .rectangle2_weight(rectangle2_weights[1771]), .rectangle3_x(rectangle3_xs[1771]), .rectangle3_y(rectangle3_ys[1771]), .rectangle3_width(rectangle3_widths[1771]), .rectangle3_height(rectangle3_heights[1771]), .rectangle3_weight(rectangle3_weights[1771]), .feature_threshold(feature_thresholds[1771]), .feature_above(feature_aboves[1771]), .feature_below(feature_belows[1771]), .scan_win_std_dev(scan_win_std_dev[1771]), .feature_accum(feature_accums[1771]));
  accum_calculator ac1772(.scan_win(scan_win1772), .rectangle1_x(rectangle1_xs[1772]), .rectangle1_y(rectangle1_ys[1772]), .rectangle1_width(rectangle1_widths[1772]), .rectangle1_height(rectangle1_heights[1772]), .rectangle1_weight(rectangle1_weights[1772]), .rectangle2_x(rectangle2_xs[1772]), .rectangle2_y(rectangle2_ys[1772]), .rectangle2_width(rectangle2_widths[1772]), .rectangle2_height(rectangle2_heights[1772]), .rectangle2_weight(rectangle2_weights[1772]), .rectangle3_x(rectangle3_xs[1772]), .rectangle3_y(rectangle3_ys[1772]), .rectangle3_width(rectangle3_widths[1772]), .rectangle3_height(rectangle3_heights[1772]), .rectangle3_weight(rectangle3_weights[1772]), .feature_threshold(feature_thresholds[1772]), .feature_above(feature_aboves[1772]), .feature_below(feature_belows[1772]), .scan_win_std_dev(scan_win_std_dev[1772]), .feature_accum(feature_accums[1772]));
  accum_calculator ac1773(.scan_win(scan_win1773), .rectangle1_x(rectangle1_xs[1773]), .rectangle1_y(rectangle1_ys[1773]), .rectangle1_width(rectangle1_widths[1773]), .rectangle1_height(rectangle1_heights[1773]), .rectangle1_weight(rectangle1_weights[1773]), .rectangle2_x(rectangle2_xs[1773]), .rectangle2_y(rectangle2_ys[1773]), .rectangle2_width(rectangle2_widths[1773]), .rectangle2_height(rectangle2_heights[1773]), .rectangle2_weight(rectangle2_weights[1773]), .rectangle3_x(rectangle3_xs[1773]), .rectangle3_y(rectangle3_ys[1773]), .rectangle3_width(rectangle3_widths[1773]), .rectangle3_height(rectangle3_heights[1773]), .rectangle3_weight(rectangle3_weights[1773]), .feature_threshold(feature_thresholds[1773]), .feature_above(feature_aboves[1773]), .feature_below(feature_belows[1773]), .scan_win_std_dev(scan_win_std_dev[1773]), .feature_accum(feature_accums[1773]));
  accum_calculator ac1774(.scan_win(scan_win1774), .rectangle1_x(rectangle1_xs[1774]), .rectangle1_y(rectangle1_ys[1774]), .rectangle1_width(rectangle1_widths[1774]), .rectangle1_height(rectangle1_heights[1774]), .rectangle1_weight(rectangle1_weights[1774]), .rectangle2_x(rectangle2_xs[1774]), .rectangle2_y(rectangle2_ys[1774]), .rectangle2_width(rectangle2_widths[1774]), .rectangle2_height(rectangle2_heights[1774]), .rectangle2_weight(rectangle2_weights[1774]), .rectangle3_x(rectangle3_xs[1774]), .rectangle3_y(rectangle3_ys[1774]), .rectangle3_width(rectangle3_widths[1774]), .rectangle3_height(rectangle3_heights[1774]), .rectangle3_weight(rectangle3_weights[1774]), .feature_threshold(feature_thresholds[1774]), .feature_above(feature_aboves[1774]), .feature_below(feature_belows[1774]), .scan_win_std_dev(scan_win_std_dev[1774]), .feature_accum(feature_accums[1774]));
  accum_calculator ac1775(.scan_win(scan_win1775), .rectangle1_x(rectangle1_xs[1775]), .rectangle1_y(rectangle1_ys[1775]), .rectangle1_width(rectangle1_widths[1775]), .rectangle1_height(rectangle1_heights[1775]), .rectangle1_weight(rectangle1_weights[1775]), .rectangle2_x(rectangle2_xs[1775]), .rectangle2_y(rectangle2_ys[1775]), .rectangle2_width(rectangle2_widths[1775]), .rectangle2_height(rectangle2_heights[1775]), .rectangle2_weight(rectangle2_weights[1775]), .rectangle3_x(rectangle3_xs[1775]), .rectangle3_y(rectangle3_ys[1775]), .rectangle3_width(rectangle3_widths[1775]), .rectangle3_height(rectangle3_heights[1775]), .rectangle3_weight(rectangle3_weights[1775]), .feature_threshold(feature_thresholds[1775]), .feature_above(feature_aboves[1775]), .feature_below(feature_belows[1775]), .scan_win_std_dev(scan_win_std_dev[1775]), .feature_accum(feature_accums[1775]));
  accum_calculator ac1776(.scan_win(scan_win1776), .rectangle1_x(rectangle1_xs[1776]), .rectangle1_y(rectangle1_ys[1776]), .rectangle1_width(rectangle1_widths[1776]), .rectangle1_height(rectangle1_heights[1776]), .rectangle1_weight(rectangle1_weights[1776]), .rectangle2_x(rectangle2_xs[1776]), .rectangle2_y(rectangle2_ys[1776]), .rectangle2_width(rectangle2_widths[1776]), .rectangle2_height(rectangle2_heights[1776]), .rectangle2_weight(rectangle2_weights[1776]), .rectangle3_x(rectangle3_xs[1776]), .rectangle3_y(rectangle3_ys[1776]), .rectangle3_width(rectangle3_widths[1776]), .rectangle3_height(rectangle3_heights[1776]), .rectangle3_weight(rectangle3_weights[1776]), .feature_threshold(feature_thresholds[1776]), .feature_above(feature_aboves[1776]), .feature_below(feature_belows[1776]), .scan_win_std_dev(scan_win_std_dev[1776]), .feature_accum(feature_accums[1776]));
  accum_calculator ac1777(.scan_win(scan_win1777), .rectangle1_x(rectangle1_xs[1777]), .rectangle1_y(rectangle1_ys[1777]), .rectangle1_width(rectangle1_widths[1777]), .rectangle1_height(rectangle1_heights[1777]), .rectangle1_weight(rectangle1_weights[1777]), .rectangle2_x(rectangle2_xs[1777]), .rectangle2_y(rectangle2_ys[1777]), .rectangle2_width(rectangle2_widths[1777]), .rectangle2_height(rectangle2_heights[1777]), .rectangle2_weight(rectangle2_weights[1777]), .rectangle3_x(rectangle3_xs[1777]), .rectangle3_y(rectangle3_ys[1777]), .rectangle3_width(rectangle3_widths[1777]), .rectangle3_height(rectangle3_heights[1777]), .rectangle3_weight(rectangle3_weights[1777]), .feature_threshold(feature_thresholds[1777]), .feature_above(feature_aboves[1777]), .feature_below(feature_belows[1777]), .scan_win_std_dev(scan_win_std_dev[1777]), .feature_accum(feature_accums[1777]));
  accum_calculator ac1778(.scan_win(scan_win1778), .rectangle1_x(rectangle1_xs[1778]), .rectangle1_y(rectangle1_ys[1778]), .rectangle1_width(rectangle1_widths[1778]), .rectangle1_height(rectangle1_heights[1778]), .rectangle1_weight(rectangle1_weights[1778]), .rectangle2_x(rectangle2_xs[1778]), .rectangle2_y(rectangle2_ys[1778]), .rectangle2_width(rectangle2_widths[1778]), .rectangle2_height(rectangle2_heights[1778]), .rectangle2_weight(rectangle2_weights[1778]), .rectangle3_x(rectangle3_xs[1778]), .rectangle3_y(rectangle3_ys[1778]), .rectangle3_width(rectangle3_widths[1778]), .rectangle3_height(rectangle3_heights[1778]), .rectangle3_weight(rectangle3_weights[1778]), .feature_threshold(feature_thresholds[1778]), .feature_above(feature_aboves[1778]), .feature_below(feature_belows[1778]), .scan_win_std_dev(scan_win_std_dev[1778]), .feature_accum(feature_accums[1778]));
  accum_calculator ac1779(.scan_win(scan_win1779), .rectangle1_x(rectangle1_xs[1779]), .rectangle1_y(rectangle1_ys[1779]), .rectangle1_width(rectangle1_widths[1779]), .rectangle1_height(rectangle1_heights[1779]), .rectangle1_weight(rectangle1_weights[1779]), .rectangle2_x(rectangle2_xs[1779]), .rectangle2_y(rectangle2_ys[1779]), .rectangle2_width(rectangle2_widths[1779]), .rectangle2_height(rectangle2_heights[1779]), .rectangle2_weight(rectangle2_weights[1779]), .rectangle3_x(rectangle3_xs[1779]), .rectangle3_y(rectangle3_ys[1779]), .rectangle3_width(rectangle3_widths[1779]), .rectangle3_height(rectangle3_heights[1779]), .rectangle3_weight(rectangle3_weights[1779]), .feature_threshold(feature_thresholds[1779]), .feature_above(feature_aboves[1779]), .feature_below(feature_belows[1779]), .scan_win_std_dev(scan_win_std_dev[1779]), .feature_accum(feature_accums[1779]));
  accum_calculator ac1780(.scan_win(scan_win1780), .rectangle1_x(rectangle1_xs[1780]), .rectangle1_y(rectangle1_ys[1780]), .rectangle1_width(rectangle1_widths[1780]), .rectangle1_height(rectangle1_heights[1780]), .rectangle1_weight(rectangle1_weights[1780]), .rectangle2_x(rectangle2_xs[1780]), .rectangle2_y(rectangle2_ys[1780]), .rectangle2_width(rectangle2_widths[1780]), .rectangle2_height(rectangle2_heights[1780]), .rectangle2_weight(rectangle2_weights[1780]), .rectangle3_x(rectangle3_xs[1780]), .rectangle3_y(rectangle3_ys[1780]), .rectangle3_width(rectangle3_widths[1780]), .rectangle3_height(rectangle3_heights[1780]), .rectangle3_weight(rectangle3_weights[1780]), .feature_threshold(feature_thresholds[1780]), .feature_above(feature_aboves[1780]), .feature_below(feature_belows[1780]), .scan_win_std_dev(scan_win_std_dev[1780]), .feature_accum(feature_accums[1780]));
  accum_calculator ac1781(.scan_win(scan_win1781), .rectangle1_x(rectangle1_xs[1781]), .rectangle1_y(rectangle1_ys[1781]), .rectangle1_width(rectangle1_widths[1781]), .rectangle1_height(rectangle1_heights[1781]), .rectangle1_weight(rectangle1_weights[1781]), .rectangle2_x(rectangle2_xs[1781]), .rectangle2_y(rectangle2_ys[1781]), .rectangle2_width(rectangle2_widths[1781]), .rectangle2_height(rectangle2_heights[1781]), .rectangle2_weight(rectangle2_weights[1781]), .rectangle3_x(rectangle3_xs[1781]), .rectangle3_y(rectangle3_ys[1781]), .rectangle3_width(rectangle3_widths[1781]), .rectangle3_height(rectangle3_heights[1781]), .rectangle3_weight(rectangle3_weights[1781]), .feature_threshold(feature_thresholds[1781]), .feature_above(feature_aboves[1781]), .feature_below(feature_belows[1781]), .scan_win_std_dev(scan_win_std_dev[1781]), .feature_accum(feature_accums[1781]));
  accum_calculator ac1782(.scan_win(scan_win1782), .rectangle1_x(rectangle1_xs[1782]), .rectangle1_y(rectangle1_ys[1782]), .rectangle1_width(rectangle1_widths[1782]), .rectangle1_height(rectangle1_heights[1782]), .rectangle1_weight(rectangle1_weights[1782]), .rectangle2_x(rectangle2_xs[1782]), .rectangle2_y(rectangle2_ys[1782]), .rectangle2_width(rectangle2_widths[1782]), .rectangle2_height(rectangle2_heights[1782]), .rectangle2_weight(rectangle2_weights[1782]), .rectangle3_x(rectangle3_xs[1782]), .rectangle3_y(rectangle3_ys[1782]), .rectangle3_width(rectangle3_widths[1782]), .rectangle3_height(rectangle3_heights[1782]), .rectangle3_weight(rectangle3_weights[1782]), .feature_threshold(feature_thresholds[1782]), .feature_above(feature_aboves[1782]), .feature_below(feature_belows[1782]), .scan_win_std_dev(scan_win_std_dev[1782]), .feature_accum(feature_accums[1782]));
  accum_calculator ac1783(.scan_win(scan_win1783), .rectangle1_x(rectangle1_xs[1783]), .rectangle1_y(rectangle1_ys[1783]), .rectangle1_width(rectangle1_widths[1783]), .rectangle1_height(rectangle1_heights[1783]), .rectangle1_weight(rectangle1_weights[1783]), .rectangle2_x(rectangle2_xs[1783]), .rectangle2_y(rectangle2_ys[1783]), .rectangle2_width(rectangle2_widths[1783]), .rectangle2_height(rectangle2_heights[1783]), .rectangle2_weight(rectangle2_weights[1783]), .rectangle3_x(rectangle3_xs[1783]), .rectangle3_y(rectangle3_ys[1783]), .rectangle3_width(rectangle3_widths[1783]), .rectangle3_height(rectangle3_heights[1783]), .rectangle3_weight(rectangle3_weights[1783]), .feature_threshold(feature_thresholds[1783]), .feature_above(feature_aboves[1783]), .feature_below(feature_belows[1783]), .scan_win_std_dev(scan_win_std_dev[1783]), .feature_accum(feature_accums[1783]));
  accum_calculator ac1784(.scan_win(scan_win1784), .rectangle1_x(rectangle1_xs[1784]), .rectangle1_y(rectangle1_ys[1784]), .rectangle1_width(rectangle1_widths[1784]), .rectangle1_height(rectangle1_heights[1784]), .rectangle1_weight(rectangle1_weights[1784]), .rectangle2_x(rectangle2_xs[1784]), .rectangle2_y(rectangle2_ys[1784]), .rectangle2_width(rectangle2_widths[1784]), .rectangle2_height(rectangle2_heights[1784]), .rectangle2_weight(rectangle2_weights[1784]), .rectangle3_x(rectangle3_xs[1784]), .rectangle3_y(rectangle3_ys[1784]), .rectangle3_width(rectangle3_widths[1784]), .rectangle3_height(rectangle3_heights[1784]), .rectangle3_weight(rectangle3_weights[1784]), .feature_threshold(feature_thresholds[1784]), .feature_above(feature_aboves[1784]), .feature_below(feature_belows[1784]), .scan_win_std_dev(scan_win_std_dev[1784]), .feature_accum(feature_accums[1784]));
  accum_calculator ac1785(.scan_win(scan_win1785), .rectangle1_x(rectangle1_xs[1785]), .rectangle1_y(rectangle1_ys[1785]), .rectangle1_width(rectangle1_widths[1785]), .rectangle1_height(rectangle1_heights[1785]), .rectangle1_weight(rectangle1_weights[1785]), .rectangle2_x(rectangle2_xs[1785]), .rectangle2_y(rectangle2_ys[1785]), .rectangle2_width(rectangle2_widths[1785]), .rectangle2_height(rectangle2_heights[1785]), .rectangle2_weight(rectangle2_weights[1785]), .rectangle3_x(rectangle3_xs[1785]), .rectangle3_y(rectangle3_ys[1785]), .rectangle3_width(rectangle3_widths[1785]), .rectangle3_height(rectangle3_heights[1785]), .rectangle3_weight(rectangle3_weights[1785]), .feature_threshold(feature_thresholds[1785]), .feature_above(feature_aboves[1785]), .feature_below(feature_belows[1785]), .scan_win_std_dev(scan_win_std_dev[1785]), .feature_accum(feature_accums[1785]));
  accum_calculator ac1786(.scan_win(scan_win1786), .rectangle1_x(rectangle1_xs[1786]), .rectangle1_y(rectangle1_ys[1786]), .rectangle1_width(rectangle1_widths[1786]), .rectangle1_height(rectangle1_heights[1786]), .rectangle1_weight(rectangle1_weights[1786]), .rectangle2_x(rectangle2_xs[1786]), .rectangle2_y(rectangle2_ys[1786]), .rectangle2_width(rectangle2_widths[1786]), .rectangle2_height(rectangle2_heights[1786]), .rectangle2_weight(rectangle2_weights[1786]), .rectangle3_x(rectangle3_xs[1786]), .rectangle3_y(rectangle3_ys[1786]), .rectangle3_width(rectangle3_widths[1786]), .rectangle3_height(rectangle3_heights[1786]), .rectangle3_weight(rectangle3_weights[1786]), .feature_threshold(feature_thresholds[1786]), .feature_above(feature_aboves[1786]), .feature_below(feature_belows[1786]), .scan_win_std_dev(scan_win_std_dev[1786]), .feature_accum(feature_accums[1786]));
  accum_calculator ac1787(.scan_win(scan_win1787), .rectangle1_x(rectangle1_xs[1787]), .rectangle1_y(rectangle1_ys[1787]), .rectangle1_width(rectangle1_widths[1787]), .rectangle1_height(rectangle1_heights[1787]), .rectangle1_weight(rectangle1_weights[1787]), .rectangle2_x(rectangle2_xs[1787]), .rectangle2_y(rectangle2_ys[1787]), .rectangle2_width(rectangle2_widths[1787]), .rectangle2_height(rectangle2_heights[1787]), .rectangle2_weight(rectangle2_weights[1787]), .rectangle3_x(rectangle3_xs[1787]), .rectangle3_y(rectangle3_ys[1787]), .rectangle3_width(rectangle3_widths[1787]), .rectangle3_height(rectangle3_heights[1787]), .rectangle3_weight(rectangle3_weights[1787]), .feature_threshold(feature_thresholds[1787]), .feature_above(feature_aboves[1787]), .feature_below(feature_belows[1787]), .scan_win_std_dev(scan_win_std_dev[1787]), .feature_accum(feature_accums[1787]));
  accum_calculator ac1788(.scan_win(scan_win1788), .rectangle1_x(rectangle1_xs[1788]), .rectangle1_y(rectangle1_ys[1788]), .rectangle1_width(rectangle1_widths[1788]), .rectangle1_height(rectangle1_heights[1788]), .rectangle1_weight(rectangle1_weights[1788]), .rectangle2_x(rectangle2_xs[1788]), .rectangle2_y(rectangle2_ys[1788]), .rectangle2_width(rectangle2_widths[1788]), .rectangle2_height(rectangle2_heights[1788]), .rectangle2_weight(rectangle2_weights[1788]), .rectangle3_x(rectangle3_xs[1788]), .rectangle3_y(rectangle3_ys[1788]), .rectangle3_width(rectangle3_widths[1788]), .rectangle3_height(rectangle3_heights[1788]), .rectangle3_weight(rectangle3_weights[1788]), .feature_threshold(feature_thresholds[1788]), .feature_above(feature_aboves[1788]), .feature_below(feature_belows[1788]), .scan_win_std_dev(scan_win_std_dev[1788]), .feature_accum(feature_accums[1788]));
  accum_calculator ac1789(.scan_win(scan_win1789), .rectangle1_x(rectangle1_xs[1789]), .rectangle1_y(rectangle1_ys[1789]), .rectangle1_width(rectangle1_widths[1789]), .rectangle1_height(rectangle1_heights[1789]), .rectangle1_weight(rectangle1_weights[1789]), .rectangle2_x(rectangle2_xs[1789]), .rectangle2_y(rectangle2_ys[1789]), .rectangle2_width(rectangle2_widths[1789]), .rectangle2_height(rectangle2_heights[1789]), .rectangle2_weight(rectangle2_weights[1789]), .rectangle3_x(rectangle3_xs[1789]), .rectangle3_y(rectangle3_ys[1789]), .rectangle3_width(rectangle3_widths[1789]), .rectangle3_height(rectangle3_heights[1789]), .rectangle3_weight(rectangle3_weights[1789]), .feature_threshold(feature_thresholds[1789]), .feature_above(feature_aboves[1789]), .feature_below(feature_belows[1789]), .scan_win_std_dev(scan_win_std_dev[1789]), .feature_accum(feature_accums[1789]));
  accum_calculator ac1790(.scan_win(scan_win1790), .rectangle1_x(rectangle1_xs[1790]), .rectangle1_y(rectangle1_ys[1790]), .rectangle1_width(rectangle1_widths[1790]), .rectangle1_height(rectangle1_heights[1790]), .rectangle1_weight(rectangle1_weights[1790]), .rectangle2_x(rectangle2_xs[1790]), .rectangle2_y(rectangle2_ys[1790]), .rectangle2_width(rectangle2_widths[1790]), .rectangle2_height(rectangle2_heights[1790]), .rectangle2_weight(rectangle2_weights[1790]), .rectangle3_x(rectangle3_xs[1790]), .rectangle3_y(rectangle3_ys[1790]), .rectangle3_width(rectangle3_widths[1790]), .rectangle3_height(rectangle3_heights[1790]), .rectangle3_weight(rectangle3_weights[1790]), .feature_threshold(feature_thresholds[1790]), .feature_above(feature_aboves[1790]), .feature_below(feature_belows[1790]), .scan_win_std_dev(scan_win_std_dev[1790]), .feature_accum(feature_accums[1790]));
  accum_calculator ac1791(.scan_win(scan_win1791), .rectangle1_x(rectangle1_xs[1791]), .rectangle1_y(rectangle1_ys[1791]), .rectangle1_width(rectangle1_widths[1791]), .rectangle1_height(rectangle1_heights[1791]), .rectangle1_weight(rectangle1_weights[1791]), .rectangle2_x(rectangle2_xs[1791]), .rectangle2_y(rectangle2_ys[1791]), .rectangle2_width(rectangle2_widths[1791]), .rectangle2_height(rectangle2_heights[1791]), .rectangle2_weight(rectangle2_weights[1791]), .rectangle3_x(rectangle3_xs[1791]), .rectangle3_y(rectangle3_ys[1791]), .rectangle3_width(rectangle3_widths[1791]), .rectangle3_height(rectangle3_heights[1791]), .rectangle3_weight(rectangle3_weights[1791]), .feature_threshold(feature_thresholds[1791]), .feature_above(feature_aboves[1791]), .feature_below(feature_belows[1791]), .scan_win_std_dev(scan_win_std_dev[1791]), .feature_accum(feature_accums[1791]));
  accum_calculator ac1792(.scan_win(scan_win1792), .rectangle1_x(rectangle1_xs[1792]), .rectangle1_y(rectangle1_ys[1792]), .rectangle1_width(rectangle1_widths[1792]), .rectangle1_height(rectangle1_heights[1792]), .rectangle1_weight(rectangle1_weights[1792]), .rectangle2_x(rectangle2_xs[1792]), .rectangle2_y(rectangle2_ys[1792]), .rectangle2_width(rectangle2_widths[1792]), .rectangle2_height(rectangle2_heights[1792]), .rectangle2_weight(rectangle2_weights[1792]), .rectangle3_x(rectangle3_xs[1792]), .rectangle3_y(rectangle3_ys[1792]), .rectangle3_width(rectangle3_widths[1792]), .rectangle3_height(rectangle3_heights[1792]), .rectangle3_weight(rectangle3_weights[1792]), .feature_threshold(feature_thresholds[1792]), .feature_above(feature_aboves[1792]), .feature_below(feature_belows[1792]), .scan_win_std_dev(scan_win_std_dev[1792]), .feature_accum(feature_accums[1792]));
  accum_calculator ac1793(.scan_win(scan_win1793), .rectangle1_x(rectangle1_xs[1793]), .rectangle1_y(rectangle1_ys[1793]), .rectangle1_width(rectangle1_widths[1793]), .rectangle1_height(rectangle1_heights[1793]), .rectangle1_weight(rectangle1_weights[1793]), .rectangle2_x(rectangle2_xs[1793]), .rectangle2_y(rectangle2_ys[1793]), .rectangle2_width(rectangle2_widths[1793]), .rectangle2_height(rectangle2_heights[1793]), .rectangle2_weight(rectangle2_weights[1793]), .rectangle3_x(rectangle3_xs[1793]), .rectangle3_y(rectangle3_ys[1793]), .rectangle3_width(rectangle3_widths[1793]), .rectangle3_height(rectangle3_heights[1793]), .rectangle3_weight(rectangle3_weights[1793]), .feature_threshold(feature_thresholds[1793]), .feature_above(feature_aboves[1793]), .feature_below(feature_belows[1793]), .scan_win_std_dev(scan_win_std_dev[1793]), .feature_accum(feature_accums[1793]));
  accum_calculator ac1794(.scan_win(scan_win1794), .rectangle1_x(rectangle1_xs[1794]), .rectangle1_y(rectangle1_ys[1794]), .rectangle1_width(rectangle1_widths[1794]), .rectangle1_height(rectangle1_heights[1794]), .rectangle1_weight(rectangle1_weights[1794]), .rectangle2_x(rectangle2_xs[1794]), .rectangle2_y(rectangle2_ys[1794]), .rectangle2_width(rectangle2_widths[1794]), .rectangle2_height(rectangle2_heights[1794]), .rectangle2_weight(rectangle2_weights[1794]), .rectangle3_x(rectangle3_xs[1794]), .rectangle3_y(rectangle3_ys[1794]), .rectangle3_width(rectangle3_widths[1794]), .rectangle3_height(rectangle3_heights[1794]), .rectangle3_weight(rectangle3_weights[1794]), .feature_threshold(feature_thresholds[1794]), .feature_above(feature_aboves[1794]), .feature_below(feature_belows[1794]), .scan_win_std_dev(scan_win_std_dev[1794]), .feature_accum(feature_accums[1794]));
  accum_calculator ac1795(.scan_win(scan_win1795), .rectangle1_x(rectangle1_xs[1795]), .rectangle1_y(rectangle1_ys[1795]), .rectangle1_width(rectangle1_widths[1795]), .rectangle1_height(rectangle1_heights[1795]), .rectangle1_weight(rectangle1_weights[1795]), .rectangle2_x(rectangle2_xs[1795]), .rectangle2_y(rectangle2_ys[1795]), .rectangle2_width(rectangle2_widths[1795]), .rectangle2_height(rectangle2_heights[1795]), .rectangle2_weight(rectangle2_weights[1795]), .rectangle3_x(rectangle3_xs[1795]), .rectangle3_y(rectangle3_ys[1795]), .rectangle3_width(rectangle3_widths[1795]), .rectangle3_height(rectangle3_heights[1795]), .rectangle3_weight(rectangle3_weights[1795]), .feature_threshold(feature_thresholds[1795]), .feature_above(feature_aboves[1795]), .feature_below(feature_belows[1795]), .scan_win_std_dev(scan_win_std_dev[1795]), .feature_accum(feature_accums[1795]));
  accum_calculator ac1796(.scan_win(scan_win1796), .rectangle1_x(rectangle1_xs[1796]), .rectangle1_y(rectangle1_ys[1796]), .rectangle1_width(rectangle1_widths[1796]), .rectangle1_height(rectangle1_heights[1796]), .rectangle1_weight(rectangle1_weights[1796]), .rectangle2_x(rectangle2_xs[1796]), .rectangle2_y(rectangle2_ys[1796]), .rectangle2_width(rectangle2_widths[1796]), .rectangle2_height(rectangle2_heights[1796]), .rectangle2_weight(rectangle2_weights[1796]), .rectangle3_x(rectangle3_xs[1796]), .rectangle3_y(rectangle3_ys[1796]), .rectangle3_width(rectangle3_widths[1796]), .rectangle3_height(rectangle3_heights[1796]), .rectangle3_weight(rectangle3_weights[1796]), .feature_threshold(feature_thresholds[1796]), .feature_above(feature_aboves[1796]), .feature_below(feature_belows[1796]), .scan_win_std_dev(scan_win_std_dev[1796]), .feature_accum(feature_accums[1796]));
  accum_calculator ac1797(.scan_win(scan_win1797), .rectangle1_x(rectangle1_xs[1797]), .rectangle1_y(rectangle1_ys[1797]), .rectangle1_width(rectangle1_widths[1797]), .rectangle1_height(rectangle1_heights[1797]), .rectangle1_weight(rectangle1_weights[1797]), .rectangle2_x(rectangle2_xs[1797]), .rectangle2_y(rectangle2_ys[1797]), .rectangle2_width(rectangle2_widths[1797]), .rectangle2_height(rectangle2_heights[1797]), .rectangle2_weight(rectangle2_weights[1797]), .rectangle3_x(rectangle3_xs[1797]), .rectangle3_y(rectangle3_ys[1797]), .rectangle3_width(rectangle3_widths[1797]), .rectangle3_height(rectangle3_heights[1797]), .rectangle3_weight(rectangle3_weights[1797]), .feature_threshold(feature_thresholds[1797]), .feature_above(feature_aboves[1797]), .feature_below(feature_belows[1797]), .scan_win_std_dev(scan_win_std_dev[1797]), .feature_accum(feature_accums[1797]));
  accum_calculator ac1798(.scan_win(scan_win1798), .rectangle1_x(rectangle1_xs[1798]), .rectangle1_y(rectangle1_ys[1798]), .rectangle1_width(rectangle1_widths[1798]), .rectangle1_height(rectangle1_heights[1798]), .rectangle1_weight(rectangle1_weights[1798]), .rectangle2_x(rectangle2_xs[1798]), .rectangle2_y(rectangle2_ys[1798]), .rectangle2_width(rectangle2_widths[1798]), .rectangle2_height(rectangle2_heights[1798]), .rectangle2_weight(rectangle2_weights[1798]), .rectangle3_x(rectangle3_xs[1798]), .rectangle3_y(rectangle3_ys[1798]), .rectangle3_width(rectangle3_widths[1798]), .rectangle3_height(rectangle3_heights[1798]), .rectangle3_weight(rectangle3_weights[1798]), .feature_threshold(feature_thresholds[1798]), .feature_above(feature_aboves[1798]), .feature_below(feature_belows[1798]), .scan_win_std_dev(scan_win_std_dev[1798]), .feature_accum(feature_accums[1798]));
  accum_calculator ac1799(.scan_win(scan_win1799), .rectangle1_x(rectangle1_xs[1799]), .rectangle1_y(rectangle1_ys[1799]), .rectangle1_width(rectangle1_widths[1799]), .rectangle1_height(rectangle1_heights[1799]), .rectangle1_weight(rectangle1_weights[1799]), .rectangle2_x(rectangle2_xs[1799]), .rectangle2_y(rectangle2_ys[1799]), .rectangle2_width(rectangle2_widths[1799]), .rectangle2_height(rectangle2_heights[1799]), .rectangle2_weight(rectangle2_weights[1799]), .rectangle3_x(rectangle3_xs[1799]), .rectangle3_y(rectangle3_ys[1799]), .rectangle3_width(rectangle3_widths[1799]), .rectangle3_height(rectangle3_heights[1799]), .rectangle3_weight(rectangle3_weights[1799]), .feature_threshold(feature_thresholds[1799]), .feature_above(feature_aboves[1799]), .feature_below(feature_belows[1799]), .scan_win_std_dev(scan_win_std_dev[1799]), .feature_accum(feature_accums[1799]));
  accum_calculator ac1800(.scan_win(scan_win1800), .rectangle1_x(rectangle1_xs[1800]), .rectangle1_y(rectangle1_ys[1800]), .rectangle1_width(rectangle1_widths[1800]), .rectangle1_height(rectangle1_heights[1800]), .rectangle1_weight(rectangle1_weights[1800]), .rectangle2_x(rectangle2_xs[1800]), .rectangle2_y(rectangle2_ys[1800]), .rectangle2_width(rectangle2_widths[1800]), .rectangle2_height(rectangle2_heights[1800]), .rectangle2_weight(rectangle2_weights[1800]), .rectangle3_x(rectangle3_xs[1800]), .rectangle3_y(rectangle3_ys[1800]), .rectangle3_width(rectangle3_widths[1800]), .rectangle3_height(rectangle3_heights[1800]), .rectangle3_weight(rectangle3_weights[1800]), .feature_threshold(feature_thresholds[1800]), .feature_above(feature_aboves[1800]), .feature_below(feature_belows[1800]), .scan_win_std_dev(scan_win_std_dev[1800]), .feature_accum(feature_accums[1800]));
  accum_calculator ac1801(.scan_win(scan_win1801), .rectangle1_x(rectangle1_xs[1801]), .rectangle1_y(rectangle1_ys[1801]), .rectangle1_width(rectangle1_widths[1801]), .rectangle1_height(rectangle1_heights[1801]), .rectangle1_weight(rectangle1_weights[1801]), .rectangle2_x(rectangle2_xs[1801]), .rectangle2_y(rectangle2_ys[1801]), .rectangle2_width(rectangle2_widths[1801]), .rectangle2_height(rectangle2_heights[1801]), .rectangle2_weight(rectangle2_weights[1801]), .rectangle3_x(rectangle3_xs[1801]), .rectangle3_y(rectangle3_ys[1801]), .rectangle3_width(rectangle3_widths[1801]), .rectangle3_height(rectangle3_heights[1801]), .rectangle3_weight(rectangle3_weights[1801]), .feature_threshold(feature_thresholds[1801]), .feature_above(feature_aboves[1801]), .feature_below(feature_belows[1801]), .scan_win_std_dev(scan_win_std_dev[1801]), .feature_accum(feature_accums[1801]));
  accum_calculator ac1802(.scan_win(scan_win1802), .rectangle1_x(rectangle1_xs[1802]), .rectangle1_y(rectangle1_ys[1802]), .rectangle1_width(rectangle1_widths[1802]), .rectangle1_height(rectangle1_heights[1802]), .rectangle1_weight(rectangle1_weights[1802]), .rectangle2_x(rectangle2_xs[1802]), .rectangle2_y(rectangle2_ys[1802]), .rectangle2_width(rectangle2_widths[1802]), .rectangle2_height(rectangle2_heights[1802]), .rectangle2_weight(rectangle2_weights[1802]), .rectangle3_x(rectangle3_xs[1802]), .rectangle3_y(rectangle3_ys[1802]), .rectangle3_width(rectangle3_widths[1802]), .rectangle3_height(rectangle3_heights[1802]), .rectangle3_weight(rectangle3_weights[1802]), .feature_threshold(feature_thresholds[1802]), .feature_above(feature_aboves[1802]), .feature_below(feature_belows[1802]), .scan_win_std_dev(scan_win_std_dev[1802]), .feature_accum(feature_accums[1802]));
  accum_calculator ac1803(.scan_win(scan_win1803), .rectangle1_x(rectangle1_xs[1803]), .rectangle1_y(rectangle1_ys[1803]), .rectangle1_width(rectangle1_widths[1803]), .rectangle1_height(rectangle1_heights[1803]), .rectangle1_weight(rectangle1_weights[1803]), .rectangle2_x(rectangle2_xs[1803]), .rectangle2_y(rectangle2_ys[1803]), .rectangle2_width(rectangle2_widths[1803]), .rectangle2_height(rectangle2_heights[1803]), .rectangle2_weight(rectangle2_weights[1803]), .rectangle3_x(rectangle3_xs[1803]), .rectangle3_y(rectangle3_ys[1803]), .rectangle3_width(rectangle3_widths[1803]), .rectangle3_height(rectangle3_heights[1803]), .rectangle3_weight(rectangle3_weights[1803]), .feature_threshold(feature_thresholds[1803]), .feature_above(feature_aboves[1803]), .feature_below(feature_belows[1803]), .scan_win_std_dev(scan_win_std_dev[1803]), .feature_accum(feature_accums[1803]));
  accum_calculator ac1804(.scan_win(scan_win1804), .rectangle1_x(rectangle1_xs[1804]), .rectangle1_y(rectangle1_ys[1804]), .rectangle1_width(rectangle1_widths[1804]), .rectangle1_height(rectangle1_heights[1804]), .rectangle1_weight(rectangle1_weights[1804]), .rectangle2_x(rectangle2_xs[1804]), .rectangle2_y(rectangle2_ys[1804]), .rectangle2_width(rectangle2_widths[1804]), .rectangle2_height(rectangle2_heights[1804]), .rectangle2_weight(rectangle2_weights[1804]), .rectangle3_x(rectangle3_xs[1804]), .rectangle3_y(rectangle3_ys[1804]), .rectangle3_width(rectangle3_widths[1804]), .rectangle3_height(rectangle3_heights[1804]), .rectangle3_weight(rectangle3_weights[1804]), .feature_threshold(feature_thresholds[1804]), .feature_above(feature_aboves[1804]), .feature_below(feature_belows[1804]), .scan_win_std_dev(scan_win_std_dev[1804]), .feature_accum(feature_accums[1804]));
  accum_calculator ac1805(.scan_win(scan_win1805), .rectangle1_x(rectangle1_xs[1805]), .rectangle1_y(rectangle1_ys[1805]), .rectangle1_width(rectangle1_widths[1805]), .rectangle1_height(rectangle1_heights[1805]), .rectangle1_weight(rectangle1_weights[1805]), .rectangle2_x(rectangle2_xs[1805]), .rectangle2_y(rectangle2_ys[1805]), .rectangle2_width(rectangle2_widths[1805]), .rectangle2_height(rectangle2_heights[1805]), .rectangle2_weight(rectangle2_weights[1805]), .rectangle3_x(rectangle3_xs[1805]), .rectangle3_y(rectangle3_ys[1805]), .rectangle3_width(rectangle3_widths[1805]), .rectangle3_height(rectangle3_heights[1805]), .rectangle3_weight(rectangle3_weights[1805]), .feature_threshold(feature_thresholds[1805]), .feature_above(feature_aboves[1805]), .feature_below(feature_belows[1805]), .scan_win_std_dev(scan_win_std_dev[1805]), .feature_accum(feature_accums[1805]));
  accum_calculator ac1806(.scan_win(scan_win1806), .rectangle1_x(rectangle1_xs[1806]), .rectangle1_y(rectangle1_ys[1806]), .rectangle1_width(rectangle1_widths[1806]), .rectangle1_height(rectangle1_heights[1806]), .rectangle1_weight(rectangle1_weights[1806]), .rectangle2_x(rectangle2_xs[1806]), .rectangle2_y(rectangle2_ys[1806]), .rectangle2_width(rectangle2_widths[1806]), .rectangle2_height(rectangle2_heights[1806]), .rectangle2_weight(rectangle2_weights[1806]), .rectangle3_x(rectangle3_xs[1806]), .rectangle3_y(rectangle3_ys[1806]), .rectangle3_width(rectangle3_widths[1806]), .rectangle3_height(rectangle3_heights[1806]), .rectangle3_weight(rectangle3_weights[1806]), .feature_threshold(feature_thresholds[1806]), .feature_above(feature_aboves[1806]), .feature_below(feature_belows[1806]), .scan_win_std_dev(scan_win_std_dev[1806]), .feature_accum(feature_accums[1806]));
  accum_calculator ac1807(.scan_win(scan_win1807), .rectangle1_x(rectangle1_xs[1807]), .rectangle1_y(rectangle1_ys[1807]), .rectangle1_width(rectangle1_widths[1807]), .rectangle1_height(rectangle1_heights[1807]), .rectangle1_weight(rectangle1_weights[1807]), .rectangle2_x(rectangle2_xs[1807]), .rectangle2_y(rectangle2_ys[1807]), .rectangle2_width(rectangle2_widths[1807]), .rectangle2_height(rectangle2_heights[1807]), .rectangle2_weight(rectangle2_weights[1807]), .rectangle3_x(rectangle3_xs[1807]), .rectangle3_y(rectangle3_ys[1807]), .rectangle3_width(rectangle3_widths[1807]), .rectangle3_height(rectangle3_heights[1807]), .rectangle3_weight(rectangle3_weights[1807]), .feature_threshold(feature_thresholds[1807]), .feature_above(feature_aboves[1807]), .feature_below(feature_belows[1807]), .scan_win_std_dev(scan_win_std_dev[1807]), .feature_accum(feature_accums[1807]));
  accum_calculator ac1808(.scan_win(scan_win1808), .rectangle1_x(rectangle1_xs[1808]), .rectangle1_y(rectangle1_ys[1808]), .rectangle1_width(rectangle1_widths[1808]), .rectangle1_height(rectangle1_heights[1808]), .rectangle1_weight(rectangle1_weights[1808]), .rectangle2_x(rectangle2_xs[1808]), .rectangle2_y(rectangle2_ys[1808]), .rectangle2_width(rectangle2_widths[1808]), .rectangle2_height(rectangle2_heights[1808]), .rectangle2_weight(rectangle2_weights[1808]), .rectangle3_x(rectangle3_xs[1808]), .rectangle3_y(rectangle3_ys[1808]), .rectangle3_width(rectangle3_widths[1808]), .rectangle3_height(rectangle3_heights[1808]), .rectangle3_weight(rectangle3_weights[1808]), .feature_threshold(feature_thresholds[1808]), .feature_above(feature_aboves[1808]), .feature_below(feature_belows[1808]), .scan_win_std_dev(scan_win_std_dev[1808]), .feature_accum(feature_accums[1808]));
  accum_calculator ac1809(.scan_win(scan_win1809), .rectangle1_x(rectangle1_xs[1809]), .rectangle1_y(rectangle1_ys[1809]), .rectangle1_width(rectangle1_widths[1809]), .rectangle1_height(rectangle1_heights[1809]), .rectangle1_weight(rectangle1_weights[1809]), .rectangle2_x(rectangle2_xs[1809]), .rectangle2_y(rectangle2_ys[1809]), .rectangle2_width(rectangle2_widths[1809]), .rectangle2_height(rectangle2_heights[1809]), .rectangle2_weight(rectangle2_weights[1809]), .rectangle3_x(rectangle3_xs[1809]), .rectangle3_y(rectangle3_ys[1809]), .rectangle3_width(rectangle3_widths[1809]), .rectangle3_height(rectangle3_heights[1809]), .rectangle3_weight(rectangle3_weights[1809]), .feature_threshold(feature_thresholds[1809]), .feature_above(feature_aboves[1809]), .feature_below(feature_belows[1809]), .scan_win_std_dev(scan_win_std_dev[1809]), .feature_accum(feature_accums[1809]));
  accum_calculator ac1810(.scan_win(scan_win1810), .rectangle1_x(rectangle1_xs[1810]), .rectangle1_y(rectangle1_ys[1810]), .rectangle1_width(rectangle1_widths[1810]), .rectangle1_height(rectangle1_heights[1810]), .rectangle1_weight(rectangle1_weights[1810]), .rectangle2_x(rectangle2_xs[1810]), .rectangle2_y(rectangle2_ys[1810]), .rectangle2_width(rectangle2_widths[1810]), .rectangle2_height(rectangle2_heights[1810]), .rectangle2_weight(rectangle2_weights[1810]), .rectangle3_x(rectangle3_xs[1810]), .rectangle3_y(rectangle3_ys[1810]), .rectangle3_width(rectangle3_widths[1810]), .rectangle3_height(rectangle3_heights[1810]), .rectangle3_weight(rectangle3_weights[1810]), .feature_threshold(feature_thresholds[1810]), .feature_above(feature_aboves[1810]), .feature_below(feature_belows[1810]), .scan_win_std_dev(scan_win_std_dev[1810]), .feature_accum(feature_accums[1810]));
  accum_calculator ac1811(.scan_win(scan_win1811), .rectangle1_x(rectangle1_xs[1811]), .rectangle1_y(rectangle1_ys[1811]), .rectangle1_width(rectangle1_widths[1811]), .rectangle1_height(rectangle1_heights[1811]), .rectangle1_weight(rectangle1_weights[1811]), .rectangle2_x(rectangle2_xs[1811]), .rectangle2_y(rectangle2_ys[1811]), .rectangle2_width(rectangle2_widths[1811]), .rectangle2_height(rectangle2_heights[1811]), .rectangle2_weight(rectangle2_weights[1811]), .rectangle3_x(rectangle3_xs[1811]), .rectangle3_y(rectangle3_ys[1811]), .rectangle3_width(rectangle3_widths[1811]), .rectangle3_height(rectangle3_heights[1811]), .rectangle3_weight(rectangle3_weights[1811]), .feature_threshold(feature_thresholds[1811]), .feature_above(feature_aboves[1811]), .feature_below(feature_belows[1811]), .scan_win_std_dev(scan_win_std_dev[1811]), .feature_accum(feature_accums[1811]));
  accum_calculator ac1812(.scan_win(scan_win1812), .rectangle1_x(rectangle1_xs[1812]), .rectangle1_y(rectangle1_ys[1812]), .rectangle1_width(rectangle1_widths[1812]), .rectangle1_height(rectangle1_heights[1812]), .rectangle1_weight(rectangle1_weights[1812]), .rectangle2_x(rectangle2_xs[1812]), .rectangle2_y(rectangle2_ys[1812]), .rectangle2_width(rectangle2_widths[1812]), .rectangle2_height(rectangle2_heights[1812]), .rectangle2_weight(rectangle2_weights[1812]), .rectangle3_x(rectangle3_xs[1812]), .rectangle3_y(rectangle3_ys[1812]), .rectangle3_width(rectangle3_widths[1812]), .rectangle3_height(rectangle3_heights[1812]), .rectangle3_weight(rectangle3_weights[1812]), .feature_threshold(feature_thresholds[1812]), .feature_above(feature_aboves[1812]), .feature_below(feature_belows[1812]), .scan_win_std_dev(scan_win_std_dev[1812]), .feature_accum(feature_accums[1812]));
  accum_calculator ac1813(.scan_win(scan_win1813), .rectangle1_x(rectangle1_xs[1813]), .rectangle1_y(rectangle1_ys[1813]), .rectangle1_width(rectangle1_widths[1813]), .rectangle1_height(rectangle1_heights[1813]), .rectangle1_weight(rectangle1_weights[1813]), .rectangle2_x(rectangle2_xs[1813]), .rectangle2_y(rectangle2_ys[1813]), .rectangle2_width(rectangle2_widths[1813]), .rectangle2_height(rectangle2_heights[1813]), .rectangle2_weight(rectangle2_weights[1813]), .rectangle3_x(rectangle3_xs[1813]), .rectangle3_y(rectangle3_ys[1813]), .rectangle3_width(rectangle3_widths[1813]), .rectangle3_height(rectangle3_heights[1813]), .rectangle3_weight(rectangle3_weights[1813]), .feature_threshold(feature_thresholds[1813]), .feature_above(feature_aboves[1813]), .feature_below(feature_belows[1813]), .scan_win_std_dev(scan_win_std_dev[1813]), .feature_accum(feature_accums[1813]));
  accum_calculator ac1814(.scan_win(scan_win1814), .rectangle1_x(rectangle1_xs[1814]), .rectangle1_y(rectangle1_ys[1814]), .rectangle1_width(rectangle1_widths[1814]), .rectangle1_height(rectangle1_heights[1814]), .rectangle1_weight(rectangle1_weights[1814]), .rectangle2_x(rectangle2_xs[1814]), .rectangle2_y(rectangle2_ys[1814]), .rectangle2_width(rectangle2_widths[1814]), .rectangle2_height(rectangle2_heights[1814]), .rectangle2_weight(rectangle2_weights[1814]), .rectangle3_x(rectangle3_xs[1814]), .rectangle3_y(rectangle3_ys[1814]), .rectangle3_width(rectangle3_widths[1814]), .rectangle3_height(rectangle3_heights[1814]), .rectangle3_weight(rectangle3_weights[1814]), .feature_threshold(feature_thresholds[1814]), .feature_above(feature_aboves[1814]), .feature_below(feature_belows[1814]), .scan_win_std_dev(scan_win_std_dev[1814]), .feature_accum(feature_accums[1814]));
  accum_calculator ac1815(.scan_win(scan_win1815), .rectangle1_x(rectangle1_xs[1815]), .rectangle1_y(rectangle1_ys[1815]), .rectangle1_width(rectangle1_widths[1815]), .rectangle1_height(rectangle1_heights[1815]), .rectangle1_weight(rectangle1_weights[1815]), .rectangle2_x(rectangle2_xs[1815]), .rectangle2_y(rectangle2_ys[1815]), .rectangle2_width(rectangle2_widths[1815]), .rectangle2_height(rectangle2_heights[1815]), .rectangle2_weight(rectangle2_weights[1815]), .rectangle3_x(rectangle3_xs[1815]), .rectangle3_y(rectangle3_ys[1815]), .rectangle3_width(rectangle3_widths[1815]), .rectangle3_height(rectangle3_heights[1815]), .rectangle3_weight(rectangle3_weights[1815]), .feature_threshold(feature_thresholds[1815]), .feature_above(feature_aboves[1815]), .feature_below(feature_belows[1815]), .scan_win_std_dev(scan_win_std_dev[1815]), .feature_accum(feature_accums[1815]));
  accum_calculator ac1816(.scan_win(scan_win1816), .rectangle1_x(rectangle1_xs[1816]), .rectangle1_y(rectangle1_ys[1816]), .rectangle1_width(rectangle1_widths[1816]), .rectangle1_height(rectangle1_heights[1816]), .rectangle1_weight(rectangle1_weights[1816]), .rectangle2_x(rectangle2_xs[1816]), .rectangle2_y(rectangle2_ys[1816]), .rectangle2_width(rectangle2_widths[1816]), .rectangle2_height(rectangle2_heights[1816]), .rectangle2_weight(rectangle2_weights[1816]), .rectangle3_x(rectangle3_xs[1816]), .rectangle3_y(rectangle3_ys[1816]), .rectangle3_width(rectangle3_widths[1816]), .rectangle3_height(rectangle3_heights[1816]), .rectangle3_weight(rectangle3_weights[1816]), .feature_threshold(feature_thresholds[1816]), .feature_above(feature_aboves[1816]), .feature_below(feature_belows[1816]), .scan_win_std_dev(scan_win_std_dev[1816]), .feature_accum(feature_accums[1816]));
  accum_calculator ac1817(.scan_win(scan_win1817), .rectangle1_x(rectangle1_xs[1817]), .rectangle1_y(rectangle1_ys[1817]), .rectangle1_width(rectangle1_widths[1817]), .rectangle1_height(rectangle1_heights[1817]), .rectangle1_weight(rectangle1_weights[1817]), .rectangle2_x(rectangle2_xs[1817]), .rectangle2_y(rectangle2_ys[1817]), .rectangle2_width(rectangle2_widths[1817]), .rectangle2_height(rectangle2_heights[1817]), .rectangle2_weight(rectangle2_weights[1817]), .rectangle3_x(rectangle3_xs[1817]), .rectangle3_y(rectangle3_ys[1817]), .rectangle3_width(rectangle3_widths[1817]), .rectangle3_height(rectangle3_heights[1817]), .rectangle3_weight(rectangle3_weights[1817]), .feature_threshold(feature_thresholds[1817]), .feature_above(feature_aboves[1817]), .feature_below(feature_belows[1817]), .scan_win_std_dev(scan_win_std_dev[1817]), .feature_accum(feature_accums[1817]));
  accum_calculator ac1818(.scan_win(scan_win1818), .rectangle1_x(rectangle1_xs[1818]), .rectangle1_y(rectangle1_ys[1818]), .rectangle1_width(rectangle1_widths[1818]), .rectangle1_height(rectangle1_heights[1818]), .rectangle1_weight(rectangle1_weights[1818]), .rectangle2_x(rectangle2_xs[1818]), .rectangle2_y(rectangle2_ys[1818]), .rectangle2_width(rectangle2_widths[1818]), .rectangle2_height(rectangle2_heights[1818]), .rectangle2_weight(rectangle2_weights[1818]), .rectangle3_x(rectangle3_xs[1818]), .rectangle3_y(rectangle3_ys[1818]), .rectangle3_width(rectangle3_widths[1818]), .rectangle3_height(rectangle3_heights[1818]), .rectangle3_weight(rectangle3_weights[1818]), .feature_threshold(feature_thresholds[1818]), .feature_above(feature_aboves[1818]), .feature_below(feature_belows[1818]), .scan_win_std_dev(scan_win_std_dev[1818]), .feature_accum(feature_accums[1818]));
  accum_calculator ac1819(.scan_win(scan_win1819), .rectangle1_x(rectangle1_xs[1819]), .rectangle1_y(rectangle1_ys[1819]), .rectangle1_width(rectangle1_widths[1819]), .rectangle1_height(rectangle1_heights[1819]), .rectangle1_weight(rectangle1_weights[1819]), .rectangle2_x(rectangle2_xs[1819]), .rectangle2_y(rectangle2_ys[1819]), .rectangle2_width(rectangle2_widths[1819]), .rectangle2_height(rectangle2_heights[1819]), .rectangle2_weight(rectangle2_weights[1819]), .rectangle3_x(rectangle3_xs[1819]), .rectangle3_y(rectangle3_ys[1819]), .rectangle3_width(rectangle3_widths[1819]), .rectangle3_height(rectangle3_heights[1819]), .rectangle3_weight(rectangle3_weights[1819]), .feature_threshold(feature_thresholds[1819]), .feature_above(feature_aboves[1819]), .feature_below(feature_belows[1819]), .scan_win_std_dev(scan_win_std_dev[1819]), .feature_accum(feature_accums[1819]));
  accum_calculator ac1820(.scan_win(scan_win1820), .rectangle1_x(rectangle1_xs[1820]), .rectangle1_y(rectangle1_ys[1820]), .rectangle1_width(rectangle1_widths[1820]), .rectangle1_height(rectangle1_heights[1820]), .rectangle1_weight(rectangle1_weights[1820]), .rectangle2_x(rectangle2_xs[1820]), .rectangle2_y(rectangle2_ys[1820]), .rectangle2_width(rectangle2_widths[1820]), .rectangle2_height(rectangle2_heights[1820]), .rectangle2_weight(rectangle2_weights[1820]), .rectangle3_x(rectangle3_xs[1820]), .rectangle3_y(rectangle3_ys[1820]), .rectangle3_width(rectangle3_widths[1820]), .rectangle3_height(rectangle3_heights[1820]), .rectangle3_weight(rectangle3_weights[1820]), .feature_threshold(feature_thresholds[1820]), .feature_above(feature_aboves[1820]), .feature_below(feature_belows[1820]), .scan_win_std_dev(scan_win_std_dev[1820]), .feature_accum(feature_accums[1820]));
  accum_calculator ac1821(.scan_win(scan_win1821), .rectangle1_x(rectangle1_xs[1821]), .rectangle1_y(rectangle1_ys[1821]), .rectangle1_width(rectangle1_widths[1821]), .rectangle1_height(rectangle1_heights[1821]), .rectangle1_weight(rectangle1_weights[1821]), .rectangle2_x(rectangle2_xs[1821]), .rectangle2_y(rectangle2_ys[1821]), .rectangle2_width(rectangle2_widths[1821]), .rectangle2_height(rectangle2_heights[1821]), .rectangle2_weight(rectangle2_weights[1821]), .rectangle3_x(rectangle3_xs[1821]), .rectangle3_y(rectangle3_ys[1821]), .rectangle3_width(rectangle3_widths[1821]), .rectangle3_height(rectangle3_heights[1821]), .rectangle3_weight(rectangle3_weights[1821]), .feature_threshold(feature_thresholds[1821]), .feature_above(feature_aboves[1821]), .feature_below(feature_belows[1821]), .scan_win_std_dev(scan_win_std_dev[1821]), .feature_accum(feature_accums[1821]));
  accum_calculator ac1822(.scan_win(scan_win1822), .rectangle1_x(rectangle1_xs[1822]), .rectangle1_y(rectangle1_ys[1822]), .rectangle1_width(rectangle1_widths[1822]), .rectangle1_height(rectangle1_heights[1822]), .rectangle1_weight(rectangle1_weights[1822]), .rectangle2_x(rectangle2_xs[1822]), .rectangle2_y(rectangle2_ys[1822]), .rectangle2_width(rectangle2_widths[1822]), .rectangle2_height(rectangle2_heights[1822]), .rectangle2_weight(rectangle2_weights[1822]), .rectangle3_x(rectangle3_xs[1822]), .rectangle3_y(rectangle3_ys[1822]), .rectangle3_width(rectangle3_widths[1822]), .rectangle3_height(rectangle3_heights[1822]), .rectangle3_weight(rectangle3_weights[1822]), .feature_threshold(feature_thresholds[1822]), .feature_above(feature_aboves[1822]), .feature_below(feature_belows[1822]), .scan_win_std_dev(scan_win_std_dev[1822]), .feature_accum(feature_accums[1822]));
  accum_calculator ac1823(.scan_win(scan_win1823), .rectangle1_x(rectangle1_xs[1823]), .rectangle1_y(rectangle1_ys[1823]), .rectangle1_width(rectangle1_widths[1823]), .rectangle1_height(rectangle1_heights[1823]), .rectangle1_weight(rectangle1_weights[1823]), .rectangle2_x(rectangle2_xs[1823]), .rectangle2_y(rectangle2_ys[1823]), .rectangle2_width(rectangle2_widths[1823]), .rectangle2_height(rectangle2_heights[1823]), .rectangle2_weight(rectangle2_weights[1823]), .rectangle3_x(rectangle3_xs[1823]), .rectangle3_y(rectangle3_ys[1823]), .rectangle3_width(rectangle3_widths[1823]), .rectangle3_height(rectangle3_heights[1823]), .rectangle3_weight(rectangle3_weights[1823]), .feature_threshold(feature_thresholds[1823]), .feature_above(feature_aboves[1823]), .feature_below(feature_belows[1823]), .scan_win_std_dev(scan_win_std_dev[1823]), .feature_accum(feature_accums[1823]));
  accum_calculator ac1824(.scan_win(scan_win1824), .rectangle1_x(rectangle1_xs[1824]), .rectangle1_y(rectangle1_ys[1824]), .rectangle1_width(rectangle1_widths[1824]), .rectangle1_height(rectangle1_heights[1824]), .rectangle1_weight(rectangle1_weights[1824]), .rectangle2_x(rectangle2_xs[1824]), .rectangle2_y(rectangle2_ys[1824]), .rectangle2_width(rectangle2_widths[1824]), .rectangle2_height(rectangle2_heights[1824]), .rectangle2_weight(rectangle2_weights[1824]), .rectangle3_x(rectangle3_xs[1824]), .rectangle3_y(rectangle3_ys[1824]), .rectangle3_width(rectangle3_widths[1824]), .rectangle3_height(rectangle3_heights[1824]), .rectangle3_weight(rectangle3_weights[1824]), .feature_threshold(feature_thresholds[1824]), .feature_above(feature_aboves[1824]), .feature_below(feature_belows[1824]), .scan_win_std_dev(scan_win_std_dev[1824]), .feature_accum(feature_accums[1824]));
  accum_calculator ac1825(.scan_win(scan_win1825), .rectangle1_x(rectangle1_xs[1825]), .rectangle1_y(rectangle1_ys[1825]), .rectangle1_width(rectangle1_widths[1825]), .rectangle1_height(rectangle1_heights[1825]), .rectangle1_weight(rectangle1_weights[1825]), .rectangle2_x(rectangle2_xs[1825]), .rectangle2_y(rectangle2_ys[1825]), .rectangle2_width(rectangle2_widths[1825]), .rectangle2_height(rectangle2_heights[1825]), .rectangle2_weight(rectangle2_weights[1825]), .rectangle3_x(rectangle3_xs[1825]), .rectangle3_y(rectangle3_ys[1825]), .rectangle3_width(rectangle3_widths[1825]), .rectangle3_height(rectangle3_heights[1825]), .rectangle3_weight(rectangle3_weights[1825]), .feature_threshold(feature_thresholds[1825]), .feature_above(feature_aboves[1825]), .feature_below(feature_belows[1825]), .scan_win_std_dev(scan_win_std_dev[1825]), .feature_accum(feature_accums[1825]));
  accum_calculator ac1826(.scan_win(scan_win1826), .rectangle1_x(rectangle1_xs[1826]), .rectangle1_y(rectangle1_ys[1826]), .rectangle1_width(rectangle1_widths[1826]), .rectangle1_height(rectangle1_heights[1826]), .rectangle1_weight(rectangle1_weights[1826]), .rectangle2_x(rectangle2_xs[1826]), .rectangle2_y(rectangle2_ys[1826]), .rectangle2_width(rectangle2_widths[1826]), .rectangle2_height(rectangle2_heights[1826]), .rectangle2_weight(rectangle2_weights[1826]), .rectangle3_x(rectangle3_xs[1826]), .rectangle3_y(rectangle3_ys[1826]), .rectangle3_width(rectangle3_widths[1826]), .rectangle3_height(rectangle3_heights[1826]), .rectangle3_weight(rectangle3_weights[1826]), .feature_threshold(feature_thresholds[1826]), .feature_above(feature_aboves[1826]), .feature_below(feature_belows[1826]), .scan_win_std_dev(scan_win_std_dev[1826]), .feature_accum(feature_accums[1826]));
  accum_calculator ac1827(.scan_win(scan_win1827), .rectangle1_x(rectangle1_xs[1827]), .rectangle1_y(rectangle1_ys[1827]), .rectangle1_width(rectangle1_widths[1827]), .rectangle1_height(rectangle1_heights[1827]), .rectangle1_weight(rectangle1_weights[1827]), .rectangle2_x(rectangle2_xs[1827]), .rectangle2_y(rectangle2_ys[1827]), .rectangle2_width(rectangle2_widths[1827]), .rectangle2_height(rectangle2_heights[1827]), .rectangle2_weight(rectangle2_weights[1827]), .rectangle3_x(rectangle3_xs[1827]), .rectangle3_y(rectangle3_ys[1827]), .rectangle3_width(rectangle3_widths[1827]), .rectangle3_height(rectangle3_heights[1827]), .rectangle3_weight(rectangle3_weights[1827]), .feature_threshold(feature_thresholds[1827]), .feature_above(feature_aboves[1827]), .feature_below(feature_belows[1827]), .scan_win_std_dev(scan_win_std_dev[1827]), .feature_accum(feature_accums[1827]));
  accum_calculator ac1828(.scan_win(scan_win1828), .rectangle1_x(rectangle1_xs[1828]), .rectangle1_y(rectangle1_ys[1828]), .rectangle1_width(rectangle1_widths[1828]), .rectangle1_height(rectangle1_heights[1828]), .rectangle1_weight(rectangle1_weights[1828]), .rectangle2_x(rectangle2_xs[1828]), .rectangle2_y(rectangle2_ys[1828]), .rectangle2_width(rectangle2_widths[1828]), .rectangle2_height(rectangle2_heights[1828]), .rectangle2_weight(rectangle2_weights[1828]), .rectangle3_x(rectangle3_xs[1828]), .rectangle3_y(rectangle3_ys[1828]), .rectangle3_width(rectangle3_widths[1828]), .rectangle3_height(rectangle3_heights[1828]), .rectangle3_weight(rectangle3_weights[1828]), .feature_threshold(feature_thresholds[1828]), .feature_above(feature_aboves[1828]), .feature_below(feature_belows[1828]), .scan_win_std_dev(scan_win_std_dev[1828]), .feature_accum(feature_accums[1828]));
  accum_calculator ac1829(.scan_win(scan_win1829), .rectangle1_x(rectangle1_xs[1829]), .rectangle1_y(rectangle1_ys[1829]), .rectangle1_width(rectangle1_widths[1829]), .rectangle1_height(rectangle1_heights[1829]), .rectangle1_weight(rectangle1_weights[1829]), .rectangle2_x(rectangle2_xs[1829]), .rectangle2_y(rectangle2_ys[1829]), .rectangle2_width(rectangle2_widths[1829]), .rectangle2_height(rectangle2_heights[1829]), .rectangle2_weight(rectangle2_weights[1829]), .rectangle3_x(rectangle3_xs[1829]), .rectangle3_y(rectangle3_ys[1829]), .rectangle3_width(rectangle3_widths[1829]), .rectangle3_height(rectangle3_heights[1829]), .rectangle3_weight(rectangle3_weights[1829]), .feature_threshold(feature_thresholds[1829]), .feature_above(feature_aboves[1829]), .feature_below(feature_belows[1829]), .scan_win_std_dev(scan_win_std_dev[1829]), .feature_accum(feature_accums[1829]));
  accum_calculator ac1830(.scan_win(scan_win1830), .rectangle1_x(rectangle1_xs[1830]), .rectangle1_y(rectangle1_ys[1830]), .rectangle1_width(rectangle1_widths[1830]), .rectangle1_height(rectangle1_heights[1830]), .rectangle1_weight(rectangle1_weights[1830]), .rectangle2_x(rectangle2_xs[1830]), .rectangle2_y(rectangle2_ys[1830]), .rectangle2_width(rectangle2_widths[1830]), .rectangle2_height(rectangle2_heights[1830]), .rectangle2_weight(rectangle2_weights[1830]), .rectangle3_x(rectangle3_xs[1830]), .rectangle3_y(rectangle3_ys[1830]), .rectangle3_width(rectangle3_widths[1830]), .rectangle3_height(rectangle3_heights[1830]), .rectangle3_weight(rectangle3_weights[1830]), .feature_threshold(feature_thresholds[1830]), .feature_above(feature_aboves[1830]), .feature_below(feature_belows[1830]), .scan_win_std_dev(scan_win_std_dev[1830]), .feature_accum(feature_accums[1830]));
  accum_calculator ac1831(.scan_win(scan_win1831), .rectangle1_x(rectangle1_xs[1831]), .rectangle1_y(rectangle1_ys[1831]), .rectangle1_width(rectangle1_widths[1831]), .rectangle1_height(rectangle1_heights[1831]), .rectangle1_weight(rectangle1_weights[1831]), .rectangle2_x(rectangle2_xs[1831]), .rectangle2_y(rectangle2_ys[1831]), .rectangle2_width(rectangle2_widths[1831]), .rectangle2_height(rectangle2_heights[1831]), .rectangle2_weight(rectangle2_weights[1831]), .rectangle3_x(rectangle3_xs[1831]), .rectangle3_y(rectangle3_ys[1831]), .rectangle3_width(rectangle3_widths[1831]), .rectangle3_height(rectangle3_heights[1831]), .rectangle3_weight(rectangle3_weights[1831]), .feature_threshold(feature_thresholds[1831]), .feature_above(feature_aboves[1831]), .feature_below(feature_belows[1831]), .scan_win_std_dev(scan_win_std_dev[1831]), .feature_accum(feature_accums[1831]));
  accum_calculator ac1832(.scan_win(scan_win1832), .rectangle1_x(rectangle1_xs[1832]), .rectangle1_y(rectangle1_ys[1832]), .rectangle1_width(rectangle1_widths[1832]), .rectangle1_height(rectangle1_heights[1832]), .rectangle1_weight(rectangle1_weights[1832]), .rectangle2_x(rectangle2_xs[1832]), .rectangle2_y(rectangle2_ys[1832]), .rectangle2_width(rectangle2_widths[1832]), .rectangle2_height(rectangle2_heights[1832]), .rectangle2_weight(rectangle2_weights[1832]), .rectangle3_x(rectangle3_xs[1832]), .rectangle3_y(rectangle3_ys[1832]), .rectangle3_width(rectangle3_widths[1832]), .rectangle3_height(rectangle3_heights[1832]), .rectangle3_weight(rectangle3_weights[1832]), .feature_threshold(feature_thresholds[1832]), .feature_above(feature_aboves[1832]), .feature_below(feature_belows[1832]), .scan_win_std_dev(scan_win_std_dev[1832]), .feature_accum(feature_accums[1832]));
  accum_calculator ac1833(.scan_win(scan_win1833), .rectangle1_x(rectangle1_xs[1833]), .rectangle1_y(rectangle1_ys[1833]), .rectangle1_width(rectangle1_widths[1833]), .rectangle1_height(rectangle1_heights[1833]), .rectangle1_weight(rectangle1_weights[1833]), .rectangle2_x(rectangle2_xs[1833]), .rectangle2_y(rectangle2_ys[1833]), .rectangle2_width(rectangle2_widths[1833]), .rectangle2_height(rectangle2_heights[1833]), .rectangle2_weight(rectangle2_weights[1833]), .rectangle3_x(rectangle3_xs[1833]), .rectangle3_y(rectangle3_ys[1833]), .rectangle3_width(rectangle3_widths[1833]), .rectangle3_height(rectangle3_heights[1833]), .rectangle3_weight(rectangle3_weights[1833]), .feature_threshold(feature_thresholds[1833]), .feature_above(feature_aboves[1833]), .feature_below(feature_belows[1833]), .scan_win_std_dev(scan_win_std_dev[1833]), .feature_accum(feature_accums[1833]));
  accum_calculator ac1834(.scan_win(scan_win1834), .rectangle1_x(rectangle1_xs[1834]), .rectangle1_y(rectangle1_ys[1834]), .rectangle1_width(rectangle1_widths[1834]), .rectangle1_height(rectangle1_heights[1834]), .rectangle1_weight(rectangle1_weights[1834]), .rectangle2_x(rectangle2_xs[1834]), .rectangle2_y(rectangle2_ys[1834]), .rectangle2_width(rectangle2_widths[1834]), .rectangle2_height(rectangle2_heights[1834]), .rectangle2_weight(rectangle2_weights[1834]), .rectangle3_x(rectangle3_xs[1834]), .rectangle3_y(rectangle3_ys[1834]), .rectangle3_width(rectangle3_widths[1834]), .rectangle3_height(rectangle3_heights[1834]), .rectangle3_weight(rectangle3_weights[1834]), .feature_threshold(feature_thresholds[1834]), .feature_above(feature_aboves[1834]), .feature_below(feature_belows[1834]), .scan_win_std_dev(scan_win_std_dev[1834]), .feature_accum(feature_accums[1834]));
  accum_calculator ac1835(.scan_win(scan_win1835), .rectangle1_x(rectangle1_xs[1835]), .rectangle1_y(rectangle1_ys[1835]), .rectangle1_width(rectangle1_widths[1835]), .rectangle1_height(rectangle1_heights[1835]), .rectangle1_weight(rectangle1_weights[1835]), .rectangle2_x(rectangle2_xs[1835]), .rectangle2_y(rectangle2_ys[1835]), .rectangle2_width(rectangle2_widths[1835]), .rectangle2_height(rectangle2_heights[1835]), .rectangle2_weight(rectangle2_weights[1835]), .rectangle3_x(rectangle3_xs[1835]), .rectangle3_y(rectangle3_ys[1835]), .rectangle3_width(rectangle3_widths[1835]), .rectangle3_height(rectangle3_heights[1835]), .rectangle3_weight(rectangle3_weights[1835]), .feature_threshold(feature_thresholds[1835]), .feature_above(feature_aboves[1835]), .feature_below(feature_belows[1835]), .scan_win_std_dev(scan_win_std_dev[1835]), .feature_accum(feature_accums[1835]));
  accum_calculator ac1836(.scan_win(scan_win1836), .rectangle1_x(rectangle1_xs[1836]), .rectangle1_y(rectangle1_ys[1836]), .rectangle1_width(rectangle1_widths[1836]), .rectangle1_height(rectangle1_heights[1836]), .rectangle1_weight(rectangle1_weights[1836]), .rectangle2_x(rectangle2_xs[1836]), .rectangle2_y(rectangle2_ys[1836]), .rectangle2_width(rectangle2_widths[1836]), .rectangle2_height(rectangle2_heights[1836]), .rectangle2_weight(rectangle2_weights[1836]), .rectangle3_x(rectangle3_xs[1836]), .rectangle3_y(rectangle3_ys[1836]), .rectangle3_width(rectangle3_widths[1836]), .rectangle3_height(rectangle3_heights[1836]), .rectangle3_weight(rectangle3_weights[1836]), .feature_threshold(feature_thresholds[1836]), .feature_above(feature_aboves[1836]), .feature_below(feature_belows[1836]), .scan_win_std_dev(scan_win_std_dev[1836]), .feature_accum(feature_accums[1836]));
  accum_calculator ac1837(.scan_win(scan_win1837), .rectangle1_x(rectangle1_xs[1837]), .rectangle1_y(rectangle1_ys[1837]), .rectangle1_width(rectangle1_widths[1837]), .rectangle1_height(rectangle1_heights[1837]), .rectangle1_weight(rectangle1_weights[1837]), .rectangle2_x(rectangle2_xs[1837]), .rectangle2_y(rectangle2_ys[1837]), .rectangle2_width(rectangle2_widths[1837]), .rectangle2_height(rectangle2_heights[1837]), .rectangle2_weight(rectangle2_weights[1837]), .rectangle3_x(rectangle3_xs[1837]), .rectangle3_y(rectangle3_ys[1837]), .rectangle3_width(rectangle3_widths[1837]), .rectangle3_height(rectangle3_heights[1837]), .rectangle3_weight(rectangle3_weights[1837]), .feature_threshold(feature_thresholds[1837]), .feature_above(feature_aboves[1837]), .feature_below(feature_belows[1837]), .scan_win_std_dev(scan_win_std_dev[1837]), .feature_accum(feature_accums[1837]));
  accum_calculator ac1838(.scan_win(scan_win1838), .rectangle1_x(rectangle1_xs[1838]), .rectangle1_y(rectangle1_ys[1838]), .rectangle1_width(rectangle1_widths[1838]), .rectangle1_height(rectangle1_heights[1838]), .rectangle1_weight(rectangle1_weights[1838]), .rectangle2_x(rectangle2_xs[1838]), .rectangle2_y(rectangle2_ys[1838]), .rectangle2_width(rectangle2_widths[1838]), .rectangle2_height(rectangle2_heights[1838]), .rectangle2_weight(rectangle2_weights[1838]), .rectangle3_x(rectangle3_xs[1838]), .rectangle3_y(rectangle3_ys[1838]), .rectangle3_width(rectangle3_widths[1838]), .rectangle3_height(rectangle3_heights[1838]), .rectangle3_weight(rectangle3_weights[1838]), .feature_threshold(feature_thresholds[1838]), .feature_above(feature_aboves[1838]), .feature_below(feature_belows[1838]), .scan_win_std_dev(scan_win_std_dev[1838]), .feature_accum(feature_accums[1838]));
  accum_calculator ac1839(.scan_win(scan_win1839), .rectangle1_x(rectangle1_xs[1839]), .rectangle1_y(rectangle1_ys[1839]), .rectangle1_width(rectangle1_widths[1839]), .rectangle1_height(rectangle1_heights[1839]), .rectangle1_weight(rectangle1_weights[1839]), .rectangle2_x(rectangle2_xs[1839]), .rectangle2_y(rectangle2_ys[1839]), .rectangle2_width(rectangle2_widths[1839]), .rectangle2_height(rectangle2_heights[1839]), .rectangle2_weight(rectangle2_weights[1839]), .rectangle3_x(rectangle3_xs[1839]), .rectangle3_y(rectangle3_ys[1839]), .rectangle3_width(rectangle3_widths[1839]), .rectangle3_height(rectangle3_heights[1839]), .rectangle3_weight(rectangle3_weights[1839]), .feature_threshold(feature_thresholds[1839]), .feature_above(feature_aboves[1839]), .feature_below(feature_belows[1839]), .scan_win_std_dev(scan_win_std_dev[1839]), .feature_accum(feature_accums[1839]));
  accum_calculator ac1840(.scan_win(scan_win1840), .rectangle1_x(rectangle1_xs[1840]), .rectangle1_y(rectangle1_ys[1840]), .rectangle1_width(rectangle1_widths[1840]), .rectangle1_height(rectangle1_heights[1840]), .rectangle1_weight(rectangle1_weights[1840]), .rectangle2_x(rectangle2_xs[1840]), .rectangle2_y(rectangle2_ys[1840]), .rectangle2_width(rectangle2_widths[1840]), .rectangle2_height(rectangle2_heights[1840]), .rectangle2_weight(rectangle2_weights[1840]), .rectangle3_x(rectangle3_xs[1840]), .rectangle3_y(rectangle3_ys[1840]), .rectangle3_width(rectangle3_widths[1840]), .rectangle3_height(rectangle3_heights[1840]), .rectangle3_weight(rectangle3_weights[1840]), .feature_threshold(feature_thresholds[1840]), .feature_above(feature_aboves[1840]), .feature_below(feature_belows[1840]), .scan_win_std_dev(scan_win_std_dev[1840]), .feature_accum(feature_accums[1840]));
  accum_calculator ac1841(.scan_win(scan_win1841), .rectangle1_x(rectangle1_xs[1841]), .rectangle1_y(rectangle1_ys[1841]), .rectangle1_width(rectangle1_widths[1841]), .rectangle1_height(rectangle1_heights[1841]), .rectangle1_weight(rectangle1_weights[1841]), .rectangle2_x(rectangle2_xs[1841]), .rectangle2_y(rectangle2_ys[1841]), .rectangle2_width(rectangle2_widths[1841]), .rectangle2_height(rectangle2_heights[1841]), .rectangle2_weight(rectangle2_weights[1841]), .rectangle3_x(rectangle3_xs[1841]), .rectangle3_y(rectangle3_ys[1841]), .rectangle3_width(rectangle3_widths[1841]), .rectangle3_height(rectangle3_heights[1841]), .rectangle3_weight(rectangle3_weights[1841]), .feature_threshold(feature_thresholds[1841]), .feature_above(feature_aboves[1841]), .feature_below(feature_belows[1841]), .scan_win_std_dev(scan_win_std_dev[1841]), .feature_accum(feature_accums[1841]));
  accum_calculator ac1842(.scan_win(scan_win1842), .rectangle1_x(rectangle1_xs[1842]), .rectangle1_y(rectangle1_ys[1842]), .rectangle1_width(rectangle1_widths[1842]), .rectangle1_height(rectangle1_heights[1842]), .rectangle1_weight(rectangle1_weights[1842]), .rectangle2_x(rectangle2_xs[1842]), .rectangle2_y(rectangle2_ys[1842]), .rectangle2_width(rectangle2_widths[1842]), .rectangle2_height(rectangle2_heights[1842]), .rectangle2_weight(rectangle2_weights[1842]), .rectangle3_x(rectangle3_xs[1842]), .rectangle3_y(rectangle3_ys[1842]), .rectangle3_width(rectangle3_widths[1842]), .rectangle3_height(rectangle3_heights[1842]), .rectangle3_weight(rectangle3_weights[1842]), .feature_threshold(feature_thresholds[1842]), .feature_above(feature_aboves[1842]), .feature_below(feature_belows[1842]), .scan_win_std_dev(scan_win_std_dev[1842]), .feature_accum(feature_accums[1842]));
  accum_calculator ac1843(.scan_win(scan_win1843), .rectangle1_x(rectangle1_xs[1843]), .rectangle1_y(rectangle1_ys[1843]), .rectangle1_width(rectangle1_widths[1843]), .rectangle1_height(rectangle1_heights[1843]), .rectangle1_weight(rectangle1_weights[1843]), .rectangle2_x(rectangle2_xs[1843]), .rectangle2_y(rectangle2_ys[1843]), .rectangle2_width(rectangle2_widths[1843]), .rectangle2_height(rectangle2_heights[1843]), .rectangle2_weight(rectangle2_weights[1843]), .rectangle3_x(rectangle3_xs[1843]), .rectangle3_y(rectangle3_ys[1843]), .rectangle3_width(rectangle3_widths[1843]), .rectangle3_height(rectangle3_heights[1843]), .rectangle3_weight(rectangle3_weights[1843]), .feature_threshold(feature_thresholds[1843]), .feature_above(feature_aboves[1843]), .feature_below(feature_belows[1843]), .scan_win_std_dev(scan_win_std_dev[1843]), .feature_accum(feature_accums[1843]));
  accum_calculator ac1844(.scan_win(scan_win1844), .rectangle1_x(rectangle1_xs[1844]), .rectangle1_y(rectangle1_ys[1844]), .rectangle1_width(rectangle1_widths[1844]), .rectangle1_height(rectangle1_heights[1844]), .rectangle1_weight(rectangle1_weights[1844]), .rectangle2_x(rectangle2_xs[1844]), .rectangle2_y(rectangle2_ys[1844]), .rectangle2_width(rectangle2_widths[1844]), .rectangle2_height(rectangle2_heights[1844]), .rectangle2_weight(rectangle2_weights[1844]), .rectangle3_x(rectangle3_xs[1844]), .rectangle3_y(rectangle3_ys[1844]), .rectangle3_width(rectangle3_widths[1844]), .rectangle3_height(rectangle3_heights[1844]), .rectangle3_weight(rectangle3_weights[1844]), .feature_threshold(feature_thresholds[1844]), .feature_above(feature_aboves[1844]), .feature_below(feature_belows[1844]), .scan_win_std_dev(scan_win_std_dev[1844]), .feature_accum(feature_accums[1844]));
  accum_calculator ac1845(.scan_win(scan_win1845), .rectangle1_x(rectangle1_xs[1845]), .rectangle1_y(rectangle1_ys[1845]), .rectangle1_width(rectangle1_widths[1845]), .rectangle1_height(rectangle1_heights[1845]), .rectangle1_weight(rectangle1_weights[1845]), .rectangle2_x(rectangle2_xs[1845]), .rectangle2_y(rectangle2_ys[1845]), .rectangle2_width(rectangle2_widths[1845]), .rectangle2_height(rectangle2_heights[1845]), .rectangle2_weight(rectangle2_weights[1845]), .rectangle3_x(rectangle3_xs[1845]), .rectangle3_y(rectangle3_ys[1845]), .rectangle3_width(rectangle3_widths[1845]), .rectangle3_height(rectangle3_heights[1845]), .rectangle3_weight(rectangle3_weights[1845]), .feature_threshold(feature_thresholds[1845]), .feature_above(feature_aboves[1845]), .feature_below(feature_belows[1845]), .scan_win_std_dev(scan_win_std_dev[1845]), .feature_accum(feature_accums[1845]));
  accum_calculator ac1846(.scan_win(scan_win1846), .rectangle1_x(rectangle1_xs[1846]), .rectangle1_y(rectangle1_ys[1846]), .rectangle1_width(rectangle1_widths[1846]), .rectangle1_height(rectangle1_heights[1846]), .rectangle1_weight(rectangle1_weights[1846]), .rectangle2_x(rectangle2_xs[1846]), .rectangle2_y(rectangle2_ys[1846]), .rectangle2_width(rectangle2_widths[1846]), .rectangle2_height(rectangle2_heights[1846]), .rectangle2_weight(rectangle2_weights[1846]), .rectangle3_x(rectangle3_xs[1846]), .rectangle3_y(rectangle3_ys[1846]), .rectangle3_width(rectangle3_widths[1846]), .rectangle3_height(rectangle3_heights[1846]), .rectangle3_weight(rectangle3_weights[1846]), .feature_threshold(feature_thresholds[1846]), .feature_above(feature_aboves[1846]), .feature_below(feature_belows[1846]), .scan_win_std_dev(scan_win_std_dev[1846]), .feature_accum(feature_accums[1846]));
  accum_calculator ac1847(.scan_win(scan_win1847), .rectangle1_x(rectangle1_xs[1847]), .rectangle1_y(rectangle1_ys[1847]), .rectangle1_width(rectangle1_widths[1847]), .rectangle1_height(rectangle1_heights[1847]), .rectangle1_weight(rectangle1_weights[1847]), .rectangle2_x(rectangle2_xs[1847]), .rectangle2_y(rectangle2_ys[1847]), .rectangle2_width(rectangle2_widths[1847]), .rectangle2_height(rectangle2_heights[1847]), .rectangle2_weight(rectangle2_weights[1847]), .rectangle3_x(rectangle3_xs[1847]), .rectangle3_y(rectangle3_ys[1847]), .rectangle3_width(rectangle3_widths[1847]), .rectangle3_height(rectangle3_heights[1847]), .rectangle3_weight(rectangle3_weights[1847]), .feature_threshold(feature_thresholds[1847]), .feature_above(feature_aboves[1847]), .feature_below(feature_belows[1847]), .scan_win_std_dev(scan_win_std_dev[1847]), .feature_accum(feature_accums[1847]));
  accum_calculator ac1848(.scan_win(scan_win1848), .rectangle1_x(rectangle1_xs[1848]), .rectangle1_y(rectangle1_ys[1848]), .rectangle1_width(rectangle1_widths[1848]), .rectangle1_height(rectangle1_heights[1848]), .rectangle1_weight(rectangle1_weights[1848]), .rectangle2_x(rectangle2_xs[1848]), .rectangle2_y(rectangle2_ys[1848]), .rectangle2_width(rectangle2_widths[1848]), .rectangle2_height(rectangle2_heights[1848]), .rectangle2_weight(rectangle2_weights[1848]), .rectangle3_x(rectangle3_xs[1848]), .rectangle3_y(rectangle3_ys[1848]), .rectangle3_width(rectangle3_widths[1848]), .rectangle3_height(rectangle3_heights[1848]), .rectangle3_weight(rectangle3_weights[1848]), .feature_threshold(feature_thresholds[1848]), .feature_above(feature_aboves[1848]), .feature_below(feature_belows[1848]), .scan_win_std_dev(scan_win_std_dev[1848]), .feature_accum(feature_accums[1848]));
  accum_calculator ac1849(.scan_win(scan_win1849), .rectangle1_x(rectangle1_xs[1849]), .rectangle1_y(rectangle1_ys[1849]), .rectangle1_width(rectangle1_widths[1849]), .rectangle1_height(rectangle1_heights[1849]), .rectangle1_weight(rectangle1_weights[1849]), .rectangle2_x(rectangle2_xs[1849]), .rectangle2_y(rectangle2_ys[1849]), .rectangle2_width(rectangle2_widths[1849]), .rectangle2_height(rectangle2_heights[1849]), .rectangle2_weight(rectangle2_weights[1849]), .rectangle3_x(rectangle3_xs[1849]), .rectangle3_y(rectangle3_ys[1849]), .rectangle3_width(rectangle3_widths[1849]), .rectangle3_height(rectangle3_heights[1849]), .rectangle3_weight(rectangle3_weights[1849]), .feature_threshold(feature_thresholds[1849]), .feature_above(feature_aboves[1849]), .feature_below(feature_belows[1849]), .scan_win_std_dev(scan_win_std_dev[1849]), .feature_accum(feature_accums[1849]));
  accum_calculator ac1850(.scan_win(scan_win1850), .rectangle1_x(rectangle1_xs[1850]), .rectangle1_y(rectangle1_ys[1850]), .rectangle1_width(rectangle1_widths[1850]), .rectangle1_height(rectangle1_heights[1850]), .rectangle1_weight(rectangle1_weights[1850]), .rectangle2_x(rectangle2_xs[1850]), .rectangle2_y(rectangle2_ys[1850]), .rectangle2_width(rectangle2_widths[1850]), .rectangle2_height(rectangle2_heights[1850]), .rectangle2_weight(rectangle2_weights[1850]), .rectangle3_x(rectangle3_xs[1850]), .rectangle3_y(rectangle3_ys[1850]), .rectangle3_width(rectangle3_widths[1850]), .rectangle3_height(rectangle3_heights[1850]), .rectangle3_weight(rectangle3_weights[1850]), .feature_threshold(feature_thresholds[1850]), .feature_above(feature_aboves[1850]), .feature_below(feature_belows[1850]), .scan_win_std_dev(scan_win_std_dev[1850]), .feature_accum(feature_accums[1850]));
  accum_calculator ac1851(.scan_win(scan_win1851), .rectangle1_x(rectangle1_xs[1851]), .rectangle1_y(rectangle1_ys[1851]), .rectangle1_width(rectangle1_widths[1851]), .rectangle1_height(rectangle1_heights[1851]), .rectangle1_weight(rectangle1_weights[1851]), .rectangle2_x(rectangle2_xs[1851]), .rectangle2_y(rectangle2_ys[1851]), .rectangle2_width(rectangle2_widths[1851]), .rectangle2_height(rectangle2_heights[1851]), .rectangle2_weight(rectangle2_weights[1851]), .rectangle3_x(rectangle3_xs[1851]), .rectangle3_y(rectangle3_ys[1851]), .rectangle3_width(rectangle3_widths[1851]), .rectangle3_height(rectangle3_heights[1851]), .rectangle3_weight(rectangle3_weights[1851]), .feature_threshold(feature_thresholds[1851]), .feature_above(feature_aboves[1851]), .feature_below(feature_belows[1851]), .scan_win_std_dev(scan_win_std_dev[1851]), .feature_accum(feature_accums[1851]));
  accum_calculator ac1852(.scan_win(scan_win1852), .rectangle1_x(rectangle1_xs[1852]), .rectangle1_y(rectangle1_ys[1852]), .rectangle1_width(rectangle1_widths[1852]), .rectangle1_height(rectangle1_heights[1852]), .rectangle1_weight(rectangle1_weights[1852]), .rectangle2_x(rectangle2_xs[1852]), .rectangle2_y(rectangle2_ys[1852]), .rectangle2_width(rectangle2_widths[1852]), .rectangle2_height(rectangle2_heights[1852]), .rectangle2_weight(rectangle2_weights[1852]), .rectangle3_x(rectangle3_xs[1852]), .rectangle3_y(rectangle3_ys[1852]), .rectangle3_width(rectangle3_widths[1852]), .rectangle3_height(rectangle3_heights[1852]), .rectangle3_weight(rectangle3_weights[1852]), .feature_threshold(feature_thresholds[1852]), .feature_above(feature_aboves[1852]), .feature_below(feature_belows[1852]), .scan_win_std_dev(scan_win_std_dev[1852]), .feature_accum(feature_accums[1852]));
  accum_calculator ac1853(.scan_win(scan_win1853), .rectangle1_x(rectangle1_xs[1853]), .rectangle1_y(rectangle1_ys[1853]), .rectangle1_width(rectangle1_widths[1853]), .rectangle1_height(rectangle1_heights[1853]), .rectangle1_weight(rectangle1_weights[1853]), .rectangle2_x(rectangle2_xs[1853]), .rectangle2_y(rectangle2_ys[1853]), .rectangle2_width(rectangle2_widths[1853]), .rectangle2_height(rectangle2_heights[1853]), .rectangle2_weight(rectangle2_weights[1853]), .rectangle3_x(rectangle3_xs[1853]), .rectangle3_y(rectangle3_ys[1853]), .rectangle3_width(rectangle3_widths[1853]), .rectangle3_height(rectangle3_heights[1853]), .rectangle3_weight(rectangle3_weights[1853]), .feature_threshold(feature_thresholds[1853]), .feature_above(feature_aboves[1853]), .feature_below(feature_belows[1853]), .scan_win_std_dev(scan_win_std_dev[1853]), .feature_accum(feature_accums[1853]));
  accum_calculator ac1854(.scan_win(scan_win1854), .rectangle1_x(rectangle1_xs[1854]), .rectangle1_y(rectangle1_ys[1854]), .rectangle1_width(rectangle1_widths[1854]), .rectangle1_height(rectangle1_heights[1854]), .rectangle1_weight(rectangle1_weights[1854]), .rectangle2_x(rectangle2_xs[1854]), .rectangle2_y(rectangle2_ys[1854]), .rectangle2_width(rectangle2_widths[1854]), .rectangle2_height(rectangle2_heights[1854]), .rectangle2_weight(rectangle2_weights[1854]), .rectangle3_x(rectangle3_xs[1854]), .rectangle3_y(rectangle3_ys[1854]), .rectangle3_width(rectangle3_widths[1854]), .rectangle3_height(rectangle3_heights[1854]), .rectangle3_weight(rectangle3_weights[1854]), .feature_threshold(feature_thresholds[1854]), .feature_above(feature_aboves[1854]), .feature_below(feature_belows[1854]), .scan_win_std_dev(scan_win_std_dev[1854]), .feature_accum(feature_accums[1854]));
  accum_calculator ac1855(.scan_win(scan_win1855), .rectangle1_x(rectangle1_xs[1855]), .rectangle1_y(rectangle1_ys[1855]), .rectangle1_width(rectangle1_widths[1855]), .rectangle1_height(rectangle1_heights[1855]), .rectangle1_weight(rectangle1_weights[1855]), .rectangle2_x(rectangle2_xs[1855]), .rectangle2_y(rectangle2_ys[1855]), .rectangle2_width(rectangle2_widths[1855]), .rectangle2_height(rectangle2_heights[1855]), .rectangle2_weight(rectangle2_weights[1855]), .rectangle3_x(rectangle3_xs[1855]), .rectangle3_y(rectangle3_ys[1855]), .rectangle3_width(rectangle3_widths[1855]), .rectangle3_height(rectangle3_heights[1855]), .rectangle3_weight(rectangle3_weights[1855]), .feature_threshold(feature_thresholds[1855]), .feature_above(feature_aboves[1855]), .feature_below(feature_belows[1855]), .scan_win_std_dev(scan_win_std_dev[1855]), .feature_accum(feature_accums[1855]));
  accum_calculator ac1856(.scan_win(scan_win1856), .rectangle1_x(rectangle1_xs[1856]), .rectangle1_y(rectangle1_ys[1856]), .rectangle1_width(rectangle1_widths[1856]), .rectangle1_height(rectangle1_heights[1856]), .rectangle1_weight(rectangle1_weights[1856]), .rectangle2_x(rectangle2_xs[1856]), .rectangle2_y(rectangle2_ys[1856]), .rectangle2_width(rectangle2_widths[1856]), .rectangle2_height(rectangle2_heights[1856]), .rectangle2_weight(rectangle2_weights[1856]), .rectangle3_x(rectangle3_xs[1856]), .rectangle3_y(rectangle3_ys[1856]), .rectangle3_width(rectangle3_widths[1856]), .rectangle3_height(rectangle3_heights[1856]), .rectangle3_weight(rectangle3_weights[1856]), .feature_threshold(feature_thresholds[1856]), .feature_above(feature_aboves[1856]), .feature_below(feature_belows[1856]), .scan_win_std_dev(scan_win_std_dev[1856]), .feature_accum(feature_accums[1856]));
  accum_calculator ac1857(.scan_win(scan_win1857), .rectangle1_x(rectangle1_xs[1857]), .rectangle1_y(rectangle1_ys[1857]), .rectangle1_width(rectangle1_widths[1857]), .rectangle1_height(rectangle1_heights[1857]), .rectangle1_weight(rectangle1_weights[1857]), .rectangle2_x(rectangle2_xs[1857]), .rectangle2_y(rectangle2_ys[1857]), .rectangle2_width(rectangle2_widths[1857]), .rectangle2_height(rectangle2_heights[1857]), .rectangle2_weight(rectangle2_weights[1857]), .rectangle3_x(rectangle3_xs[1857]), .rectangle3_y(rectangle3_ys[1857]), .rectangle3_width(rectangle3_widths[1857]), .rectangle3_height(rectangle3_heights[1857]), .rectangle3_weight(rectangle3_weights[1857]), .feature_threshold(feature_thresholds[1857]), .feature_above(feature_aboves[1857]), .feature_below(feature_belows[1857]), .scan_win_std_dev(scan_win_std_dev[1857]), .feature_accum(feature_accums[1857]));
  accum_calculator ac1858(.scan_win(scan_win1858), .rectangle1_x(rectangle1_xs[1858]), .rectangle1_y(rectangle1_ys[1858]), .rectangle1_width(rectangle1_widths[1858]), .rectangle1_height(rectangle1_heights[1858]), .rectangle1_weight(rectangle1_weights[1858]), .rectangle2_x(rectangle2_xs[1858]), .rectangle2_y(rectangle2_ys[1858]), .rectangle2_width(rectangle2_widths[1858]), .rectangle2_height(rectangle2_heights[1858]), .rectangle2_weight(rectangle2_weights[1858]), .rectangle3_x(rectangle3_xs[1858]), .rectangle3_y(rectangle3_ys[1858]), .rectangle3_width(rectangle3_widths[1858]), .rectangle3_height(rectangle3_heights[1858]), .rectangle3_weight(rectangle3_weights[1858]), .feature_threshold(feature_thresholds[1858]), .feature_above(feature_aboves[1858]), .feature_below(feature_belows[1858]), .scan_win_std_dev(scan_win_std_dev[1858]), .feature_accum(feature_accums[1858]));
  accum_calculator ac1859(.scan_win(scan_win1859), .rectangle1_x(rectangle1_xs[1859]), .rectangle1_y(rectangle1_ys[1859]), .rectangle1_width(rectangle1_widths[1859]), .rectangle1_height(rectangle1_heights[1859]), .rectangle1_weight(rectangle1_weights[1859]), .rectangle2_x(rectangle2_xs[1859]), .rectangle2_y(rectangle2_ys[1859]), .rectangle2_width(rectangle2_widths[1859]), .rectangle2_height(rectangle2_heights[1859]), .rectangle2_weight(rectangle2_weights[1859]), .rectangle3_x(rectangle3_xs[1859]), .rectangle3_y(rectangle3_ys[1859]), .rectangle3_width(rectangle3_widths[1859]), .rectangle3_height(rectangle3_heights[1859]), .rectangle3_weight(rectangle3_weights[1859]), .feature_threshold(feature_thresholds[1859]), .feature_above(feature_aboves[1859]), .feature_below(feature_belows[1859]), .scan_win_std_dev(scan_win_std_dev[1859]), .feature_accum(feature_accums[1859]));
  accum_calculator ac1860(.scan_win(scan_win1860), .rectangle1_x(rectangle1_xs[1860]), .rectangle1_y(rectangle1_ys[1860]), .rectangle1_width(rectangle1_widths[1860]), .rectangle1_height(rectangle1_heights[1860]), .rectangle1_weight(rectangle1_weights[1860]), .rectangle2_x(rectangle2_xs[1860]), .rectangle2_y(rectangle2_ys[1860]), .rectangle2_width(rectangle2_widths[1860]), .rectangle2_height(rectangle2_heights[1860]), .rectangle2_weight(rectangle2_weights[1860]), .rectangle3_x(rectangle3_xs[1860]), .rectangle3_y(rectangle3_ys[1860]), .rectangle3_width(rectangle3_widths[1860]), .rectangle3_height(rectangle3_heights[1860]), .rectangle3_weight(rectangle3_weights[1860]), .feature_threshold(feature_thresholds[1860]), .feature_above(feature_aboves[1860]), .feature_below(feature_belows[1860]), .scan_win_std_dev(scan_win_std_dev[1860]), .feature_accum(feature_accums[1860]));
  accum_calculator ac1861(.scan_win(scan_win1861), .rectangle1_x(rectangle1_xs[1861]), .rectangle1_y(rectangle1_ys[1861]), .rectangle1_width(rectangle1_widths[1861]), .rectangle1_height(rectangle1_heights[1861]), .rectangle1_weight(rectangle1_weights[1861]), .rectangle2_x(rectangle2_xs[1861]), .rectangle2_y(rectangle2_ys[1861]), .rectangle2_width(rectangle2_widths[1861]), .rectangle2_height(rectangle2_heights[1861]), .rectangle2_weight(rectangle2_weights[1861]), .rectangle3_x(rectangle3_xs[1861]), .rectangle3_y(rectangle3_ys[1861]), .rectangle3_width(rectangle3_widths[1861]), .rectangle3_height(rectangle3_heights[1861]), .rectangle3_weight(rectangle3_weights[1861]), .feature_threshold(feature_thresholds[1861]), .feature_above(feature_aboves[1861]), .feature_below(feature_belows[1861]), .scan_win_std_dev(scan_win_std_dev[1861]), .feature_accum(feature_accums[1861]));
  accum_calculator ac1862(.scan_win(scan_win1862), .rectangle1_x(rectangle1_xs[1862]), .rectangle1_y(rectangle1_ys[1862]), .rectangle1_width(rectangle1_widths[1862]), .rectangle1_height(rectangle1_heights[1862]), .rectangle1_weight(rectangle1_weights[1862]), .rectangle2_x(rectangle2_xs[1862]), .rectangle2_y(rectangle2_ys[1862]), .rectangle2_width(rectangle2_widths[1862]), .rectangle2_height(rectangle2_heights[1862]), .rectangle2_weight(rectangle2_weights[1862]), .rectangle3_x(rectangle3_xs[1862]), .rectangle3_y(rectangle3_ys[1862]), .rectangle3_width(rectangle3_widths[1862]), .rectangle3_height(rectangle3_heights[1862]), .rectangle3_weight(rectangle3_weights[1862]), .feature_threshold(feature_thresholds[1862]), .feature_above(feature_aboves[1862]), .feature_below(feature_belows[1862]), .scan_win_std_dev(scan_win_std_dev[1862]), .feature_accum(feature_accums[1862]));
  accum_calculator ac1863(.scan_win(scan_win1863), .rectangle1_x(rectangle1_xs[1863]), .rectangle1_y(rectangle1_ys[1863]), .rectangle1_width(rectangle1_widths[1863]), .rectangle1_height(rectangle1_heights[1863]), .rectangle1_weight(rectangle1_weights[1863]), .rectangle2_x(rectangle2_xs[1863]), .rectangle2_y(rectangle2_ys[1863]), .rectangle2_width(rectangle2_widths[1863]), .rectangle2_height(rectangle2_heights[1863]), .rectangle2_weight(rectangle2_weights[1863]), .rectangle3_x(rectangle3_xs[1863]), .rectangle3_y(rectangle3_ys[1863]), .rectangle3_width(rectangle3_widths[1863]), .rectangle3_height(rectangle3_heights[1863]), .rectangle3_weight(rectangle3_weights[1863]), .feature_threshold(feature_thresholds[1863]), .feature_above(feature_aboves[1863]), .feature_below(feature_belows[1863]), .scan_win_std_dev(scan_win_std_dev[1863]), .feature_accum(feature_accums[1863]));
  accum_calculator ac1864(.scan_win(scan_win1864), .rectangle1_x(rectangle1_xs[1864]), .rectangle1_y(rectangle1_ys[1864]), .rectangle1_width(rectangle1_widths[1864]), .rectangle1_height(rectangle1_heights[1864]), .rectangle1_weight(rectangle1_weights[1864]), .rectangle2_x(rectangle2_xs[1864]), .rectangle2_y(rectangle2_ys[1864]), .rectangle2_width(rectangle2_widths[1864]), .rectangle2_height(rectangle2_heights[1864]), .rectangle2_weight(rectangle2_weights[1864]), .rectangle3_x(rectangle3_xs[1864]), .rectangle3_y(rectangle3_ys[1864]), .rectangle3_width(rectangle3_widths[1864]), .rectangle3_height(rectangle3_heights[1864]), .rectangle3_weight(rectangle3_weights[1864]), .feature_threshold(feature_thresholds[1864]), .feature_above(feature_aboves[1864]), .feature_below(feature_belows[1864]), .scan_win_std_dev(scan_win_std_dev[1864]), .feature_accum(feature_accums[1864]));
  accum_calculator ac1865(.scan_win(scan_win1865), .rectangle1_x(rectangle1_xs[1865]), .rectangle1_y(rectangle1_ys[1865]), .rectangle1_width(rectangle1_widths[1865]), .rectangle1_height(rectangle1_heights[1865]), .rectangle1_weight(rectangle1_weights[1865]), .rectangle2_x(rectangle2_xs[1865]), .rectangle2_y(rectangle2_ys[1865]), .rectangle2_width(rectangle2_widths[1865]), .rectangle2_height(rectangle2_heights[1865]), .rectangle2_weight(rectangle2_weights[1865]), .rectangle3_x(rectangle3_xs[1865]), .rectangle3_y(rectangle3_ys[1865]), .rectangle3_width(rectangle3_widths[1865]), .rectangle3_height(rectangle3_heights[1865]), .rectangle3_weight(rectangle3_weights[1865]), .feature_threshold(feature_thresholds[1865]), .feature_above(feature_aboves[1865]), .feature_below(feature_belows[1865]), .scan_win_std_dev(scan_win_std_dev[1865]), .feature_accum(feature_accums[1865]));
  accum_calculator ac1866(.scan_win(scan_win1866), .rectangle1_x(rectangle1_xs[1866]), .rectangle1_y(rectangle1_ys[1866]), .rectangle1_width(rectangle1_widths[1866]), .rectangle1_height(rectangle1_heights[1866]), .rectangle1_weight(rectangle1_weights[1866]), .rectangle2_x(rectangle2_xs[1866]), .rectangle2_y(rectangle2_ys[1866]), .rectangle2_width(rectangle2_widths[1866]), .rectangle2_height(rectangle2_heights[1866]), .rectangle2_weight(rectangle2_weights[1866]), .rectangle3_x(rectangle3_xs[1866]), .rectangle3_y(rectangle3_ys[1866]), .rectangle3_width(rectangle3_widths[1866]), .rectangle3_height(rectangle3_heights[1866]), .rectangle3_weight(rectangle3_weights[1866]), .feature_threshold(feature_thresholds[1866]), .feature_above(feature_aboves[1866]), .feature_below(feature_belows[1866]), .scan_win_std_dev(scan_win_std_dev[1866]), .feature_accum(feature_accums[1866]));
  accum_calculator ac1867(.scan_win(scan_win1867), .rectangle1_x(rectangle1_xs[1867]), .rectangle1_y(rectangle1_ys[1867]), .rectangle1_width(rectangle1_widths[1867]), .rectangle1_height(rectangle1_heights[1867]), .rectangle1_weight(rectangle1_weights[1867]), .rectangle2_x(rectangle2_xs[1867]), .rectangle2_y(rectangle2_ys[1867]), .rectangle2_width(rectangle2_widths[1867]), .rectangle2_height(rectangle2_heights[1867]), .rectangle2_weight(rectangle2_weights[1867]), .rectangle3_x(rectangle3_xs[1867]), .rectangle3_y(rectangle3_ys[1867]), .rectangle3_width(rectangle3_widths[1867]), .rectangle3_height(rectangle3_heights[1867]), .rectangle3_weight(rectangle3_weights[1867]), .feature_threshold(feature_thresholds[1867]), .feature_above(feature_aboves[1867]), .feature_below(feature_belows[1867]), .scan_win_std_dev(scan_win_std_dev[1867]), .feature_accum(feature_accums[1867]));
  accum_calculator ac1868(.scan_win(scan_win1868), .rectangle1_x(rectangle1_xs[1868]), .rectangle1_y(rectangle1_ys[1868]), .rectangle1_width(rectangle1_widths[1868]), .rectangle1_height(rectangle1_heights[1868]), .rectangle1_weight(rectangle1_weights[1868]), .rectangle2_x(rectangle2_xs[1868]), .rectangle2_y(rectangle2_ys[1868]), .rectangle2_width(rectangle2_widths[1868]), .rectangle2_height(rectangle2_heights[1868]), .rectangle2_weight(rectangle2_weights[1868]), .rectangle3_x(rectangle3_xs[1868]), .rectangle3_y(rectangle3_ys[1868]), .rectangle3_width(rectangle3_widths[1868]), .rectangle3_height(rectangle3_heights[1868]), .rectangle3_weight(rectangle3_weights[1868]), .feature_threshold(feature_thresholds[1868]), .feature_above(feature_aboves[1868]), .feature_below(feature_belows[1868]), .scan_win_std_dev(scan_win_std_dev[1868]), .feature_accum(feature_accums[1868]));
  accum_calculator ac1869(.scan_win(scan_win1869), .rectangle1_x(rectangle1_xs[1869]), .rectangle1_y(rectangle1_ys[1869]), .rectangle1_width(rectangle1_widths[1869]), .rectangle1_height(rectangle1_heights[1869]), .rectangle1_weight(rectangle1_weights[1869]), .rectangle2_x(rectangle2_xs[1869]), .rectangle2_y(rectangle2_ys[1869]), .rectangle2_width(rectangle2_widths[1869]), .rectangle2_height(rectangle2_heights[1869]), .rectangle2_weight(rectangle2_weights[1869]), .rectangle3_x(rectangle3_xs[1869]), .rectangle3_y(rectangle3_ys[1869]), .rectangle3_width(rectangle3_widths[1869]), .rectangle3_height(rectangle3_heights[1869]), .rectangle3_weight(rectangle3_weights[1869]), .feature_threshold(feature_thresholds[1869]), .feature_above(feature_aboves[1869]), .feature_below(feature_belows[1869]), .scan_win_std_dev(scan_win_std_dev[1869]), .feature_accum(feature_accums[1869]));
  accum_calculator ac1870(.scan_win(scan_win1870), .rectangle1_x(rectangle1_xs[1870]), .rectangle1_y(rectangle1_ys[1870]), .rectangle1_width(rectangle1_widths[1870]), .rectangle1_height(rectangle1_heights[1870]), .rectangle1_weight(rectangle1_weights[1870]), .rectangle2_x(rectangle2_xs[1870]), .rectangle2_y(rectangle2_ys[1870]), .rectangle2_width(rectangle2_widths[1870]), .rectangle2_height(rectangle2_heights[1870]), .rectangle2_weight(rectangle2_weights[1870]), .rectangle3_x(rectangle3_xs[1870]), .rectangle3_y(rectangle3_ys[1870]), .rectangle3_width(rectangle3_widths[1870]), .rectangle3_height(rectangle3_heights[1870]), .rectangle3_weight(rectangle3_weights[1870]), .feature_threshold(feature_thresholds[1870]), .feature_above(feature_aboves[1870]), .feature_below(feature_belows[1870]), .scan_win_std_dev(scan_win_std_dev[1870]), .feature_accum(feature_accums[1870]));
  accum_calculator ac1871(.scan_win(scan_win1871), .rectangle1_x(rectangle1_xs[1871]), .rectangle1_y(rectangle1_ys[1871]), .rectangle1_width(rectangle1_widths[1871]), .rectangle1_height(rectangle1_heights[1871]), .rectangle1_weight(rectangle1_weights[1871]), .rectangle2_x(rectangle2_xs[1871]), .rectangle2_y(rectangle2_ys[1871]), .rectangle2_width(rectangle2_widths[1871]), .rectangle2_height(rectangle2_heights[1871]), .rectangle2_weight(rectangle2_weights[1871]), .rectangle3_x(rectangle3_xs[1871]), .rectangle3_y(rectangle3_ys[1871]), .rectangle3_width(rectangle3_widths[1871]), .rectangle3_height(rectangle3_heights[1871]), .rectangle3_weight(rectangle3_weights[1871]), .feature_threshold(feature_thresholds[1871]), .feature_above(feature_aboves[1871]), .feature_below(feature_belows[1871]), .scan_win_std_dev(scan_win_std_dev[1871]), .feature_accum(feature_accums[1871]));
  accum_calculator ac1872(.scan_win(scan_win1872), .rectangle1_x(rectangle1_xs[1872]), .rectangle1_y(rectangle1_ys[1872]), .rectangle1_width(rectangle1_widths[1872]), .rectangle1_height(rectangle1_heights[1872]), .rectangle1_weight(rectangle1_weights[1872]), .rectangle2_x(rectangle2_xs[1872]), .rectangle2_y(rectangle2_ys[1872]), .rectangle2_width(rectangle2_widths[1872]), .rectangle2_height(rectangle2_heights[1872]), .rectangle2_weight(rectangle2_weights[1872]), .rectangle3_x(rectangle3_xs[1872]), .rectangle3_y(rectangle3_ys[1872]), .rectangle3_width(rectangle3_widths[1872]), .rectangle3_height(rectangle3_heights[1872]), .rectangle3_weight(rectangle3_weights[1872]), .feature_threshold(feature_thresholds[1872]), .feature_above(feature_aboves[1872]), .feature_below(feature_belows[1872]), .scan_win_std_dev(scan_win_std_dev[1872]), .feature_accum(feature_accums[1872]));
  accum_calculator ac1873(.scan_win(scan_win1873), .rectangle1_x(rectangle1_xs[1873]), .rectangle1_y(rectangle1_ys[1873]), .rectangle1_width(rectangle1_widths[1873]), .rectangle1_height(rectangle1_heights[1873]), .rectangle1_weight(rectangle1_weights[1873]), .rectangle2_x(rectangle2_xs[1873]), .rectangle2_y(rectangle2_ys[1873]), .rectangle2_width(rectangle2_widths[1873]), .rectangle2_height(rectangle2_heights[1873]), .rectangle2_weight(rectangle2_weights[1873]), .rectangle3_x(rectangle3_xs[1873]), .rectangle3_y(rectangle3_ys[1873]), .rectangle3_width(rectangle3_widths[1873]), .rectangle3_height(rectangle3_heights[1873]), .rectangle3_weight(rectangle3_weights[1873]), .feature_threshold(feature_thresholds[1873]), .feature_above(feature_aboves[1873]), .feature_below(feature_belows[1873]), .scan_win_std_dev(scan_win_std_dev[1873]), .feature_accum(feature_accums[1873]));
  accum_calculator ac1874(.scan_win(scan_win1874), .rectangle1_x(rectangle1_xs[1874]), .rectangle1_y(rectangle1_ys[1874]), .rectangle1_width(rectangle1_widths[1874]), .rectangle1_height(rectangle1_heights[1874]), .rectangle1_weight(rectangle1_weights[1874]), .rectangle2_x(rectangle2_xs[1874]), .rectangle2_y(rectangle2_ys[1874]), .rectangle2_width(rectangle2_widths[1874]), .rectangle2_height(rectangle2_heights[1874]), .rectangle2_weight(rectangle2_weights[1874]), .rectangle3_x(rectangle3_xs[1874]), .rectangle3_y(rectangle3_ys[1874]), .rectangle3_width(rectangle3_widths[1874]), .rectangle3_height(rectangle3_heights[1874]), .rectangle3_weight(rectangle3_weights[1874]), .feature_threshold(feature_thresholds[1874]), .feature_above(feature_aboves[1874]), .feature_below(feature_belows[1874]), .scan_win_std_dev(scan_win_std_dev[1874]), .feature_accum(feature_accums[1874]));
  accum_calculator ac1875(.scan_win(scan_win1875), .rectangle1_x(rectangle1_xs[1875]), .rectangle1_y(rectangle1_ys[1875]), .rectangle1_width(rectangle1_widths[1875]), .rectangle1_height(rectangle1_heights[1875]), .rectangle1_weight(rectangle1_weights[1875]), .rectangle2_x(rectangle2_xs[1875]), .rectangle2_y(rectangle2_ys[1875]), .rectangle2_width(rectangle2_widths[1875]), .rectangle2_height(rectangle2_heights[1875]), .rectangle2_weight(rectangle2_weights[1875]), .rectangle3_x(rectangle3_xs[1875]), .rectangle3_y(rectangle3_ys[1875]), .rectangle3_width(rectangle3_widths[1875]), .rectangle3_height(rectangle3_heights[1875]), .rectangle3_weight(rectangle3_weights[1875]), .feature_threshold(feature_thresholds[1875]), .feature_above(feature_aboves[1875]), .feature_below(feature_belows[1875]), .scan_win_std_dev(scan_win_std_dev[1875]), .feature_accum(feature_accums[1875]));
  accum_calculator ac1876(.scan_win(scan_win1876), .rectangle1_x(rectangle1_xs[1876]), .rectangle1_y(rectangle1_ys[1876]), .rectangle1_width(rectangle1_widths[1876]), .rectangle1_height(rectangle1_heights[1876]), .rectangle1_weight(rectangle1_weights[1876]), .rectangle2_x(rectangle2_xs[1876]), .rectangle2_y(rectangle2_ys[1876]), .rectangle2_width(rectangle2_widths[1876]), .rectangle2_height(rectangle2_heights[1876]), .rectangle2_weight(rectangle2_weights[1876]), .rectangle3_x(rectangle3_xs[1876]), .rectangle3_y(rectangle3_ys[1876]), .rectangle3_width(rectangle3_widths[1876]), .rectangle3_height(rectangle3_heights[1876]), .rectangle3_weight(rectangle3_weights[1876]), .feature_threshold(feature_thresholds[1876]), .feature_above(feature_aboves[1876]), .feature_below(feature_belows[1876]), .scan_win_std_dev(scan_win_std_dev[1876]), .feature_accum(feature_accums[1876]));
  accum_calculator ac1877(.scan_win(scan_win1877), .rectangle1_x(rectangle1_xs[1877]), .rectangle1_y(rectangle1_ys[1877]), .rectangle1_width(rectangle1_widths[1877]), .rectangle1_height(rectangle1_heights[1877]), .rectangle1_weight(rectangle1_weights[1877]), .rectangle2_x(rectangle2_xs[1877]), .rectangle2_y(rectangle2_ys[1877]), .rectangle2_width(rectangle2_widths[1877]), .rectangle2_height(rectangle2_heights[1877]), .rectangle2_weight(rectangle2_weights[1877]), .rectangle3_x(rectangle3_xs[1877]), .rectangle3_y(rectangle3_ys[1877]), .rectangle3_width(rectangle3_widths[1877]), .rectangle3_height(rectangle3_heights[1877]), .rectangle3_weight(rectangle3_weights[1877]), .feature_threshold(feature_thresholds[1877]), .feature_above(feature_aboves[1877]), .feature_below(feature_belows[1877]), .scan_win_std_dev(scan_win_std_dev[1877]), .feature_accum(feature_accums[1877]));
  accum_calculator ac1878(.scan_win(scan_win1878), .rectangle1_x(rectangle1_xs[1878]), .rectangle1_y(rectangle1_ys[1878]), .rectangle1_width(rectangle1_widths[1878]), .rectangle1_height(rectangle1_heights[1878]), .rectangle1_weight(rectangle1_weights[1878]), .rectangle2_x(rectangle2_xs[1878]), .rectangle2_y(rectangle2_ys[1878]), .rectangle2_width(rectangle2_widths[1878]), .rectangle2_height(rectangle2_heights[1878]), .rectangle2_weight(rectangle2_weights[1878]), .rectangle3_x(rectangle3_xs[1878]), .rectangle3_y(rectangle3_ys[1878]), .rectangle3_width(rectangle3_widths[1878]), .rectangle3_height(rectangle3_heights[1878]), .rectangle3_weight(rectangle3_weights[1878]), .feature_threshold(feature_thresholds[1878]), .feature_above(feature_aboves[1878]), .feature_below(feature_belows[1878]), .scan_win_std_dev(scan_win_std_dev[1878]), .feature_accum(feature_accums[1878]));
  accum_calculator ac1879(.scan_win(scan_win1879), .rectangle1_x(rectangle1_xs[1879]), .rectangle1_y(rectangle1_ys[1879]), .rectangle1_width(rectangle1_widths[1879]), .rectangle1_height(rectangle1_heights[1879]), .rectangle1_weight(rectangle1_weights[1879]), .rectangle2_x(rectangle2_xs[1879]), .rectangle2_y(rectangle2_ys[1879]), .rectangle2_width(rectangle2_widths[1879]), .rectangle2_height(rectangle2_heights[1879]), .rectangle2_weight(rectangle2_weights[1879]), .rectangle3_x(rectangle3_xs[1879]), .rectangle3_y(rectangle3_ys[1879]), .rectangle3_width(rectangle3_widths[1879]), .rectangle3_height(rectangle3_heights[1879]), .rectangle3_weight(rectangle3_weights[1879]), .feature_threshold(feature_thresholds[1879]), .feature_above(feature_aboves[1879]), .feature_below(feature_belows[1879]), .scan_win_std_dev(scan_win_std_dev[1879]), .feature_accum(feature_accums[1879]));
  accum_calculator ac1880(.scan_win(scan_win1880), .rectangle1_x(rectangle1_xs[1880]), .rectangle1_y(rectangle1_ys[1880]), .rectangle1_width(rectangle1_widths[1880]), .rectangle1_height(rectangle1_heights[1880]), .rectangle1_weight(rectangle1_weights[1880]), .rectangle2_x(rectangle2_xs[1880]), .rectangle2_y(rectangle2_ys[1880]), .rectangle2_width(rectangle2_widths[1880]), .rectangle2_height(rectangle2_heights[1880]), .rectangle2_weight(rectangle2_weights[1880]), .rectangle3_x(rectangle3_xs[1880]), .rectangle3_y(rectangle3_ys[1880]), .rectangle3_width(rectangle3_widths[1880]), .rectangle3_height(rectangle3_heights[1880]), .rectangle3_weight(rectangle3_weights[1880]), .feature_threshold(feature_thresholds[1880]), .feature_above(feature_aboves[1880]), .feature_below(feature_belows[1880]), .scan_win_std_dev(scan_win_std_dev[1880]), .feature_accum(feature_accums[1880]));
  accum_calculator ac1881(.scan_win(scan_win1881), .rectangle1_x(rectangle1_xs[1881]), .rectangle1_y(rectangle1_ys[1881]), .rectangle1_width(rectangle1_widths[1881]), .rectangle1_height(rectangle1_heights[1881]), .rectangle1_weight(rectangle1_weights[1881]), .rectangle2_x(rectangle2_xs[1881]), .rectangle2_y(rectangle2_ys[1881]), .rectangle2_width(rectangle2_widths[1881]), .rectangle2_height(rectangle2_heights[1881]), .rectangle2_weight(rectangle2_weights[1881]), .rectangle3_x(rectangle3_xs[1881]), .rectangle3_y(rectangle3_ys[1881]), .rectangle3_width(rectangle3_widths[1881]), .rectangle3_height(rectangle3_heights[1881]), .rectangle3_weight(rectangle3_weights[1881]), .feature_threshold(feature_thresholds[1881]), .feature_above(feature_aboves[1881]), .feature_below(feature_belows[1881]), .scan_win_std_dev(scan_win_std_dev[1881]), .feature_accum(feature_accums[1881]));
  accum_calculator ac1882(.scan_win(scan_win1882), .rectangle1_x(rectangle1_xs[1882]), .rectangle1_y(rectangle1_ys[1882]), .rectangle1_width(rectangle1_widths[1882]), .rectangle1_height(rectangle1_heights[1882]), .rectangle1_weight(rectangle1_weights[1882]), .rectangle2_x(rectangle2_xs[1882]), .rectangle2_y(rectangle2_ys[1882]), .rectangle2_width(rectangle2_widths[1882]), .rectangle2_height(rectangle2_heights[1882]), .rectangle2_weight(rectangle2_weights[1882]), .rectangle3_x(rectangle3_xs[1882]), .rectangle3_y(rectangle3_ys[1882]), .rectangle3_width(rectangle3_widths[1882]), .rectangle3_height(rectangle3_heights[1882]), .rectangle3_weight(rectangle3_weights[1882]), .feature_threshold(feature_thresholds[1882]), .feature_above(feature_aboves[1882]), .feature_below(feature_belows[1882]), .scan_win_std_dev(scan_win_std_dev[1882]), .feature_accum(feature_accums[1882]));
  accum_calculator ac1883(.scan_win(scan_win1883), .rectangle1_x(rectangle1_xs[1883]), .rectangle1_y(rectangle1_ys[1883]), .rectangle1_width(rectangle1_widths[1883]), .rectangle1_height(rectangle1_heights[1883]), .rectangle1_weight(rectangle1_weights[1883]), .rectangle2_x(rectangle2_xs[1883]), .rectangle2_y(rectangle2_ys[1883]), .rectangle2_width(rectangle2_widths[1883]), .rectangle2_height(rectangle2_heights[1883]), .rectangle2_weight(rectangle2_weights[1883]), .rectangle3_x(rectangle3_xs[1883]), .rectangle3_y(rectangle3_ys[1883]), .rectangle3_width(rectangle3_widths[1883]), .rectangle3_height(rectangle3_heights[1883]), .rectangle3_weight(rectangle3_weights[1883]), .feature_threshold(feature_thresholds[1883]), .feature_above(feature_aboves[1883]), .feature_below(feature_belows[1883]), .scan_win_std_dev(scan_win_std_dev[1883]), .feature_accum(feature_accums[1883]));
  accum_calculator ac1884(.scan_win(scan_win1884), .rectangle1_x(rectangle1_xs[1884]), .rectangle1_y(rectangle1_ys[1884]), .rectangle1_width(rectangle1_widths[1884]), .rectangle1_height(rectangle1_heights[1884]), .rectangle1_weight(rectangle1_weights[1884]), .rectangle2_x(rectangle2_xs[1884]), .rectangle2_y(rectangle2_ys[1884]), .rectangle2_width(rectangle2_widths[1884]), .rectangle2_height(rectangle2_heights[1884]), .rectangle2_weight(rectangle2_weights[1884]), .rectangle3_x(rectangle3_xs[1884]), .rectangle3_y(rectangle3_ys[1884]), .rectangle3_width(rectangle3_widths[1884]), .rectangle3_height(rectangle3_heights[1884]), .rectangle3_weight(rectangle3_weights[1884]), .feature_threshold(feature_thresholds[1884]), .feature_above(feature_aboves[1884]), .feature_below(feature_belows[1884]), .scan_win_std_dev(scan_win_std_dev[1884]), .feature_accum(feature_accums[1884]));
  accum_calculator ac1885(.scan_win(scan_win1885), .rectangle1_x(rectangle1_xs[1885]), .rectangle1_y(rectangle1_ys[1885]), .rectangle1_width(rectangle1_widths[1885]), .rectangle1_height(rectangle1_heights[1885]), .rectangle1_weight(rectangle1_weights[1885]), .rectangle2_x(rectangle2_xs[1885]), .rectangle2_y(rectangle2_ys[1885]), .rectangle2_width(rectangle2_widths[1885]), .rectangle2_height(rectangle2_heights[1885]), .rectangle2_weight(rectangle2_weights[1885]), .rectangle3_x(rectangle3_xs[1885]), .rectangle3_y(rectangle3_ys[1885]), .rectangle3_width(rectangle3_widths[1885]), .rectangle3_height(rectangle3_heights[1885]), .rectangle3_weight(rectangle3_weights[1885]), .feature_threshold(feature_thresholds[1885]), .feature_above(feature_aboves[1885]), .feature_below(feature_belows[1885]), .scan_win_std_dev(scan_win_std_dev[1885]), .feature_accum(feature_accums[1885]));
  accum_calculator ac1886(.scan_win(scan_win1886), .rectangle1_x(rectangle1_xs[1886]), .rectangle1_y(rectangle1_ys[1886]), .rectangle1_width(rectangle1_widths[1886]), .rectangle1_height(rectangle1_heights[1886]), .rectangle1_weight(rectangle1_weights[1886]), .rectangle2_x(rectangle2_xs[1886]), .rectangle2_y(rectangle2_ys[1886]), .rectangle2_width(rectangle2_widths[1886]), .rectangle2_height(rectangle2_heights[1886]), .rectangle2_weight(rectangle2_weights[1886]), .rectangle3_x(rectangle3_xs[1886]), .rectangle3_y(rectangle3_ys[1886]), .rectangle3_width(rectangle3_widths[1886]), .rectangle3_height(rectangle3_heights[1886]), .rectangle3_weight(rectangle3_weights[1886]), .feature_threshold(feature_thresholds[1886]), .feature_above(feature_aboves[1886]), .feature_below(feature_belows[1886]), .scan_win_std_dev(scan_win_std_dev[1886]), .feature_accum(feature_accums[1886]));
  accum_calculator ac1887(.scan_win(scan_win1887), .rectangle1_x(rectangle1_xs[1887]), .rectangle1_y(rectangle1_ys[1887]), .rectangle1_width(rectangle1_widths[1887]), .rectangle1_height(rectangle1_heights[1887]), .rectangle1_weight(rectangle1_weights[1887]), .rectangle2_x(rectangle2_xs[1887]), .rectangle2_y(rectangle2_ys[1887]), .rectangle2_width(rectangle2_widths[1887]), .rectangle2_height(rectangle2_heights[1887]), .rectangle2_weight(rectangle2_weights[1887]), .rectangle3_x(rectangle3_xs[1887]), .rectangle3_y(rectangle3_ys[1887]), .rectangle3_width(rectangle3_widths[1887]), .rectangle3_height(rectangle3_heights[1887]), .rectangle3_weight(rectangle3_weights[1887]), .feature_threshold(feature_thresholds[1887]), .feature_above(feature_aboves[1887]), .feature_below(feature_belows[1887]), .scan_win_std_dev(scan_win_std_dev[1887]), .feature_accum(feature_accums[1887]));
  accum_calculator ac1888(.scan_win(scan_win1888), .rectangle1_x(rectangle1_xs[1888]), .rectangle1_y(rectangle1_ys[1888]), .rectangle1_width(rectangle1_widths[1888]), .rectangle1_height(rectangle1_heights[1888]), .rectangle1_weight(rectangle1_weights[1888]), .rectangle2_x(rectangle2_xs[1888]), .rectangle2_y(rectangle2_ys[1888]), .rectangle2_width(rectangle2_widths[1888]), .rectangle2_height(rectangle2_heights[1888]), .rectangle2_weight(rectangle2_weights[1888]), .rectangle3_x(rectangle3_xs[1888]), .rectangle3_y(rectangle3_ys[1888]), .rectangle3_width(rectangle3_widths[1888]), .rectangle3_height(rectangle3_heights[1888]), .rectangle3_weight(rectangle3_weights[1888]), .feature_threshold(feature_thresholds[1888]), .feature_above(feature_aboves[1888]), .feature_below(feature_belows[1888]), .scan_win_std_dev(scan_win_std_dev[1888]), .feature_accum(feature_accums[1888]));
  accum_calculator ac1889(.scan_win(scan_win1889), .rectangle1_x(rectangle1_xs[1889]), .rectangle1_y(rectangle1_ys[1889]), .rectangle1_width(rectangle1_widths[1889]), .rectangle1_height(rectangle1_heights[1889]), .rectangle1_weight(rectangle1_weights[1889]), .rectangle2_x(rectangle2_xs[1889]), .rectangle2_y(rectangle2_ys[1889]), .rectangle2_width(rectangle2_widths[1889]), .rectangle2_height(rectangle2_heights[1889]), .rectangle2_weight(rectangle2_weights[1889]), .rectangle3_x(rectangle3_xs[1889]), .rectangle3_y(rectangle3_ys[1889]), .rectangle3_width(rectangle3_widths[1889]), .rectangle3_height(rectangle3_heights[1889]), .rectangle3_weight(rectangle3_weights[1889]), .feature_threshold(feature_thresholds[1889]), .feature_above(feature_aboves[1889]), .feature_below(feature_belows[1889]), .scan_win_std_dev(scan_win_std_dev[1889]), .feature_accum(feature_accums[1889]));
  accum_calculator ac1890(.scan_win(scan_win1890), .rectangle1_x(rectangle1_xs[1890]), .rectangle1_y(rectangle1_ys[1890]), .rectangle1_width(rectangle1_widths[1890]), .rectangle1_height(rectangle1_heights[1890]), .rectangle1_weight(rectangle1_weights[1890]), .rectangle2_x(rectangle2_xs[1890]), .rectangle2_y(rectangle2_ys[1890]), .rectangle2_width(rectangle2_widths[1890]), .rectangle2_height(rectangle2_heights[1890]), .rectangle2_weight(rectangle2_weights[1890]), .rectangle3_x(rectangle3_xs[1890]), .rectangle3_y(rectangle3_ys[1890]), .rectangle3_width(rectangle3_widths[1890]), .rectangle3_height(rectangle3_heights[1890]), .rectangle3_weight(rectangle3_weights[1890]), .feature_threshold(feature_thresholds[1890]), .feature_above(feature_aboves[1890]), .feature_below(feature_belows[1890]), .scan_win_std_dev(scan_win_std_dev[1890]), .feature_accum(feature_accums[1890]));
  accum_calculator ac1891(.scan_win(scan_win1891), .rectangle1_x(rectangle1_xs[1891]), .rectangle1_y(rectangle1_ys[1891]), .rectangle1_width(rectangle1_widths[1891]), .rectangle1_height(rectangle1_heights[1891]), .rectangle1_weight(rectangle1_weights[1891]), .rectangle2_x(rectangle2_xs[1891]), .rectangle2_y(rectangle2_ys[1891]), .rectangle2_width(rectangle2_widths[1891]), .rectangle2_height(rectangle2_heights[1891]), .rectangle2_weight(rectangle2_weights[1891]), .rectangle3_x(rectangle3_xs[1891]), .rectangle3_y(rectangle3_ys[1891]), .rectangle3_width(rectangle3_widths[1891]), .rectangle3_height(rectangle3_heights[1891]), .rectangle3_weight(rectangle3_weights[1891]), .feature_threshold(feature_thresholds[1891]), .feature_above(feature_aboves[1891]), .feature_below(feature_belows[1891]), .scan_win_std_dev(scan_win_std_dev[1891]), .feature_accum(feature_accums[1891]));
  accum_calculator ac1892(.scan_win(scan_win1892), .rectangle1_x(rectangle1_xs[1892]), .rectangle1_y(rectangle1_ys[1892]), .rectangle1_width(rectangle1_widths[1892]), .rectangle1_height(rectangle1_heights[1892]), .rectangle1_weight(rectangle1_weights[1892]), .rectangle2_x(rectangle2_xs[1892]), .rectangle2_y(rectangle2_ys[1892]), .rectangle2_width(rectangle2_widths[1892]), .rectangle2_height(rectangle2_heights[1892]), .rectangle2_weight(rectangle2_weights[1892]), .rectangle3_x(rectangle3_xs[1892]), .rectangle3_y(rectangle3_ys[1892]), .rectangle3_width(rectangle3_widths[1892]), .rectangle3_height(rectangle3_heights[1892]), .rectangle3_weight(rectangle3_weights[1892]), .feature_threshold(feature_thresholds[1892]), .feature_above(feature_aboves[1892]), .feature_below(feature_belows[1892]), .scan_win_std_dev(scan_win_std_dev[1892]), .feature_accum(feature_accums[1892]));
  accum_calculator ac1893(.scan_win(scan_win1893), .rectangle1_x(rectangle1_xs[1893]), .rectangle1_y(rectangle1_ys[1893]), .rectangle1_width(rectangle1_widths[1893]), .rectangle1_height(rectangle1_heights[1893]), .rectangle1_weight(rectangle1_weights[1893]), .rectangle2_x(rectangle2_xs[1893]), .rectangle2_y(rectangle2_ys[1893]), .rectangle2_width(rectangle2_widths[1893]), .rectangle2_height(rectangle2_heights[1893]), .rectangle2_weight(rectangle2_weights[1893]), .rectangle3_x(rectangle3_xs[1893]), .rectangle3_y(rectangle3_ys[1893]), .rectangle3_width(rectangle3_widths[1893]), .rectangle3_height(rectangle3_heights[1893]), .rectangle3_weight(rectangle3_weights[1893]), .feature_threshold(feature_thresholds[1893]), .feature_above(feature_aboves[1893]), .feature_below(feature_belows[1893]), .scan_win_std_dev(scan_win_std_dev[1893]), .feature_accum(feature_accums[1893]));
  accum_calculator ac1894(.scan_win(scan_win1894), .rectangle1_x(rectangle1_xs[1894]), .rectangle1_y(rectangle1_ys[1894]), .rectangle1_width(rectangle1_widths[1894]), .rectangle1_height(rectangle1_heights[1894]), .rectangle1_weight(rectangle1_weights[1894]), .rectangle2_x(rectangle2_xs[1894]), .rectangle2_y(rectangle2_ys[1894]), .rectangle2_width(rectangle2_widths[1894]), .rectangle2_height(rectangle2_heights[1894]), .rectangle2_weight(rectangle2_weights[1894]), .rectangle3_x(rectangle3_xs[1894]), .rectangle3_y(rectangle3_ys[1894]), .rectangle3_width(rectangle3_widths[1894]), .rectangle3_height(rectangle3_heights[1894]), .rectangle3_weight(rectangle3_weights[1894]), .feature_threshold(feature_thresholds[1894]), .feature_above(feature_aboves[1894]), .feature_below(feature_belows[1894]), .scan_win_std_dev(scan_win_std_dev[1894]), .feature_accum(feature_accums[1894]));
  accum_calculator ac1895(.scan_win(scan_win1895), .rectangle1_x(rectangle1_xs[1895]), .rectangle1_y(rectangle1_ys[1895]), .rectangle1_width(rectangle1_widths[1895]), .rectangle1_height(rectangle1_heights[1895]), .rectangle1_weight(rectangle1_weights[1895]), .rectangle2_x(rectangle2_xs[1895]), .rectangle2_y(rectangle2_ys[1895]), .rectangle2_width(rectangle2_widths[1895]), .rectangle2_height(rectangle2_heights[1895]), .rectangle2_weight(rectangle2_weights[1895]), .rectangle3_x(rectangle3_xs[1895]), .rectangle3_y(rectangle3_ys[1895]), .rectangle3_width(rectangle3_widths[1895]), .rectangle3_height(rectangle3_heights[1895]), .rectangle3_weight(rectangle3_weights[1895]), .feature_threshold(feature_thresholds[1895]), .feature_above(feature_aboves[1895]), .feature_below(feature_belows[1895]), .scan_win_std_dev(scan_win_std_dev[1895]), .feature_accum(feature_accums[1895]));
  accum_calculator ac1896(.scan_win(scan_win1896), .rectangle1_x(rectangle1_xs[1896]), .rectangle1_y(rectangle1_ys[1896]), .rectangle1_width(rectangle1_widths[1896]), .rectangle1_height(rectangle1_heights[1896]), .rectangle1_weight(rectangle1_weights[1896]), .rectangle2_x(rectangle2_xs[1896]), .rectangle2_y(rectangle2_ys[1896]), .rectangle2_width(rectangle2_widths[1896]), .rectangle2_height(rectangle2_heights[1896]), .rectangle2_weight(rectangle2_weights[1896]), .rectangle3_x(rectangle3_xs[1896]), .rectangle3_y(rectangle3_ys[1896]), .rectangle3_width(rectangle3_widths[1896]), .rectangle3_height(rectangle3_heights[1896]), .rectangle3_weight(rectangle3_weights[1896]), .feature_threshold(feature_thresholds[1896]), .feature_above(feature_aboves[1896]), .feature_below(feature_belows[1896]), .scan_win_std_dev(scan_win_std_dev[1896]), .feature_accum(feature_accums[1896]));
  accum_calculator ac1897(.scan_win(scan_win1897), .rectangle1_x(rectangle1_xs[1897]), .rectangle1_y(rectangle1_ys[1897]), .rectangle1_width(rectangle1_widths[1897]), .rectangle1_height(rectangle1_heights[1897]), .rectangle1_weight(rectangle1_weights[1897]), .rectangle2_x(rectangle2_xs[1897]), .rectangle2_y(rectangle2_ys[1897]), .rectangle2_width(rectangle2_widths[1897]), .rectangle2_height(rectangle2_heights[1897]), .rectangle2_weight(rectangle2_weights[1897]), .rectangle3_x(rectangle3_xs[1897]), .rectangle3_y(rectangle3_ys[1897]), .rectangle3_width(rectangle3_widths[1897]), .rectangle3_height(rectangle3_heights[1897]), .rectangle3_weight(rectangle3_weights[1897]), .feature_threshold(feature_thresholds[1897]), .feature_above(feature_aboves[1897]), .feature_below(feature_belows[1897]), .scan_win_std_dev(scan_win_std_dev[1897]), .feature_accum(feature_accums[1897]));
  accum_calculator ac1898(.scan_win(scan_win1898), .rectangle1_x(rectangle1_xs[1898]), .rectangle1_y(rectangle1_ys[1898]), .rectangle1_width(rectangle1_widths[1898]), .rectangle1_height(rectangle1_heights[1898]), .rectangle1_weight(rectangle1_weights[1898]), .rectangle2_x(rectangle2_xs[1898]), .rectangle2_y(rectangle2_ys[1898]), .rectangle2_width(rectangle2_widths[1898]), .rectangle2_height(rectangle2_heights[1898]), .rectangle2_weight(rectangle2_weights[1898]), .rectangle3_x(rectangle3_xs[1898]), .rectangle3_y(rectangle3_ys[1898]), .rectangle3_width(rectangle3_widths[1898]), .rectangle3_height(rectangle3_heights[1898]), .rectangle3_weight(rectangle3_weights[1898]), .feature_threshold(feature_thresholds[1898]), .feature_above(feature_aboves[1898]), .feature_below(feature_belows[1898]), .scan_win_std_dev(scan_win_std_dev[1898]), .feature_accum(feature_accums[1898]));
  accum_calculator ac1899(.scan_win(scan_win1899), .rectangle1_x(rectangle1_xs[1899]), .rectangle1_y(rectangle1_ys[1899]), .rectangle1_width(rectangle1_widths[1899]), .rectangle1_height(rectangle1_heights[1899]), .rectangle1_weight(rectangle1_weights[1899]), .rectangle2_x(rectangle2_xs[1899]), .rectangle2_y(rectangle2_ys[1899]), .rectangle2_width(rectangle2_widths[1899]), .rectangle2_height(rectangle2_heights[1899]), .rectangle2_weight(rectangle2_weights[1899]), .rectangle3_x(rectangle3_xs[1899]), .rectangle3_y(rectangle3_ys[1899]), .rectangle3_width(rectangle3_widths[1899]), .rectangle3_height(rectangle3_heights[1899]), .rectangle3_weight(rectangle3_weights[1899]), .feature_threshold(feature_thresholds[1899]), .feature_above(feature_aboves[1899]), .feature_below(feature_belows[1899]), .scan_win_std_dev(scan_win_std_dev[1899]), .feature_accum(feature_accums[1899]));
  accum_calculator ac1900(.scan_win(scan_win1900), .rectangle1_x(rectangle1_xs[1900]), .rectangle1_y(rectangle1_ys[1900]), .rectangle1_width(rectangle1_widths[1900]), .rectangle1_height(rectangle1_heights[1900]), .rectangle1_weight(rectangle1_weights[1900]), .rectangle2_x(rectangle2_xs[1900]), .rectangle2_y(rectangle2_ys[1900]), .rectangle2_width(rectangle2_widths[1900]), .rectangle2_height(rectangle2_heights[1900]), .rectangle2_weight(rectangle2_weights[1900]), .rectangle3_x(rectangle3_xs[1900]), .rectangle3_y(rectangle3_ys[1900]), .rectangle3_width(rectangle3_widths[1900]), .rectangle3_height(rectangle3_heights[1900]), .rectangle3_weight(rectangle3_weights[1900]), .feature_threshold(feature_thresholds[1900]), .feature_above(feature_aboves[1900]), .feature_below(feature_belows[1900]), .scan_win_std_dev(scan_win_std_dev[1900]), .feature_accum(feature_accums[1900]));
  accum_calculator ac1901(.scan_win(scan_win1901), .rectangle1_x(rectangle1_xs[1901]), .rectangle1_y(rectangle1_ys[1901]), .rectangle1_width(rectangle1_widths[1901]), .rectangle1_height(rectangle1_heights[1901]), .rectangle1_weight(rectangle1_weights[1901]), .rectangle2_x(rectangle2_xs[1901]), .rectangle2_y(rectangle2_ys[1901]), .rectangle2_width(rectangle2_widths[1901]), .rectangle2_height(rectangle2_heights[1901]), .rectangle2_weight(rectangle2_weights[1901]), .rectangle3_x(rectangle3_xs[1901]), .rectangle3_y(rectangle3_ys[1901]), .rectangle3_width(rectangle3_widths[1901]), .rectangle3_height(rectangle3_heights[1901]), .rectangle3_weight(rectangle3_weights[1901]), .feature_threshold(feature_thresholds[1901]), .feature_above(feature_aboves[1901]), .feature_below(feature_belows[1901]), .scan_win_std_dev(scan_win_std_dev[1901]), .feature_accum(feature_accums[1901]));
  accum_calculator ac1902(.scan_win(scan_win1902), .rectangle1_x(rectangle1_xs[1902]), .rectangle1_y(rectangle1_ys[1902]), .rectangle1_width(rectangle1_widths[1902]), .rectangle1_height(rectangle1_heights[1902]), .rectangle1_weight(rectangle1_weights[1902]), .rectangle2_x(rectangle2_xs[1902]), .rectangle2_y(rectangle2_ys[1902]), .rectangle2_width(rectangle2_widths[1902]), .rectangle2_height(rectangle2_heights[1902]), .rectangle2_weight(rectangle2_weights[1902]), .rectangle3_x(rectangle3_xs[1902]), .rectangle3_y(rectangle3_ys[1902]), .rectangle3_width(rectangle3_widths[1902]), .rectangle3_height(rectangle3_heights[1902]), .rectangle3_weight(rectangle3_weights[1902]), .feature_threshold(feature_thresholds[1902]), .feature_above(feature_aboves[1902]), .feature_below(feature_belows[1902]), .scan_win_std_dev(scan_win_std_dev[1902]), .feature_accum(feature_accums[1902]));
  accum_calculator ac1903(.scan_win(scan_win1903), .rectangle1_x(rectangle1_xs[1903]), .rectangle1_y(rectangle1_ys[1903]), .rectangle1_width(rectangle1_widths[1903]), .rectangle1_height(rectangle1_heights[1903]), .rectangle1_weight(rectangle1_weights[1903]), .rectangle2_x(rectangle2_xs[1903]), .rectangle2_y(rectangle2_ys[1903]), .rectangle2_width(rectangle2_widths[1903]), .rectangle2_height(rectangle2_heights[1903]), .rectangle2_weight(rectangle2_weights[1903]), .rectangle3_x(rectangle3_xs[1903]), .rectangle3_y(rectangle3_ys[1903]), .rectangle3_width(rectangle3_widths[1903]), .rectangle3_height(rectangle3_heights[1903]), .rectangle3_weight(rectangle3_weights[1903]), .feature_threshold(feature_thresholds[1903]), .feature_above(feature_aboves[1903]), .feature_below(feature_belows[1903]), .scan_win_std_dev(scan_win_std_dev[1903]), .feature_accum(feature_accums[1903]));
  accum_calculator ac1904(.scan_win(scan_win1904), .rectangle1_x(rectangle1_xs[1904]), .rectangle1_y(rectangle1_ys[1904]), .rectangle1_width(rectangle1_widths[1904]), .rectangle1_height(rectangle1_heights[1904]), .rectangle1_weight(rectangle1_weights[1904]), .rectangle2_x(rectangle2_xs[1904]), .rectangle2_y(rectangle2_ys[1904]), .rectangle2_width(rectangle2_widths[1904]), .rectangle2_height(rectangle2_heights[1904]), .rectangle2_weight(rectangle2_weights[1904]), .rectangle3_x(rectangle3_xs[1904]), .rectangle3_y(rectangle3_ys[1904]), .rectangle3_width(rectangle3_widths[1904]), .rectangle3_height(rectangle3_heights[1904]), .rectangle3_weight(rectangle3_weights[1904]), .feature_threshold(feature_thresholds[1904]), .feature_above(feature_aboves[1904]), .feature_below(feature_belows[1904]), .scan_win_std_dev(scan_win_std_dev[1904]), .feature_accum(feature_accums[1904]));
  accum_calculator ac1905(.scan_win(scan_win1905), .rectangle1_x(rectangle1_xs[1905]), .rectangle1_y(rectangle1_ys[1905]), .rectangle1_width(rectangle1_widths[1905]), .rectangle1_height(rectangle1_heights[1905]), .rectangle1_weight(rectangle1_weights[1905]), .rectangle2_x(rectangle2_xs[1905]), .rectangle2_y(rectangle2_ys[1905]), .rectangle2_width(rectangle2_widths[1905]), .rectangle2_height(rectangle2_heights[1905]), .rectangle2_weight(rectangle2_weights[1905]), .rectangle3_x(rectangle3_xs[1905]), .rectangle3_y(rectangle3_ys[1905]), .rectangle3_width(rectangle3_widths[1905]), .rectangle3_height(rectangle3_heights[1905]), .rectangle3_weight(rectangle3_weights[1905]), .feature_threshold(feature_thresholds[1905]), .feature_above(feature_aboves[1905]), .feature_below(feature_belows[1905]), .scan_win_std_dev(scan_win_std_dev[1905]), .feature_accum(feature_accums[1905]));
  accum_calculator ac1906(.scan_win(scan_win1906), .rectangle1_x(rectangle1_xs[1906]), .rectangle1_y(rectangle1_ys[1906]), .rectangle1_width(rectangle1_widths[1906]), .rectangle1_height(rectangle1_heights[1906]), .rectangle1_weight(rectangle1_weights[1906]), .rectangle2_x(rectangle2_xs[1906]), .rectangle2_y(rectangle2_ys[1906]), .rectangle2_width(rectangle2_widths[1906]), .rectangle2_height(rectangle2_heights[1906]), .rectangle2_weight(rectangle2_weights[1906]), .rectangle3_x(rectangle3_xs[1906]), .rectangle3_y(rectangle3_ys[1906]), .rectangle3_width(rectangle3_widths[1906]), .rectangle3_height(rectangle3_heights[1906]), .rectangle3_weight(rectangle3_weights[1906]), .feature_threshold(feature_thresholds[1906]), .feature_above(feature_aboves[1906]), .feature_below(feature_belows[1906]), .scan_win_std_dev(scan_win_std_dev[1906]), .feature_accum(feature_accums[1906]));
  accum_calculator ac1907(.scan_win(scan_win1907), .rectangle1_x(rectangle1_xs[1907]), .rectangle1_y(rectangle1_ys[1907]), .rectangle1_width(rectangle1_widths[1907]), .rectangle1_height(rectangle1_heights[1907]), .rectangle1_weight(rectangle1_weights[1907]), .rectangle2_x(rectangle2_xs[1907]), .rectangle2_y(rectangle2_ys[1907]), .rectangle2_width(rectangle2_widths[1907]), .rectangle2_height(rectangle2_heights[1907]), .rectangle2_weight(rectangle2_weights[1907]), .rectangle3_x(rectangle3_xs[1907]), .rectangle3_y(rectangle3_ys[1907]), .rectangle3_width(rectangle3_widths[1907]), .rectangle3_height(rectangle3_heights[1907]), .rectangle3_weight(rectangle3_weights[1907]), .feature_threshold(feature_thresholds[1907]), .feature_above(feature_aboves[1907]), .feature_below(feature_belows[1907]), .scan_win_std_dev(scan_win_std_dev[1907]), .feature_accum(feature_accums[1907]));
  accum_calculator ac1908(.scan_win(scan_win1908), .rectangle1_x(rectangle1_xs[1908]), .rectangle1_y(rectangle1_ys[1908]), .rectangle1_width(rectangle1_widths[1908]), .rectangle1_height(rectangle1_heights[1908]), .rectangle1_weight(rectangle1_weights[1908]), .rectangle2_x(rectangle2_xs[1908]), .rectangle2_y(rectangle2_ys[1908]), .rectangle2_width(rectangle2_widths[1908]), .rectangle2_height(rectangle2_heights[1908]), .rectangle2_weight(rectangle2_weights[1908]), .rectangle3_x(rectangle3_xs[1908]), .rectangle3_y(rectangle3_ys[1908]), .rectangle3_width(rectangle3_widths[1908]), .rectangle3_height(rectangle3_heights[1908]), .rectangle3_weight(rectangle3_weights[1908]), .feature_threshold(feature_thresholds[1908]), .feature_above(feature_aboves[1908]), .feature_below(feature_belows[1908]), .scan_win_std_dev(scan_win_std_dev[1908]), .feature_accum(feature_accums[1908]));
  accum_calculator ac1909(.scan_win(scan_win1909), .rectangle1_x(rectangle1_xs[1909]), .rectangle1_y(rectangle1_ys[1909]), .rectangle1_width(rectangle1_widths[1909]), .rectangle1_height(rectangle1_heights[1909]), .rectangle1_weight(rectangle1_weights[1909]), .rectangle2_x(rectangle2_xs[1909]), .rectangle2_y(rectangle2_ys[1909]), .rectangle2_width(rectangle2_widths[1909]), .rectangle2_height(rectangle2_heights[1909]), .rectangle2_weight(rectangle2_weights[1909]), .rectangle3_x(rectangle3_xs[1909]), .rectangle3_y(rectangle3_ys[1909]), .rectangle3_width(rectangle3_widths[1909]), .rectangle3_height(rectangle3_heights[1909]), .rectangle3_weight(rectangle3_weights[1909]), .feature_threshold(feature_thresholds[1909]), .feature_above(feature_aboves[1909]), .feature_below(feature_belows[1909]), .scan_win_std_dev(scan_win_std_dev[1909]), .feature_accum(feature_accums[1909]));
  accum_calculator ac1910(.scan_win(scan_win1910), .rectangle1_x(rectangle1_xs[1910]), .rectangle1_y(rectangle1_ys[1910]), .rectangle1_width(rectangle1_widths[1910]), .rectangle1_height(rectangle1_heights[1910]), .rectangle1_weight(rectangle1_weights[1910]), .rectangle2_x(rectangle2_xs[1910]), .rectangle2_y(rectangle2_ys[1910]), .rectangle2_width(rectangle2_widths[1910]), .rectangle2_height(rectangle2_heights[1910]), .rectangle2_weight(rectangle2_weights[1910]), .rectangle3_x(rectangle3_xs[1910]), .rectangle3_y(rectangle3_ys[1910]), .rectangle3_width(rectangle3_widths[1910]), .rectangle3_height(rectangle3_heights[1910]), .rectangle3_weight(rectangle3_weights[1910]), .feature_threshold(feature_thresholds[1910]), .feature_above(feature_aboves[1910]), .feature_below(feature_belows[1910]), .scan_win_std_dev(scan_win_std_dev[1910]), .feature_accum(feature_accums[1910]));
  accum_calculator ac1911(.scan_win(scan_win1911), .rectangle1_x(rectangle1_xs[1911]), .rectangle1_y(rectangle1_ys[1911]), .rectangle1_width(rectangle1_widths[1911]), .rectangle1_height(rectangle1_heights[1911]), .rectangle1_weight(rectangle1_weights[1911]), .rectangle2_x(rectangle2_xs[1911]), .rectangle2_y(rectangle2_ys[1911]), .rectangle2_width(rectangle2_widths[1911]), .rectangle2_height(rectangle2_heights[1911]), .rectangle2_weight(rectangle2_weights[1911]), .rectangle3_x(rectangle3_xs[1911]), .rectangle3_y(rectangle3_ys[1911]), .rectangle3_width(rectangle3_widths[1911]), .rectangle3_height(rectangle3_heights[1911]), .rectangle3_weight(rectangle3_weights[1911]), .feature_threshold(feature_thresholds[1911]), .feature_above(feature_aboves[1911]), .feature_below(feature_belows[1911]), .scan_win_std_dev(scan_win_std_dev[1911]), .feature_accum(feature_accums[1911]));
  accum_calculator ac1912(.scan_win(scan_win1912), .rectangle1_x(rectangle1_xs[1912]), .rectangle1_y(rectangle1_ys[1912]), .rectangle1_width(rectangle1_widths[1912]), .rectangle1_height(rectangle1_heights[1912]), .rectangle1_weight(rectangle1_weights[1912]), .rectangle2_x(rectangle2_xs[1912]), .rectangle2_y(rectangle2_ys[1912]), .rectangle2_width(rectangle2_widths[1912]), .rectangle2_height(rectangle2_heights[1912]), .rectangle2_weight(rectangle2_weights[1912]), .rectangle3_x(rectangle3_xs[1912]), .rectangle3_y(rectangle3_ys[1912]), .rectangle3_width(rectangle3_widths[1912]), .rectangle3_height(rectangle3_heights[1912]), .rectangle3_weight(rectangle3_weights[1912]), .feature_threshold(feature_thresholds[1912]), .feature_above(feature_aboves[1912]), .feature_below(feature_belows[1912]), .scan_win_std_dev(scan_win_std_dev[1912]), .feature_accum(feature_accums[1912]));
  accum_calculator ac1913(.scan_win(scan_win1913), .rectangle1_x(rectangle1_xs[1913]), .rectangle1_y(rectangle1_ys[1913]), .rectangle1_width(rectangle1_widths[1913]), .rectangle1_height(rectangle1_heights[1913]), .rectangle1_weight(rectangle1_weights[1913]), .rectangle2_x(rectangle2_xs[1913]), .rectangle2_y(rectangle2_ys[1913]), .rectangle2_width(rectangle2_widths[1913]), .rectangle2_height(rectangle2_heights[1913]), .rectangle2_weight(rectangle2_weights[1913]), .rectangle3_x(rectangle3_xs[1913]), .rectangle3_y(rectangle3_ys[1913]), .rectangle3_width(rectangle3_widths[1913]), .rectangle3_height(rectangle3_heights[1913]), .rectangle3_weight(rectangle3_weights[1913]), .feature_threshold(feature_thresholds[1913]), .feature_above(feature_aboves[1913]), .feature_below(feature_belows[1913]), .scan_win_std_dev(scan_win_std_dev[1913]), .feature_accum(feature_accums[1913]));
  accum_calculator ac1914(.scan_win(scan_win1914), .rectangle1_x(rectangle1_xs[1914]), .rectangle1_y(rectangle1_ys[1914]), .rectangle1_width(rectangle1_widths[1914]), .rectangle1_height(rectangle1_heights[1914]), .rectangle1_weight(rectangle1_weights[1914]), .rectangle2_x(rectangle2_xs[1914]), .rectangle2_y(rectangle2_ys[1914]), .rectangle2_width(rectangle2_widths[1914]), .rectangle2_height(rectangle2_heights[1914]), .rectangle2_weight(rectangle2_weights[1914]), .rectangle3_x(rectangle3_xs[1914]), .rectangle3_y(rectangle3_ys[1914]), .rectangle3_width(rectangle3_widths[1914]), .rectangle3_height(rectangle3_heights[1914]), .rectangle3_weight(rectangle3_weights[1914]), .feature_threshold(feature_thresholds[1914]), .feature_above(feature_aboves[1914]), .feature_below(feature_belows[1914]), .scan_win_std_dev(scan_win_std_dev[1914]), .feature_accum(feature_accums[1914]));
  accum_calculator ac1915(.scan_win(scan_win1915), .rectangle1_x(rectangle1_xs[1915]), .rectangle1_y(rectangle1_ys[1915]), .rectangle1_width(rectangle1_widths[1915]), .rectangle1_height(rectangle1_heights[1915]), .rectangle1_weight(rectangle1_weights[1915]), .rectangle2_x(rectangle2_xs[1915]), .rectangle2_y(rectangle2_ys[1915]), .rectangle2_width(rectangle2_widths[1915]), .rectangle2_height(rectangle2_heights[1915]), .rectangle2_weight(rectangle2_weights[1915]), .rectangle3_x(rectangle3_xs[1915]), .rectangle3_y(rectangle3_ys[1915]), .rectangle3_width(rectangle3_widths[1915]), .rectangle3_height(rectangle3_heights[1915]), .rectangle3_weight(rectangle3_weights[1915]), .feature_threshold(feature_thresholds[1915]), .feature_above(feature_aboves[1915]), .feature_below(feature_belows[1915]), .scan_win_std_dev(scan_win_std_dev[1915]), .feature_accum(feature_accums[1915]));
  accum_calculator ac1916(.scan_win(scan_win1916), .rectangle1_x(rectangle1_xs[1916]), .rectangle1_y(rectangle1_ys[1916]), .rectangle1_width(rectangle1_widths[1916]), .rectangle1_height(rectangle1_heights[1916]), .rectangle1_weight(rectangle1_weights[1916]), .rectangle2_x(rectangle2_xs[1916]), .rectangle2_y(rectangle2_ys[1916]), .rectangle2_width(rectangle2_widths[1916]), .rectangle2_height(rectangle2_heights[1916]), .rectangle2_weight(rectangle2_weights[1916]), .rectangle3_x(rectangle3_xs[1916]), .rectangle3_y(rectangle3_ys[1916]), .rectangle3_width(rectangle3_widths[1916]), .rectangle3_height(rectangle3_heights[1916]), .rectangle3_weight(rectangle3_weights[1916]), .feature_threshold(feature_thresholds[1916]), .feature_above(feature_aboves[1916]), .feature_below(feature_belows[1916]), .scan_win_std_dev(scan_win_std_dev[1916]), .feature_accum(feature_accums[1916]));
  accum_calculator ac1917(.scan_win(scan_win1917), .rectangle1_x(rectangle1_xs[1917]), .rectangle1_y(rectangle1_ys[1917]), .rectangle1_width(rectangle1_widths[1917]), .rectangle1_height(rectangle1_heights[1917]), .rectangle1_weight(rectangle1_weights[1917]), .rectangle2_x(rectangle2_xs[1917]), .rectangle2_y(rectangle2_ys[1917]), .rectangle2_width(rectangle2_widths[1917]), .rectangle2_height(rectangle2_heights[1917]), .rectangle2_weight(rectangle2_weights[1917]), .rectangle3_x(rectangle3_xs[1917]), .rectangle3_y(rectangle3_ys[1917]), .rectangle3_width(rectangle3_widths[1917]), .rectangle3_height(rectangle3_heights[1917]), .rectangle3_weight(rectangle3_weights[1917]), .feature_threshold(feature_thresholds[1917]), .feature_above(feature_aboves[1917]), .feature_below(feature_belows[1917]), .scan_win_std_dev(scan_win_std_dev[1917]), .feature_accum(feature_accums[1917]));
  accum_calculator ac1918(.scan_win(scan_win1918), .rectangle1_x(rectangle1_xs[1918]), .rectangle1_y(rectangle1_ys[1918]), .rectangle1_width(rectangle1_widths[1918]), .rectangle1_height(rectangle1_heights[1918]), .rectangle1_weight(rectangle1_weights[1918]), .rectangle2_x(rectangle2_xs[1918]), .rectangle2_y(rectangle2_ys[1918]), .rectangle2_width(rectangle2_widths[1918]), .rectangle2_height(rectangle2_heights[1918]), .rectangle2_weight(rectangle2_weights[1918]), .rectangle3_x(rectangle3_xs[1918]), .rectangle3_y(rectangle3_ys[1918]), .rectangle3_width(rectangle3_widths[1918]), .rectangle3_height(rectangle3_heights[1918]), .rectangle3_weight(rectangle3_weights[1918]), .feature_threshold(feature_thresholds[1918]), .feature_above(feature_aboves[1918]), .feature_below(feature_belows[1918]), .scan_win_std_dev(scan_win_std_dev[1918]), .feature_accum(feature_accums[1918]));
  accum_calculator ac1919(.scan_win(scan_win1919), .rectangle1_x(rectangle1_xs[1919]), .rectangle1_y(rectangle1_ys[1919]), .rectangle1_width(rectangle1_widths[1919]), .rectangle1_height(rectangle1_heights[1919]), .rectangle1_weight(rectangle1_weights[1919]), .rectangle2_x(rectangle2_xs[1919]), .rectangle2_y(rectangle2_ys[1919]), .rectangle2_width(rectangle2_widths[1919]), .rectangle2_height(rectangle2_heights[1919]), .rectangle2_weight(rectangle2_weights[1919]), .rectangle3_x(rectangle3_xs[1919]), .rectangle3_y(rectangle3_ys[1919]), .rectangle3_width(rectangle3_widths[1919]), .rectangle3_height(rectangle3_heights[1919]), .rectangle3_weight(rectangle3_weights[1919]), .feature_threshold(feature_thresholds[1919]), .feature_above(feature_aboves[1919]), .feature_below(feature_belows[1919]), .scan_win_std_dev(scan_win_std_dev[1919]), .feature_accum(feature_accums[1919]));
  accum_calculator ac1920(.scan_win(scan_win1920), .rectangle1_x(rectangle1_xs[1920]), .rectangle1_y(rectangle1_ys[1920]), .rectangle1_width(rectangle1_widths[1920]), .rectangle1_height(rectangle1_heights[1920]), .rectangle1_weight(rectangle1_weights[1920]), .rectangle2_x(rectangle2_xs[1920]), .rectangle2_y(rectangle2_ys[1920]), .rectangle2_width(rectangle2_widths[1920]), .rectangle2_height(rectangle2_heights[1920]), .rectangle2_weight(rectangle2_weights[1920]), .rectangle3_x(rectangle3_xs[1920]), .rectangle3_y(rectangle3_ys[1920]), .rectangle3_width(rectangle3_widths[1920]), .rectangle3_height(rectangle3_heights[1920]), .rectangle3_weight(rectangle3_weights[1920]), .feature_threshold(feature_thresholds[1920]), .feature_above(feature_aboves[1920]), .feature_below(feature_belows[1920]), .scan_win_std_dev(scan_win_std_dev[1920]), .feature_accum(feature_accums[1920]));
  accum_calculator ac1921(.scan_win(scan_win1921), .rectangle1_x(rectangle1_xs[1921]), .rectangle1_y(rectangle1_ys[1921]), .rectangle1_width(rectangle1_widths[1921]), .rectangle1_height(rectangle1_heights[1921]), .rectangle1_weight(rectangle1_weights[1921]), .rectangle2_x(rectangle2_xs[1921]), .rectangle2_y(rectangle2_ys[1921]), .rectangle2_width(rectangle2_widths[1921]), .rectangle2_height(rectangle2_heights[1921]), .rectangle2_weight(rectangle2_weights[1921]), .rectangle3_x(rectangle3_xs[1921]), .rectangle3_y(rectangle3_ys[1921]), .rectangle3_width(rectangle3_widths[1921]), .rectangle3_height(rectangle3_heights[1921]), .rectangle3_weight(rectangle3_weights[1921]), .feature_threshold(feature_thresholds[1921]), .feature_above(feature_aboves[1921]), .feature_below(feature_belows[1921]), .scan_win_std_dev(scan_win_std_dev[1921]), .feature_accum(feature_accums[1921]));
  accum_calculator ac1922(.scan_win(scan_win1922), .rectangle1_x(rectangle1_xs[1922]), .rectangle1_y(rectangle1_ys[1922]), .rectangle1_width(rectangle1_widths[1922]), .rectangle1_height(rectangle1_heights[1922]), .rectangle1_weight(rectangle1_weights[1922]), .rectangle2_x(rectangle2_xs[1922]), .rectangle2_y(rectangle2_ys[1922]), .rectangle2_width(rectangle2_widths[1922]), .rectangle2_height(rectangle2_heights[1922]), .rectangle2_weight(rectangle2_weights[1922]), .rectangle3_x(rectangle3_xs[1922]), .rectangle3_y(rectangle3_ys[1922]), .rectangle3_width(rectangle3_widths[1922]), .rectangle3_height(rectangle3_heights[1922]), .rectangle3_weight(rectangle3_weights[1922]), .feature_threshold(feature_thresholds[1922]), .feature_above(feature_aboves[1922]), .feature_below(feature_belows[1922]), .scan_win_std_dev(scan_win_std_dev[1922]), .feature_accum(feature_accums[1922]));
  accum_calculator ac1923(.scan_win(scan_win1923), .rectangle1_x(rectangle1_xs[1923]), .rectangle1_y(rectangle1_ys[1923]), .rectangle1_width(rectangle1_widths[1923]), .rectangle1_height(rectangle1_heights[1923]), .rectangle1_weight(rectangle1_weights[1923]), .rectangle2_x(rectangle2_xs[1923]), .rectangle2_y(rectangle2_ys[1923]), .rectangle2_width(rectangle2_widths[1923]), .rectangle2_height(rectangle2_heights[1923]), .rectangle2_weight(rectangle2_weights[1923]), .rectangle3_x(rectangle3_xs[1923]), .rectangle3_y(rectangle3_ys[1923]), .rectangle3_width(rectangle3_widths[1923]), .rectangle3_height(rectangle3_heights[1923]), .rectangle3_weight(rectangle3_weights[1923]), .feature_threshold(feature_thresholds[1923]), .feature_above(feature_aboves[1923]), .feature_below(feature_belows[1923]), .scan_win_std_dev(scan_win_std_dev[1923]), .feature_accum(feature_accums[1923]));
  accum_calculator ac1924(.scan_win(scan_win1924), .rectangle1_x(rectangle1_xs[1924]), .rectangle1_y(rectangle1_ys[1924]), .rectangle1_width(rectangle1_widths[1924]), .rectangle1_height(rectangle1_heights[1924]), .rectangle1_weight(rectangle1_weights[1924]), .rectangle2_x(rectangle2_xs[1924]), .rectangle2_y(rectangle2_ys[1924]), .rectangle2_width(rectangle2_widths[1924]), .rectangle2_height(rectangle2_heights[1924]), .rectangle2_weight(rectangle2_weights[1924]), .rectangle3_x(rectangle3_xs[1924]), .rectangle3_y(rectangle3_ys[1924]), .rectangle3_width(rectangle3_widths[1924]), .rectangle3_height(rectangle3_heights[1924]), .rectangle3_weight(rectangle3_weights[1924]), .feature_threshold(feature_thresholds[1924]), .feature_above(feature_aboves[1924]), .feature_below(feature_belows[1924]), .scan_win_std_dev(scan_win_std_dev[1924]), .feature_accum(feature_accums[1924]));
  accum_calculator ac1925(.scan_win(scan_win1925), .rectangle1_x(rectangle1_xs[1925]), .rectangle1_y(rectangle1_ys[1925]), .rectangle1_width(rectangle1_widths[1925]), .rectangle1_height(rectangle1_heights[1925]), .rectangle1_weight(rectangle1_weights[1925]), .rectangle2_x(rectangle2_xs[1925]), .rectangle2_y(rectangle2_ys[1925]), .rectangle2_width(rectangle2_widths[1925]), .rectangle2_height(rectangle2_heights[1925]), .rectangle2_weight(rectangle2_weights[1925]), .rectangle3_x(rectangle3_xs[1925]), .rectangle3_y(rectangle3_ys[1925]), .rectangle3_width(rectangle3_widths[1925]), .rectangle3_height(rectangle3_heights[1925]), .rectangle3_weight(rectangle3_weights[1925]), .feature_threshold(feature_thresholds[1925]), .feature_above(feature_aboves[1925]), .feature_below(feature_belows[1925]), .scan_win_std_dev(scan_win_std_dev[1925]), .feature_accum(feature_accums[1925]));
  accum_calculator ac1926(.scan_win(scan_win1926), .rectangle1_x(rectangle1_xs[1926]), .rectangle1_y(rectangle1_ys[1926]), .rectangle1_width(rectangle1_widths[1926]), .rectangle1_height(rectangle1_heights[1926]), .rectangle1_weight(rectangle1_weights[1926]), .rectangle2_x(rectangle2_xs[1926]), .rectangle2_y(rectangle2_ys[1926]), .rectangle2_width(rectangle2_widths[1926]), .rectangle2_height(rectangle2_heights[1926]), .rectangle2_weight(rectangle2_weights[1926]), .rectangle3_x(rectangle3_xs[1926]), .rectangle3_y(rectangle3_ys[1926]), .rectangle3_width(rectangle3_widths[1926]), .rectangle3_height(rectangle3_heights[1926]), .rectangle3_weight(rectangle3_weights[1926]), .feature_threshold(feature_thresholds[1926]), .feature_above(feature_aboves[1926]), .feature_below(feature_belows[1926]), .scan_win_std_dev(scan_win_std_dev[1926]), .feature_accum(feature_accums[1926]));
  accum_calculator ac1927(.scan_win(scan_win1927), .rectangle1_x(rectangle1_xs[1927]), .rectangle1_y(rectangle1_ys[1927]), .rectangle1_width(rectangle1_widths[1927]), .rectangle1_height(rectangle1_heights[1927]), .rectangle1_weight(rectangle1_weights[1927]), .rectangle2_x(rectangle2_xs[1927]), .rectangle2_y(rectangle2_ys[1927]), .rectangle2_width(rectangle2_widths[1927]), .rectangle2_height(rectangle2_heights[1927]), .rectangle2_weight(rectangle2_weights[1927]), .rectangle3_x(rectangle3_xs[1927]), .rectangle3_y(rectangle3_ys[1927]), .rectangle3_width(rectangle3_widths[1927]), .rectangle3_height(rectangle3_heights[1927]), .rectangle3_weight(rectangle3_weights[1927]), .feature_threshold(feature_thresholds[1927]), .feature_above(feature_aboves[1927]), .feature_below(feature_belows[1927]), .scan_win_std_dev(scan_win_std_dev[1927]), .feature_accum(feature_accums[1927]));
  accum_calculator ac1928(.scan_win(scan_win1928), .rectangle1_x(rectangle1_xs[1928]), .rectangle1_y(rectangle1_ys[1928]), .rectangle1_width(rectangle1_widths[1928]), .rectangle1_height(rectangle1_heights[1928]), .rectangle1_weight(rectangle1_weights[1928]), .rectangle2_x(rectangle2_xs[1928]), .rectangle2_y(rectangle2_ys[1928]), .rectangle2_width(rectangle2_widths[1928]), .rectangle2_height(rectangle2_heights[1928]), .rectangle2_weight(rectangle2_weights[1928]), .rectangle3_x(rectangle3_xs[1928]), .rectangle3_y(rectangle3_ys[1928]), .rectangle3_width(rectangle3_widths[1928]), .rectangle3_height(rectangle3_heights[1928]), .rectangle3_weight(rectangle3_weights[1928]), .feature_threshold(feature_thresholds[1928]), .feature_above(feature_aboves[1928]), .feature_below(feature_belows[1928]), .scan_win_std_dev(scan_win_std_dev[1928]), .feature_accum(feature_accums[1928]));
  accum_calculator ac1929(.scan_win(scan_win1929), .rectangle1_x(rectangle1_xs[1929]), .rectangle1_y(rectangle1_ys[1929]), .rectangle1_width(rectangle1_widths[1929]), .rectangle1_height(rectangle1_heights[1929]), .rectangle1_weight(rectangle1_weights[1929]), .rectangle2_x(rectangle2_xs[1929]), .rectangle2_y(rectangle2_ys[1929]), .rectangle2_width(rectangle2_widths[1929]), .rectangle2_height(rectangle2_heights[1929]), .rectangle2_weight(rectangle2_weights[1929]), .rectangle3_x(rectangle3_xs[1929]), .rectangle3_y(rectangle3_ys[1929]), .rectangle3_width(rectangle3_widths[1929]), .rectangle3_height(rectangle3_heights[1929]), .rectangle3_weight(rectangle3_weights[1929]), .feature_threshold(feature_thresholds[1929]), .feature_above(feature_aboves[1929]), .feature_below(feature_belows[1929]), .scan_win_std_dev(scan_win_std_dev[1929]), .feature_accum(feature_accums[1929]));
  accum_calculator ac1930(.scan_win(scan_win1930), .rectangle1_x(rectangle1_xs[1930]), .rectangle1_y(rectangle1_ys[1930]), .rectangle1_width(rectangle1_widths[1930]), .rectangle1_height(rectangle1_heights[1930]), .rectangle1_weight(rectangle1_weights[1930]), .rectangle2_x(rectangle2_xs[1930]), .rectangle2_y(rectangle2_ys[1930]), .rectangle2_width(rectangle2_widths[1930]), .rectangle2_height(rectangle2_heights[1930]), .rectangle2_weight(rectangle2_weights[1930]), .rectangle3_x(rectangle3_xs[1930]), .rectangle3_y(rectangle3_ys[1930]), .rectangle3_width(rectangle3_widths[1930]), .rectangle3_height(rectangle3_heights[1930]), .rectangle3_weight(rectangle3_weights[1930]), .feature_threshold(feature_thresholds[1930]), .feature_above(feature_aboves[1930]), .feature_below(feature_belows[1930]), .scan_win_std_dev(scan_win_std_dev[1930]), .feature_accum(feature_accums[1930]));
  accum_calculator ac1931(.scan_win(scan_win1931), .rectangle1_x(rectangle1_xs[1931]), .rectangle1_y(rectangle1_ys[1931]), .rectangle1_width(rectangle1_widths[1931]), .rectangle1_height(rectangle1_heights[1931]), .rectangle1_weight(rectangle1_weights[1931]), .rectangle2_x(rectangle2_xs[1931]), .rectangle2_y(rectangle2_ys[1931]), .rectangle2_width(rectangle2_widths[1931]), .rectangle2_height(rectangle2_heights[1931]), .rectangle2_weight(rectangle2_weights[1931]), .rectangle3_x(rectangle3_xs[1931]), .rectangle3_y(rectangle3_ys[1931]), .rectangle3_width(rectangle3_widths[1931]), .rectangle3_height(rectangle3_heights[1931]), .rectangle3_weight(rectangle3_weights[1931]), .feature_threshold(feature_thresholds[1931]), .feature_above(feature_aboves[1931]), .feature_below(feature_belows[1931]), .scan_win_std_dev(scan_win_std_dev[1931]), .feature_accum(feature_accums[1931]));
  accum_calculator ac1932(.scan_win(scan_win1932), .rectangle1_x(rectangle1_xs[1932]), .rectangle1_y(rectangle1_ys[1932]), .rectangle1_width(rectangle1_widths[1932]), .rectangle1_height(rectangle1_heights[1932]), .rectangle1_weight(rectangle1_weights[1932]), .rectangle2_x(rectangle2_xs[1932]), .rectangle2_y(rectangle2_ys[1932]), .rectangle2_width(rectangle2_widths[1932]), .rectangle2_height(rectangle2_heights[1932]), .rectangle2_weight(rectangle2_weights[1932]), .rectangle3_x(rectangle3_xs[1932]), .rectangle3_y(rectangle3_ys[1932]), .rectangle3_width(rectangle3_widths[1932]), .rectangle3_height(rectangle3_heights[1932]), .rectangle3_weight(rectangle3_weights[1932]), .feature_threshold(feature_thresholds[1932]), .feature_above(feature_aboves[1932]), .feature_below(feature_belows[1932]), .scan_win_std_dev(scan_win_std_dev[1932]), .feature_accum(feature_accums[1932]));
  accum_calculator ac1933(.scan_win(scan_win1933), .rectangle1_x(rectangle1_xs[1933]), .rectangle1_y(rectangle1_ys[1933]), .rectangle1_width(rectangle1_widths[1933]), .rectangle1_height(rectangle1_heights[1933]), .rectangle1_weight(rectangle1_weights[1933]), .rectangle2_x(rectangle2_xs[1933]), .rectangle2_y(rectangle2_ys[1933]), .rectangle2_width(rectangle2_widths[1933]), .rectangle2_height(rectangle2_heights[1933]), .rectangle2_weight(rectangle2_weights[1933]), .rectangle3_x(rectangle3_xs[1933]), .rectangle3_y(rectangle3_ys[1933]), .rectangle3_width(rectangle3_widths[1933]), .rectangle3_height(rectangle3_heights[1933]), .rectangle3_weight(rectangle3_weights[1933]), .feature_threshold(feature_thresholds[1933]), .feature_above(feature_aboves[1933]), .feature_below(feature_belows[1933]), .scan_win_std_dev(scan_win_std_dev[1933]), .feature_accum(feature_accums[1933]));
  accum_calculator ac1934(.scan_win(scan_win1934), .rectangle1_x(rectangle1_xs[1934]), .rectangle1_y(rectangle1_ys[1934]), .rectangle1_width(rectangle1_widths[1934]), .rectangle1_height(rectangle1_heights[1934]), .rectangle1_weight(rectangle1_weights[1934]), .rectangle2_x(rectangle2_xs[1934]), .rectangle2_y(rectangle2_ys[1934]), .rectangle2_width(rectangle2_widths[1934]), .rectangle2_height(rectangle2_heights[1934]), .rectangle2_weight(rectangle2_weights[1934]), .rectangle3_x(rectangle3_xs[1934]), .rectangle3_y(rectangle3_ys[1934]), .rectangle3_width(rectangle3_widths[1934]), .rectangle3_height(rectangle3_heights[1934]), .rectangle3_weight(rectangle3_weights[1934]), .feature_threshold(feature_thresholds[1934]), .feature_above(feature_aboves[1934]), .feature_below(feature_belows[1934]), .scan_win_std_dev(scan_win_std_dev[1934]), .feature_accum(feature_accums[1934]));
  accum_calculator ac1935(.scan_win(scan_win1935), .rectangle1_x(rectangle1_xs[1935]), .rectangle1_y(rectangle1_ys[1935]), .rectangle1_width(rectangle1_widths[1935]), .rectangle1_height(rectangle1_heights[1935]), .rectangle1_weight(rectangle1_weights[1935]), .rectangle2_x(rectangle2_xs[1935]), .rectangle2_y(rectangle2_ys[1935]), .rectangle2_width(rectangle2_widths[1935]), .rectangle2_height(rectangle2_heights[1935]), .rectangle2_weight(rectangle2_weights[1935]), .rectangle3_x(rectangle3_xs[1935]), .rectangle3_y(rectangle3_ys[1935]), .rectangle3_width(rectangle3_widths[1935]), .rectangle3_height(rectangle3_heights[1935]), .rectangle3_weight(rectangle3_weights[1935]), .feature_threshold(feature_thresholds[1935]), .feature_above(feature_aboves[1935]), .feature_below(feature_belows[1935]), .scan_win_std_dev(scan_win_std_dev[1935]), .feature_accum(feature_accums[1935]));
  accum_calculator ac1936(.scan_win(scan_win1936), .rectangle1_x(rectangle1_xs[1936]), .rectangle1_y(rectangle1_ys[1936]), .rectangle1_width(rectangle1_widths[1936]), .rectangle1_height(rectangle1_heights[1936]), .rectangle1_weight(rectangle1_weights[1936]), .rectangle2_x(rectangle2_xs[1936]), .rectangle2_y(rectangle2_ys[1936]), .rectangle2_width(rectangle2_widths[1936]), .rectangle2_height(rectangle2_heights[1936]), .rectangle2_weight(rectangle2_weights[1936]), .rectangle3_x(rectangle3_xs[1936]), .rectangle3_y(rectangle3_ys[1936]), .rectangle3_width(rectangle3_widths[1936]), .rectangle3_height(rectangle3_heights[1936]), .rectangle3_weight(rectangle3_weights[1936]), .feature_threshold(feature_thresholds[1936]), .feature_above(feature_aboves[1936]), .feature_below(feature_belows[1936]), .scan_win_std_dev(scan_win_std_dev[1936]), .feature_accum(feature_accums[1936]));
  accum_calculator ac1937(.scan_win(scan_win1937), .rectangle1_x(rectangle1_xs[1937]), .rectangle1_y(rectangle1_ys[1937]), .rectangle1_width(rectangle1_widths[1937]), .rectangle1_height(rectangle1_heights[1937]), .rectangle1_weight(rectangle1_weights[1937]), .rectangle2_x(rectangle2_xs[1937]), .rectangle2_y(rectangle2_ys[1937]), .rectangle2_width(rectangle2_widths[1937]), .rectangle2_height(rectangle2_heights[1937]), .rectangle2_weight(rectangle2_weights[1937]), .rectangle3_x(rectangle3_xs[1937]), .rectangle3_y(rectangle3_ys[1937]), .rectangle3_width(rectangle3_widths[1937]), .rectangle3_height(rectangle3_heights[1937]), .rectangle3_weight(rectangle3_weights[1937]), .feature_threshold(feature_thresholds[1937]), .feature_above(feature_aboves[1937]), .feature_below(feature_belows[1937]), .scan_win_std_dev(scan_win_std_dev[1937]), .feature_accum(feature_accums[1937]));
  accum_calculator ac1938(.scan_win(scan_win1938), .rectangle1_x(rectangle1_xs[1938]), .rectangle1_y(rectangle1_ys[1938]), .rectangle1_width(rectangle1_widths[1938]), .rectangle1_height(rectangle1_heights[1938]), .rectangle1_weight(rectangle1_weights[1938]), .rectangle2_x(rectangle2_xs[1938]), .rectangle2_y(rectangle2_ys[1938]), .rectangle2_width(rectangle2_widths[1938]), .rectangle2_height(rectangle2_heights[1938]), .rectangle2_weight(rectangle2_weights[1938]), .rectangle3_x(rectangle3_xs[1938]), .rectangle3_y(rectangle3_ys[1938]), .rectangle3_width(rectangle3_widths[1938]), .rectangle3_height(rectangle3_heights[1938]), .rectangle3_weight(rectangle3_weights[1938]), .feature_threshold(feature_thresholds[1938]), .feature_above(feature_aboves[1938]), .feature_below(feature_belows[1938]), .scan_win_std_dev(scan_win_std_dev[1938]), .feature_accum(feature_accums[1938]));
  accum_calculator ac1939(.scan_win(scan_win1939), .rectangle1_x(rectangle1_xs[1939]), .rectangle1_y(rectangle1_ys[1939]), .rectangle1_width(rectangle1_widths[1939]), .rectangle1_height(rectangle1_heights[1939]), .rectangle1_weight(rectangle1_weights[1939]), .rectangle2_x(rectangle2_xs[1939]), .rectangle2_y(rectangle2_ys[1939]), .rectangle2_width(rectangle2_widths[1939]), .rectangle2_height(rectangle2_heights[1939]), .rectangle2_weight(rectangle2_weights[1939]), .rectangle3_x(rectangle3_xs[1939]), .rectangle3_y(rectangle3_ys[1939]), .rectangle3_width(rectangle3_widths[1939]), .rectangle3_height(rectangle3_heights[1939]), .rectangle3_weight(rectangle3_weights[1939]), .feature_threshold(feature_thresholds[1939]), .feature_above(feature_aboves[1939]), .feature_below(feature_belows[1939]), .scan_win_std_dev(scan_win_std_dev[1939]), .feature_accum(feature_accums[1939]));
  accum_calculator ac1940(.scan_win(scan_win1940), .rectangle1_x(rectangle1_xs[1940]), .rectangle1_y(rectangle1_ys[1940]), .rectangle1_width(rectangle1_widths[1940]), .rectangle1_height(rectangle1_heights[1940]), .rectangle1_weight(rectangle1_weights[1940]), .rectangle2_x(rectangle2_xs[1940]), .rectangle2_y(rectangle2_ys[1940]), .rectangle2_width(rectangle2_widths[1940]), .rectangle2_height(rectangle2_heights[1940]), .rectangle2_weight(rectangle2_weights[1940]), .rectangle3_x(rectangle3_xs[1940]), .rectangle3_y(rectangle3_ys[1940]), .rectangle3_width(rectangle3_widths[1940]), .rectangle3_height(rectangle3_heights[1940]), .rectangle3_weight(rectangle3_weights[1940]), .feature_threshold(feature_thresholds[1940]), .feature_above(feature_aboves[1940]), .feature_below(feature_belows[1940]), .scan_win_std_dev(scan_win_std_dev[1940]), .feature_accum(feature_accums[1940]));
  accum_calculator ac1941(.scan_win(scan_win1941), .rectangle1_x(rectangle1_xs[1941]), .rectangle1_y(rectangle1_ys[1941]), .rectangle1_width(rectangle1_widths[1941]), .rectangle1_height(rectangle1_heights[1941]), .rectangle1_weight(rectangle1_weights[1941]), .rectangle2_x(rectangle2_xs[1941]), .rectangle2_y(rectangle2_ys[1941]), .rectangle2_width(rectangle2_widths[1941]), .rectangle2_height(rectangle2_heights[1941]), .rectangle2_weight(rectangle2_weights[1941]), .rectangle3_x(rectangle3_xs[1941]), .rectangle3_y(rectangle3_ys[1941]), .rectangle3_width(rectangle3_widths[1941]), .rectangle3_height(rectangle3_heights[1941]), .rectangle3_weight(rectangle3_weights[1941]), .feature_threshold(feature_thresholds[1941]), .feature_above(feature_aboves[1941]), .feature_below(feature_belows[1941]), .scan_win_std_dev(scan_win_std_dev[1941]), .feature_accum(feature_accums[1941]));
  accum_calculator ac1942(.scan_win(scan_win1942), .rectangle1_x(rectangle1_xs[1942]), .rectangle1_y(rectangle1_ys[1942]), .rectangle1_width(rectangle1_widths[1942]), .rectangle1_height(rectangle1_heights[1942]), .rectangle1_weight(rectangle1_weights[1942]), .rectangle2_x(rectangle2_xs[1942]), .rectangle2_y(rectangle2_ys[1942]), .rectangle2_width(rectangle2_widths[1942]), .rectangle2_height(rectangle2_heights[1942]), .rectangle2_weight(rectangle2_weights[1942]), .rectangle3_x(rectangle3_xs[1942]), .rectangle3_y(rectangle3_ys[1942]), .rectangle3_width(rectangle3_widths[1942]), .rectangle3_height(rectangle3_heights[1942]), .rectangle3_weight(rectangle3_weights[1942]), .feature_threshold(feature_thresholds[1942]), .feature_above(feature_aboves[1942]), .feature_below(feature_belows[1942]), .scan_win_std_dev(scan_win_std_dev[1942]), .feature_accum(feature_accums[1942]));
  accum_calculator ac1943(.scan_win(scan_win1943), .rectangle1_x(rectangle1_xs[1943]), .rectangle1_y(rectangle1_ys[1943]), .rectangle1_width(rectangle1_widths[1943]), .rectangle1_height(rectangle1_heights[1943]), .rectangle1_weight(rectangle1_weights[1943]), .rectangle2_x(rectangle2_xs[1943]), .rectangle2_y(rectangle2_ys[1943]), .rectangle2_width(rectangle2_widths[1943]), .rectangle2_height(rectangle2_heights[1943]), .rectangle2_weight(rectangle2_weights[1943]), .rectangle3_x(rectangle3_xs[1943]), .rectangle3_y(rectangle3_ys[1943]), .rectangle3_width(rectangle3_widths[1943]), .rectangle3_height(rectangle3_heights[1943]), .rectangle3_weight(rectangle3_weights[1943]), .feature_threshold(feature_thresholds[1943]), .feature_above(feature_aboves[1943]), .feature_below(feature_belows[1943]), .scan_win_std_dev(scan_win_std_dev[1943]), .feature_accum(feature_accums[1943]));
  accum_calculator ac1944(.scan_win(scan_win1944), .rectangle1_x(rectangle1_xs[1944]), .rectangle1_y(rectangle1_ys[1944]), .rectangle1_width(rectangle1_widths[1944]), .rectangle1_height(rectangle1_heights[1944]), .rectangle1_weight(rectangle1_weights[1944]), .rectangle2_x(rectangle2_xs[1944]), .rectangle2_y(rectangle2_ys[1944]), .rectangle2_width(rectangle2_widths[1944]), .rectangle2_height(rectangle2_heights[1944]), .rectangle2_weight(rectangle2_weights[1944]), .rectangle3_x(rectangle3_xs[1944]), .rectangle3_y(rectangle3_ys[1944]), .rectangle3_width(rectangle3_widths[1944]), .rectangle3_height(rectangle3_heights[1944]), .rectangle3_weight(rectangle3_weights[1944]), .feature_threshold(feature_thresholds[1944]), .feature_above(feature_aboves[1944]), .feature_below(feature_belows[1944]), .scan_win_std_dev(scan_win_std_dev[1944]), .feature_accum(feature_accums[1944]));
  accum_calculator ac1945(.scan_win(scan_win1945), .rectangle1_x(rectangle1_xs[1945]), .rectangle1_y(rectangle1_ys[1945]), .rectangle1_width(rectangle1_widths[1945]), .rectangle1_height(rectangle1_heights[1945]), .rectangle1_weight(rectangle1_weights[1945]), .rectangle2_x(rectangle2_xs[1945]), .rectangle2_y(rectangle2_ys[1945]), .rectangle2_width(rectangle2_widths[1945]), .rectangle2_height(rectangle2_heights[1945]), .rectangle2_weight(rectangle2_weights[1945]), .rectangle3_x(rectangle3_xs[1945]), .rectangle3_y(rectangle3_ys[1945]), .rectangle3_width(rectangle3_widths[1945]), .rectangle3_height(rectangle3_heights[1945]), .rectangle3_weight(rectangle3_weights[1945]), .feature_threshold(feature_thresholds[1945]), .feature_above(feature_aboves[1945]), .feature_below(feature_belows[1945]), .scan_win_std_dev(scan_win_std_dev[1945]), .feature_accum(feature_accums[1945]));
  accum_calculator ac1946(.scan_win(scan_win1946), .rectangle1_x(rectangle1_xs[1946]), .rectangle1_y(rectangle1_ys[1946]), .rectangle1_width(rectangle1_widths[1946]), .rectangle1_height(rectangle1_heights[1946]), .rectangle1_weight(rectangle1_weights[1946]), .rectangle2_x(rectangle2_xs[1946]), .rectangle2_y(rectangle2_ys[1946]), .rectangle2_width(rectangle2_widths[1946]), .rectangle2_height(rectangle2_heights[1946]), .rectangle2_weight(rectangle2_weights[1946]), .rectangle3_x(rectangle3_xs[1946]), .rectangle3_y(rectangle3_ys[1946]), .rectangle3_width(rectangle3_widths[1946]), .rectangle3_height(rectangle3_heights[1946]), .rectangle3_weight(rectangle3_weights[1946]), .feature_threshold(feature_thresholds[1946]), .feature_above(feature_aboves[1946]), .feature_below(feature_belows[1946]), .scan_win_std_dev(scan_win_std_dev[1946]), .feature_accum(feature_accums[1946]));
  accum_calculator ac1947(.scan_win(scan_win1947), .rectangle1_x(rectangle1_xs[1947]), .rectangle1_y(rectangle1_ys[1947]), .rectangle1_width(rectangle1_widths[1947]), .rectangle1_height(rectangle1_heights[1947]), .rectangle1_weight(rectangle1_weights[1947]), .rectangle2_x(rectangle2_xs[1947]), .rectangle2_y(rectangle2_ys[1947]), .rectangle2_width(rectangle2_widths[1947]), .rectangle2_height(rectangle2_heights[1947]), .rectangle2_weight(rectangle2_weights[1947]), .rectangle3_x(rectangle3_xs[1947]), .rectangle3_y(rectangle3_ys[1947]), .rectangle3_width(rectangle3_widths[1947]), .rectangle3_height(rectangle3_heights[1947]), .rectangle3_weight(rectangle3_weights[1947]), .feature_threshold(feature_thresholds[1947]), .feature_above(feature_aboves[1947]), .feature_below(feature_belows[1947]), .scan_win_std_dev(scan_win_std_dev[1947]), .feature_accum(feature_accums[1947]));
  accum_calculator ac1948(.scan_win(scan_win1948), .rectangle1_x(rectangle1_xs[1948]), .rectangle1_y(rectangle1_ys[1948]), .rectangle1_width(rectangle1_widths[1948]), .rectangle1_height(rectangle1_heights[1948]), .rectangle1_weight(rectangle1_weights[1948]), .rectangle2_x(rectangle2_xs[1948]), .rectangle2_y(rectangle2_ys[1948]), .rectangle2_width(rectangle2_widths[1948]), .rectangle2_height(rectangle2_heights[1948]), .rectangle2_weight(rectangle2_weights[1948]), .rectangle3_x(rectangle3_xs[1948]), .rectangle3_y(rectangle3_ys[1948]), .rectangle3_width(rectangle3_widths[1948]), .rectangle3_height(rectangle3_heights[1948]), .rectangle3_weight(rectangle3_weights[1948]), .feature_threshold(feature_thresholds[1948]), .feature_above(feature_aboves[1948]), .feature_below(feature_belows[1948]), .scan_win_std_dev(scan_win_std_dev[1948]), .feature_accum(feature_accums[1948]));
  accum_calculator ac1949(.scan_win(scan_win1949), .rectangle1_x(rectangle1_xs[1949]), .rectangle1_y(rectangle1_ys[1949]), .rectangle1_width(rectangle1_widths[1949]), .rectangle1_height(rectangle1_heights[1949]), .rectangle1_weight(rectangle1_weights[1949]), .rectangle2_x(rectangle2_xs[1949]), .rectangle2_y(rectangle2_ys[1949]), .rectangle2_width(rectangle2_widths[1949]), .rectangle2_height(rectangle2_heights[1949]), .rectangle2_weight(rectangle2_weights[1949]), .rectangle3_x(rectangle3_xs[1949]), .rectangle3_y(rectangle3_ys[1949]), .rectangle3_width(rectangle3_widths[1949]), .rectangle3_height(rectangle3_heights[1949]), .rectangle3_weight(rectangle3_weights[1949]), .feature_threshold(feature_thresholds[1949]), .feature_above(feature_aboves[1949]), .feature_below(feature_belows[1949]), .scan_win_std_dev(scan_win_std_dev[1949]), .feature_accum(feature_accums[1949]));
  accum_calculator ac1950(.scan_win(scan_win1950), .rectangle1_x(rectangle1_xs[1950]), .rectangle1_y(rectangle1_ys[1950]), .rectangle1_width(rectangle1_widths[1950]), .rectangle1_height(rectangle1_heights[1950]), .rectangle1_weight(rectangle1_weights[1950]), .rectangle2_x(rectangle2_xs[1950]), .rectangle2_y(rectangle2_ys[1950]), .rectangle2_width(rectangle2_widths[1950]), .rectangle2_height(rectangle2_heights[1950]), .rectangle2_weight(rectangle2_weights[1950]), .rectangle3_x(rectangle3_xs[1950]), .rectangle3_y(rectangle3_ys[1950]), .rectangle3_width(rectangle3_widths[1950]), .rectangle3_height(rectangle3_heights[1950]), .rectangle3_weight(rectangle3_weights[1950]), .feature_threshold(feature_thresholds[1950]), .feature_above(feature_aboves[1950]), .feature_below(feature_belows[1950]), .scan_win_std_dev(scan_win_std_dev[1950]), .feature_accum(feature_accums[1950]));
  accum_calculator ac1951(.scan_win(scan_win1951), .rectangle1_x(rectangle1_xs[1951]), .rectangle1_y(rectangle1_ys[1951]), .rectangle1_width(rectangle1_widths[1951]), .rectangle1_height(rectangle1_heights[1951]), .rectangle1_weight(rectangle1_weights[1951]), .rectangle2_x(rectangle2_xs[1951]), .rectangle2_y(rectangle2_ys[1951]), .rectangle2_width(rectangle2_widths[1951]), .rectangle2_height(rectangle2_heights[1951]), .rectangle2_weight(rectangle2_weights[1951]), .rectangle3_x(rectangle3_xs[1951]), .rectangle3_y(rectangle3_ys[1951]), .rectangle3_width(rectangle3_widths[1951]), .rectangle3_height(rectangle3_heights[1951]), .rectangle3_weight(rectangle3_weights[1951]), .feature_threshold(feature_thresholds[1951]), .feature_above(feature_aboves[1951]), .feature_below(feature_belows[1951]), .scan_win_std_dev(scan_win_std_dev[1951]), .feature_accum(feature_accums[1951]));
  accum_calculator ac1952(.scan_win(scan_win1952), .rectangle1_x(rectangle1_xs[1952]), .rectangle1_y(rectangle1_ys[1952]), .rectangle1_width(rectangle1_widths[1952]), .rectangle1_height(rectangle1_heights[1952]), .rectangle1_weight(rectangle1_weights[1952]), .rectangle2_x(rectangle2_xs[1952]), .rectangle2_y(rectangle2_ys[1952]), .rectangle2_width(rectangle2_widths[1952]), .rectangle2_height(rectangle2_heights[1952]), .rectangle2_weight(rectangle2_weights[1952]), .rectangle3_x(rectangle3_xs[1952]), .rectangle3_y(rectangle3_ys[1952]), .rectangle3_width(rectangle3_widths[1952]), .rectangle3_height(rectangle3_heights[1952]), .rectangle3_weight(rectangle3_weights[1952]), .feature_threshold(feature_thresholds[1952]), .feature_above(feature_aboves[1952]), .feature_below(feature_belows[1952]), .scan_win_std_dev(scan_win_std_dev[1952]), .feature_accum(feature_accums[1952]));
  accum_calculator ac1953(.scan_win(scan_win1953), .rectangle1_x(rectangle1_xs[1953]), .rectangle1_y(rectangle1_ys[1953]), .rectangle1_width(rectangle1_widths[1953]), .rectangle1_height(rectangle1_heights[1953]), .rectangle1_weight(rectangle1_weights[1953]), .rectangle2_x(rectangle2_xs[1953]), .rectangle2_y(rectangle2_ys[1953]), .rectangle2_width(rectangle2_widths[1953]), .rectangle2_height(rectangle2_heights[1953]), .rectangle2_weight(rectangle2_weights[1953]), .rectangle3_x(rectangle3_xs[1953]), .rectangle3_y(rectangle3_ys[1953]), .rectangle3_width(rectangle3_widths[1953]), .rectangle3_height(rectangle3_heights[1953]), .rectangle3_weight(rectangle3_weights[1953]), .feature_threshold(feature_thresholds[1953]), .feature_above(feature_aboves[1953]), .feature_below(feature_belows[1953]), .scan_win_std_dev(scan_win_std_dev[1953]), .feature_accum(feature_accums[1953]));
  accum_calculator ac1954(.scan_win(scan_win1954), .rectangle1_x(rectangle1_xs[1954]), .rectangle1_y(rectangle1_ys[1954]), .rectangle1_width(rectangle1_widths[1954]), .rectangle1_height(rectangle1_heights[1954]), .rectangle1_weight(rectangle1_weights[1954]), .rectangle2_x(rectangle2_xs[1954]), .rectangle2_y(rectangle2_ys[1954]), .rectangle2_width(rectangle2_widths[1954]), .rectangle2_height(rectangle2_heights[1954]), .rectangle2_weight(rectangle2_weights[1954]), .rectangle3_x(rectangle3_xs[1954]), .rectangle3_y(rectangle3_ys[1954]), .rectangle3_width(rectangle3_widths[1954]), .rectangle3_height(rectangle3_heights[1954]), .rectangle3_weight(rectangle3_weights[1954]), .feature_threshold(feature_thresholds[1954]), .feature_above(feature_aboves[1954]), .feature_below(feature_belows[1954]), .scan_win_std_dev(scan_win_std_dev[1954]), .feature_accum(feature_accums[1954]));
  accum_calculator ac1955(.scan_win(scan_win1955), .rectangle1_x(rectangle1_xs[1955]), .rectangle1_y(rectangle1_ys[1955]), .rectangle1_width(rectangle1_widths[1955]), .rectangle1_height(rectangle1_heights[1955]), .rectangle1_weight(rectangle1_weights[1955]), .rectangle2_x(rectangle2_xs[1955]), .rectangle2_y(rectangle2_ys[1955]), .rectangle2_width(rectangle2_widths[1955]), .rectangle2_height(rectangle2_heights[1955]), .rectangle2_weight(rectangle2_weights[1955]), .rectangle3_x(rectangle3_xs[1955]), .rectangle3_y(rectangle3_ys[1955]), .rectangle3_width(rectangle3_widths[1955]), .rectangle3_height(rectangle3_heights[1955]), .rectangle3_weight(rectangle3_weights[1955]), .feature_threshold(feature_thresholds[1955]), .feature_above(feature_aboves[1955]), .feature_below(feature_belows[1955]), .scan_win_std_dev(scan_win_std_dev[1955]), .feature_accum(feature_accums[1955]));
  accum_calculator ac1956(.scan_win(scan_win1956), .rectangle1_x(rectangle1_xs[1956]), .rectangle1_y(rectangle1_ys[1956]), .rectangle1_width(rectangle1_widths[1956]), .rectangle1_height(rectangle1_heights[1956]), .rectangle1_weight(rectangle1_weights[1956]), .rectangle2_x(rectangle2_xs[1956]), .rectangle2_y(rectangle2_ys[1956]), .rectangle2_width(rectangle2_widths[1956]), .rectangle2_height(rectangle2_heights[1956]), .rectangle2_weight(rectangle2_weights[1956]), .rectangle3_x(rectangle3_xs[1956]), .rectangle3_y(rectangle3_ys[1956]), .rectangle3_width(rectangle3_widths[1956]), .rectangle3_height(rectangle3_heights[1956]), .rectangle3_weight(rectangle3_weights[1956]), .feature_threshold(feature_thresholds[1956]), .feature_above(feature_aboves[1956]), .feature_below(feature_belows[1956]), .scan_win_std_dev(scan_win_std_dev[1956]), .feature_accum(feature_accums[1956]));
  accum_calculator ac1957(.scan_win(scan_win1957), .rectangle1_x(rectangle1_xs[1957]), .rectangle1_y(rectangle1_ys[1957]), .rectangle1_width(rectangle1_widths[1957]), .rectangle1_height(rectangle1_heights[1957]), .rectangle1_weight(rectangle1_weights[1957]), .rectangle2_x(rectangle2_xs[1957]), .rectangle2_y(rectangle2_ys[1957]), .rectangle2_width(rectangle2_widths[1957]), .rectangle2_height(rectangle2_heights[1957]), .rectangle2_weight(rectangle2_weights[1957]), .rectangle3_x(rectangle3_xs[1957]), .rectangle3_y(rectangle3_ys[1957]), .rectangle3_width(rectangle3_widths[1957]), .rectangle3_height(rectangle3_heights[1957]), .rectangle3_weight(rectangle3_weights[1957]), .feature_threshold(feature_thresholds[1957]), .feature_above(feature_aboves[1957]), .feature_below(feature_belows[1957]), .scan_win_std_dev(scan_win_std_dev[1957]), .feature_accum(feature_accums[1957]));
  accum_calculator ac1958(.scan_win(scan_win1958), .rectangle1_x(rectangle1_xs[1958]), .rectangle1_y(rectangle1_ys[1958]), .rectangle1_width(rectangle1_widths[1958]), .rectangle1_height(rectangle1_heights[1958]), .rectangle1_weight(rectangle1_weights[1958]), .rectangle2_x(rectangle2_xs[1958]), .rectangle2_y(rectangle2_ys[1958]), .rectangle2_width(rectangle2_widths[1958]), .rectangle2_height(rectangle2_heights[1958]), .rectangle2_weight(rectangle2_weights[1958]), .rectangle3_x(rectangle3_xs[1958]), .rectangle3_y(rectangle3_ys[1958]), .rectangle3_width(rectangle3_widths[1958]), .rectangle3_height(rectangle3_heights[1958]), .rectangle3_weight(rectangle3_weights[1958]), .feature_threshold(feature_thresholds[1958]), .feature_above(feature_aboves[1958]), .feature_below(feature_belows[1958]), .scan_win_std_dev(scan_win_std_dev[1958]), .feature_accum(feature_accums[1958]));
  accum_calculator ac1959(.scan_win(scan_win1959), .rectangle1_x(rectangle1_xs[1959]), .rectangle1_y(rectangle1_ys[1959]), .rectangle1_width(rectangle1_widths[1959]), .rectangle1_height(rectangle1_heights[1959]), .rectangle1_weight(rectangle1_weights[1959]), .rectangle2_x(rectangle2_xs[1959]), .rectangle2_y(rectangle2_ys[1959]), .rectangle2_width(rectangle2_widths[1959]), .rectangle2_height(rectangle2_heights[1959]), .rectangle2_weight(rectangle2_weights[1959]), .rectangle3_x(rectangle3_xs[1959]), .rectangle3_y(rectangle3_ys[1959]), .rectangle3_width(rectangle3_widths[1959]), .rectangle3_height(rectangle3_heights[1959]), .rectangle3_weight(rectangle3_weights[1959]), .feature_threshold(feature_thresholds[1959]), .feature_above(feature_aboves[1959]), .feature_below(feature_belows[1959]), .scan_win_std_dev(scan_win_std_dev[1959]), .feature_accum(feature_accums[1959]));
  accum_calculator ac1960(.scan_win(scan_win1960), .rectangle1_x(rectangle1_xs[1960]), .rectangle1_y(rectangle1_ys[1960]), .rectangle1_width(rectangle1_widths[1960]), .rectangle1_height(rectangle1_heights[1960]), .rectangle1_weight(rectangle1_weights[1960]), .rectangle2_x(rectangle2_xs[1960]), .rectangle2_y(rectangle2_ys[1960]), .rectangle2_width(rectangle2_widths[1960]), .rectangle2_height(rectangle2_heights[1960]), .rectangle2_weight(rectangle2_weights[1960]), .rectangle3_x(rectangle3_xs[1960]), .rectangle3_y(rectangle3_ys[1960]), .rectangle3_width(rectangle3_widths[1960]), .rectangle3_height(rectangle3_heights[1960]), .rectangle3_weight(rectangle3_weights[1960]), .feature_threshold(feature_thresholds[1960]), .feature_above(feature_aboves[1960]), .feature_below(feature_belows[1960]), .scan_win_std_dev(scan_win_std_dev[1960]), .feature_accum(feature_accums[1960]));
  accum_calculator ac1961(.scan_win(scan_win1961), .rectangle1_x(rectangle1_xs[1961]), .rectangle1_y(rectangle1_ys[1961]), .rectangle1_width(rectangle1_widths[1961]), .rectangle1_height(rectangle1_heights[1961]), .rectangle1_weight(rectangle1_weights[1961]), .rectangle2_x(rectangle2_xs[1961]), .rectangle2_y(rectangle2_ys[1961]), .rectangle2_width(rectangle2_widths[1961]), .rectangle2_height(rectangle2_heights[1961]), .rectangle2_weight(rectangle2_weights[1961]), .rectangle3_x(rectangle3_xs[1961]), .rectangle3_y(rectangle3_ys[1961]), .rectangle3_width(rectangle3_widths[1961]), .rectangle3_height(rectangle3_heights[1961]), .rectangle3_weight(rectangle3_weights[1961]), .feature_threshold(feature_thresholds[1961]), .feature_above(feature_aboves[1961]), .feature_below(feature_belows[1961]), .scan_win_std_dev(scan_win_std_dev[1961]), .feature_accum(feature_accums[1961]));
  accum_calculator ac1962(.scan_win(scan_win1962), .rectangle1_x(rectangle1_xs[1962]), .rectangle1_y(rectangle1_ys[1962]), .rectangle1_width(rectangle1_widths[1962]), .rectangle1_height(rectangle1_heights[1962]), .rectangle1_weight(rectangle1_weights[1962]), .rectangle2_x(rectangle2_xs[1962]), .rectangle2_y(rectangle2_ys[1962]), .rectangle2_width(rectangle2_widths[1962]), .rectangle2_height(rectangle2_heights[1962]), .rectangle2_weight(rectangle2_weights[1962]), .rectangle3_x(rectangle3_xs[1962]), .rectangle3_y(rectangle3_ys[1962]), .rectangle3_width(rectangle3_widths[1962]), .rectangle3_height(rectangle3_heights[1962]), .rectangle3_weight(rectangle3_weights[1962]), .feature_threshold(feature_thresholds[1962]), .feature_above(feature_aboves[1962]), .feature_below(feature_belows[1962]), .scan_win_std_dev(scan_win_std_dev[1962]), .feature_accum(feature_accums[1962]));
  accum_calculator ac1963(.scan_win(scan_win1963), .rectangle1_x(rectangle1_xs[1963]), .rectangle1_y(rectangle1_ys[1963]), .rectangle1_width(rectangle1_widths[1963]), .rectangle1_height(rectangle1_heights[1963]), .rectangle1_weight(rectangle1_weights[1963]), .rectangle2_x(rectangle2_xs[1963]), .rectangle2_y(rectangle2_ys[1963]), .rectangle2_width(rectangle2_widths[1963]), .rectangle2_height(rectangle2_heights[1963]), .rectangle2_weight(rectangle2_weights[1963]), .rectangle3_x(rectangle3_xs[1963]), .rectangle3_y(rectangle3_ys[1963]), .rectangle3_width(rectangle3_widths[1963]), .rectangle3_height(rectangle3_heights[1963]), .rectangle3_weight(rectangle3_weights[1963]), .feature_threshold(feature_thresholds[1963]), .feature_above(feature_aboves[1963]), .feature_below(feature_belows[1963]), .scan_win_std_dev(scan_win_std_dev[1963]), .feature_accum(feature_accums[1963]));
  accum_calculator ac1964(.scan_win(scan_win1964), .rectangle1_x(rectangle1_xs[1964]), .rectangle1_y(rectangle1_ys[1964]), .rectangle1_width(rectangle1_widths[1964]), .rectangle1_height(rectangle1_heights[1964]), .rectangle1_weight(rectangle1_weights[1964]), .rectangle2_x(rectangle2_xs[1964]), .rectangle2_y(rectangle2_ys[1964]), .rectangle2_width(rectangle2_widths[1964]), .rectangle2_height(rectangle2_heights[1964]), .rectangle2_weight(rectangle2_weights[1964]), .rectangle3_x(rectangle3_xs[1964]), .rectangle3_y(rectangle3_ys[1964]), .rectangle3_width(rectangle3_widths[1964]), .rectangle3_height(rectangle3_heights[1964]), .rectangle3_weight(rectangle3_weights[1964]), .feature_threshold(feature_thresholds[1964]), .feature_above(feature_aboves[1964]), .feature_below(feature_belows[1964]), .scan_win_std_dev(scan_win_std_dev[1964]), .feature_accum(feature_accums[1964]));
  accum_calculator ac1965(.scan_win(scan_win1965), .rectangle1_x(rectangle1_xs[1965]), .rectangle1_y(rectangle1_ys[1965]), .rectangle1_width(rectangle1_widths[1965]), .rectangle1_height(rectangle1_heights[1965]), .rectangle1_weight(rectangle1_weights[1965]), .rectangle2_x(rectangle2_xs[1965]), .rectangle2_y(rectangle2_ys[1965]), .rectangle2_width(rectangle2_widths[1965]), .rectangle2_height(rectangle2_heights[1965]), .rectangle2_weight(rectangle2_weights[1965]), .rectangle3_x(rectangle3_xs[1965]), .rectangle3_y(rectangle3_ys[1965]), .rectangle3_width(rectangle3_widths[1965]), .rectangle3_height(rectangle3_heights[1965]), .rectangle3_weight(rectangle3_weights[1965]), .feature_threshold(feature_thresholds[1965]), .feature_above(feature_aboves[1965]), .feature_below(feature_belows[1965]), .scan_win_std_dev(scan_win_std_dev[1965]), .feature_accum(feature_accums[1965]));
  accum_calculator ac1966(.scan_win(scan_win1966), .rectangle1_x(rectangle1_xs[1966]), .rectangle1_y(rectangle1_ys[1966]), .rectangle1_width(rectangle1_widths[1966]), .rectangle1_height(rectangle1_heights[1966]), .rectangle1_weight(rectangle1_weights[1966]), .rectangle2_x(rectangle2_xs[1966]), .rectangle2_y(rectangle2_ys[1966]), .rectangle2_width(rectangle2_widths[1966]), .rectangle2_height(rectangle2_heights[1966]), .rectangle2_weight(rectangle2_weights[1966]), .rectangle3_x(rectangle3_xs[1966]), .rectangle3_y(rectangle3_ys[1966]), .rectangle3_width(rectangle3_widths[1966]), .rectangle3_height(rectangle3_heights[1966]), .rectangle3_weight(rectangle3_weights[1966]), .feature_threshold(feature_thresholds[1966]), .feature_above(feature_aboves[1966]), .feature_below(feature_belows[1966]), .scan_win_std_dev(scan_win_std_dev[1966]), .feature_accum(feature_accums[1966]));
  accum_calculator ac1967(.scan_win(scan_win1967), .rectangle1_x(rectangle1_xs[1967]), .rectangle1_y(rectangle1_ys[1967]), .rectangle1_width(rectangle1_widths[1967]), .rectangle1_height(rectangle1_heights[1967]), .rectangle1_weight(rectangle1_weights[1967]), .rectangle2_x(rectangle2_xs[1967]), .rectangle2_y(rectangle2_ys[1967]), .rectangle2_width(rectangle2_widths[1967]), .rectangle2_height(rectangle2_heights[1967]), .rectangle2_weight(rectangle2_weights[1967]), .rectangle3_x(rectangle3_xs[1967]), .rectangle3_y(rectangle3_ys[1967]), .rectangle3_width(rectangle3_widths[1967]), .rectangle3_height(rectangle3_heights[1967]), .rectangle3_weight(rectangle3_weights[1967]), .feature_threshold(feature_thresholds[1967]), .feature_above(feature_aboves[1967]), .feature_below(feature_belows[1967]), .scan_win_std_dev(scan_win_std_dev[1967]), .feature_accum(feature_accums[1967]));
  accum_calculator ac1968(.scan_win(scan_win1968), .rectangle1_x(rectangle1_xs[1968]), .rectangle1_y(rectangle1_ys[1968]), .rectangle1_width(rectangle1_widths[1968]), .rectangle1_height(rectangle1_heights[1968]), .rectangle1_weight(rectangle1_weights[1968]), .rectangle2_x(rectangle2_xs[1968]), .rectangle2_y(rectangle2_ys[1968]), .rectangle2_width(rectangle2_widths[1968]), .rectangle2_height(rectangle2_heights[1968]), .rectangle2_weight(rectangle2_weights[1968]), .rectangle3_x(rectangle3_xs[1968]), .rectangle3_y(rectangle3_ys[1968]), .rectangle3_width(rectangle3_widths[1968]), .rectangle3_height(rectangle3_heights[1968]), .rectangle3_weight(rectangle3_weights[1968]), .feature_threshold(feature_thresholds[1968]), .feature_above(feature_aboves[1968]), .feature_below(feature_belows[1968]), .scan_win_std_dev(scan_win_std_dev[1968]), .feature_accum(feature_accums[1968]));
  accum_calculator ac1969(.scan_win(scan_win1969), .rectangle1_x(rectangle1_xs[1969]), .rectangle1_y(rectangle1_ys[1969]), .rectangle1_width(rectangle1_widths[1969]), .rectangle1_height(rectangle1_heights[1969]), .rectangle1_weight(rectangle1_weights[1969]), .rectangle2_x(rectangle2_xs[1969]), .rectangle2_y(rectangle2_ys[1969]), .rectangle2_width(rectangle2_widths[1969]), .rectangle2_height(rectangle2_heights[1969]), .rectangle2_weight(rectangle2_weights[1969]), .rectangle3_x(rectangle3_xs[1969]), .rectangle3_y(rectangle3_ys[1969]), .rectangle3_width(rectangle3_widths[1969]), .rectangle3_height(rectangle3_heights[1969]), .rectangle3_weight(rectangle3_weights[1969]), .feature_threshold(feature_thresholds[1969]), .feature_above(feature_aboves[1969]), .feature_below(feature_belows[1969]), .scan_win_std_dev(scan_win_std_dev[1969]), .feature_accum(feature_accums[1969]));
  accum_calculator ac1970(.scan_win(scan_win1970), .rectangle1_x(rectangle1_xs[1970]), .rectangle1_y(rectangle1_ys[1970]), .rectangle1_width(rectangle1_widths[1970]), .rectangle1_height(rectangle1_heights[1970]), .rectangle1_weight(rectangle1_weights[1970]), .rectangle2_x(rectangle2_xs[1970]), .rectangle2_y(rectangle2_ys[1970]), .rectangle2_width(rectangle2_widths[1970]), .rectangle2_height(rectangle2_heights[1970]), .rectangle2_weight(rectangle2_weights[1970]), .rectangle3_x(rectangle3_xs[1970]), .rectangle3_y(rectangle3_ys[1970]), .rectangle3_width(rectangle3_widths[1970]), .rectangle3_height(rectangle3_heights[1970]), .rectangle3_weight(rectangle3_weights[1970]), .feature_threshold(feature_thresholds[1970]), .feature_above(feature_aboves[1970]), .feature_below(feature_belows[1970]), .scan_win_std_dev(scan_win_std_dev[1970]), .feature_accum(feature_accums[1970]));
  accum_calculator ac1971(.scan_win(scan_win1971), .rectangle1_x(rectangle1_xs[1971]), .rectangle1_y(rectangle1_ys[1971]), .rectangle1_width(rectangle1_widths[1971]), .rectangle1_height(rectangle1_heights[1971]), .rectangle1_weight(rectangle1_weights[1971]), .rectangle2_x(rectangle2_xs[1971]), .rectangle2_y(rectangle2_ys[1971]), .rectangle2_width(rectangle2_widths[1971]), .rectangle2_height(rectangle2_heights[1971]), .rectangle2_weight(rectangle2_weights[1971]), .rectangle3_x(rectangle3_xs[1971]), .rectangle3_y(rectangle3_ys[1971]), .rectangle3_width(rectangle3_widths[1971]), .rectangle3_height(rectangle3_heights[1971]), .rectangle3_weight(rectangle3_weights[1971]), .feature_threshold(feature_thresholds[1971]), .feature_above(feature_aboves[1971]), .feature_below(feature_belows[1971]), .scan_win_std_dev(scan_win_std_dev[1971]), .feature_accum(feature_accums[1971]));
  accum_calculator ac1972(.scan_win(scan_win1972), .rectangle1_x(rectangle1_xs[1972]), .rectangle1_y(rectangle1_ys[1972]), .rectangle1_width(rectangle1_widths[1972]), .rectangle1_height(rectangle1_heights[1972]), .rectangle1_weight(rectangle1_weights[1972]), .rectangle2_x(rectangle2_xs[1972]), .rectangle2_y(rectangle2_ys[1972]), .rectangle2_width(rectangle2_widths[1972]), .rectangle2_height(rectangle2_heights[1972]), .rectangle2_weight(rectangle2_weights[1972]), .rectangle3_x(rectangle3_xs[1972]), .rectangle3_y(rectangle3_ys[1972]), .rectangle3_width(rectangle3_widths[1972]), .rectangle3_height(rectangle3_heights[1972]), .rectangle3_weight(rectangle3_weights[1972]), .feature_threshold(feature_thresholds[1972]), .feature_above(feature_aboves[1972]), .feature_below(feature_belows[1972]), .scan_win_std_dev(scan_win_std_dev[1972]), .feature_accum(feature_accums[1972]));
  accum_calculator ac1973(.scan_win(scan_win1973), .rectangle1_x(rectangle1_xs[1973]), .rectangle1_y(rectangle1_ys[1973]), .rectangle1_width(rectangle1_widths[1973]), .rectangle1_height(rectangle1_heights[1973]), .rectangle1_weight(rectangle1_weights[1973]), .rectangle2_x(rectangle2_xs[1973]), .rectangle2_y(rectangle2_ys[1973]), .rectangle2_width(rectangle2_widths[1973]), .rectangle2_height(rectangle2_heights[1973]), .rectangle2_weight(rectangle2_weights[1973]), .rectangle3_x(rectangle3_xs[1973]), .rectangle3_y(rectangle3_ys[1973]), .rectangle3_width(rectangle3_widths[1973]), .rectangle3_height(rectangle3_heights[1973]), .rectangle3_weight(rectangle3_weights[1973]), .feature_threshold(feature_thresholds[1973]), .feature_above(feature_aboves[1973]), .feature_below(feature_belows[1973]), .scan_win_std_dev(scan_win_std_dev[1973]), .feature_accum(feature_accums[1973]));
  accum_calculator ac1974(.scan_win(scan_win1974), .rectangle1_x(rectangle1_xs[1974]), .rectangle1_y(rectangle1_ys[1974]), .rectangle1_width(rectangle1_widths[1974]), .rectangle1_height(rectangle1_heights[1974]), .rectangle1_weight(rectangle1_weights[1974]), .rectangle2_x(rectangle2_xs[1974]), .rectangle2_y(rectangle2_ys[1974]), .rectangle2_width(rectangle2_widths[1974]), .rectangle2_height(rectangle2_heights[1974]), .rectangle2_weight(rectangle2_weights[1974]), .rectangle3_x(rectangle3_xs[1974]), .rectangle3_y(rectangle3_ys[1974]), .rectangle3_width(rectangle3_widths[1974]), .rectangle3_height(rectangle3_heights[1974]), .rectangle3_weight(rectangle3_weights[1974]), .feature_threshold(feature_thresholds[1974]), .feature_above(feature_aboves[1974]), .feature_below(feature_belows[1974]), .scan_win_std_dev(scan_win_std_dev[1974]), .feature_accum(feature_accums[1974]));
  accum_calculator ac1975(.scan_win(scan_win1975), .rectangle1_x(rectangle1_xs[1975]), .rectangle1_y(rectangle1_ys[1975]), .rectangle1_width(rectangle1_widths[1975]), .rectangle1_height(rectangle1_heights[1975]), .rectangle1_weight(rectangle1_weights[1975]), .rectangle2_x(rectangle2_xs[1975]), .rectangle2_y(rectangle2_ys[1975]), .rectangle2_width(rectangle2_widths[1975]), .rectangle2_height(rectangle2_heights[1975]), .rectangle2_weight(rectangle2_weights[1975]), .rectangle3_x(rectangle3_xs[1975]), .rectangle3_y(rectangle3_ys[1975]), .rectangle3_width(rectangle3_widths[1975]), .rectangle3_height(rectangle3_heights[1975]), .rectangle3_weight(rectangle3_weights[1975]), .feature_threshold(feature_thresholds[1975]), .feature_above(feature_aboves[1975]), .feature_below(feature_belows[1975]), .scan_win_std_dev(scan_win_std_dev[1975]), .feature_accum(feature_accums[1975]));
  accum_calculator ac1976(.scan_win(scan_win1976), .rectangle1_x(rectangle1_xs[1976]), .rectangle1_y(rectangle1_ys[1976]), .rectangle1_width(rectangle1_widths[1976]), .rectangle1_height(rectangle1_heights[1976]), .rectangle1_weight(rectangle1_weights[1976]), .rectangle2_x(rectangle2_xs[1976]), .rectangle2_y(rectangle2_ys[1976]), .rectangle2_width(rectangle2_widths[1976]), .rectangle2_height(rectangle2_heights[1976]), .rectangle2_weight(rectangle2_weights[1976]), .rectangle3_x(rectangle3_xs[1976]), .rectangle3_y(rectangle3_ys[1976]), .rectangle3_width(rectangle3_widths[1976]), .rectangle3_height(rectangle3_heights[1976]), .rectangle3_weight(rectangle3_weights[1976]), .feature_threshold(feature_thresholds[1976]), .feature_above(feature_aboves[1976]), .feature_below(feature_belows[1976]), .scan_win_std_dev(scan_win_std_dev[1976]), .feature_accum(feature_accums[1976]));
  accum_calculator ac1977(.scan_win(scan_win1977), .rectangle1_x(rectangle1_xs[1977]), .rectangle1_y(rectangle1_ys[1977]), .rectangle1_width(rectangle1_widths[1977]), .rectangle1_height(rectangle1_heights[1977]), .rectangle1_weight(rectangle1_weights[1977]), .rectangle2_x(rectangle2_xs[1977]), .rectangle2_y(rectangle2_ys[1977]), .rectangle2_width(rectangle2_widths[1977]), .rectangle2_height(rectangle2_heights[1977]), .rectangle2_weight(rectangle2_weights[1977]), .rectangle3_x(rectangle3_xs[1977]), .rectangle3_y(rectangle3_ys[1977]), .rectangle3_width(rectangle3_widths[1977]), .rectangle3_height(rectangle3_heights[1977]), .rectangle3_weight(rectangle3_weights[1977]), .feature_threshold(feature_thresholds[1977]), .feature_above(feature_aboves[1977]), .feature_below(feature_belows[1977]), .scan_win_std_dev(scan_win_std_dev[1977]), .feature_accum(feature_accums[1977]));
  accum_calculator ac1978(.scan_win(scan_win1978), .rectangle1_x(rectangle1_xs[1978]), .rectangle1_y(rectangle1_ys[1978]), .rectangle1_width(rectangle1_widths[1978]), .rectangle1_height(rectangle1_heights[1978]), .rectangle1_weight(rectangle1_weights[1978]), .rectangle2_x(rectangle2_xs[1978]), .rectangle2_y(rectangle2_ys[1978]), .rectangle2_width(rectangle2_widths[1978]), .rectangle2_height(rectangle2_heights[1978]), .rectangle2_weight(rectangle2_weights[1978]), .rectangle3_x(rectangle3_xs[1978]), .rectangle3_y(rectangle3_ys[1978]), .rectangle3_width(rectangle3_widths[1978]), .rectangle3_height(rectangle3_heights[1978]), .rectangle3_weight(rectangle3_weights[1978]), .feature_threshold(feature_thresholds[1978]), .feature_above(feature_aboves[1978]), .feature_below(feature_belows[1978]), .scan_win_std_dev(scan_win_std_dev[1978]), .feature_accum(feature_accums[1978]));
  accum_calculator ac1979(.scan_win(scan_win1979), .rectangle1_x(rectangle1_xs[1979]), .rectangle1_y(rectangle1_ys[1979]), .rectangle1_width(rectangle1_widths[1979]), .rectangle1_height(rectangle1_heights[1979]), .rectangle1_weight(rectangle1_weights[1979]), .rectangle2_x(rectangle2_xs[1979]), .rectangle2_y(rectangle2_ys[1979]), .rectangle2_width(rectangle2_widths[1979]), .rectangle2_height(rectangle2_heights[1979]), .rectangle2_weight(rectangle2_weights[1979]), .rectangle3_x(rectangle3_xs[1979]), .rectangle3_y(rectangle3_ys[1979]), .rectangle3_width(rectangle3_widths[1979]), .rectangle3_height(rectangle3_heights[1979]), .rectangle3_weight(rectangle3_weights[1979]), .feature_threshold(feature_thresholds[1979]), .feature_above(feature_aboves[1979]), .feature_below(feature_belows[1979]), .scan_win_std_dev(scan_win_std_dev[1979]), .feature_accum(feature_accums[1979]));
  accum_calculator ac1980(.scan_win(scan_win1980), .rectangle1_x(rectangle1_xs[1980]), .rectangle1_y(rectangle1_ys[1980]), .rectangle1_width(rectangle1_widths[1980]), .rectangle1_height(rectangle1_heights[1980]), .rectangle1_weight(rectangle1_weights[1980]), .rectangle2_x(rectangle2_xs[1980]), .rectangle2_y(rectangle2_ys[1980]), .rectangle2_width(rectangle2_widths[1980]), .rectangle2_height(rectangle2_heights[1980]), .rectangle2_weight(rectangle2_weights[1980]), .rectangle3_x(rectangle3_xs[1980]), .rectangle3_y(rectangle3_ys[1980]), .rectangle3_width(rectangle3_widths[1980]), .rectangle3_height(rectangle3_heights[1980]), .rectangle3_weight(rectangle3_weights[1980]), .feature_threshold(feature_thresholds[1980]), .feature_above(feature_aboves[1980]), .feature_below(feature_belows[1980]), .scan_win_std_dev(scan_win_std_dev[1980]), .feature_accum(feature_accums[1980]));
  accum_calculator ac1981(.scan_win(scan_win1981), .rectangle1_x(rectangle1_xs[1981]), .rectangle1_y(rectangle1_ys[1981]), .rectangle1_width(rectangle1_widths[1981]), .rectangle1_height(rectangle1_heights[1981]), .rectangle1_weight(rectangle1_weights[1981]), .rectangle2_x(rectangle2_xs[1981]), .rectangle2_y(rectangle2_ys[1981]), .rectangle2_width(rectangle2_widths[1981]), .rectangle2_height(rectangle2_heights[1981]), .rectangle2_weight(rectangle2_weights[1981]), .rectangle3_x(rectangle3_xs[1981]), .rectangle3_y(rectangle3_ys[1981]), .rectangle3_width(rectangle3_widths[1981]), .rectangle3_height(rectangle3_heights[1981]), .rectangle3_weight(rectangle3_weights[1981]), .feature_threshold(feature_thresholds[1981]), .feature_above(feature_aboves[1981]), .feature_below(feature_belows[1981]), .scan_win_std_dev(scan_win_std_dev[1981]), .feature_accum(feature_accums[1981]));
  accum_calculator ac1982(.scan_win(scan_win1982), .rectangle1_x(rectangle1_xs[1982]), .rectangle1_y(rectangle1_ys[1982]), .rectangle1_width(rectangle1_widths[1982]), .rectangle1_height(rectangle1_heights[1982]), .rectangle1_weight(rectangle1_weights[1982]), .rectangle2_x(rectangle2_xs[1982]), .rectangle2_y(rectangle2_ys[1982]), .rectangle2_width(rectangle2_widths[1982]), .rectangle2_height(rectangle2_heights[1982]), .rectangle2_weight(rectangle2_weights[1982]), .rectangle3_x(rectangle3_xs[1982]), .rectangle3_y(rectangle3_ys[1982]), .rectangle3_width(rectangle3_widths[1982]), .rectangle3_height(rectangle3_heights[1982]), .rectangle3_weight(rectangle3_weights[1982]), .feature_threshold(feature_thresholds[1982]), .feature_above(feature_aboves[1982]), .feature_below(feature_belows[1982]), .scan_win_std_dev(scan_win_std_dev[1982]), .feature_accum(feature_accums[1982]));
  accum_calculator ac1983(.scan_win(scan_win1983), .rectangle1_x(rectangle1_xs[1983]), .rectangle1_y(rectangle1_ys[1983]), .rectangle1_width(rectangle1_widths[1983]), .rectangle1_height(rectangle1_heights[1983]), .rectangle1_weight(rectangle1_weights[1983]), .rectangle2_x(rectangle2_xs[1983]), .rectangle2_y(rectangle2_ys[1983]), .rectangle2_width(rectangle2_widths[1983]), .rectangle2_height(rectangle2_heights[1983]), .rectangle2_weight(rectangle2_weights[1983]), .rectangle3_x(rectangle3_xs[1983]), .rectangle3_y(rectangle3_ys[1983]), .rectangle3_width(rectangle3_widths[1983]), .rectangle3_height(rectangle3_heights[1983]), .rectangle3_weight(rectangle3_weights[1983]), .feature_threshold(feature_thresholds[1983]), .feature_above(feature_aboves[1983]), .feature_below(feature_belows[1983]), .scan_win_std_dev(scan_win_std_dev[1983]), .feature_accum(feature_accums[1983]));
  accum_calculator ac1984(.scan_win(scan_win1984), .rectangle1_x(rectangle1_xs[1984]), .rectangle1_y(rectangle1_ys[1984]), .rectangle1_width(rectangle1_widths[1984]), .rectangle1_height(rectangle1_heights[1984]), .rectangle1_weight(rectangle1_weights[1984]), .rectangle2_x(rectangle2_xs[1984]), .rectangle2_y(rectangle2_ys[1984]), .rectangle2_width(rectangle2_widths[1984]), .rectangle2_height(rectangle2_heights[1984]), .rectangle2_weight(rectangle2_weights[1984]), .rectangle3_x(rectangle3_xs[1984]), .rectangle3_y(rectangle3_ys[1984]), .rectangle3_width(rectangle3_widths[1984]), .rectangle3_height(rectangle3_heights[1984]), .rectangle3_weight(rectangle3_weights[1984]), .feature_threshold(feature_thresholds[1984]), .feature_above(feature_aboves[1984]), .feature_below(feature_belows[1984]), .scan_win_std_dev(scan_win_std_dev[1984]), .feature_accum(feature_accums[1984]));
  accum_calculator ac1985(.scan_win(scan_win1985), .rectangle1_x(rectangle1_xs[1985]), .rectangle1_y(rectangle1_ys[1985]), .rectangle1_width(rectangle1_widths[1985]), .rectangle1_height(rectangle1_heights[1985]), .rectangle1_weight(rectangle1_weights[1985]), .rectangle2_x(rectangle2_xs[1985]), .rectangle2_y(rectangle2_ys[1985]), .rectangle2_width(rectangle2_widths[1985]), .rectangle2_height(rectangle2_heights[1985]), .rectangle2_weight(rectangle2_weights[1985]), .rectangle3_x(rectangle3_xs[1985]), .rectangle3_y(rectangle3_ys[1985]), .rectangle3_width(rectangle3_widths[1985]), .rectangle3_height(rectangle3_heights[1985]), .rectangle3_weight(rectangle3_weights[1985]), .feature_threshold(feature_thresholds[1985]), .feature_above(feature_aboves[1985]), .feature_below(feature_belows[1985]), .scan_win_std_dev(scan_win_std_dev[1985]), .feature_accum(feature_accums[1985]));
  accum_calculator ac1986(.scan_win(scan_win1986), .rectangle1_x(rectangle1_xs[1986]), .rectangle1_y(rectangle1_ys[1986]), .rectangle1_width(rectangle1_widths[1986]), .rectangle1_height(rectangle1_heights[1986]), .rectangle1_weight(rectangle1_weights[1986]), .rectangle2_x(rectangle2_xs[1986]), .rectangle2_y(rectangle2_ys[1986]), .rectangle2_width(rectangle2_widths[1986]), .rectangle2_height(rectangle2_heights[1986]), .rectangle2_weight(rectangle2_weights[1986]), .rectangle3_x(rectangle3_xs[1986]), .rectangle3_y(rectangle3_ys[1986]), .rectangle3_width(rectangle3_widths[1986]), .rectangle3_height(rectangle3_heights[1986]), .rectangle3_weight(rectangle3_weights[1986]), .feature_threshold(feature_thresholds[1986]), .feature_above(feature_aboves[1986]), .feature_below(feature_belows[1986]), .scan_win_std_dev(scan_win_std_dev[1986]), .feature_accum(feature_accums[1986]));
  accum_calculator ac1987(.scan_win(scan_win1987), .rectangle1_x(rectangle1_xs[1987]), .rectangle1_y(rectangle1_ys[1987]), .rectangle1_width(rectangle1_widths[1987]), .rectangle1_height(rectangle1_heights[1987]), .rectangle1_weight(rectangle1_weights[1987]), .rectangle2_x(rectangle2_xs[1987]), .rectangle2_y(rectangle2_ys[1987]), .rectangle2_width(rectangle2_widths[1987]), .rectangle2_height(rectangle2_heights[1987]), .rectangle2_weight(rectangle2_weights[1987]), .rectangle3_x(rectangle3_xs[1987]), .rectangle3_y(rectangle3_ys[1987]), .rectangle3_width(rectangle3_widths[1987]), .rectangle3_height(rectangle3_heights[1987]), .rectangle3_weight(rectangle3_weights[1987]), .feature_threshold(feature_thresholds[1987]), .feature_above(feature_aboves[1987]), .feature_below(feature_belows[1987]), .scan_win_std_dev(scan_win_std_dev[1987]), .feature_accum(feature_accums[1987]));
  accum_calculator ac1988(.scan_win(scan_win1988), .rectangle1_x(rectangle1_xs[1988]), .rectangle1_y(rectangle1_ys[1988]), .rectangle1_width(rectangle1_widths[1988]), .rectangle1_height(rectangle1_heights[1988]), .rectangle1_weight(rectangle1_weights[1988]), .rectangle2_x(rectangle2_xs[1988]), .rectangle2_y(rectangle2_ys[1988]), .rectangle2_width(rectangle2_widths[1988]), .rectangle2_height(rectangle2_heights[1988]), .rectangle2_weight(rectangle2_weights[1988]), .rectangle3_x(rectangle3_xs[1988]), .rectangle3_y(rectangle3_ys[1988]), .rectangle3_width(rectangle3_widths[1988]), .rectangle3_height(rectangle3_heights[1988]), .rectangle3_weight(rectangle3_weights[1988]), .feature_threshold(feature_thresholds[1988]), .feature_above(feature_aboves[1988]), .feature_below(feature_belows[1988]), .scan_win_std_dev(scan_win_std_dev[1988]), .feature_accum(feature_accums[1988]));
  accum_calculator ac1989(.scan_win(scan_win1989), .rectangle1_x(rectangle1_xs[1989]), .rectangle1_y(rectangle1_ys[1989]), .rectangle1_width(rectangle1_widths[1989]), .rectangle1_height(rectangle1_heights[1989]), .rectangle1_weight(rectangle1_weights[1989]), .rectangle2_x(rectangle2_xs[1989]), .rectangle2_y(rectangle2_ys[1989]), .rectangle2_width(rectangle2_widths[1989]), .rectangle2_height(rectangle2_heights[1989]), .rectangle2_weight(rectangle2_weights[1989]), .rectangle3_x(rectangle3_xs[1989]), .rectangle3_y(rectangle3_ys[1989]), .rectangle3_width(rectangle3_widths[1989]), .rectangle3_height(rectangle3_heights[1989]), .rectangle3_weight(rectangle3_weights[1989]), .feature_threshold(feature_thresholds[1989]), .feature_above(feature_aboves[1989]), .feature_below(feature_belows[1989]), .scan_win_std_dev(scan_win_std_dev[1989]), .feature_accum(feature_accums[1989]));
  accum_calculator ac1990(.scan_win(scan_win1990), .rectangle1_x(rectangle1_xs[1990]), .rectangle1_y(rectangle1_ys[1990]), .rectangle1_width(rectangle1_widths[1990]), .rectangle1_height(rectangle1_heights[1990]), .rectangle1_weight(rectangle1_weights[1990]), .rectangle2_x(rectangle2_xs[1990]), .rectangle2_y(rectangle2_ys[1990]), .rectangle2_width(rectangle2_widths[1990]), .rectangle2_height(rectangle2_heights[1990]), .rectangle2_weight(rectangle2_weights[1990]), .rectangle3_x(rectangle3_xs[1990]), .rectangle3_y(rectangle3_ys[1990]), .rectangle3_width(rectangle3_widths[1990]), .rectangle3_height(rectangle3_heights[1990]), .rectangle3_weight(rectangle3_weights[1990]), .feature_threshold(feature_thresholds[1990]), .feature_above(feature_aboves[1990]), .feature_below(feature_belows[1990]), .scan_win_std_dev(scan_win_std_dev[1990]), .feature_accum(feature_accums[1990]));
  accum_calculator ac1991(.scan_win(scan_win1991), .rectangle1_x(rectangle1_xs[1991]), .rectangle1_y(rectangle1_ys[1991]), .rectangle1_width(rectangle1_widths[1991]), .rectangle1_height(rectangle1_heights[1991]), .rectangle1_weight(rectangle1_weights[1991]), .rectangle2_x(rectangle2_xs[1991]), .rectangle2_y(rectangle2_ys[1991]), .rectangle2_width(rectangle2_widths[1991]), .rectangle2_height(rectangle2_heights[1991]), .rectangle2_weight(rectangle2_weights[1991]), .rectangle3_x(rectangle3_xs[1991]), .rectangle3_y(rectangle3_ys[1991]), .rectangle3_width(rectangle3_widths[1991]), .rectangle3_height(rectangle3_heights[1991]), .rectangle3_weight(rectangle3_weights[1991]), .feature_threshold(feature_thresholds[1991]), .feature_above(feature_aboves[1991]), .feature_below(feature_belows[1991]), .scan_win_std_dev(scan_win_std_dev[1991]), .feature_accum(feature_accums[1991]));
  accum_calculator ac1992(.scan_win(scan_win1992), .rectangle1_x(rectangle1_xs[1992]), .rectangle1_y(rectangle1_ys[1992]), .rectangle1_width(rectangle1_widths[1992]), .rectangle1_height(rectangle1_heights[1992]), .rectangle1_weight(rectangle1_weights[1992]), .rectangle2_x(rectangle2_xs[1992]), .rectangle2_y(rectangle2_ys[1992]), .rectangle2_width(rectangle2_widths[1992]), .rectangle2_height(rectangle2_heights[1992]), .rectangle2_weight(rectangle2_weights[1992]), .rectangle3_x(rectangle3_xs[1992]), .rectangle3_y(rectangle3_ys[1992]), .rectangle3_width(rectangle3_widths[1992]), .rectangle3_height(rectangle3_heights[1992]), .rectangle3_weight(rectangle3_weights[1992]), .feature_threshold(feature_thresholds[1992]), .feature_above(feature_aboves[1992]), .feature_below(feature_belows[1992]), .scan_win_std_dev(scan_win_std_dev[1992]), .feature_accum(feature_accums[1992]));
  accum_calculator ac1993(.scan_win(scan_win1993), .rectangle1_x(rectangle1_xs[1993]), .rectangle1_y(rectangle1_ys[1993]), .rectangle1_width(rectangle1_widths[1993]), .rectangle1_height(rectangle1_heights[1993]), .rectangle1_weight(rectangle1_weights[1993]), .rectangle2_x(rectangle2_xs[1993]), .rectangle2_y(rectangle2_ys[1993]), .rectangle2_width(rectangle2_widths[1993]), .rectangle2_height(rectangle2_heights[1993]), .rectangle2_weight(rectangle2_weights[1993]), .rectangle3_x(rectangle3_xs[1993]), .rectangle3_y(rectangle3_ys[1993]), .rectangle3_width(rectangle3_widths[1993]), .rectangle3_height(rectangle3_heights[1993]), .rectangle3_weight(rectangle3_weights[1993]), .feature_threshold(feature_thresholds[1993]), .feature_above(feature_aboves[1993]), .feature_below(feature_belows[1993]), .scan_win_std_dev(scan_win_std_dev[1993]), .feature_accum(feature_accums[1993]));
  accum_calculator ac1994(.scan_win(scan_win1994), .rectangle1_x(rectangle1_xs[1994]), .rectangle1_y(rectangle1_ys[1994]), .rectangle1_width(rectangle1_widths[1994]), .rectangle1_height(rectangle1_heights[1994]), .rectangle1_weight(rectangle1_weights[1994]), .rectangle2_x(rectangle2_xs[1994]), .rectangle2_y(rectangle2_ys[1994]), .rectangle2_width(rectangle2_widths[1994]), .rectangle2_height(rectangle2_heights[1994]), .rectangle2_weight(rectangle2_weights[1994]), .rectangle3_x(rectangle3_xs[1994]), .rectangle3_y(rectangle3_ys[1994]), .rectangle3_width(rectangle3_widths[1994]), .rectangle3_height(rectangle3_heights[1994]), .rectangle3_weight(rectangle3_weights[1994]), .feature_threshold(feature_thresholds[1994]), .feature_above(feature_aboves[1994]), .feature_below(feature_belows[1994]), .scan_win_std_dev(scan_win_std_dev[1994]), .feature_accum(feature_accums[1994]));
  accum_calculator ac1995(.scan_win(scan_win1995), .rectangle1_x(rectangle1_xs[1995]), .rectangle1_y(rectangle1_ys[1995]), .rectangle1_width(rectangle1_widths[1995]), .rectangle1_height(rectangle1_heights[1995]), .rectangle1_weight(rectangle1_weights[1995]), .rectangle2_x(rectangle2_xs[1995]), .rectangle2_y(rectangle2_ys[1995]), .rectangle2_width(rectangle2_widths[1995]), .rectangle2_height(rectangle2_heights[1995]), .rectangle2_weight(rectangle2_weights[1995]), .rectangle3_x(rectangle3_xs[1995]), .rectangle3_y(rectangle3_ys[1995]), .rectangle3_width(rectangle3_widths[1995]), .rectangle3_height(rectangle3_heights[1995]), .rectangle3_weight(rectangle3_weights[1995]), .feature_threshold(feature_thresholds[1995]), .feature_above(feature_aboves[1995]), .feature_below(feature_belows[1995]), .scan_win_std_dev(scan_win_std_dev[1995]), .feature_accum(feature_accums[1995]));
  accum_calculator ac1996(.scan_win(scan_win1996), .rectangle1_x(rectangle1_xs[1996]), .rectangle1_y(rectangle1_ys[1996]), .rectangle1_width(rectangle1_widths[1996]), .rectangle1_height(rectangle1_heights[1996]), .rectangle1_weight(rectangle1_weights[1996]), .rectangle2_x(rectangle2_xs[1996]), .rectangle2_y(rectangle2_ys[1996]), .rectangle2_width(rectangle2_widths[1996]), .rectangle2_height(rectangle2_heights[1996]), .rectangle2_weight(rectangle2_weights[1996]), .rectangle3_x(rectangle3_xs[1996]), .rectangle3_y(rectangle3_ys[1996]), .rectangle3_width(rectangle3_widths[1996]), .rectangle3_height(rectangle3_heights[1996]), .rectangle3_weight(rectangle3_weights[1996]), .feature_threshold(feature_thresholds[1996]), .feature_above(feature_aboves[1996]), .feature_below(feature_belows[1996]), .scan_win_std_dev(scan_win_std_dev[1996]), .feature_accum(feature_accums[1996]));
  accum_calculator ac1997(.scan_win(scan_win1997), .rectangle1_x(rectangle1_xs[1997]), .rectangle1_y(rectangle1_ys[1997]), .rectangle1_width(rectangle1_widths[1997]), .rectangle1_height(rectangle1_heights[1997]), .rectangle1_weight(rectangle1_weights[1997]), .rectangle2_x(rectangle2_xs[1997]), .rectangle2_y(rectangle2_ys[1997]), .rectangle2_width(rectangle2_widths[1997]), .rectangle2_height(rectangle2_heights[1997]), .rectangle2_weight(rectangle2_weights[1997]), .rectangle3_x(rectangle3_xs[1997]), .rectangle3_y(rectangle3_ys[1997]), .rectangle3_width(rectangle3_widths[1997]), .rectangle3_height(rectangle3_heights[1997]), .rectangle3_weight(rectangle3_weights[1997]), .feature_threshold(feature_thresholds[1997]), .feature_above(feature_aboves[1997]), .feature_below(feature_belows[1997]), .scan_win_std_dev(scan_win_std_dev[1997]), .feature_accum(feature_accums[1997]));
  accum_calculator ac1998(.scan_win(scan_win1998), .rectangle1_x(rectangle1_xs[1998]), .rectangle1_y(rectangle1_ys[1998]), .rectangle1_width(rectangle1_widths[1998]), .rectangle1_height(rectangle1_heights[1998]), .rectangle1_weight(rectangle1_weights[1998]), .rectangle2_x(rectangle2_xs[1998]), .rectangle2_y(rectangle2_ys[1998]), .rectangle2_width(rectangle2_widths[1998]), .rectangle2_height(rectangle2_heights[1998]), .rectangle2_weight(rectangle2_weights[1998]), .rectangle3_x(rectangle3_xs[1998]), .rectangle3_y(rectangle3_ys[1998]), .rectangle3_width(rectangle3_widths[1998]), .rectangle3_height(rectangle3_heights[1998]), .rectangle3_weight(rectangle3_weights[1998]), .feature_threshold(feature_thresholds[1998]), .feature_above(feature_aboves[1998]), .feature_below(feature_belows[1998]), .scan_win_std_dev(scan_win_std_dev[1998]), .feature_accum(feature_accums[1998]));
  accum_calculator ac1999(.scan_win(scan_win1999), .rectangle1_x(rectangle1_xs[1999]), .rectangle1_y(rectangle1_ys[1999]), .rectangle1_width(rectangle1_widths[1999]), .rectangle1_height(rectangle1_heights[1999]), .rectangle1_weight(rectangle1_weights[1999]), .rectangle2_x(rectangle2_xs[1999]), .rectangle2_y(rectangle2_ys[1999]), .rectangle2_width(rectangle2_widths[1999]), .rectangle2_height(rectangle2_heights[1999]), .rectangle2_weight(rectangle2_weights[1999]), .rectangle3_x(rectangle3_xs[1999]), .rectangle3_y(rectangle3_ys[1999]), .rectangle3_width(rectangle3_widths[1999]), .rectangle3_height(rectangle3_heights[1999]), .rectangle3_weight(rectangle3_weights[1999]), .feature_threshold(feature_thresholds[1999]), .feature_above(feature_aboves[1999]), .feature_below(feature_belows[1999]), .scan_win_std_dev(scan_win_std_dev[1999]), .feature_accum(feature_accums[1999]));
  accum_calculator ac2000(.scan_win(scan_win2000), .rectangle1_x(rectangle1_xs[2000]), .rectangle1_y(rectangle1_ys[2000]), .rectangle1_width(rectangle1_widths[2000]), .rectangle1_height(rectangle1_heights[2000]), .rectangle1_weight(rectangle1_weights[2000]), .rectangle2_x(rectangle2_xs[2000]), .rectangle2_y(rectangle2_ys[2000]), .rectangle2_width(rectangle2_widths[2000]), .rectangle2_height(rectangle2_heights[2000]), .rectangle2_weight(rectangle2_weights[2000]), .rectangle3_x(rectangle3_xs[2000]), .rectangle3_y(rectangle3_ys[2000]), .rectangle3_width(rectangle3_widths[2000]), .rectangle3_height(rectangle3_heights[2000]), .rectangle3_weight(rectangle3_weights[2000]), .feature_threshold(feature_thresholds[2000]), .feature_above(feature_aboves[2000]), .feature_below(feature_belows[2000]), .scan_win_std_dev(scan_win_std_dev[2000]), .feature_accum(feature_accums[2000]));
  accum_calculator ac2001(.scan_win(scan_win2001), .rectangle1_x(rectangle1_xs[2001]), .rectangle1_y(rectangle1_ys[2001]), .rectangle1_width(rectangle1_widths[2001]), .rectangle1_height(rectangle1_heights[2001]), .rectangle1_weight(rectangle1_weights[2001]), .rectangle2_x(rectangle2_xs[2001]), .rectangle2_y(rectangle2_ys[2001]), .rectangle2_width(rectangle2_widths[2001]), .rectangle2_height(rectangle2_heights[2001]), .rectangle2_weight(rectangle2_weights[2001]), .rectangle3_x(rectangle3_xs[2001]), .rectangle3_y(rectangle3_ys[2001]), .rectangle3_width(rectangle3_widths[2001]), .rectangle3_height(rectangle3_heights[2001]), .rectangle3_weight(rectangle3_weights[2001]), .feature_threshold(feature_thresholds[2001]), .feature_above(feature_aboves[2001]), .feature_below(feature_belows[2001]), .scan_win_std_dev(scan_win_std_dev[2001]), .feature_accum(feature_accums[2001]));
  accum_calculator ac2002(.scan_win(scan_win2002), .rectangle1_x(rectangle1_xs[2002]), .rectangle1_y(rectangle1_ys[2002]), .rectangle1_width(rectangle1_widths[2002]), .rectangle1_height(rectangle1_heights[2002]), .rectangle1_weight(rectangle1_weights[2002]), .rectangle2_x(rectangle2_xs[2002]), .rectangle2_y(rectangle2_ys[2002]), .rectangle2_width(rectangle2_widths[2002]), .rectangle2_height(rectangle2_heights[2002]), .rectangle2_weight(rectangle2_weights[2002]), .rectangle3_x(rectangle3_xs[2002]), .rectangle3_y(rectangle3_ys[2002]), .rectangle3_width(rectangle3_widths[2002]), .rectangle3_height(rectangle3_heights[2002]), .rectangle3_weight(rectangle3_weights[2002]), .feature_threshold(feature_thresholds[2002]), .feature_above(feature_aboves[2002]), .feature_below(feature_belows[2002]), .scan_win_std_dev(scan_win_std_dev[2002]), .feature_accum(feature_accums[2002]));
  accum_calculator ac2003(.scan_win(scan_win2003), .rectangle1_x(rectangle1_xs[2003]), .rectangle1_y(rectangle1_ys[2003]), .rectangle1_width(rectangle1_widths[2003]), .rectangle1_height(rectangle1_heights[2003]), .rectangle1_weight(rectangle1_weights[2003]), .rectangle2_x(rectangle2_xs[2003]), .rectangle2_y(rectangle2_ys[2003]), .rectangle2_width(rectangle2_widths[2003]), .rectangle2_height(rectangle2_heights[2003]), .rectangle2_weight(rectangle2_weights[2003]), .rectangle3_x(rectangle3_xs[2003]), .rectangle3_y(rectangle3_ys[2003]), .rectangle3_width(rectangle3_widths[2003]), .rectangle3_height(rectangle3_heights[2003]), .rectangle3_weight(rectangle3_weights[2003]), .feature_threshold(feature_thresholds[2003]), .feature_above(feature_aboves[2003]), .feature_below(feature_belows[2003]), .scan_win_std_dev(scan_win_std_dev[2003]), .feature_accum(feature_accums[2003]));
  accum_calculator ac2004(.scan_win(scan_win2004), .rectangle1_x(rectangle1_xs[2004]), .rectangle1_y(rectangle1_ys[2004]), .rectangle1_width(rectangle1_widths[2004]), .rectangle1_height(rectangle1_heights[2004]), .rectangle1_weight(rectangle1_weights[2004]), .rectangle2_x(rectangle2_xs[2004]), .rectangle2_y(rectangle2_ys[2004]), .rectangle2_width(rectangle2_widths[2004]), .rectangle2_height(rectangle2_heights[2004]), .rectangle2_weight(rectangle2_weights[2004]), .rectangle3_x(rectangle3_xs[2004]), .rectangle3_y(rectangle3_ys[2004]), .rectangle3_width(rectangle3_widths[2004]), .rectangle3_height(rectangle3_heights[2004]), .rectangle3_weight(rectangle3_weights[2004]), .feature_threshold(feature_thresholds[2004]), .feature_above(feature_aboves[2004]), .feature_below(feature_belows[2004]), .scan_win_std_dev(scan_win_std_dev[2004]), .feature_accum(feature_accums[2004]));
  accum_calculator ac2005(.scan_win(scan_win2005), .rectangle1_x(rectangle1_xs[2005]), .rectangle1_y(rectangle1_ys[2005]), .rectangle1_width(rectangle1_widths[2005]), .rectangle1_height(rectangle1_heights[2005]), .rectangle1_weight(rectangle1_weights[2005]), .rectangle2_x(rectangle2_xs[2005]), .rectangle2_y(rectangle2_ys[2005]), .rectangle2_width(rectangle2_widths[2005]), .rectangle2_height(rectangle2_heights[2005]), .rectangle2_weight(rectangle2_weights[2005]), .rectangle3_x(rectangle3_xs[2005]), .rectangle3_y(rectangle3_ys[2005]), .rectangle3_width(rectangle3_widths[2005]), .rectangle3_height(rectangle3_heights[2005]), .rectangle3_weight(rectangle3_weights[2005]), .feature_threshold(feature_thresholds[2005]), .feature_above(feature_aboves[2005]), .feature_below(feature_belows[2005]), .scan_win_std_dev(scan_win_std_dev[2005]), .feature_accum(feature_accums[2005]));
  accum_calculator ac2006(.scan_win(scan_win2006), .rectangle1_x(rectangle1_xs[2006]), .rectangle1_y(rectangle1_ys[2006]), .rectangle1_width(rectangle1_widths[2006]), .rectangle1_height(rectangle1_heights[2006]), .rectangle1_weight(rectangle1_weights[2006]), .rectangle2_x(rectangle2_xs[2006]), .rectangle2_y(rectangle2_ys[2006]), .rectangle2_width(rectangle2_widths[2006]), .rectangle2_height(rectangle2_heights[2006]), .rectangle2_weight(rectangle2_weights[2006]), .rectangle3_x(rectangle3_xs[2006]), .rectangle3_y(rectangle3_ys[2006]), .rectangle3_width(rectangle3_widths[2006]), .rectangle3_height(rectangle3_heights[2006]), .rectangle3_weight(rectangle3_weights[2006]), .feature_threshold(feature_thresholds[2006]), .feature_above(feature_aboves[2006]), .feature_below(feature_belows[2006]), .scan_win_std_dev(scan_win_std_dev[2006]), .feature_accum(feature_accums[2006]));
  accum_calculator ac2007(.scan_win(scan_win2007), .rectangle1_x(rectangle1_xs[2007]), .rectangle1_y(rectangle1_ys[2007]), .rectangle1_width(rectangle1_widths[2007]), .rectangle1_height(rectangle1_heights[2007]), .rectangle1_weight(rectangle1_weights[2007]), .rectangle2_x(rectangle2_xs[2007]), .rectangle2_y(rectangle2_ys[2007]), .rectangle2_width(rectangle2_widths[2007]), .rectangle2_height(rectangle2_heights[2007]), .rectangle2_weight(rectangle2_weights[2007]), .rectangle3_x(rectangle3_xs[2007]), .rectangle3_y(rectangle3_ys[2007]), .rectangle3_width(rectangle3_widths[2007]), .rectangle3_height(rectangle3_heights[2007]), .rectangle3_weight(rectangle3_weights[2007]), .feature_threshold(feature_thresholds[2007]), .feature_above(feature_aboves[2007]), .feature_below(feature_belows[2007]), .scan_win_std_dev(scan_win_std_dev[2007]), .feature_accum(feature_accums[2007]));
  accum_calculator ac2008(.scan_win(scan_win2008), .rectangle1_x(rectangle1_xs[2008]), .rectangle1_y(rectangle1_ys[2008]), .rectangle1_width(rectangle1_widths[2008]), .rectangle1_height(rectangle1_heights[2008]), .rectangle1_weight(rectangle1_weights[2008]), .rectangle2_x(rectangle2_xs[2008]), .rectangle2_y(rectangle2_ys[2008]), .rectangle2_width(rectangle2_widths[2008]), .rectangle2_height(rectangle2_heights[2008]), .rectangle2_weight(rectangle2_weights[2008]), .rectangle3_x(rectangle3_xs[2008]), .rectangle3_y(rectangle3_ys[2008]), .rectangle3_width(rectangle3_widths[2008]), .rectangle3_height(rectangle3_heights[2008]), .rectangle3_weight(rectangle3_weights[2008]), .feature_threshold(feature_thresholds[2008]), .feature_above(feature_aboves[2008]), .feature_below(feature_belows[2008]), .scan_win_std_dev(scan_win_std_dev[2008]), .feature_accum(feature_accums[2008]));
  accum_calculator ac2009(.scan_win(scan_win2009), .rectangle1_x(rectangle1_xs[2009]), .rectangle1_y(rectangle1_ys[2009]), .rectangle1_width(rectangle1_widths[2009]), .rectangle1_height(rectangle1_heights[2009]), .rectangle1_weight(rectangle1_weights[2009]), .rectangle2_x(rectangle2_xs[2009]), .rectangle2_y(rectangle2_ys[2009]), .rectangle2_width(rectangle2_widths[2009]), .rectangle2_height(rectangle2_heights[2009]), .rectangle2_weight(rectangle2_weights[2009]), .rectangle3_x(rectangle3_xs[2009]), .rectangle3_y(rectangle3_ys[2009]), .rectangle3_width(rectangle3_widths[2009]), .rectangle3_height(rectangle3_heights[2009]), .rectangle3_weight(rectangle3_weights[2009]), .feature_threshold(feature_thresholds[2009]), .feature_above(feature_aboves[2009]), .feature_below(feature_belows[2009]), .scan_win_std_dev(scan_win_std_dev[2009]), .feature_accum(feature_accums[2009]));
  accum_calculator ac2010(.scan_win(scan_win2010), .rectangle1_x(rectangle1_xs[2010]), .rectangle1_y(rectangle1_ys[2010]), .rectangle1_width(rectangle1_widths[2010]), .rectangle1_height(rectangle1_heights[2010]), .rectangle1_weight(rectangle1_weights[2010]), .rectangle2_x(rectangle2_xs[2010]), .rectangle2_y(rectangle2_ys[2010]), .rectangle2_width(rectangle2_widths[2010]), .rectangle2_height(rectangle2_heights[2010]), .rectangle2_weight(rectangle2_weights[2010]), .rectangle3_x(rectangle3_xs[2010]), .rectangle3_y(rectangle3_ys[2010]), .rectangle3_width(rectangle3_widths[2010]), .rectangle3_height(rectangle3_heights[2010]), .rectangle3_weight(rectangle3_weights[2010]), .feature_threshold(feature_thresholds[2010]), .feature_above(feature_aboves[2010]), .feature_below(feature_belows[2010]), .scan_win_std_dev(scan_win_std_dev[2010]), .feature_accum(feature_accums[2010]));
  accum_calculator ac2011(.scan_win(scan_win2011), .rectangle1_x(rectangle1_xs[2011]), .rectangle1_y(rectangle1_ys[2011]), .rectangle1_width(rectangle1_widths[2011]), .rectangle1_height(rectangle1_heights[2011]), .rectangle1_weight(rectangle1_weights[2011]), .rectangle2_x(rectangle2_xs[2011]), .rectangle2_y(rectangle2_ys[2011]), .rectangle2_width(rectangle2_widths[2011]), .rectangle2_height(rectangle2_heights[2011]), .rectangle2_weight(rectangle2_weights[2011]), .rectangle3_x(rectangle3_xs[2011]), .rectangle3_y(rectangle3_ys[2011]), .rectangle3_width(rectangle3_widths[2011]), .rectangle3_height(rectangle3_heights[2011]), .rectangle3_weight(rectangle3_weights[2011]), .feature_threshold(feature_thresholds[2011]), .feature_above(feature_aboves[2011]), .feature_below(feature_belows[2011]), .scan_win_std_dev(scan_win_std_dev[2011]), .feature_accum(feature_accums[2011]));
  accum_calculator ac2012(.scan_win(scan_win2012), .rectangle1_x(rectangle1_xs[2012]), .rectangle1_y(rectangle1_ys[2012]), .rectangle1_width(rectangle1_widths[2012]), .rectangle1_height(rectangle1_heights[2012]), .rectangle1_weight(rectangle1_weights[2012]), .rectangle2_x(rectangle2_xs[2012]), .rectangle2_y(rectangle2_ys[2012]), .rectangle2_width(rectangle2_widths[2012]), .rectangle2_height(rectangle2_heights[2012]), .rectangle2_weight(rectangle2_weights[2012]), .rectangle3_x(rectangle3_xs[2012]), .rectangle3_y(rectangle3_ys[2012]), .rectangle3_width(rectangle3_widths[2012]), .rectangle3_height(rectangle3_heights[2012]), .rectangle3_weight(rectangle3_weights[2012]), .feature_threshold(feature_thresholds[2012]), .feature_above(feature_aboves[2012]), .feature_below(feature_belows[2012]), .scan_win_std_dev(scan_win_std_dev[2012]), .feature_accum(feature_accums[2012]));
  accum_calculator ac2013(.scan_win(scan_win2013), .rectangle1_x(rectangle1_xs[2013]), .rectangle1_y(rectangle1_ys[2013]), .rectangle1_width(rectangle1_widths[2013]), .rectangle1_height(rectangle1_heights[2013]), .rectangle1_weight(rectangle1_weights[2013]), .rectangle2_x(rectangle2_xs[2013]), .rectangle2_y(rectangle2_ys[2013]), .rectangle2_width(rectangle2_widths[2013]), .rectangle2_height(rectangle2_heights[2013]), .rectangle2_weight(rectangle2_weights[2013]), .rectangle3_x(rectangle3_xs[2013]), .rectangle3_y(rectangle3_ys[2013]), .rectangle3_width(rectangle3_widths[2013]), .rectangle3_height(rectangle3_heights[2013]), .rectangle3_weight(rectangle3_weights[2013]), .feature_threshold(feature_thresholds[2013]), .feature_above(feature_aboves[2013]), .feature_below(feature_belows[2013]), .scan_win_std_dev(scan_win_std_dev[2013]), .feature_accum(feature_accums[2013]));
  accum_calculator ac2014(.scan_win(scan_win2014), .rectangle1_x(rectangle1_xs[2014]), .rectangle1_y(rectangle1_ys[2014]), .rectangle1_width(rectangle1_widths[2014]), .rectangle1_height(rectangle1_heights[2014]), .rectangle1_weight(rectangle1_weights[2014]), .rectangle2_x(rectangle2_xs[2014]), .rectangle2_y(rectangle2_ys[2014]), .rectangle2_width(rectangle2_widths[2014]), .rectangle2_height(rectangle2_heights[2014]), .rectangle2_weight(rectangle2_weights[2014]), .rectangle3_x(rectangle3_xs[2014]), .rectangle3_y(rectangle3_ys[2014]), .rectangle3_width(rectangle3_widths[2014]), .rectangle3_height(rectangle3_heights[2014]), .rectangle3_weight(rectangle3_weights[2014]), .feature_threshold(feature_thresholds[2014]), .feature_above(feature_aboves[2014]), .feature_below(feature_belows[2014]), .scan_win_std_dev(scan_win_std_dev[2014]), .feature_accum(feature_accums[2014]));
  accum_calculator ac2015(.scan_win(scan_win2015), .rectangle1_x(rectangle1_xs[2015]), .rectangle1_y(rectangle1_ys[2015]), .rectangle1_width(rectangle1_widths[2015]), .rectangle1_height(rectangle1_heights[2015]), .rectangle1_weight(rectangle1_weights[2015]), .rectangle2_x(rectangle2_xs[2015]), .rectangle2_y(rectangle2_ys[2015]), .rectangle2_width(rectangle2_widths[2015]), .rectangle2_height(rectangle2_heights[2015]), .rectangle2_weight(rectangle2_weights[2015]), .rectangle3_x(rectangle3_xs[2015]), .rectangle3_y(rectangle3_ys[2015]), .rectangle3_width(rectangle3_widths[2015]), .rectangle3_height(rectangle3_heights[2015]), .rectangle3_weight(rectangle3_weights[2015]), .feature_threshold(feature_thresholds[2015]), .feature_above(feature_aboves[2015]), .feature_below(feature_belows[2015]), .scan_win_std_dev(scan_win_std_dev[2015]), .feature_accum(feature_accums[2015]));
  accum_calculator ac2016(.scan_win(scan_win2016), .rectangle1_x(rectangle1_xs[2016]), .rectangle1_y(rectangle1_ys[2016]), .rectangle1_width(rectangle1_widths[2016]), .rectangle1_height(rectangle1_heights[2016]), .rectangle1_weight(rectangle1_weights[2016]), .rectangle2_x(rectangle2_xs[2016]), .rectangle2_y(rectangle2_ys[2016]), .rectangle2_width(rectangle2_widths[2016]), .rectangle2_height(rectangle2_heights[2016]), .rectangle2_weight(rectangle2_weights[2016]), .rectangle3_x(rectangle3_xs[2016]), .rectangle3_y(rectangle3_ys[2016]), .rectangle3_width(rectangle3_widths[2016]), .rectangle3_height(rectangle3_heights[2016]), .rectangle3_weight(rectangle3_weights[2016]), .feature_threshold(feature_thresholds[2016]), .feature_above(feature_aboves[2016]), .feature_below(feature_belows[2016]), .scan_win_std_dev(scan_win_std_dev[2016]), .feature_accum(feature_accums[2016]));
  accum_calculator ac2017(.scan_win(scan_win2017), .rectangle1_x(rectangle1_xs[2017]), .rectangle1_y(rectangle1_ys[2017]), .rectangle1_width(rectangle1_widths[2017]), .rectangle1_height(rectangle1_heights[2017]), .rectangle1_weight(rectangle1_weights[2017]), .rectangle2_x(rectangle2_xs[2017]), .rectangle2_y(rectangle2_ys[2017]), .rectangle2_width(rectangle2_widths[2017]), .rectangle2_height(rectangle2_heights[2017]), .rectangle2_weight(rectangle2_weights[2017]), .rectangle3_x(rectangle3_xs[2017]), .rectangle3_y(rectangle3_ys[2017]), .rectangle3_width(rectangle3_widths[2017]), .rectangle3_height(rectangle3_heights[2017]), .rectangle3_weight(rectangle3_weights[2017]), .feature_threshold(feature_thresholds[2017]), .feature_above(feature_aboves[2017]), .feature_below(feature_belows[2017]), .scan_win_std_dev(scan_win_std_dev[2017]), .feature_accum(feature_accums[2017]));
  accum_calculator ac2018(.scan_win(scan_win2018), .rectangle1_x(rectangle1_xs[2018]), .rectangle1_y(rectangle1_ys[2018]), .rectangle1_width(rectangle1_widths[2018]), .rectangle1_height(rectangle1_heights[2018]), .rectangle1_weight(rectangle1_weights[2018]), .rectangle2_x(rectangle2_xs[2018]), .rectangle2_y(rectangle2_ys[2018]), .rectangle2_width(rectangle2_widths[2018]), .rectangle2_height(rectangle2_heights[2018]), .rectangle2_weight(rectangle2_weights[2018]), .rectangle3_x(rectangle3_xs[2018]), .rectangle3_y(rectangle3_ys[2018]), .rectangle3_width(rectangle3_widths[2018]), .rectangle3_height(rectangle3_heights[2018]), .rectangle3_weight(rectangle3_weights[2018]), .feature_threshold(feature_thresholds[2018]), .feature_above(feature_aboves[2018]), .feature_below(feature_belows[2018]), .scan_win_std_dev(scan_win_std_dev[2018]), .feature_accum(feature_accums[2018]));
  accum_calculator ac2019(.scan_win(scan_win2019), .rectangle1_x(rectangle1_xs[2019]), .rectangle1_y(rectangle1_ys[2019]), .rectangle1_width(rectangle1_widths[2019]), .rectangle1_height(rectangle1_heights[2019]), .rectangle1_weight(rectangle1_weights[2019]), .rectangle2_x(rectangle2_xs[2019]), .rectangle2_y(rectangle2_ys[2019]), .rectangle2_width(rectangle2_widths[2019]), .rectangle2_height(rectangle2_heights[2019]), .rectangle2_weight(rectangle2_weights[2019]), .rectangle3_x(rectangle3_xs[2019]), .rectangle3_y(rectangle3_ys[2019]), .rectangle3_width(rectangle3_widths[2019]), .rectangle3_height(rectangle3_heights[2019]), .rectangle3_weight(rectangle3_weights[2019]), .feature_threshold(feature_thresholds[2019]), .feature_above(feature_aboves[2019]), .feature_below(feature_belows[2019]), .scan_win_std_dev(scan_win_std_dev[2019]), .feature_accum(feature_accums[2019]));
  accum_calculator ac2020(.scan_win(scan_win2020), .rectangle1_x(rectangle1_xs[2020]), .rectangle1_y(rectangle1_ys[2020]), .rectangle1_width(rectangle1_widths[2020]), .rectangle1_height(rectangle1_heights[2020]), .rectangle1_weight(rectangle1_weights[2020]), .rectangle2_x(rectangle2_xs[2020]), .rectangle2_y(rectangle2_ys[2020]), .rectangle2_width(rectangle2_widths[2020]), .rectangle2_height(rectangle2_heights[2020]), .rectangle2_weight(rectangle2_weights[2020]), .rectangle3_x(rectangle3_xs[2020]), .rectangle3_y(rectangle3_ys[2020]), .rectangle3_width(rectangle3_widths[2020]), .rectangle3_height(rectangle3_heights[2020]), .rectangle3_weight(rectangle3_weights[2020]), .feature_threshold(feature_thresholds[2020]), .feature_above(feature_aboves[2020]), .feature_below(feature_belows[2020]), .scan_win_std_dev(scan_win_std_dev[2020]), .feature_accum(feature_accums[2020]));
  accum_calculator ac2021(.scan_win(scan_win2021), .rectangle1_x(rectangle1_xs[2021]), .rectangle1_y(rectangle1_ys[2021]), .rectangle1_width(rectangle1_widths[2021]), .rectangle1_height(rectangle1_heights[2021]), .rectangle1_weight(rectangle1_weights[2021]), .rectangle2_x(rectangle2_xs[2021]), .rectangle2_y(rectangle2_ys[2021]), .rectangle2_width(rectangle2_widths[2021]), .rectangle2_height(rectangle2_heights[2021]), .rectangle2_weight(rectangle2_weights[2021]), .rectangle3_x(rectangle3_xs[2021]), .rectangle3_y(rectangle3_ys[2021]), .rectangle3_width(rectangle3_widths[2021]), .rectangle3_height(rectangle3_heights[2021]), .rectangle3_weight(rectangle3_weights[2021]), .feature_threshold(feature_thresholds[2021]), .feature_above(feature_aboves[2021]), .feature_below(feature_belows[2021]), .scan_win_std_dev(scan_win_std_dev[2021]), .feature_accum(feature_accums[2021]));
  accum_calculator ac2022(.scan_win(scan_win2022), .rectangle1_x(rectangle1_xs[2022]), .rectangle1_y(rectangle1_ys[2022]), .rectangle1_width(rectangle1_widths[2022]), .rectangle1_height(rectangle1_heights[2022]), .rectangle1_weight(rectangle1_weights[2022]), .rectangle2_x(rectangle2_xs[2022]), .rectangle2_y(rectangle2_ys[2022]), .rectangle2_width(rectangle2_widths[2022]), .rectangle2_height(rectangle2_heights[2022]), .rectangle2_weight(rectangle2_weights[2022]), .rectangle3_x(rectangle3_xs[2022]), .rectangle3_y(rectangle3_ys[2022]), .rectangle3_width(rectangle3_widths[2022]), .rectangle3_height(rectangle3_heights[2022]), .rectangle3_weight(rectangle3_weights[2022]), .feature_threshold(feature_thresholds[2022]), .feature_above(feature_aboves[2022]), .feature_below(feature_belows[2022]), .scan_win_std_dev(scan_win_std_dev[2022]), .feature_accum(feature_accums[2022]));
  accum_calculator ac2023(.scan_win(scan_win2023), .rectangle1_x(rectangle1_xs[2023]), .rectangle1_y(rectangle1_ys[2023]), .rectangle1_width(rectangle1_widths[2023]), .rectangle1_height(rectangle1_heights[2023]), .rectangle1_weight(rectangle1_weights[2023]), .rectangle2_x(rectangle2_xs[2023]), .rectangle2_y(rectangle2_ys[2023]), .rectangle2_width(rectangle2_widths[2023]), .rectangle2_height(rectangle2_heights[2023]), .rectangle2_weight(rectangle2_weights[2023]), .rectangle3_x(rectangle3_xs[2023]), .rectangle3_y(rectangle3_ys[2023]), .rectangle3_width(rectangle3_widths[2023]), .rectangle3_height(rectangle3_heights[2023]), .rectangle3_weight(rectangle3_weights[2023]), .feature_threshold(feature_thresholds[2023]), .feature_above(feature_aboves[2023]), .feature_below(feature_belows[2023]), .scan_win_std_dev(scan_win_std_dev[2023]), .feature_accum(feature_accums[2023]));
  accum_calculator ac2024(.scan_win(scan_win2024), .rectangle1_x(rectangle1_xs[2024]), .rectangle1_y(rectangle1_ys[2024]), .rectangle1_width(rectangle1_widths[2024]), .rectangle1_height(rectangle1_heights[2024]), .rectangle1_weight(rectangle1_weights[2024]), .rectangle2_x(rectangle2_xs[2024]), .rectangle2_y(rectangle2_ys[2024]), .rectangle2_width(rectangle2_widths[2024]), .rectangle2_height(rectangle2_heights[2024]), .rectangle2_weight(rectangle2_weights[2024]), .rectangle3_x(rectangle3_xs[2024]), .rectangle3_y(rectangle3_ys[2024]), .rectangle3_width(rectangle3_widths[2024]), .rectangle3_height(rectangle3_heights[2024]), .rectangle3_weight(rectangle3_weights[2024]), .feature_threshold(feature_thresholds[2024]), .feature_above(feature_aboves[2024]), .feature_below(feature_belows[2024]), .scan_win_std_dev(scan_win_std_dev[2024]), .feature_accum(feature_accums[2024]));
  accum_calculator ac2025(.scan_win(scan_win2025), .rectangle1_x(rectangle1_xs[2025]), .rectangle1_y(rectangle1_ys[2025]), .rectangle1_width(rectangle1_widths[2025]), .rectangle1_height(rectangle1_heights[2025]), .rectangle1_weight(rectangle1_weights[2025]), .rectangle2_x(rectangle2_xs[2025]), .rectangle2_y(rectangle2_ys[2025]), .rectangle2_width(rectangle2_widths[2025]), .rectangle2_height(rectangle2_heights[2025]), .rectangle2_weight(rectangle2_weights[2025]), .rectangle3_x(rectangle3_xs[2025]), .rectangle3_y(rectangle3_ys[2025]), .rectangle3_width(rectangle3_widths[2025]), .rectangle3_height(rectangle3_heights[2025]), .rectangle3_weight(rectangle3_weights[2025]), .feature_threshold(feature_thresholds[2025]), .feature_above(feature_aboves[2025]), .feature_below(feature_belows[2025]), .scan_win_std_dev(scan_win_std_dev[2025]), .feature_accum(feature_accums[2025]));
  accum_calculator ac2026(.scan_win(scan_win2026), .rectangle1_x(rectangle1_xs[2026]), .rectangle1_y(rectangle1_ys[2026]), .rectangle1_width(rectangle1_widths[2026]), .rectangle1_height(rectangle1_heights[2026]), .rectangle1_weight(rectangle1_weights[2026]), .rectangle2_x(rectangle2_xs[2026]), .rectangle2_y(rectangle2_ys[2026]), .rectangle2_width(rectangle2_widths[2026]), .rectangle2_height(rectangle2_heights[2026]), .rectangle2_weight(rectangle2_weights[2026]), .rectangle3_x(rectangle3_xs[2026]), .rectangle3_y(rectangle3_ys[2026]), .rectangle3_width(rectangle3_widths[2026]), .rectangle3_height(rectangle3_heights[2026]), .rectangle3_weight(rectangle3_weights[2026]), .feature_threshold(feature_thresholds[2026]), .feature_above(feature_aboves[2026]), .feature_below(feature_belows[2026]), .scan_win_std_dev(scan_win_std_dev[2026]), .feature_accum(feature_accums[2026]));
  accum_calculator ac2027(.scan_win(scan_win2027), .rectangle1_x(rectangle1_xs[2027]), .rectangle1_y(rectangle1_ys[2027]), .rectangle1_width(rectangle1_widths[2027]), .rectangle1_height(rectangle1_heights[2027]), .rectangle1_weight(rectangle1_weights[2027]), .rectangle2_x(rectangle2_xs[2027]), .rectangle2_y(rectangle2_ys[2027]), .rectangle2_width(rectangle2_widths[2027]), .rectangle2_height(rectangle2_heights[2027]), .rectangle2_weight(rectangle2_weights[2027]), .rectangle3_x(rectangle3_xs[2027]), .rectangle3_y(rectangle3_ys[2027]), .rectangle3_width(rectangle3_widths[2027]), .rectangle3_height(rectangle3_heights[2027]), .rectangle3_weight(rectangle3_weights[2027]), .feature_threshold(feature_thresholds[2027]), .feature_above(feature_aboves[2027]), .feature_below(feature_belows[2027]), .scan_win_std_dev(scan_win_std_dev[2027]), .feature_accum(feature_accums[2027]));
  accum_calculator ac2028(.scan_win(scan_win2028), .rectangle1_x(rectangle1_xs[2028]), .rectangle1_y(rectangle1_ys[2028]), .rectangle1_width(rectangle1_widths[2028]), .rectangle1_height(rectangle1_heights[2028]), .rectangle1_weight(rectangle1_weights[2028]), .rectangle2_x(rectangle2_xs[2028]), .rectangle2_y(rectangle2_ys[2028]), .rectangle2_width(rectangle2_widths[2028]), .rectangle2_height(rectangle2_heights[2028]), .rectangle2_weight(rectangle2_weights[2028]), .rectangle3_x(rectangle3_xs[2028]), .rectangle3_y(rectangle3_ys[2028]), .rectangle3_width(rectangle3_widths[2028]), .rectangle3_height(rectangle3_heights[2028]), .rectangle3_weight(rectangle3_weights[2028]), .feature_threshold(feature_thresholds[2028]), .feature_above(feature_aboves[2028]), .feature_below(feature_belows[2028]), .scan_win_std_dev(scan_win_std_dev[2028]), .feature_accum(feature_accums[2028]));
  accum_calculator ac2029(.scan_win(scan_win2029), .rectangle1_x(rectangle1_xs[2029]), .rectangle1_y(rectangle1_ys[2029]), .rectangle1_width(rectangle1_widths[2029]), .rectangle1_height(rectangle1_heights[2029]), .rectangle1_weight(rectangle1_weights[2029]), .rectangle2_x(rectangle2_xs[2029]), .rectangle2_y(rectangle2_ys[2029]), .rectangle2_width(rectangle2_widths[2029]), .rectangle2_height(rectangle2_heights[2029]), .rectangle2_weight(rectangle2_weights[2029]), .rectangle3_x(rectangle3_xs[2029]), .rectangle3_y(rectangle3_ys[2029]), .rectangle3_width(rectangle3_widths[2029]), .rectangle3_height(rectangle3_heights[2029]), .rectangle3_weight(rectangle3_weights[2029]), .feature_threshold(feature_thresholds[2029]), .feature_above(feature_aboves[2029]), .feature_below(feature_belows[2029]), .scan_win_std_dev(scan_win_std_dev[2029]), .feature_accum(feature_accums[2029]));
  accum_calculator ac2030(.scan_win(scan_win2030), .rectangle1_x(rectangle1_xs[2030]), .rectangle1_y(rectangle1_ys[2030]), .rectangle1_width(rectangle1_widths[2030]), .rectangle1_height(rectangle1_heights[2030]), .rectangle1_weight(rectangle1_weights[2030]), .rectangle2_x(rectangle2_xs[2030]), .rectangle2_y(rectangle2_ys[2030]), .rectangle2_width(rectangle2_widths[2030]), .rectangle2_height(rectangle2_heights[2030]), .rectangle2_weight(rectangle2_weights[2030]), .rectangle3_x(rectangle3_xs[2030]), .rectangle3_y(rectangle3_ys[2030]), .rectangle3_width(rectangle3_widths[2030]), .rectangle3_height(rectangle3_heights[2030]), .rectangle3_weight(rectangle3_weights[2030]), .feature_threshold(feature_thresholds[2030]), .feature_above(feature_aboves[2030]), .feature_below(feature_belows[2030]), .scan_win_std_dev(scan_win_std_dev[2030]), .feature_accum(feature_accums[2030]));
  accum_calculator ac2031(.scan_win(scan_win2031), .rectangle1_x(rectangle1_xs[2031]), .rectangle1_y(rectangle1_ys[2031]), .rectangle1_width(rectangle1_widths[2031]), .rectangle1_height(rectangle1_heights[2031]), .rectangle1_weight(rectangle1_weights[2031]), .rectangle2_x(rectangle2_xs[2031]), .rectangle2_y(rectangle2_ys[2031]), .rectangle2_width(rectangle2_widths[2031]), .rectangle2_height(rectangle2_heights[2031]), .rectangle2_weight(rectangle2_weights[2031]), .rectangle3_x(rectangle3_xs[2031]), .rectangle3_y(rectangle3_ys[2031]), .rectangle3_width(rectangle3_widths[2031]), .rectangle3_height(rectangle3_heights[2031]), .rectangle3_weight(rectangle3_weights[2031]), .feature_threshold(feature_thresholds[2031]), .feature_above(feature_aboves[2031]), .feature_below(feature_belows[2031]), .scan_win_std_dev(scan_win_std_dev[2031]), .feature_accum(feature_accums[2031]));
  accum_calculator ac2032(.scan_win(scan_win2032), .rectangle1_x(rectangle1_xs[2032]), .rectangle1_y(rectangle1_ys[2032]), .rectangle1_width(rectangle1_widths[2032]), .rectangle1_height(rectangle1_heights[2032]), .rectangle1_weight(rectangle1_weights[2032]), .rectangle2_x(rectangle2_xs[2032]), .rectangle2_y(rectangle2_ys[2032]), .rectangle2_width(rectangle2_widths[2032]), .rectangle2_height(rectangle2_heights[2032]), .rectangle2_weight(rectangle2_weights[2032]), .rectangle3_x(rectangle3_xs[2032]), .rectangle3_y(rectangle3_ys[2032]), .rectangle3_width(rectangle3_widths[2032]), .rectangle3_height(rectangle3_heights[2032]), .rectangle3_weight(rectangle3_weights[2032]), .feature_threshold(feature_thresholds[2032]), .feature_above(feature_aboves[2032]), .feature_below(feature_belows[2032]), .scan_win_std_dev(scan_win_std_dev[2032]), .feature_accum(feature_accums[2032]));
  accum_calculator ac2033(.scan_win(scan_win2033), .rectangle1_x(rectangle1_xs[2033]), .rectangle1_y(rectangle1_ys[2033]), .rectangle1_width(rectangle1_widths[2033]), .rectangle1_height(rectangle1_heights[2033]), .rectangle1_weight(rectangle1_weights[2033]), .rectangle2_x(rectangle2_xs[2033]), .rectangle2_y(rectangle2_ys[2033]), .rectangle2_width(rectangle2_widths[2033]), .rectangle2_height(rectangle2_heights[2033]), .rectangle2_weight(rectangle2_weights[2033]), .rectangle3_x(rectangle3_xs[2033]), .rectangle3_y(rectangle3_ys[2033]), .rectangle3_width(rectangle3_widths[2033]), .rectangle3_height(rectangle3_heights[2033]), .rectangle3_weight(rectangle3_weights[2033]), .feature_threshold(feature_thresholds[2033]), .feature_above(feature_aboves[2033]), .feature_below(feature_belows[2033]), .scan_win_std_dev(scan_win_std_dev[2033]), .feature_accum(feature_accums[2033]));
  accum_calculator ac2034(.scan_win(scan_win2034), .rectangle1_x(rectangle1_xs[2034]), .rectangle1_y(rectangle1_ys[2034]), .rectangle1_width(rectangle1_widths[2034]), .rectangle1_height(rectangle1_heights[2034]), .rectangle1_weight(rectangle1_weights[2034]), .rectangle2_x(rectangle2_xs[2034]), .rectangle2_y(rectangle2_ys[2034]), .rectangle2_width(rectangle2_widths[2034]), .rectangle2_height(rectangle2_heights[2034]), .rectangle2_weight(rectangle2_weights[2034]), .rectangle3_x(rectangle3_xs[2034]), .rectangle3_y(rectangle3_ys[2034]), .rectangle3_width(rectangle3_widths[2034]), .rectangle3_height(rectangle3_heights[2034]), .rectangle3_weight(rectangle3_weights[2034]), .feature_threshold(feature_thresholds[2034]), .feature_above(feature_aboves[2034]), .feature_below(feature_belows[2034]), .scan_win_std_dev(scan_win_std_dev[2034]), .feature_accum(feature_accums[2034]));
  accum_calculator ac2035(.scan_win(scan_win2035), .rectangle1_x(rectangle1_xs[2035]), .rectangle1_y(rectangle1_ys[2035]), .rectangle1_width(rectangle1_widths[2035]), .rectangle1_height(rectangle1_heights[2035]), .rectangle1_weight(rectangle1_weights[2035]), .rectangle2_x(rectangle2_xs[2035]), .rectangle2_y(rectangle2_ys[2035]), .rectangle2_width(rectangle2_widths[2035]), .rectangle2_height(rectangle2_heights[2035]), .rectangle2_weight(rectangle2_weights[2035]), .rectangle3_x(rectangle3_xs[2035]), .rectangle3_y(rectangle3_ys[2035]), .rectangle3_width(rectangle3_widths[2035]), .rectangle3_height(rectangle3_heights[2035]), .rectangle3_weight(rectangle3_weights[2035]), .feature_threshold(feature_thresholds[2035]), .feature_above(feature_aboves[2035]), .feature_below(feature_belows[2035]), .scan_win_std_dev(scan_win_std_dev[2035]), .feature_accum(feature_accums[2035]));
  accum_calculator ac2036(.scan_win(scan_win2036), .rectangle1_x(rectangle1_xs[2036]), .rectangle1_y(rectangle1_ys[2036]), .rectangle1_width(rectangle1_widths[2036]), .rectangle1_height(rectangle1_heights[2036]), .rectangle1_weight(rectangle1_weights[2036]), .rectangle2_x(rectangle2_xs[2036]), .rectangle2_y(rectangle2_ys[2036]), .rectangle2_width(rectangle2_widths[2036]), .rectangle2_height(rectangle2_heights[2036]), .rectangle2_weight(rectangle2_weights[2036]), .rectangle3_x(rectangle3_xs[2036]), .rectangle3_y(rectangle3_ys[2036]), .rectangle3_width(rectangle3_widths[2036]), .rectangle3_height(rectangle3_heights[2036]), .rectangle3_weight(rectangle3_weights[2036]), .feature_threshold(feature_thresholds[2036]), .feature_above(feature_aboves[2036]), .feature_below(feature_belows[2036]), .scan_win_std_dev(scan_win_std_dev[2036]), .feature_accum(feature_accums[2036]));
  accum_calculator ac2037(.scan_win(scan_win2037), .rectangle1_x(rectangle1_xs[2037]), .rectangle1_y(rectangle1_ys[2037]), .rectangle1_width(rectangle1_widths[2037]), .rectangle1_height(rectangle1_heights[2037]), .rectangle1_weight(rectangle1_weights[2037]), .rectangle2_x(rectangle2_xs[2037]), .rectangle2_y(rectangle2_ys[2037]), .rectangle2_width(rectangle2_widths[2037]), .rectangle2_height(rectangle2_heights[2037]), .rectangle2_weight(rectangle2_weights[2037]), .rectangle3_x(rectangle3_xs[2037]), .rectangle3_y(rectangle3_ys[2037]), .rectangle3_width(rectangle3_widths[2037]), .rectangle3_height(rectangle3_heights[2037]), .rectangle3_weight(rectangle3_weights[2037]), .feature_threshold(feature_thresholds[2037]), .feature_above(feature_aboves[2037]), .feature_below(feature_belows[2037]), .scan_win_std_dev(scan_win_std_dev[2037]), .feature_accum(feature_accums[2037]));
  accum_calculator ac2038(.scan_win(scan_win2038), .rectangle1_x(rectangle1_xs[2038]), .rectangle1_y(rectangle1_ys[2038]), .rectangle1_width(rectangle1_widths[2038]), .rectangle1_height(rectangle1_heights[2038]), .rectangle1_weight(rectangle1_weights[2038]), .rectangle2_x(rectangle2_xs[2038]), .rectangle2_y(rectangle2_ys[2038]), .rectangle2_width(rectangle2_widths[2038]), .rectangle2_height(rectangle2_heights[2038]), .rectangle2_weight(rectangle2_weights[2038]), .rectangle3_x(rectangle3_xs[2038]), .rectangle3_y(rectangle3_ys[2038]), .rectangle3_width(rectangle3_widths[2038]), .rectangle3_height(rectangle3_heights[2038]), .rectangle3_weight(rectangle3_weights[2038]), .feature_threshold(feature_thresholds[2038]), .feature_above(feature_aboves[2038]), .feature_below(feature_belows[2038]), .scan_win_std_dev(scan_win_std_dev[2038]), .feature_accum(feature_accums[2038]));
  accum_calculator ac2039(.scan_win(scan_win2039), .rectangle1_x(rectangle1_xs[2039]), .rectangle1_y(rectangle1_ys[2039]), .rectangle1_width(rectangle1_widths[2039]), .rectangle1_height(rectangle1_heights[2039]), .rectangle1_weight(rectangle1_weights[2039]), .rectangle2_x(rectangle2_xs[2039]), .rectangle2_y(rectangle2_ys[2039]), .rectangle2_width(rectangle2_widths[2039]), .rectangle2_height(rectangle2_heights[2039]), .rectangle2_weight(rectangle2_weights[2039]), .rectangle3_x(rectangle3_xs[2039]), .rectangle3_y(rectangle3_ys[2039]), .rectangle3_width(rectangle3_widths[2039]), .rectangle3_height(rectangle3_heights[2039]), .rectangle3_weight(rectangle3_weights[2039]), .feature_threshold(feature_thresholds[2039]), .feature_above(feature_aboves[2039]), .feature_below(feature_belows[2039]), .scan_win_std_dev(scan_win_std_dev[2039]), .feature_accum(feature_accums[2039]));
  accum_calculator ac2040(.scan_win(scan_win2040), .rectangle1_x(rectangle1_xs[2040]), .rectangle1_y(rectangle1_ys[2040]), .rectangle1_width(rectangle1_widths[2040]), .rectangle1_height(rectangle1_heights[2040]), .rectangle1_weight(rectangle1_weights[2040]), .rectangle2_x(rectangle2_xs[2040]), .rectangle2_y(rectangle2_ys[2040]), .rectangle2_width(rectangle2_widths[2040]), .rectangle2_height(rectangle2_heights[2040]), .rectangle2_weight(rectangle2_weights[2040]), .rectangle3_x(rectangle3_xs[2040]), .rectangle3_y(rectangle3_ys[2040]), .rectangle3_width(rectangle3_widths[2040]), .rectangle3_height(rectangle3_heights[2040]), .rectangle3_weight(rectangle3_weights[2040]), .feature_threshold(feature_thresholds[2040]), .feature_above(feature_aboves[2040]), .feature_below(feature_belows[2040]), .scan_win_std_dev(scan_win_std_dev[2040]), .feature_accum(feature_accums[2040]));
  accum_calculator ac2041(.scan_win(scan_win2041), .rectangle1_x(rectangle1_xs[2041]), .rectangle1_y(rectangle1_ys[2041]), .rectangle1_width(rectangle1_widths[2041]), .rectangle1_height(rectangle1_heights[2041]), .rectangle1_weight(rectangle1_weights[2041]), .rectangle2_x(rectangle2_xs[2041]), .rectangle2_y(rectangle2_ys[2041]), .rectangle2_width(rectangle2_widths[2041]), .rectangle2_height(rectangle2_heights[2041]), .rectangle2_weight(rectangle2_weights[2041]), .rectangle3_x(rectangle3_xs[2041]), .rectangle3_y(rectangle3_ys[2041]), .rectangle3_width(rectangle3_widths[2041]), .rectangle3_height(rectangle3_heights[2041]), .rectangle3_weight(rectangle3_weights[2041]), .feature_threshold(feature_thresholds[2041]), .feature_above(feature_aboves[2041]), .feature_below(feature_belows[2041]), .scan_win_std_dev(scan_win_std_dev[2041]), .feature_accum(feature_accums[2041]));
  accum_calculator ac2042(.scan_win(scan_win2042), .rectangle1_x(rectangle1_xs[2042]), .rectangle1_y(rectangle1_ys[2042]), .rectangle1_width(rectangle1_widths[2042]), .rectangle1_height(rectangle1_heights[2042]), .rectangle1_weight(rectangle1_weights[2042]), .rectangle2_x(rectangle2_xs[2042]), .rectangle2_y(rectangle2_ys[2042]), .rectangle2_width(rectangle2_widths[2042]), .rectangle2_height(rectangle2_heights[2042]), .rectangle2_weight(rectangle2_weights[2042]), .rectangle3_x(rectangle3_xs[2042]), .rectangle3_y(rectangle3_ys[2042]), .rectangle3_width(rectangle3_widths[2042]), .rectangle3_height(rectangle3_heights[2042]), .rectangle3_weight(rectangle3_weights[2042]), .feature_threshold(feature_thresholds[2042]), .feature_above(feature_aboves[2042]), .feature_below(feature_belows[2042]), .scan_win_std_dev(scan_win_std_dev[2042]), .feature_accum(feature_accums[2042]));
  accum_calculator ac2043(.scan_win(scan_win2043), .rectangle1_x(rectangle1_xs[2043]), .rectangle1_y(rectangle1_ys[2043]), .rectangle1_width(rectangle1_widths[2043]), .rectangle1_height(rectangle1_heights[2043]), .rectangle1_weight(rectangle1_weights[2043]), .rectangle2_x(rectangle2_xs[2043]), .rectangle2_y(rectangle2_ys[2043]), .rectangle2_width(rectangle2_widths[2043]), .rectangle2_height(rectangle2_heights[2043]), .rectangle2_weight(rectangle2_weights[2043]), .rectangle3_x(rectangle3_xs[2043]), .rectangle3_y(rectangle3_ys[2043]), .rectangle3_width(rectangle3_widths[2043]), .rectangle3_height(rectangle3_heights[2043]), .rectangle3_weight(rectangle3_weights[2043]), .feature_threshold(feature_thresholds[2043]), .feature_above(feature_aboves[2043]), .feature_below(feature_belows[2043]), .scan_win_std_dev(scan_win_std_dev[2043]), .feature_accum(feature_accums[2043]));
  accum_calculator ac2044(.scan_win(scan_win2044), .rectangle1_x(rectangle1_xs[2044]), .rectangle1_y(rectangle1_ys[2044]), .rectangle1_width(rectangle1_widths[2044]), .rectangle1_height(rectangle1_heights[2044]), .rectangle1_weight(rectangle1_weights[2044]), .rectangle2_x(rectangle2_xs[2044]), .rectangle2_y(rectangle2_ys[2044]), .rectangle2_width(rectangle2_widths[2044]), .rectangle2_height(rectangle2_heights[2044]), .rectangle2_weight(rectangle2_weights[2044]), .rectangle3_x(rectangle3_xs[2044]), .rectangle3_y(rectangle3_ys[2044]), .rectangle3_width(rectangle3_widths[2044]), .rectangle3_height(rectangle3_heights[2044]), .rectangle3_weight(rectangle3_weights[2044]), .feature_threshold(feature_thresholds[2044]), .feature_above(feature_aboves[2044]), .feature_below(feature_belows[2044]), .scan_win_std_dev(scan_win_std_dev[2044]), .feature_accum(feature_accums[2044]));
  accum_calculator ac2045(.scan_win(scan_win2045), .rectangle1_x(rectangle1_xs[2045]), .rectangle1_y(rectangle1_ys[2045]), .rectangle1_width(rectangle1_widths[2045]), .rectangle1_height(rectangle1_heights[2045]), .rectangle1_weight(rectangle1_weights[2045]), .rectangle2_x(rectangle2_xs[2045]), .rectangle2_y(rectangle2_ys[2045]), .rectangle2_width(rectangle2_widths[2045]), .rectangle2_height(rectangle2_heights[2045]), .rectangle2_weight(rectangle2_weights[2045]), .rectangle3_x(rectangle3_xs[2045]), .rectangle3_y(rectangle3_ys[2045]), .rectangle3_width(rectangle3_widths[2045]), .rectangle3_height(rectangle3_heights[2045]), .rectangle3_weight(rectangle3_weights[2045]), .feature_threshold(feature_thresholds[2045]), .feature_above(feature_aboves[2045]), .feature_below(feature_belows[2045]), .scan_win_std_dev(scan_win_std_dev[2045]), .feature_accum(feature_accums[2045]));
  accum_calculator ac2046(.scan_win(scan_win2046), .rectangle1_x(rectangle1_xs[2046]), .rectangle1_y(rectangle1_ys[2046]), .rectangle1_width(rectangle1_widths[2046]), .rectangle1_height(rectangle1_heights[2046]), .rectangle1_weight(rectangle1_weights[2046]), .rectangle2_x(rectangle2_xs[2046]), .rectangle2_y(rectangle2_ys[2046]), .rectangle2_width(rectangle2_widths[2046]), .rectangle2_height(rectangle2_heights[2046]), .rectangle2_weight(rectangle2_weights[2046]), .rectangle3_x(rectangle3_xs[2046]), .rectangle3_y(rectangle3_ys[2046]), .rectangle3_width(rectangle3_widths[2046]), .rectangle3_height(rectangle3_heights[2046]), .rectangle3_weight(rectangle3_weights[2046]), .feature_threshold(feature_thresholds[2046]), .feature_above(feature_aboves[2046]), .feature_below(feature_belows[2046]), .scan_win_std_dev(scan_win_std_dev[2046]), .feature_accum(feature_accums[2046]));
  accum_calculator ac2047(.scan_win(scan_win2047), .rectangle1_x(rectangle1_xs[2047]), .rectangle1_y(rectangle1_ys[2047]), .rectangle1_width(rectangle1_widths[2047]), .rectangle1_height(rectangle1_heights[2047]), .rectangle1_weight(rectangle1_weights[2047]), .rectangle2_x(rectangle2_xs[2047]), .rectangle2_y(rectangle2_ys[2047]), .rectangle2_width(rectangle2_widths[2047]), .rectangle2_height(rectangle2_heights[2047]), .rectangle2_weight(rectangle2_weights[2047]), .rectangle3_x(rectangle3_xs[2047]), .rectangle3_y(rectangle3_ys[2047]), .rectangle3_width(rectangle3_widths[2047]), .rectangle3_height(rectangle3_heights[2047]), .rectangle3_weight(rectangle3_weights[2047]), .feature_threshold(feature_thresholds[2047]), .feature_above(feature_aboves[2047]), .feature_below(feature_belows[2047]), .scan_win_std_dev(scan_win_std_dev[2047]), .feature_accum(feature_accums[2047]));
  accum_calculator ac2048(.scan_win(scan_win2048), .rectangle1_x(rectangle1_xs[2048]), .rectangle1_y(rectangle1_ys[2048]), .rectangle1_width(rectangle1_widths[2048]), .rectangle1_height(rectangle1_heights[2048]), .rectangle1_weight(rectangle1_weights[2048]), .rectangle2_x(rectangle2_xs[2048]), .rectangle2_y(rectangle2_ys[2048]), .rectangle2_width(rectangle2_widths[2048]), .rectangle2_height(rectangle2_heights[2048]), .rectangle2_weight(rectangle2_weights[2048]), .rectangle3_x(rectangle3_xs[2048]), .rectangle3_y(rectangle3_ys[2048]), .rectangle3_width(rectangle3_widths[2048]), .rectangle3_height(rectangle3_heights[2048]), .rectangle3_weight(rectangle3_weights[2048]), .feature_threshold(feature_thresholds[2048]), .feature_above(feature_aboves[2048]), .feature_below(feature_belows[2048]), .scan_win_std_dev(scan_win_std_dev[2048]), .feature_accum(feature_accums[2048]));
  accum_calculator ac2049(.scan_win(scan_win2049), .rectangle1_x(rectangle1_xs[2049]), .rectangle1_y(rectangle1_ys[2049]), .rectangle1_width(rectangle1_widths[2049]), .rectangle1_height(rectangle1_heights[2049]), .rectangle1_weight(rectangle1_weights[2049]), .rectangle2_x(rectangle2_xs[2049]), .rectangle2_y(rectangle2_ys[2049]), .rectangle2_width(rectangle2_widths[2049]), .rectangle2_height(rectangle2_heights[2049]), .rectangle2_weight(rectangle2_weights[2049]), .rectangle3_x(rectangle3_xs[2049]), .rectangle3_y(rectangle3_ys[2049]), .rectangle3_width(rectangle3_widths[2049]), .rectangle3_height(rectangle3_heights[2049]), .rectangle3_weight(rectangle3_weights[2049]), .feature_threshold(feature_thresholds[2049]), .feature_above(feature_aboves[2049]), .feature_below(feature_belows[2049]), .scan_win_std_dev(scan_win_std_dev[2049]), .feature_accum(feature_accums[2049]));
  accum_calculator ac2050(.scan_win(scan_win2050), .rectangle1_x(rectangle1_xs[2050]), .rectangle1_y(rectangle1_ys[2050]), .rectangle1_width(rectangle1_widths[2050]), .rectangle1_height(rectangle1_heights[2050]), .rectangle1_weight(rectangle1_weights[2050]), .rectangle2_x(rectangle2_xs[2050]), .rectangle2_y(rectangle2_ys[2050]), .rectangle2_width(rectangle2_widths[2050]), .rectangle2_height(rectangle2_heights[2050]), .rectangle2_weight(rectangle2_weights[2050]), .rectangle3_x(rectangle3_xs[2050]), .rectangle3_y(rectangle3_ys[2050]), .rectangle3_width(rectangle3_widths[2050]), .rectangle3_height(rectangle3_heights[2050]), .rectangle3_weight(rectangle3_weights[2050]), .feature_threshold(feature_thresholds[2050]), .feature_above(feature_aboves[2050]), .feature_below(feature_belows[2050]), .scan_win_std_dev(scan_win_std_dev[2050]), .feature_accum(feature_accums[2050]));
  accum_calculator ac2051(.scan_win(scan_win2051), .rectangle1_x(rectangle1_xs[2051]), .rectangle1_y(rectangle1_ys[2051]), .rectangle1_width(rectangle1_widths[2051]), .rectangle1_height(rectangle1_heights[2051]), .rectangle1_weight(rectangle1_weights[2051]), .rectangle2_x(rectangle2_xs[2051]), .rectangle2_y(rectangle2_ys[2051]), .rectangle2_width(rectangle2_widths[2051]), .rectangle2_height(rectangle2_heights[2051]), .rectangle2_weight(rectangle2_weights[2051]), .rectangle3_x(rectangle3_xs[2051]), .rectangle3_y(rectangle3_ys[2051]), .rectangle3_width(rectangle3_widths[2051]), .rectangle3_height(rectangle3_heights[2051]), .rectangle3_weight(rectangle3_weights[2051]), .feature_threshold(feature_thresholds[2051]), .feature_above(feature_aboves[2051]), .feature_below(feature_belows[2051]), .scan_win_std_dev(scan_win_std_dev[2051]), .feature_accum(feature_accums[2051]));
  accum_calculator ac2052(.scan_win(scan_win2052), .rectangle1_x(rectangle1_xs[2052]), .rectangle1_y(rectangle1_ys[2052]), .rectangle1_width(rectangle1_widths[2052]), .rectangle1_height(rectangle1_heights[2052]), .rectangle1_weight(rectangle1_weights[2052]), .rectangle2_x(rectangle2_xs[2052]), .rectangle2_y(rectangle2_ys[2052]), .rectangle2_width(rectangle2_widths[2052]), .rectangle2_height(rectangle2_heights[2052]), .rectangle2_weight(rectangle2_weights[2052]), .rectangle3_x(rectangle3_xs[2052]), .rectangle3_y(rectangle3_ys[2052]), .rectangle3_width(rectangle3_widths[2052]), .rectangle3_height(rectangle3_heights[2052]), .rectangle3_weight(rectangle3_weights[2052]), .feature_threshold(feature_thresholds[2052]), .feature_above(feature_aboves[2052]), .feature_below(feature_belows[2052]), .scan_win_std_dev(scan_win_std_dev[2052]), .feature_accum(feature_accums[2052]));
  accum_calculator ac2053(.scan_win(scan_win2053), .rectangle1_x(rectangle1_xs[2053]), .rectangle1_y(rectangle1_ys[2053]), .rectangle1_width(rectangle1_widths[2053]), .rectangle1_height(rectangle1_heights[2053]), .rectangle1_weight(rectangle1_weights[2053]), .rectangle2_x(rectangle2_xs[2053]), .rectangle2_y(rectangle2_ys[2053]), .rectangle2_width(rectangle2_widths[2053]), .rectangle2_height(rectangle2_heights[2053]), .rectangle2_weight(rectangle2_weights[2053]), .rectangle3_x(rectangle3_xs[2053]), .rectangle3_y(rectangle3_ys[2053]), .rectangle3_width(rectangle3_widths[2053]), .rectangle3_height(rectangle3_heights[2053]), .rectangle3_weight(rectangle3_weights[2053]), .feature_threshold(feature_thresholds[2053]), .feature_above(feature_aboves[2053]), .feature_below(feature_belows[2053]), .scan_win_std_dev(scan_win_std_dev[2053]), .feature_accum(feature_accums[2053]));
  accum_calculator ac2054(.scan_win(scan_win2054), .rectangle1_x(rectangle1_xs[2054]), .rectangle1_y(rectangle1_ys[2054]), .rectangle1_width(rectangle1_widths[2054]), .rectangle1_height(rectangle1_heights[2054]), .rectangle1_weight(rectangle1_weights[2054]), .rectangle2_x(rectangle2_xs[2054]), .rectangle2_y(rectangle2_ys[2054]), .rectangle2_width(rectangle2_widths[2054]), .rectangle2_height(rectangle2_heights[2054]), .rectangle2_weight(rectangle2_weights[2054]), .rectangle3_x(rectangle3_xs[2054]), .rectangle3_y(rectangle3_ys[2054]), .rectangle3_width(rectangle3_widths[2054]), .rectangle3_height(rectangle3_heights[2054]), .rectangle3_weight(rectangle3_weights[2054]), .feature_threshold(feature_thresholds[2054]), .feature_above(feature_aboves[2054]), .feature_below(feature_belows[2054]), .scan_win_std_dev(scan_win_std_dev[2054]), .feature_accum(feature_accums[2054]));
  accum_calculator ac2055(.scan_win(scan_win2055), .rectangle1_x(rectangle1_xs[2055]), .rectangle1_y(rectangle1_ys[2055]), .rectangle1_width(rectangle1_widths[2055]), .rectangle1_height(rectangle1_heights[2055]), .rectangle1_weight(rectangle1_weights[2055]), .rectangle2_x(rectangle2_xs[2055]), .rectangle2_y(rectangle2_ys[2055]), .rectangle2_width(rectangle2_widths[2055]), .rectangle2_height(rectangle2_heights[2055]), .rectangle2_weight(rectangle2_weights[2055]), .rectangle3_x(rectangle3_xs[2055]), .rectangle3_y(rectangle3_ys[2055]), .rectangle3_width(rectangle3_widths[2055]), .rectangle3_height(rectangle3_heights[2055]), .rectangle3_weight(rectangle3_weights[2055]), .feature_threshold(feature_thresholds[2055]), .feature_above(feature_aboves[2055]), .feature_below(feature_belows[2055]), .scan_win_std_dev(scan_win_std_dev[2055]), .feature_accum(feature_accums[2055]));
  accum_calculator ac2056(.scan_win(scan_win2056), .rectangle1_x(rectangle1_xs[2056]), .rectangle1_y(rectangle1_ys[2056]), .rectangle1_width(rectangle1_widths[2056]), .rectangle1_height(rectangle1_heights[2056]), .rectangle1_weight(rectangle1_weights[2056]), .rectangle2_x(rectangle2_xs[2056]), .rectangle2_y(rectangle2_ys[2056]), .rectangle2_width(rectangle2_widths[2056]), .rectangle2_height(rectangle2_heights[2056]), .rectangle2_weight(rectangle2_weights[2056]), .rectangle3_x(rectangle3_xs[2056]), .rectangle3_y(rectangle3_ys[2056]), .rectangle3_width(rectangle3_widths[2056]), .rectangle3_height(rectangle3_heights[2056]), .rectangle3_weight(rectangle3_weights[2056]), .feature_threshold(feature_thresholds[2056]), .feature_above(feature_aboves[2056]), .feature_below(feature_belows[2056]), .scan_win_std_dev(scan_win_std_dev[2056]), .feature_accum(feature_accums[2056]));
  accum_calculator ac2057(.scan_win(scan_win2057), .rectangle1_x(rectangle1_xs[2057]), .rectangle1_y(rectangle1_ys[2057]), .rectangle1_width(rectangle1_widths[2057]), .rectangle1_height(rectangle1_heights[2057]), .rectangle1_weight(rectangle1_weights[2057]), .rectangle2_x(rectangle2_xs[2057]), .rectangle2_y(rectangle2_ys[2057]), .rectangle2_width(rectangle2_widths[2057]), .rectangle2_height(rectangle2_heights[2057]), .rectangle2_weight(rectangle2_weights[2057]), .rectangle3_x(rectangle3_xs[2057]), .rectangle3_y(rectangle3_ys[2057]), .rectangle3_width(rectangle3_widths[2057]), .rectangle3_height(rectangle3_heights[2057]), .rectangle3_weight(rectangle3_weights[2057]), .feature_threshold(feature_thresholds[2057]), .feature_above(feature_aboves[2057]), .feature_below(feature_belows[2057]), .scan_win_std_dev(scan_win_std_dev[2057]), .feature_accum(feature_accums[2057]));
  accum_calculator ac2058(.scan_win(scan_win2058), .rectangle1_x(rectangle1_xs[2058]), .rectangle1_y(rectangle1_ys[2058]), .rectangle1_width(rectangle1_widths[2058]), .rectangle1_height(rectangle1_heights[2058]), .rectangle1_weight(rectangle1_weights[2058]), .rectangle2_x(rectangle2_xs[2058]), .rectangle2_y(rectangle2_ys[2058]), .rectangle2_width(rectangle2_widths[2058]), .rectangle2_height(rectangle2_heights[2058]), .rectangle2_weight(rectangle2_weights[2058]), .rectangle3_x(rectangle3_xs[2058]), .rectangle3_y(rectangle3_ys[2058]), .rectangle3_width(rectangle3_widths[2058]), .rectangle3_height(rectangle3_heights[2058]), .rectangle3_weight(rectangle3_weights[2058]), .feature_threshold(feature_thresholds[2058]), .feature_above(feature_aboves[2058]), .feature_below(feature_belows[2058]), .scan_win_std_dev(scan_win_std_dev[2058]), .feature_accum(feature_accums[2058]));
  accum_calculator ac2059(.scan_win(scan_win2059), .rectangle1_x(rectangle1_xs[2059]), .rectangle1_y(rectangle1_ys[2059]), .rectangle1_width(rectangle1_widths[2059]), .rectangle1_height(rectangle1_heights[2059]), .rectangle1_weight(rectangle1_weights[2059]), .rectangle2_x(rectangle2_xs[2059]), .rectangle2_y(rectangle2_ys[2059]), .rectangle2_width(rectangle2_widths[2059]), .rectangle2_height(rectangle2_heights[2059]), .rectangle2_weight(rectangle2_weights[2059]), .rectangle3_x(rectangle3_xs[2059]), .rectangle3_y(rectangle3_ys[2059]), .rectangle3_width(rectangle3_widths[2059]), .rectangle3_height(rectangle3_heights[2059]), .rectangle3_weight(rectangle3_weights[2059]), .feature_threshold(feature_thresholds[2059]), .feature_above(feature_aboves[2059]), .feature_below(feature_belows[2059]), .scan_win_std_dev(scan_win_std_dev[2059]), .feature_accum(feature_accums[2059]));
  accum_calculator ac2060(.scan_win(scan_win2060), .rectangle1_x(rectangle1_xs[2060]), .rectangle1_y(rectangle1_ys[2060]), .rectangle1_width(rectangle1_widths[2060]), .rectangle1_height(rectangle1_heights[2060]), .rectangle1_weight(rectangle1_weights[2060]), .rectangle2_x(rectangle2_xs[2060]), .rectangle2_y(rectangle2_ys[2060]), .rectangle2_width(rectangle2_widths[2060]), .rectangle2_height(rectangle2_heights[2060]), .rectangle2_weight(rectangle2_weights[2060]), .rectangle3_x(rectangle3_xs[2060]), .rectangle3_y(rectangle3_ys[2060]), .rectangle3_width(rectangle3_widths[2060]), .rectangle3_height(rectangle3_heights[2060]), .rectangle3_weight(rectangle3_weights[2060]), .feature_threshold(feature_thresholds[2060]), .feature_above(feature_aboves[2060]), .feature_below(feature_belows[2060]), .scan_win_std_dev(scan_win_std_dev[2060]), .feature_accum(feature_accums[2060]));
  accum_calculator ac2061(.scan_win(scan_win2061), .rectangle1_x(rectangle1_xs[2061]), .rectangle1_y(rectangle1_ys[2061]), .rectangle1_width(rectangle1_widths[2061]), .rectangle1_height(rectangle1_heights[2061]), .rectangle1_weight(rectangle1_weights[2061]), .rectangle2_x(rectangle2_xs[2061]), .rectangle2_y(rectangle2_ys[2061]), .rectangle2_width(rectangle2_widths[2061]), .rectangle2_height(rectangle2_heights[2061]), .rectangle2_weight(rectangle2_weights[2061]), .rectangle3_x(rectangle3_xs[2061]), .rectangle3_y(rectangle3_ys[2061]), .rectangle3_width(rectangle3_widths[2061]), .rectangle3_height(rectangle3_heights[2061]), .rectangle3_weight(rectangle3_weights[2061]), .feature_threshold(feature_thresholds[2061]), .feature_above(feature_aboves[2061]), .feature_below(feature_belows[2061]), .scan_win_std_dev(scan_win_std_dev[2061]), .feature_accum(feature_accums[2061]));
  accum_calculator ac2062(.scan_win(scan_win2062), .rectangle1_x(rectangle1_xs[2062]), .rectangle1_y(rectangle1_ys[2062]), .rectangle1_width(rectangle1_widths[2062]), .rectangle1_height(rectangle1_heights[2062]), .rectangle1_weight(rectangle1_weights[2062]), .rectangle2_x(rectangle2_xs[2062]), .rectangle2_y(rectangle2_ys[2062]), .rectangle2_width(rectangle2_widths[2062]), .rectangle2_height(rectangle2_heights[2062]), .rectangle2_weight(rectangle2_weights[2062]), .rectangle3_x(rectangle3_xs[2062]), .rectangle3_y(rectangle3_ys[2062]), .rectangle3_width(rectangle3_widths[2062]), .rectangle3_height(rectangle3_heights[2062]), .rectangle3_weight(rectangle3_weights[2062]), .feature_threshold(feature_thresholds[2062]), .feature_above(feature_aboves[2062]), .feature_below(feature_belows[2062]), .scan_win_std_dev(scan_win_std_dev[2062]), .feature_accum(feature_accums[2062]));
  accum_calculator ac2063(.scan_win(scan_win2063), .rectangle1_x(rectangle1_xs[2063]), .rectangle1_y(rectangle1_ys[2063]), .rectangle1_width(rectangle1_widths[2063]), .rectangle1_height(rectangle1_heights[2063]), .rectangle1_weight(rectangle1_weights[2063]), .rectangle2_x(rectangle2_xs[2063]), .rectangle2_y(rectangle2_ys[2063]), .rectangle2_width(rectangle2_widths[2063]), .rectangle2_height(rectangle2_heights[2063]), .rectangle2_weight(rectangle2_weights[2063]), .rectangle3_x(rectangle3_xs[2063]), .rectangle3_y(rectangle3_ys[2063]), .rectangle3_width(rectangle3_widths[2063]), .rectangle3_height(rectangle3_heights[2063]), .rectangle3_weight(rectangle3_weights[2063]), .feature_threshold(feature_thresholds[2063]), .feature_above(feature_aboves[2063]), .feature_below(feature_belows[2063]), .scan_win_std_dev(scan_win_std_dev[2063]), .feature_accum(feature_accums[2063]));
  accum_calculator ac2064(.scan_win(scan_win2064), .rectangle1_x(rectangle1_xs[2064]), .rectangle1_y(rectangle1_ys[2064]), .rectangle1_width(rectangle1_widths[2064]), .rectangle1_height(rectangle1_heights[2064]), .rectangle1_weight(rectangle1_weights[2064]), .rectangle2_x(rectangle2_xs[2064]), .rectangle2_y(rectangle2_ys[2064]), .rectangle2_width(rectangle2_widths[2064]), .rectangle2_height(rectangle2_heights[2064]), .rectangle2_weight(rectangle2_weights[2064]), .rectangle3_x(rectangle3_xs[2064]), .rectangle3_y(rectangle3_ys[2064]), .rectangle3_width(rectangle3_widths[2064]), .rectangle3_height(rectangle3_heights[2064]), .rectangle3_weight(rectangle3_weights[2064]), .feature_threshold(feature_thresholds[2064]), .feature_above(feature_aboves[2064]), .feature_below(feature_belows[2064]), .scan_win_std_dev(scan_win_std_dev[2064]), .feature_accum(feature_accums[2064]));
  accum_calculator ac2065(.scan_win(scan_win2065), .rectangle1_x(rectangle1_xs[2065]), .rectangle1_y(rectangle1_ys[2065]), .rectangle1_width(rectangle1_widths[2065]), .rectangle1_height(rectangle1_heights[2065]), .rectangle1_weight(rectangle1_weights[2065]), .rectangle2_x(rectangle2_xs[2065]), .rectangle2_y(rectangle2_ys[2065]), .rectangle2_width(rectangle2_widths[2065]), .rectangle2_height(rectangle2_heights[2065]), .rectangle2_weight(rectangle2_weights[2065]), .rectangle3_x(rectangle3_xs[2065]), .rectangle3_y(rectangle3_ys[2065]), .rectangle3_width(rectangle3_widths[2065]), .rectangle3_height(rectangle3_heights[2065]), .rectangle3_weight(rectangle3_weights[2065]), .feature_threshold(feature_thresholds[2065]), .feature_above(feature_aboves[2065]), .feature_below(feature_belows[2065]), .scan_win_std_dev(scan_win_std_dev[2065]), .feature_accum(feature_accums[2065]));
  accum_calculator ac2066(.scan_win(scan_win2066), .rectangle1_x(rectangle1_xs[2066]), .rectangle1_y(rectangle1_ys[2066]), .rectangle1_width(rectangle1_widths[2066]), .rectangle1_height(rectangle1_heights[2066]), .rectangle1_weight(rectangle1_weights[2066]), .rectangle2_x(rectangle2_xs[2066]), .rectangle2_y(rectangle2_ys[2066]), .rectangle2_width(rectangle2_widths[2066]), .rectangle2_height(rectangle2_heights[2066]), .rectangle2_weight(rectangle2_weights[2066]), .rectangle3_x(rectangle3_xs[2066]), .rectangle3_y(rectangle3_ys[2066]), .rectangle3_width(rectangle3_widths[2066]), .rectangle3_height(rectangle3_heights[2066]), .rectangle3_weight(rectangle3_weights[2066]), .feature_threshold(feature_thresholds[2066]), .feature_above(feature_aboves[2066]), .feature_below(feature_belows[2066]), .scan_win_std_dev(scan_win_std_dev[2066]), .feature_accum(feature_accums[2066]));
  accum_calculator ac2067(.scan_win(scan_win2067), .rectangle1_x(rectangle1_xs[2067]), .rectangle1_y(rectangle1_ys[2067]), .rectangle1_width(rectangle1_widths[2067]), .rectangle1_height(rectangle1_heights[2067]), .rectangle1_weight(rectangle1_weights[2067]), .rectangle2_x(rectangle2_xs[2067]), .rectangle2_y(rectangle2_ys[2067]), .rectangle2_width(rectangle2_widths[2067]), .rectangle2_height(rectangle2_heights[2067]), .rectangle2_weight(rectangle2_weights[2067]), .rectangle3_x(rectangle3_xs[2067]), .rectangle3_y(rectangle3_ys[2067]), .rectangle3_width(rectangle3_widths[2067]), .rectangle3_height(rectangle3_heights[2067]), .rectangle3_weight(rectangle3_weights[2067]), .feature_threshold(feature_thresholds[2067]), .feature_above(feature_aboves[2067]), .feature_below(feature_belows[2067]), .scan_win_std_dev(scan_win_std_dev[2067]), .feature_accum(feature_accums[2067]));
  accum_calculator ac2068(.scan_win(scan_win2068), .rectangle1_x(rectangle1_xs[2068]), .rectangle1_y(rectangle1_ys[2068]), .rectangle1_width(rectangle1_widths[2068]), .rectangle1_height(rectangle1_heights[2068]), .rectangle1_weight(rectangle1_weights[2068]), .rectangle2_x(rectangle2_xs[2068]), .rectangle2_y(rectangle2_ys[2068]), .rectangle2_width(rectangle2_widths[2068]), .rectangle2_height(rectangle2_heights[2068]), .rectangle2_weight(rectangle2_weights[2068]), .rectangle3_x(rectangle3_xs[2068]), .rectangle3_y(rectangle3_ys[2068]), .rectangle3_width(rectangle3_widths[2068]), .rectangle3_height(rectangle3_heights[2068]), .rectangle3_weight(rectangle3_weights[2068]), .feature_threshold(feature_thresholds[2068]), .feature_above(feature_aboves[2068]), .feature_below(feature_belows[2068]), .scan_win_std_dev(scan_win_std_dev[2068]), .feature_accum(feature_accums[2068]));
  accum_calculator ac2069(.scan_win(scan_win2069), .rectangle1_x(rectangle1_xs[2069]), .rectangle1_y(rectangle1_ys[2069]), .rectangle1_width(rectangle1_widths[2069]), .rectangle1_height(rectangle1_heights[2069]), .rectangle1_weight(rectangle1_weights[2069]), .rectangle2_x(rectangle2_xs[2069]), .rectangle2_y(rectangle2_ys[2069]), .rectangle2_width(rectangle2_widths[2069]), .rectangle2_height(rectangle2_heights[2069]), .rectangle2_weight(rectangle2_weights[2069]), .rectangle3_x(rectangle3_xs[2069]), .rectangle3_y(rectangle3_ys[2069]), .rectangle3_width(rectangle3_widths[2069]), .rectangle3_height(rectangle3_heights[2069]), .rectangle3_weight(rectangle3_weights[2069]), .feature_threshold(feature_thresholds[2069]), .feature_above(feature_aboves[2069]), .feature_below(feature_belows[2069]), .scan_win_std_dev(scan_win_std_dev[2069]), .feature_accum(feature_accums[2069]));
  accum_calculator ac2070(.scan_win(scan_win2070), .rectangle1_x(rectangle1_xs[2070]), .rectangle1_y(rectangle1_ys[2070]), .rectangle1_width(rectangle1_widths[2070]), .rectangle1_height(rectangle1_heights[2070]), .rectangle1_weight(rectangle1_weights[2070]), .rectangle2_x(rectangle2_xs[2070]), .rectangle2_y(rectangle2_ys[2070]), .rectangle2_width(rectangle2_widths[2070]), .rectangle2_height(rectangle2_heights[2070]), .rectangle2_weight(rectangle2_weights[2070]), .rectangle3_x(rectangle3_xs[2070]), .rectangle3_y(rectangle3_ys[2070]), .rectangle3_width(rectangle3_widths[2070]), .rectangle3_height(rectangle3_heights[2070]), .rectangle3_weight(rectangle3_weights[2070]), .feature_threshold(feature_thresholds[2070]), .feature_above(feature_aboves[2070]), .feature_below(feature_belows[2070]), .scan_win_std_dev(scan_win_std_dev[2070]), .feature_accum(feature_accums[2070]));
  accum_calculator ac2071(.scan_win(scan_win2071), .rectangle1_x(rectangle1_xs[2071]), .rectangle1_y(rectangle1_ys[2071]), .rectangle1_width(rectangle1_widths[2071]), .rectangle1_height(rectangle1_heights[2071]), .rectangle1_weight(rectangle1_weights[2071]), .rectangle2_x(rectangle2_xs[2071]), .rectangle2_y(rectangle2_ys[2071]), .rectangle2_width(rectangle2_widths[2071]), .rectangle2_height(rectangle2_heights[2071]), .rectangle2_weight(rectangle2_weights[2071]), .rectangle3_x(rectangle3_xs[2071]), .rectangle3_y(rectangle3_ys[2071]), .rectangle3_width(rectangle3_widths[2071]), .rectangle3_height(rectangle3_heights[2071]), .rectangle3_weight(rectangle3_weights[2071]), .feature_threshold(feature_thresholds[2071]), .feature_above(feature_aboves[2071]), .feature_below(feature_belows[2071]), .scan_win_std_dev(scan_win_std_dev[2071]), .feature_accum(feature_accums[2071]));
  accum_calculator ac2072(.scan_win(scan_win2072), .rectangle1_x(rectangle1_xs[2072]), .rectangle1_y(rectangle1_ys[2072]), .rectangle1_width(rectangle1_widths[2072]), .rectangle1_height(rectangle1_heights[2072]), .rectangle1_weight(rectangle1_weights[2072]), .rectangle2_x(rectangle2_xs[2072]), .rectangle2_y(rectangle2_ys[2072]), .rectangle2_width(rectangle2_widths[2072]), .rectangle2_height(rectangle2_heights[2072]), .rectangle2_weight(rectangle2_weights[2072]), .rectangle3_x(rectangle3_xs[2072]), .rectangle3_y(rectangle3_ys[2072]), .rectangle3_width(rectangle3_widths[2072]), .rectangle3_height(rectangle3_heights[2072]), .rectangle3_weight(rectangle3_weights[2072]), .feature_threshold(feature_thresholds[2072]), .feature_above(feature_aboves[2072]), .feature_below(feature_belows[2072]), .scan_win_std_dev(scan_win_std_dev[2072]), .feature_accum(feature_accums[2072]));
  accum_calculator ac2073(.scan_win(scan_win2073), .rectangle1_x(rectangle1_xs[2073]), .rectangle1_y(rectangle1_ys[2073]), .rectangle1_width(rectangle1_widths[2073]), .rectangle1_height(rectangle1_heights[2073]), .rectangle1_weight(rectangle1_weights[2073]), .rectangle2_x(rectangle2_xs[2073]), .rectangle2_y(rectangle2_ys[2073]), .rectangle2_width(rectangle2_widths[2073]), .rectangle2_height(rectangle2_heights[2073]), .rectangle2_weight(rectangle2_weights[2073]), .rectangle3_x(rectangle3_xs[2073]), .rectangle3_y(rectangle3_ys[2073]), .rectangle3_width(rectangle3_widths[2073]), .rectangle3_height(rectangle3_heights[2073]), .rectangle3_weight(rectangle3_weights[2073]), .feature_threshold(feature_thresholds[2073]), .feature_above(feature_aboves[2073]), .feature_below(feature_belows[2073]), .scan_win_std_dev(scan_win_std_dev[2073]), .feature_accum(feature_accums[2073]));
  accum_calculator ac2074(.scan_win(scan_win2074), .rectangle1_x(rectangle1_xs[2074]), .rectangle1_y(rectangle1_ys[2074]), .rectangle1_width(rectangle1_widths[2074]), .rectangle1_height(rectangle1_heights[2074]), .rectangle1_weight(rectangle1_weights[2074]), .rectangle2_x(rectangle2_xs[2074]), .rectangle2_y(rectangle2_ys[2074]), .rectangle2_width(rectangle2_widths[2074]), .rectangle2_height(rectangle2_heights[2074]), .rectangle2_weight(rectangle2_weights[2074]), .rectangle3_x(rectangle3_xs[2074]), .rectangle3_y(rectangle3_ys[2074]), .rectangle3_width(rectangle3_widths[2074]), .rectangle3_height(rectangle3_heights[2074]), .rectangle3_weight(rectangle3_weights[2074]), .feature_threshold(feature_thresholds[2074]), .feature_above(feature_aboves[2074]), .feature_below(feature_belows[2074]), .scan_win_std_dev(scan_win_std_dev[2074]), .feature_accum(feature_accums[2074]));
  accum_calculator ac2075(.scan_win(scan_win2075), .rectangle1_x(rectangle1_xs[2075]), .rectangle1_y(rectangle1_ys[2075]), .rectangle1_width(rectangle1_widths[2075]), .rectangle1_height(rectangle1_heights[2075]), .rectangle1_weight(rectangle1_weights[2075]), .rectangle2_x(rectangle2_xs[2075]), .rectangle2_y(rectangle2_ys[2075]), .rectangle2_width(rectangle2_widths[2075]), .rectangle2_height(rectangle2_heights[2075]), .rectangle2_weight(rectangle2_weights[2075]), .rectangle3_x(rectangle3_xs[2075]), .rectangle3_y(rectangle3_ys[2075]), .rectangle3_width(rectangle3_widths[2075]), .rectangle3_height(rectangle3_heights[2075]), .rectangle3_weight(rectangle3_weights[2075]), .feature_threshold(feature_thresholds[2075]), .feature_above(feature_aboves[2075]), .feature_below(feature_belows[2075]), .scan_win_std_dev(scan_win_std_dev[2075]), .feature_accum(feature_accums[2075]));
  accum_calculator ac2076(.scan_win(scan_win2076), .rectangle1_x(rectangle1_xs[2076]), .rectangle1_y(rectangle1_ys[2076]), .rectangle1_width(rectangle1_widths[2076]), .rectangle1_height(rectangle1_heights[2076]), .rectangle1_weight(rectangle1_weights[2076]), .rectangle2_x(rectangle2_xs[2076]), .rectangle2_y(rectangle2_ys[2076]), .rectangle2_width(rectangle2_widths[2076]), .rectangle2_height(rectangle2_heights[2076]), .rectangle2_weight(rectangle2_weights[2076]), .rectangle3_x(rectangle3_xs[2076]), .rectangle3_y(rectangle3_ys[2076]), .rectangle3_width(rectangle3_widths[2076]), .rectangle3_height(rectangle3_heights[2076]), .rectangle3_weight(rectangle3_weights[2076]), .feature_threshold(feature_thresholds[2076]), .feature_above(feature_aboves[2076]), .feature_below(feature_belows[2076]), .scan_win_std_dev(scan_win_std_dev[2076]), .feature_accum(feature_accums[2076]));
  accum_calculator ac2077(.scan_win(scan_win2077), .rectangle1_x(rectangle1_xs[2077]), .rectangle1_y(rectangle1_ys[2077]), .rectangle1_width(rectangle1_widths[2077]), .rectangle1_height(rectangle1_heights[2077]), .rectangle1_weight(rectangle1_weights[2077]), .rectangle2_x(rectangle2_xs[2077]), .rectangle2_y(rectangle2_ys[2077]), .rectangle2_width(rectangle2_widths[2077]), .rectangle2_height(rectangle2_heights[2077]), .rectangle2_weight(rectangle2_weights[2077]), .rectangle3_x(rectangle3_xs[2077]), .rectangle3_y(rectangle3_ys[2077]), .rectangle3_width(rectangle3_widths[2077]), .rectangle3_height(rectangle3_heights[2077]), .rectangle3_weight(rectangle3_weights[2077]), .feature_threshold(feature_thresholds[2077]), .feature_above(feature_aboves[2077]), .feature_below(feature_belows[2077]), .scan_win_std_dev(scan_win_std_dev[2077]), .feature_accum(feature_accums[2077]));
  accum_calculator ac2078(.scan_win(scan_win2078), .rectangle1_x(rectangle1_xs[2078]), .rectangle1_y(rectangle1_ys[2078]), .rectangle1_width(rectangle1_widths[2078]), .rectangle1_height(rectangle1_heights[2078]), .rectangle1_weight(rectangle1_weights[2078]), .rectangle2_x(rectangle2_xs[2078]), .rectangle2_y(rectangle2_ys[2078]), .rectangle2_width(rectangle2_widths[2078]), .rectangle2_height(rectangle2_heights[2078]), .rectangle2_weight(rectangle2_weights[2078]), .rectangle3_x(rectangle3_xs[2078]), .rectangle3_y(rectangle3_ys[2078]), .rectangle3_width(rectangle3_widths[2078]), .rectangle3_height(rectangle3_heights[2078]), .rectangle3_weight(rectangle3_weights[2078]), .feature_threshold(feature_thresholds[2078]), .feature_above(feature_aboves[2078]), .feature_below(feature_belows[2078]), .scan_win_std_dev(scan_win_std_dev[2078]), .feature_accum(feature_accums[2078]));
  accum_calculator ac2079(.scan_win(scan_win2079), .rectangle1_x(rectangle1_xs[2079]), .rectangle1_y(rectangle1_ys[2079]), .rectangle1_width(rectangle1_widths[2079]), .rectangle1_height(rectangle1_heights[2079]), .rectangle1_weight(rectangle1_weights[2079]), .rectangle2_x(rectangle2_xs[2079]), .rectangle2_y(rectangle2_ys[2079]), .rectangle2_width(rectangle2_widths[2079]), .rectangle2_height(rectangle2_heights[2079]), .rectangle2_weight(rectangle2_weights[2079]), .rectangle3_x(rectangle3_xs[2079]), .rectangle3_y(rectangle3_ys[2079]), .rectangle3_width(rectangle3_widths[2079]), .rectangle3_height(rectangle3_heights[2079]), .rectangle3_weight(rectangle3_weights[2079]), .feature_threshold(feature_thresholds[2079]), .feature_above(feature_aboves[2079]), .feature_below(feature_belows[2079]), .scan_win_std_dev(scan_win_std_dev[2079]), .feature_accum(feature_accums[2079]));
  accum_calculator ac2080(.scan_win(scan_win2080), .rectangle1_x(rectangle1_xs[2080]), .rectangle1_y(rectangle1_ys[2080]), .rectangle1_width(rectangle1_widths[2080]), .rectangle1_height(rectangle1_heights[2080]), .rectangle1_weight(rectangle1_weights[2080]), .rectangle2_x(rectangle2_xs[2080]), .rectangle2_y(rectangle2_ys[2080]), .rectangle2_width(rectangle2_widths[2080]), .rectangle2_height(rectangle2_heights[2080]), .rectangle2_weight(rectangle2_weights[2080]), .rectangle3_x(rectangle3_xs[2080]), .rectangle3_y(rectangle3_ys[2080]), .rectangle3_width(rectangle3_widths[2080]), .rectangle3_height(rectangle3_heights[2080]), .rectangle3_weight(rectangle3_weights[2080]), .feature_threshold(feature_thresholds[2080]), .feature_above(feature_aboves[2080]), .feature_below(feature_belows[2080]), .scan_win_std_dev(scan_win_std_dev[2080]), .feature_accum(feature_accums[2080]));
  accum_calculator ac2081(.scan_win(scan_win2081), .rectangle1_x(rectangle1_xs[2081]), .rectangle1_y(rectangle1_ys[2081]), .rectangle1_width(rectangle1_widths[2081]), .rectangle1_height(rectangle1_heights[2081]), .rectangle1_weight(rectangle1_weights[2081]), .rectangle2_x(rectangle2_xs[2081]), .rectangle2_y(rectangle2_ys[2081]), .rectangle2_width(rectangle2_widths[2081]), .rectangle2_height(rectangle2_heights[2081]), .rectangle2_weight(rectangle2_weights[2081]), .rectangle3_x(rectangle3_xs[2081]), .rectangle3_y(rectangle3_ys[2081]), .rectangle3_width(rectangle3_widths[2081]), .rectangle3_height(rectangle3_heights[2081]), .rectangle3_weight(rectangle3_weights[2081]), .feature_threshold(feature_thresholds[2081]), .feature_above(feature_aboves[2081]), .feature_below(feature_belows[2081]), .scan_win_std_dev(scan_win_std_dev[2081]), .feature_accum(feature_accums[2081]));
  accum_calculator ac2082(.scan_win(scan_win2082), .rectangle1_x(rectangle1_xs[2082]), .rectangle1_y(rectangle1_ys[2082]), .rectangle1_width(rectangle1_widths[2082]), .rectangle1_height(rectangle1_heights[2082]), .rectangle1_weight(rectangle1_weights[2082]), .rectangle2_x(rectangle2_xs[2082]), .rectangle2_y(rectangle2_ys[2082]), .rectangle2_width(rectangle2_widths[2082]), .rectangle2_height(rectangle2_heights[2082]), .rectangle2_weight(rectangle2_weights[2082]), .rectangle3_x(rectangle3_xs[2082]), .rectangle3_y(rectangle3_ys[2082]), .rectangle3_width(rectangle3_widths[2082]), .rectangle3_height(rectangle3_heights[2082]), .rectangle3_weight(rectangle3_weights[2082]), .feature_threshold(feature_thresholds[2082]), .feature_above(feature_aboves[2082]), .feature_below(feature_belows[2082]), .scan_win_std_dev(scan_win_std_dev[2082]), .feature_accum(feature_accums[2082]));
  accum_calculator ac2083(.scan_win(scan_win2083), .rectangle1_x(rectangle1_xs[2083]), .rectangle1_y(rectangle1_ys[2083]), .rectangle1_width(rectangle1_widths[2083]), .rectangle1_height(rectangle1_heights[2083]), .rectangle1_weight(rectangle1_weights[2083]), .rectangle2_x(rectangle2_xs[2083]), .rectangle2_y(rectangle2_ys[2083]), .rectangle2_width(rectangle2_widths[2083]), .rectangle2_height(rectangle2_heights[2083]), .rectangle2_weight(rectangle2_weights[2083]), .rectangle3_x(rectangle3_xs[2083]), .rectangle3_y(rectangle3_ys[2083]), .rectangle3_width(rectangle3_widths[2083]), .rectangle3_height(rectangle3_heights[2083]), .rectangle3_weight(rectangle3_weights[2083]), .feature_threshold(feature_thresholds[2083]), .feature_above(feature_aboves[2083]), .feature_below(feature_belows[2083]), .scan_win_std_dev(scan_win_std_dev[2083]), .feature_accum(feature_accums[2083]));
  accum_calculator ac2084(.scan_win(scan_win2084), .rectangle1_x(rectangle1_xs[2084]), .rectangle1_y(rectangle1_ys[2084]), .rectangle1_width(rectangle1_widths[2084]), .rectangle1_height(rectangle1_heights[2084]), .rectangle1_weight(rectangle1_weights[2084]), .rectangle2_x(rectangle2_xs[2084]), .rectangle2_y(rectangle2_ys[2084]), .rectangle2_width(rectangle2_widths[2084]), .rectangle2_height(rectangle2_heights[2084]), .rectangle2_weight(rectangle2_weights[2084]), .rectangle3_x(rectangle3_xs[2084]), .rectangle3_y(rectangle3_ys[2084]), .rectangle3_width(rectangle3_widths[2084]), .rectangle3_height(rectangle3_heights[2084]), .rectangle3_weight(rectangle3_weights[2084]), .feature_threshold(feature_thresholds[2084]), .feature_above(feature_aboves[2084]), .feature_below(feature_belows[2084]), .scan_win_std_dev(scan_win_std_dev[2084]), .feature_accum(feature_accums[2084]));
  accum_calculator ac2085(.scan_win(scan_win2085), .rectangle1_x(rectangle1_xs[2085]), .rectangle1_y(rectangle1_ys[2085]), .rectangle1_width(rectangle1_widths[2085]), .rectangle1_height(rectangle1_heights[2085]), .rectangle1_weight(rectangle1_weights[2085]), .rectangle2_x(rectangle2_xs[2085]), .rectangle2_y(rectangle2_ys[2085]), .rectangle2_width(rectangle2_widths[2085]), .rectangle2_height(rectangle2_heights[2085]), .rectangle2_weight(rectangle2_weights[2085]), .rectangle3_x(rectangle3_xs[2085]), .rectangle3_y(rectangle3_ys[2085]), .rectangle3_width(rectangle3_widths[2085]), .rectangle3_height(rectangle3_heights[2085]), .rectangle3_weight(rectangle3_weights[2085]), .feature_threshold(feature_thresholds[2085]), .feature_above(feature_aboves[2085]), .feature_below(feature_belows[2085]), .scan_win_std_dev(scan_win_std_dev[2085]), .feature_accum(feature_accums[2085]));
  accum_calculator ac2086(.scan_win(scan_win2086), .rectangle1_x(rectangle1_xs[2086]), .rectangle1_y(rectangle1_ys[2086]), .rectangle1_width(rectangle1_widths[2086]), .rectangle1_height(rectangle1_heights[2086]), .rectangle1_weight(rectangle1_weights[2086]), .rectangle2_x(rectangle2_xs[2086]), .rectangle2_y(rectangle2_ys[2086]), .rectangle2_width(rectangle2_widths[2086]), .rectangle2_height(rectangle2_heights[2086]), .rectangle2_weight(rectangle2_weights[2086]), .rectangle3_x(rectangle3_xs[2086]), .rectangle3_y(rectangle3_ys[2086]), .rectangle3_width(rectangle3_widths[2086]), .rectangle3_height(rectangle3_heights[2086]), .rectangle3_weight(rectangle3_weights[2086]), .feature_threshold(feature_thresholds[2086]), .feature_above(feature_aboves[2086]), .feature_below(feature_belows[2086]), .scan_win_std_dev(scan_win_std_dev[2086]), .feature_accum(feature_accums[2086]));
  accum_calculator ac2087(.scan_win(scan_win2087), .rectangle1_x(rectangle1_xs[2087]), .rectangle1_y(rectangle1_ys[2087]), .rectangle1_width(rectangle1_widths[2087]), .rectangle1_height(rectangle1_heights[2087]), .rectangle1_weight(rectangle1_weights[2087]), .rectangle2_x(rectangle2_xs[2087]), .rectangle2_y(rectangle2_ys[2087]), .rectangle2_width(rectangle2_widths[2087]), .rectangle2_height(rectangle2_heights[2087]), .rectangle2_weight(rectangle2_weights[2087]), .rectangle3_x(rectangle3_xs[2087]), .rectangle3_y(rectangle3_ys[2087]), .rectangle3_width(rectangle3_widths[2087]), .rectangle3_height(rectangle3_heights[2087]), .rectangle3_weight(rectangle3_weights[2087]), .feature_threshold(feature_thresholds[2087]), .feature_above(feature_aboves[2087]), .feature_below(feature_belows[2087]), .scan_win_std_dev(scan_win_std_dev[2087]), .feature_accum(feature_accums[2087]));
  accum_calculator ac2088(.scan_win(scan_win2088), .rectangle1_x(rectangle1_xs[2088]), .rectangle1_y(rectangle1_ys[2088]), .rectangle1_width(rectangle1_widths[2088]), .rectangle1_height(rectangle1_heights[2088]), .rectangle1_weight(rectangle1_weights[2088]), .rectangle2_x(rectangle2_xs[2088]), .rectangle2_y(rectangle2_ys[2088]), .rectangle2_width(rectangle2_widths[2088]), .rectangle2_height(rectangle2_heights[2088]), .rectangle2_weight(rectangle2_weights[2088]), .rectangle3_x(rectangle3_xs[2088]), .rectangle3_y(rectangle3_ys[2088]), .rectangle3_width(rectangle3_widths[2088]), .rectangle3_height(rectangle3_heights[2088]), .rectangle3_weight(rectangle3_weights[2088]), .feature_threshold(feature_thresholds[2088]), .feature_above(feature_aboves[2088]), .feature_below(feature_belows[2088]), .scan_win_std_dev(scan_win_std_dev[2088]), .feature_accum(feature_accums[2088]));
  accum_calculator ac2089(.scan_win(scan_win2089), .rectangle1_x(rectangle1_xs[2089]), .rectangle1_y(rectangle1_ys[2089]), .rectangle1_width(rectangle1_widths[2089]), .rectangle1_height(rectangle1_heights[2089]), .rectangle1_weight(rectangle1_weights[2089]), .rectangle2_x(rectangle2_xs[2089]), .rectangle2_y(rectangle2_ys[2089]), .rectangle2_width(rectangle2_widths[2089]), .rectangle2_height(rectangle2_heights[2089]), .rectangle2_weight(rectangle2_weights[2089]), .rectangle3_x(rectangle3_xs[2089]), .rectangle3_y(rectangle3_ys[2089]), .rectangle3_width(rectangle3_widths[2089]), .rectangle3_height(rectangle3_heights[2089]), .rectangle3_weight(rectangle3_weights[2089]), .feature_threshold(feature_thresholds[2089]), .feature_above(feature_aboves[2089]), .feature_below(feature_belows[2089]), .scan_win_std_dev(scan_win_std_dev[2089]), .feature_accum(feature_accums[2089]));
  accum_calculator ac2090(.scan_win(scan_win2090), .rectangle1_x(rectangle1_xs[2090]), .rectangle1_y(rectangle1_ys[2090]), .rectangle1_width(rectangle1_widths[2090]), .rectangle1_height(rectangle1_heights[2090]), .rectangle1_weight(rectangle1_weights[2090]), .rectangle2_x(rectangle2_xs[2090]), .rectangle2_y(rectangle2_ys[2090]), .rectangle2_width(rectangle2_widths[2090]), .rectangle2_height(rectangle2_heights[2090]), .rectangle2_weight(rectangle2_weights[2090]), .rectangle3_x(rectangle3_xs[2090]), .rectangle3_y(rectangle3_ys[2090]), .rectangle3_width(rectangle3_widths[2090]), .rectangle3_height(rectangle3_heights[2090]), .rectangle3_weight(rectangle3_weights[2090]), .feature_threshold(feature_thresholds[2090]), .feature_above(feature_aboves[2090]), .feature_below(feature_belows[2090]), .scan_win_std_dev(scan_win_std_dev[2090]), .feature_accum(feature_accums[2090]));
  accum_calculator ac2091(.scan_win(scan_win2091), .rectangle1_x(rectangle1_xs[2091]), .rectangle1_y(rectangle1_ys[2091]), .rectangle1_width(rectangle1_widths[2091]), .rectangle1_height(rectangle1_heights[2091]), .rectangle1_weight(rectangle1_weights[2091]), .rectangle2_x(rectangle2_xs[2091]), .rectangle2_y(rectangle2_ys[2091]), .rectangle2_width(rectangle2_widths[2091]), .rectangle2_height(rectangle2_heights[2091]), .rectangle2_weight(rectangle2_weights[2091]), .rectangle3_x(rectangle3_xs[2091]), .rectangle3_y(rectangle3_ys[2091]), .rectangle3_width(rectangle3_widths[2091]), .rectangle3_height(rectangle3_heights[2091]), .rectangle3_weight(rectangle3_weights[2091]), .feature_threshold(feature_thresholds[2091]), .feature_above(feature_aboves[2091]), .feature_below(feature_belows[2091]), .scan_win_std_dev(scan_win_std_dev[2091]), .feature_accum(feature_accums[2091]));
  accum_calculator ac2092(.scan_win(scan_win2092), .rectangle1_x(rectangle1_xs[2092]), .rectangle1_y(rectangle1_ys[2092]), .rectangle1_width(rectangle1_widths[2092]), .rectangle1_height(rectangle1_heights[2092]), .rectangle1_weight(rectangle1_weights[2092]), .rectangle2_x(rectangle2_xs[2092]), .rectangle2_y(rectangle2_ys[2092]), .rectangle2_width(rectangle2_widths[2092]), .rectangle2_height(rectangle2_heights[2092]), .rectangle2_weight(rectangle2_weights[2092]), .rectangle3_x(rectangle3_xs[2092]), .rectangle3_y(rectangle3_ys[2092]), .rectangle3_width(rectangle3_widths[2092]), .rectangle3_height(rectangle3_heights[2092]), .rectangle3_weight(rectangle3_weights[2092]), .feature_threshold(feature_thresholds[2092]), .feature_above(feature_aboves[2092]), .feature_below(feature_belows[2092]), .scan_win_std_dev(scan_win_std_dev[2092]), .feature_accum(feature_accums[2092]));
  accum_calculator ac2093(.scan_win(scan_win2093), .rectangle1_x(rectangle1_xs[2093]), .rectangle1_y(rectangle1_ys[2093]), .rectangle1_width(rectangle1_widths[2093]), .rectangle1_height(rectangle1_heights[2093]), .rectangle1_weight(rectangle1_weights[2093]), .rectangle2_x(rectangle2_xs[2093]), .rectangle2_y(rectangle2_ys[2093]), .rectangle2_width(rectangle2_widths[2093]), .rectangle2_height(rectangle2_heights[2093]), .rectangle2_weight(rectangle2_weights[2093]), .rectangle3_x(rectangle3_xs[2093]), .rectangle3_y(rectangle3_ys[2093]), .rectangle3_width(rectangle3_widths[2093]), .rectangle3_height(rectangle3_heights[2093]), .rectangle3_weight(rectangle3_weights[2093]), .feature_threshold(feature_thresholds[2093]), .feature_above(feature_aboves[2093]), .feature_below(feature_belows[2093]), .scan_win_std_dev(scan_win_std_dev[2093]), .feature_accum(feature_accums[2093]));
  accum_calculator ac2094(.scan_win(scan_win2094), .rectangle1_x(rectangle1_xs[2094]), .rectangle1_y(rectangle1_ys[2094]), .rectangle1_width(rectangle1_widths[2094]), .rectangle1_height(rectangle1_heights[2094]), .rectangle1_weight(rectangle1_weights[2094]), .rectangle2_x(rectangle2_xs[2094]), .rectangle2_y(rectangle2_ys[2094]), .rectangle2_width(rectangle2_widths[2094]), .rectangle2_height(rectangle2_heights[2094]), .rectangle2_weight(rectangle2_weights[2094]), .rectangle3_x(rectangle3_xs[2094]), .rectangle3_y(rectangle3_ys[2094]), .rectangle3_width(rectangle3_widths[2094]), .rectangle3_height(rectangle3_heights[2094]), .rectangle3_weight(rectangle3_weights[2094]), .feature_threshold(feature_thresholds[2094]), .feature_above(feature_aboves[2094]), .feature_below(feature_belows[2094]), .scan_win_std_dev(scan_win_std_dev[2094]), .feature_accum(feature_accums[2094]));
  accum_calculator ac2095(.scan_win(scan_win2095), .rectangle1_x(rectangle1_xs[2095]), .rectangle1_y(rectangle1_ys[2095]), .rectangle1_width(rectangle1_widths[2095]), .rectangle1_height(rectangle1_heights[2095]), .rectangle1_weight(rectangle1_weights[2095]), .rectangle2_x(rectangle2_xs[2095]), .rectangle2_y(rectangle2_ys[2095]), .rectangle2_width(rectangle2_widths[2095]), .rectangle2_height(rectangle2_heights[2095]), .rectangle2_weight(rectangle2_weights[2095]), .rectangle3_x(rectangle3_xs[2095]), .rectangle3_y(rectangle3_ys[2095]), .rectangle3_width(rectangle3_widths[2095]), .rectangle3_height(rectangle3_heights[2095]), .rectangle3_weight(rectangle3_weights[2095]), .feature_threshold(feature_thresholds[2095]), .feature_above(feature_aboves[2095]), .feature_below(feature_belows[2095]), .scan_win_std_dev(scan_win_std_dev[2095]), .feature_accum(feature_accums[2095]));
  accum_calculator ac2096(.scan_win(scan_win2096), .rectangle1_x(rectangle1_xs[2096]), .rectangle1_y(rectangle1_ys[2096]), .rectangle1_width(rectangle1_widths[2096]), .rectangle1_height(rectangle1_heights[2096]), .rectangle1_weight(rectangle1_weights[2096]), .rectangle2_x(rectangle2_xs[2096]), .rectangle2_y(rectangle2_ys[2096]), .rectangle2_width(rectangle2_widths[2096]), .rectangle2_height(rectangle2_heights[2096]), .rectangle2_weight(rectangle2_weights[2096]), .rectangle3_x(rectangle3_xs[2096]), .rectangle3_y(rectangle3_ys[2096]), .rectangle3_width(rectangle3_widths[2096]), .rectangle3_height(rectangle3_heights[2096]), .rectangle3_weight(rectangle3_weights[2096]), .feature_threshold(feature_thresholds[2096]), .feature_above(feature_aboves[2096]), .feature_below(feature_belows[2096]), .scan_win_std_dev(scan_win_std_dev[2096]), .feature_accum(feature_accums[2096]));
  accum_calculator ac2097(.scan_win(scan_win2097), .rectangle1_x(rectangle1_xs[2097]), .rectangle1_y(rectangle1_ys[2097]), .rectangle1_width(rectangle1_widths[2097]), .rectangle1_height(rectangle1_heights[2097]), .rectangle1_weight(rectangle1_weights[2097]), .rectangle2_x(rectangle2_xs[2097]), .rectangle2_y(rectangle2_ys[2097]), .rectangle2_width(rectangle2_widths[2097]), .rectangle2_height(rectangle2_heights[2097]), .rectangle2_weight(rectangle2_weights[2097]), .rectangle3_x(rectangle3_xs[2097]), .rectangle3_y(rectangle3_ys[2097]), .rectangle3_width(rectangle3_widths[2097]), .rectangle3_height(rectangle3_heights[2097]), .rectangle3_weight(rectangle3_weights[2097]), .feature_threshold(feature_thresholds[2097]), .feature_above(feature_aboves[2097]), .feature_below(feature_belows[2097]), .scan_win_std_dev(scan_win_std_dev[2097]), .feature_accum(feature_accums[2097]));
  accum_calculator ac2098(.scan_win(scan_win2098), .rectangle1_x(rectangle1_xs[2098]), .rectangle1_y(rectangle1_ys[2098]), .rectangle1_width(rectangle1_widths[2098]), .rectangle1_height(rectangle1_heights[2098]), .rectangle1_weight(rectangle1_weights[2098]), .rectangle2_x(rectangle2_xs[2098]), .rectangle2_y(rectangle2_ys[2098]), .rectangle2_width(rectangle2_widths[2098]), .rectangle2_height(rectangle2_heights[2098]), .rectangle2_weight(rectangle2_weights[2098]), .rectangle3_x(rectangle3_xs[2098]), .rectangle3_y(rectangle3_ys[2098]), .rectangle3_width(rectangle3_widths[2098]), .rectangle3_height(rectangle3_heights[2098]), .rectangle3_weight(rectangle3_weights[2098]), .feature_threshold(feature_thresholds[2098]), .feature_above(feature_aboves[2098]), .feature_below(feature_belows[2098]), .scan_win_std_dev(scan_win_std_dev[2098]), .feature_accum(feature_accums[2098]));
  accum_calculator ac2099(.scan_win(scan_win2099), .rectangle1_x(rectangle1_xs[2099]), .rectangle1_y(rectangle1_ys[2099]), .rectangle1_width(rectangle1_widths[2099]), .rectangle1_height(rectangle1_heights[2099]), .rectangle1_weight(rectangle1_weights[2099]), .rectangle2_x(rectangle2_xs[2099]), .rectangle2_y(rectangle2_ys[2099]), .rectangle2_width(rectangle2_widths[2099]), .rectangle2_height(rectangle2_heights[2099]), .rectangle2_weight(rectangle2_weights[2099]), .rectangle3_x(rectangle3_xs[2099]), .rectangle3_y(rectangle3_ys[2099]), .rectangle3_width(rectangle3_widths[2099]), .rectangle3_height(rectangle3_heights[2099]), .rectangle3_weight(rectangle3_weights[2099]), .feature_threshold(feature_thresholds[2099]), .feature_above(feature_aboves[2099]), .feature_below(feature_belows[2099]), .scan_win_std_dev(scan_win_std_dev[2099]), .feature_accum(feature_accums[2099]));
  accum_calculator ac2100(.scan_win(scan_win2100), .rectangle1_x(rectangle1_xs[2100]), .rectangle1_y(rectangle1_ys[2100]), .rectangle1_width(rectangle1_widths[2100]), .rectangle1_height(rectangle1_heights[2100]), .rectangle1_weight(rectangle1_weights[2100]), .rectangle2_x(rectangle2_xs[2100]), .rectangle2_y(rectangle2_ys[2100]), .rectangle2_width(rectangle2_widths[2100]), .rectangle2_height(rectangle2_heights[2100]), .rectangle2_weight(rectangle2_weights[2100]), .rectangle3_x(rectangle3_xs[2100]), .rectangle3_y(rectangle3_ys[2100]), .rectangle3_width(rectangle3_widths[2100]), .rectangle3_height(rectangle3_heights[2100]), .rectangle3_weight(rectangle3_weights[2100]), .feature_threshold(feature_thresholds[2100]), .feature_above(feature_aboves[2100]), .feature_below(feature_belows[2100]), .scan_win_std_dev(scan_win_std_dev[2100]), .feature_accum(feature_accums[2100]));
  accum_calculator ac2101(.scan_win(scan_win2101), .rectangle1_x(rectangle1_xs[2101]), .rectangle1_y(rectangle1_ys[2101]), .rectangle1_width(rectangle1_widths[2101]), .rectangle1_height(rectangle1_heights[2101]), .rectangle1_weight(rectangle1_weights[2101]), .rectangle2_x(rectangle2_xs[2101]), .rectangle2_y(rectangle2_ys[2101]), .rectangle2_width(rectangle2_widths[2101]), .rectangle2_height(rectangle2_heights[2101]), .rectangle2_weight(rectangle2_weights[2101]), .rectangle3_x(rectangle3_xs[2101]), .rectangle3_y(rectangle3_ys[2101]), .rectangle3_width(rectangle3_widths[2101]), .rectangle3_height(rectangle3_heights[2101]), .rectangle3_weight(rectangle3_weights[2101]), .feature_threshold(feature_thresholds[2101]), .feature_above(feature_aboves[2101]), .feature_below(feature_belows[2101]), .scan_win_std_dev(scan_win_std_dev[2101]), .feature_accum(feature_accums[2101]));
  accum_calculator ac2102(.scan_win(scan_win2102), .rectangle1_x(rectangle1_xs[2102]), .rectangle1_y(rectangle1_ys[2102]), .rectangle1_width(rectangle1_widths[2102]), .rectangle1_height(rectangle1_heights[2102]), .rectangle1_weight(rectangle1_weights[2102]), .rectangle2_x(rectangle2_xs[2102]), .rectangle2_y(rectangle2_ys[2102]), .rectangle2_width(rectangle2_widths[2102]), .rectangle2_height(rectangle2_heights[2102]), .rectangle2_weight(rectangle2_weights[2102]), .rectangle3_x(rectangle3_xs[2102]), .rectangle3_y(rectangle3_ys[2102]), .rectangle3_width(rectangle3_widths[2102]), .rectangle3_height(rectangle3_heights[2102]), .rectangle3_weight(rectangle3_weights[2102]), .feature_threshold(feature_thresholds[2102]), .feature_above(feature_aboves[2102]), .feature_below(feature_belows[2102]), .scan_win_std_dev(scan_win_std_dev[2102]), .feature_accum(feature_accums[2102]));
  accum_calculator ac2103(.scan_win(scan_win2103), .rectangle1_x(rectangle1_xs[2103]), .rectangle1_y(rectangle1_ys[2103]), .rectangle1_width(rectangle1_widths[2103]), .rectangle1_height(rectangle1_heights[2103]), .rectangle1_weight(rectangle1_weights[2103]), .rectangle2_x(rectangle2_xs[2103]), .rectangle2_y(rectangle2_ys[2103]), .rectangle2_width(rectangle2_widths[2103]), .rectangle2_height(rectangle2_heights[2103]), .rectangle2_weight(rectangle2_weights[2103]), .rectangle3_x(rectangle3_xs[2103]), .rectangle3_y(rectangle3_ys[2103]), .rectangle3_width(rectangle3_widths[2103]), .rectangle3_height(rectangle3_heights[2103]), .rectangle3_weight(rectangle3_weights[2103]), .feature_threshold(feature_thresholds[2103]), .feature_above(feature_aboves[2103]), .feature_below(feature_belows[2103]), .scan_win_std_dev(scan_win_std_dev[2103]), .feature_accum(feature_accums[2103]));
  accum_calculator ac2104(.scan_win(scan_win2104), .rectangle1_x(rectangle1_xs[2104]), .rectangle1_y(rectangle1_ys[2104]), .rectangle1_width(rectangle1_widths[2104]), .rectangle1_height(rectangle1_heights[2104]), .rectangle1_weight(rectangle1_weights[2104]), .rectangle2_x(rectangle2_xs[2104]), .rectangle2_y(rectangle2_ys[2104]), .rectangle2_width(rectangle2_widths[2104]), .rectangle2_height(rectangle2_heights[2104]), .rectangle2_weight(rectangle2_weights[2104]), .rectangle3_x(rectangle3_xs[2104]), .rectangle3_y(rectangle3_ys[2104]), .rectangle3_width(rectangle3_widths[2104]), .rectangle3_height(rectangle3_heights[2104]), .rectangle3_weight(rectangle3_weights[2104]), .feature_threshold(feature_thresholds[2104]), .feature_above(feature_aboves[2104]), .feature_below(feature_belows[2104]), .scan_win_std_dev(scan_win_std_dev[2104]), .feature_accum(feature_accums[2104]));
  accum_calculator ac2105(.scan_win(scan_win2105), .rectangle1_x(rectangle1_xs[2105]), .rectangle1_y(rectangle1_ys[2105]), .rectangle1_width(rectangle1_widths[2105]), .rectangle1_height(rectangle1_heights[2105]), .rectangle1_weight(rectangle1_weights[2105]), .rectangle2_x(rectangle2_xs[2105]), .rectangle2_y(rectangle2_ys[2105]), .rectangle2_width(rectangle2_widths[2105]), .rectangle2_height(rectangle2_heights[2105]), .rectangle2_weight(rectangle2_weights[2105]), .rectangle3_x(rectangle3_xs[2105]), .rectangle3_y(rectangle3_ys[2105]), .rectangle3_width(rectangle3_widths[2105]), .rectangle3_height(rectangle3_heights[2105]), .rectangle3_weight(rectangle3_weights[2105]), .feature_threshold(feature_thresholds[2105]), .feature_above(feature_aboves[2105]), .feature_below(feature_belows[2105]), .scan_win_std_dev(scan_win_std_dev[2105]), .feature_accum(feature_accums[2105]));
  accum_calculator ac2106(.scan_win(scan_win2106), .rectangle1_x(rectangle1_xs[2106]), .rectangle1_y(rectangle1_ys[2106]), .rectangle1_width(rectangle1_widths[2106]), .rectangle1_height(rectangle1_heights[2106]), .rectangle1_weight(rectangle1_weights[2106]), .rectangle2_x(rectangle2_xs[2106]), .rectangle2_y(rectangle2_ys[2106]), .rectangle2_width(rectangle2_widths[2106]), .rectangle2_height(rectangle2_heights[2106]), .rectangle2_weight(rectangle2_weights[2106]), .rectangle3_x(rectangle3_xs[2106]), .rectangle3_y(rectangle3_ys[2106]), .rectangle3_width(rectangle3_widths[2106]), .rectangle3_height(rectangle3_heights[2106]), .rectangle3_weight(rectangle3_weights[2106]), .feature_threshold(feature_thresholds[2106]), .feature_above(feature_aboves[2106]), .feature_below(feature_belows[2106]), .scan_win_std_dev(scan_win_std_dev[2106]), .feature_accum(feature_accums[2106]));
  accum_calculator ac2107(.scan_win(scan_win2107), .rectangle1_x(rectangle1_xs[2107]), .rectangle1_y(rectangle1_ys[2107]), .rectangle1_width(rectangle1_widths[2107]), .rectangle1_height(rectangle1_heights[2107]), .rectangle1_weight(rectangle1_weights[2107]), .rectangle2_x(rectangle2_xs[2107]), .rectangle2_y(rectangle2_ys[2107]), .rectangle2_width(rectangle2_widths[2107]), .rectangle2_height(rectangle2_heights[2107]), .rectangle2_weight(rectangle2_weights[2107]), .rectangle3_x(rectangle3_xs[2107]), .rectangle3_y(rectangle3_ys[2107]), .rectangle3_width(rectangle3_widths[2107]), .rectangle3_height(rectangle3_heights[2107]), .rectangle3_weight(rectangle3_weights[2107]), .feature_threshold(feature_thresholds[2107]), .feature_above(feature_aboves[2107]), .feature_below(feature_belows[2107]), .scan_win_std_dev(scan_win_std_dev[2107]), .feature_accum(feature_accums[2107]));
  accum_calculator ac2108(.scan_win(scan_win2108), .rectangle1_x(rectangle1_xs[2108]), .rectangle1_y(rectangle1_ys[2108]), .rectangle1_width(rectangle1_widths[2108]), .rectangle1_height(rectangle1_heights[2108]), .rectangle1_weight(rectangle1_weights[2108]), .rectangle2_x(rectangle2_xs[2108]), .rectangle2_y(rectangle2_ys[2108]), .rectangle2_width(rectangle2_widths[2108]), .rectangle2_height(rectangle2_heights[2108]), .rectangle2_weight(rectangle2_weights[2108]), .rectangle3_x(rectangle3_xs[2108]), .rectangle3_y(rectangle3_ys[2108]), .rectangle3_width(rectangle3_widths[2108]), .rectangle3_height(rectangle3_heights[2108]), .rectangle3_weight(rectangle3_weights[2108]), .feature_threshold(feature_thresholds[2108]), .feature_above(feature_aboves[2108]), .feature_below(feature_belows[2108]), .scan_win_std_dev(scan_win_std_dev[2108]), .feature_accum(feature_accums[2108]));
  accum_calculator ac2109(.scan_win(scan_win2109), .rectangle1_x(rectangle1_xs[2109]), .rectangle1_y(rectangle1_ys[2109]), .rectangle1_width(rectangle1_widths[2109]), .rectangle1_height(rectangle1_heights[2109]), .rectangle1_weight(rectangle1_weights[2109]), .rectangle2_x(rectangle2_xs[2109]), .rectangle2_y(rectangle2_ys[2109]), .rectangle2_width(rectangle2_widths[2109]), .rectangle2_height(rectangle2_heights[2109]), .rectangle2_weight(rectangle2_weights[2109]), .rectangle3_x(rectangle3_xs[2109]), .rectangle3_y(rectangle3_ys[2109]), .rectangle3_width(rectangle3_widths[2109]), .rectangle3_height(rectangle3_heights[2109]), .rectangle3_weight(rectangle3_weights[2109]), .feature_threshold(feature_thresholds[2109]), .feature_above(feature_aboves[2109]), .feature_below(feature_belows[2109]), .scan_win_std_dev(scan_win_std_dev[2109]), .feature_accum(feature_accums[2109]));
  accum_calculator ac2110(.scan_win(scan_win2110), .rectangle1_x(rectangle1_xs[2110]), .rectangle1_y(rectangle1_ys[2110]), .rectangle1_width(rectangle1_widths[2110]), .rectangle1_height(rectangle1_heights[2110]), .rectangle1_weight(rectangle1_weights[2110]), .rectangle2_x(rectangle2_xs[2110]), .rectangle2_y(rectangle2_ys[2110]), .rectangle2_width(rectangle2_widths[2110]), .rectangle2_height(rectangle2_heights[2110]), .rectangle2_weight(rectangle2_weights[2110]), .rectangle3_x(rectangle3_xs[2110]), .rectangle3_y(rectangle3_ys[2110]), .rectangle3_width(rectangle3_widths[2110]), .rectangle3_height(rectangle3_heights[2110]), .rectangle3_weight(rectangle3_weights[2110]), .feature_threshold(feature_thresholds[2110]), .feature_above(feature_aboves[2110]), .feature_below(feature_belows[2110]), .scan_win_std_dev(scan_win_std_dev[2110]), .feature_accum(feature_accums[2110]));
  accum_calculator ac2111(.scan_win(scan_win2111), .rectangle1_x(rectangle1_xs[2111]), .rectangle1_y(rectangle1_ys[2111]), .rectangle1_width(rectangle1_widths[2111]), .rectangle1_height(rectangle1_heights[2111]), .rectangle1_weight(rectangle1_weights[2111]), .rectangle2_x(rectangle2_xs[2111]), .rectangle2_y(rectangle2_ys[2111]), .rectangle2_width(rectangle2_widths[2111]), .rectangle2_height(rectangle2_heights[2111]), .rectangle2_weight(rectangle2_weights[2111]), .rectangle3_x(rectangle3_xs[2111]), .rectangle3_y(rectangle3_ys[2111]), .rectangle3_width(rectangle3_widths[2111]), .rectangle3_height(rectangle3_heights[2111]), .rectangle3_weight(rectangle3_weights[2111]), .feature_threshold(feature_thresholds[2111]), .feature_above(feature_aboves[2111]), .feature_below(feature_belows[2111]), .scan_win_std_dev(scan_win_std_dev[2111]), .feature_accum(feature_accums[2111]));
  accum_calculator ac2112(.scan_win(scan_win2112), .rectangle1_x(rectangle1_xs[2112]), .rectangle1_y(rectangle1_ys[2112]), .rectangle1_width(rectangle1_widths[2112]), .rectangle1_height(rectangle1_heights[2112]), .rectangle1_weight(rectangle1_weights[2112]), .rectangle2_x(rectangle2_xs[2112]), .rectangle2_y(rectangle2_ys[2112]), .rectangle2_width(rectangle2_widths[2112]), .rectangle2_height(rectangle2_heights[2112]), .rectangle2_weight(rectangle2_weights[2112]), .rectangle3_x(rectangle3_xs[2112]), .rectangle3_y(rectangle3_ys[2112]), .rectangle3_width(rectangle3_widths[2112]), .rectangle3_height(rectangle3_heights[2112]), .rectangle3_weight(rectangle3_weights[2112]), .feature_threshold(feature_thresholds[2112]), .feature_above(feature_aboves[2112]), .feature_below(feature_belows[2112]), .scan_win_std_dev(scan_win_std_dev[2112]), .feature_accum(feature_accums[2112]));
  accum_calculator ac2113(.scan_win(scan_win2113), .rectangle1_x(rectangle1_xs[2113]), .rectangle1_y(rectangle1_ys[2113]), .rectangle1_width(rectangle1_widths[2113]), .rectangle1_height(rectangle1_heights[2113]), .rectangle1_weight(rectangle1_weights[2113]), .rectangle2_x(rectangle2_xs[2113]), .rectangle2_y(rectangle2_ys[2113]), .rectangle2_width(rectangle2_widths[2113]), .rectangle2_height(rectangle2_heights[2113]), .rectangle2_weight(rectangle2_weights[2113]), .rectangle3_x(rectangle3_xs[2113]), .rectangle3_y(rectangle3_ys[2113]), .rectangle3_width(rectangle3_widths[2113]), .rectangle3_height(rectangle3_heights[2113]), .rectangle3_weight(rectangle3_weights[2113]), .feature_threshold(feature_thresholds[2113]), .feature_above(feature_aboves[2113]), .feature_below(feature_belows[2113]), .scan_win_std_dev(scan_win_std_dev[2113]), .feature_accum(feature_accums[2113]));
  accum_calculator ac2114(.scan_win(scan_win2114), .rectangle1_x(rectangle1_xs[2114]), .rectangle1_y(rectangle1_ys[2114]), .rectangle1_width(rectangle1_widths[2114]), .rectangle1_height(rectangle1_heights[2114]), .rectangle1_weight(rectangle1_weights[2114]), .rectangle2_x(rectangle2_xs[2114]), .rectangle2_y(rectangle2_ys[2114]), .rectangle2_width(rectangle2_widths[2114]), .rectangle2_height(rectangle2_heights[2114]), .rectangle2_weight(rectangle2_weights[2114]), .rectangle3_x(rectangle3_xs[2114]), .rectangle3_y(rectangle3_ys[2114]), .rectangle3_width(rectangle3_widths[2114]), .rectangle3_height(rectangle3_heights[2114]), .rectangle3_weight(rectangle3_weights[2114]), .feature_threshold(feature_thresholds[2114]), .feature_above(feature_aboves[2114]), .feature_below(feature_belows[2114]), .scan_win_std_dev(scan_win_std_dev[2114]), .feature_accum(feature_accums[2114]));
  accum_calculator ac2115(.scan_win(scan_win2115), .rectangle1_x(rectangle1_xs[2115]), .rectangle1_y(rectangle1_ys[2115]), .rectangle1_width(rectangle1_widths[2115]), .rectangle1_height(rectangle1_heights[2115]), .rectangle1_weight(rectangle1_weights[2115]), .rectangle2_x(rectangle2_xs[2115]), .rectangle2_y(rectangle2_ys[2115]), .rectangle2_width(rectangle2_widths[2115]), .rectangle2_height(rectangle2_heights[2115]), .rectangle2_weight(rectangle2_weights[2115]), .rectangle3_x(rectangle3_xs[2115]), .rectangle3_y(rectangle3_ys[2115]), .rectangle3_width(rectangle3_widths[2115]), .rectangle3_height(rectangle3_heights[2115]), .rectangle3_weight(rectangle3_weights[2115]), .feature_threshold(feature_thresholds[2115]), .feature_above(feature_aboves[2115]), .feature_below(feature_belows[2115]), .scan_win_std_dev(scan_win_std_dev[2115]), .feature_accum(feature_accums[2115]));
  accum_calculator ac2116(.scan_win(scan_win2116), .rectangle1_x(rectangle1_xs[2116]), .rectangle1_y(rectangle1_ys[2116]), .rectangle1_width(rectangle1_widths[2116]), .rectangle1_height(rectangle1_heights[2116]), .rectangle1_weight(rectangle1_weights[2116]), .rectangle2_x(rectangle2_xs[2116]), .rectangle2_y(rectangle2_ys[2116]), .rectangle2_width(rectangle2_widths[2116]), .rectangle2_height(rectangle2_heights[2116]), .rectangle2_weight(rectangle2_weights[2116]), .rectangle3_x(rectangle3_xs[2116]), .rectangle3_y(rectangle3_ys[2116]), .rectangle3_width(rectangle3_widths[2116]), .rectangle3_height(rectangle3_heights[2116]), .rectangle3_weight(rectangle3_weights[2116]), .feature_threshold(feature_thresholds[2116]), .feature_above(feature_aboves[2116]), .feature_below(feature_belows[2116]), .scan_win_std_dev(scan_win_std_dev[2116]), .feature_accum(feature_accums[2116]));
  accum_calculator ac2117(.scan_win(scan_win2117), .rectangle1_x(rectangle1_xs[2117]), .rectangle1_y(rectangle1_ys[2117]), .rectangle1_width(rectangle1_widths[2117]), .rectangle1_height(rectangle1_heights[2117]), .rectangle1_weight(rectangle1_weights[2117]), .rectangle2_x(rectangle2_xs[2117]), .rectangle2_y(rectangle2_ys[2117]), .rectangle2_width(rectangle2_widths[2117]), .rectangle2_height(rectangle2_heights[2117]), .rectangle2_weight(rectangle2_weights[2117]), .rectangle3_x(rectangle3_xs[2117]), .rectangle3_y(rectangle3_ys[2117]), .rectangle3_width(rectangle3_widths[2117]), .rectangle3_height(rectangle3_heights[2117]), .rectangle3_weight(rectangle3_weights[2117]), .feature_threshold(feature_thresholds[2117]), .feature_above(feature_aboves[2117]), .feature_below(feature_belows[2117]), .scan_win_std_dev(scan_win_std_dev[2117]), .feature_accum(feature_accums[2117]));
  accum_calculator ac2118(.scan_win(scan_win2118), .rectangle1_x(rectangle1_xs[2118]), .rectangle1_y(rectangle1_ys[2118]), .rectangle1_width(rectangle1_widths[2118]), .rectangle1_height(rectangle1_heights[2118]), .rectangle1_weight(rectangle1_weights[2118]), .rectangle2_x(rectangle2_xs[2118]), .rectangle2_y(rectangle2_ys[2118]), .rectangle2_width(rectangle2_widths[2118]), .rectangle2_height(rectangle2_heights[2118]), .rectangle2_weight(rectangle2_weights[2118]), .rectangle3_x(rectangle3_xs[2118]), .rectangle3_y(rectangle3_ys[2118]), .rectangle3_width(rectangle3_widths[2118]), .rectangle3_height(rectangle3_heights[2118]), .rectangle3_weight(rectangle3_weights[2118]), .feature_threshold(feature_thresholds[2118]), .feature_above(feature_aboves[2118]), .feature_below(feature_belows[2118]), .scan_win_std_dev(scan_win_std_dev[2118]), .feature_accum(feature_accums[2118]));
  accum_calculator ac2119(.scan_win(scan_win2119), .rectangle1_x(rectangle1_xs[2119]), .rectangle1_y(rectangle1_ys[2119]), .rectangle1_width(rectangle1_widths[2119]), .rectangle1_height(rectangle1_heights[2119]), .rectangle1_weight(rectangle1_weights[2119]), .rectangle2_x(rectangle2_xs[2119]), .rectangle2_y(rectangle2_ys[2119]), .rectangle2_width(rectangle2_widths[2119]), .rectangle2_height(rectangle2_heights[2119]), .rectangle2_weight(rectangle2_weights[2119]), .rectangle3_x(rectangle3_xs[2119]), .rectangle3_y(rectangle3_ys[2119]), .rectangle3_width(rectangle3_widths[2119]), .rectangle3_height(rectangle3_heights[2119]), .rectangle3_weight(rectangle3_weights[2119]), .feature_threshold(feature_thresholds[2119]), .feature_above(feature_aboves[2119]), .feature_below(feature_belows[2119]), .scan_win_std_dev(scan_win_std_dev[2119]), .feature_accum(feature_accums[2119]));
  accum_calculator ac2120(.scan_win(scan_win2120), .rectangle1_x(rectangle1_xs[2120]), .rectangle1_y(rectangle1_ys[2120]), .rectangle1_width(rectangle1_widths[2120]), .rectangle1_height(rectangle1_heights[2120]), .rectangle1_weight(rectangle1_weights[2120]), .rectangle2_x(rectangle2_xs[2120]), .rectangle2_y(rectangle2_ys[2120]), .rectangle2_width(rectangle2_widths[2120]), .rectangle2_height(rectangle2_heights[2120]), .rectangle2_weight(rectangle2_weights[2120]), .rectangle3_x(rectangle3_xs[2120]), .rectangle3_y(rectangle3_ys[2120]), .rectangle3_width(rectangle3_widths[2120]), .rectangle3_height(rectangle3_heights[2120]), .rectangle3_weight(rectangle3_weights[2120]), .feature_threshold(feature_thresholds[2120]), .feature_above(feature_aboves[2120]), .feature_below(feature_belows[2120]), .scan_win_std_dev(scan_win_std_dev[2120]), .feature_accum(feature_accums[2120]));
  accum_calculator ac2121(.scan_win(scan_win2121), .rectangle1_x(rectangle1_xs[2121]), .rectangle1_y(rectangle1_ys[2121]), .rectangle1_width(rectangle1_widths[2121]), .rectangle1_height(rectangle1_heights[2121]), .rectangle1_weight(rectangle1_weights[2121]), .rectangle2_x(rectangle2_xs[2121]), .rectangle2_y(rectangle2_ys[2121]), .rectangle2_width(rectangle2_widths[2121]), .rectangle2_height(rectangle2_heights[2121]), .rectangle2_weight(rectangle2_weights[2121]), .rectangle3_x(rectangle3_xs[2121]), .rectangle3_y(rectangle3_ys[2121]), .rectangle3_width(rectangle3_widths[2121]), .rectangle3_height(rectangle3_heights[2121]), .rectangle3_weight(rectangle3_weights[2121]), .feature_threshold(feature_thresholds[2121]), .feature_above(feature_aboves[2121]), .feature_below(feature_belows[2121]), .scan_win_std_dev(scan_win_std_dev[2121]), .feature_accum(feature_accums[2121]));
  accum_calculator ac2122(.scan_win(scan_win2122), .rectangle1_x(rectangle1_xs[2122]), .rectangle1_y(rectangle1_ys[2122]), .rectangle1_width(rectangle1_widths[2122]), .rectangle1_height(rectangle1_heights[2122]), .rectangle1_weight(rectangle1_weights[2122]), .rectangle2_x(rectangle2_xs[2122]), .rectangle2_y(rectangle2_ys[2122]), .rectangle2_width(rectangle2_widths[2122]), .rectangle2_height(rectangle2_heights[2122]), .rectangle2_weight(rectangle2_weights[2122]), .rectangle3_x(rectangle3_xs[2122]), .rectangle3_y(rectangle3_ys[2122]), .rectangle3_width(rectangle3_widths[2122]), .rectangle3_height(rectangle3_heights[2122]), .rectangle3_weight(rectangle3_weights[2122]), .feature_threshold(feature_thresholds[2122]), .feature_above(feature_aboves[2122]), .feature_below(feature_belows[2122]), .scan_win_std_dev(scan_win_std_dev[2122]), .feature_accum(feature_accums[2122]));
  accum_calculator ac2123(.scan_win(scan_win2123), .rectangle1_x(rectangle1_xs[2123]), .rectangle1_y(rectangle1_ys[2123]), .rectangle1_width(rectangle1_widths[2123]), .rectangle1_height(rectangle1_heights[2123]), .rectangle1_weight(rectangle1_weights[2123]), .rectangle2_x(rectangle2_xs[2123]), .rectangle2_y(rectangle2_ys[2123]), .rectangle2_width(rectangle2_widths[2123]), .rectangle2_height(rectangle2_heights[2123]), .rectangle2_weight(rectangle2_weights[2123]), .rectangle3_x(rectangle3_xs[2123]), .rectangle3_y(rectangle3_ys[2123]), .rectangle3_width(rectangle3_widths[2123]), .rectangle3_height(rectangle3_heights[2123]), .rectangle3_weight(rectangle3_weights[2123]), .feature_threshold(feature_thresholds[2123]), .feature_above(feature_aboves[2123]), .feature_below(feature_belows[2123]), .scan_win_std_dev(scan_win_std_dev[2123]), .feature_accum(feature_accums[2123]));
  accum_calculator ac2124(.scan_win(scan_win2124), .rectangle1_x(rectangle1_xs[2124]), .rectangle1_y(rectangle1_ys[2124]), .rectangle1_width(rectangle1_widths[2124]), .rectangle1_height(rectangle1_heights[2124]), .rectangle1_weight(rectangle1_weights[2124]), .rectangle2_x(rectangle2_xs[2124]), .rectangle2_y(rectangle2_ys[2124]), .rectangle2_width(rectangle2_widths[2124]), .rectangle2_height(rectangle2_heights[2124]), .rectangle2_weight(rectangle2_weights[2124]), .rectangle3_x(rectangle3_xs[2124]), .rectangle3_y(rectangle3_ys[2124]), .rectangle3_width(rectangle3_widths[2124]), .rectangle3_height(rectangle3_heights[2124]), .rectangle3_weight(rectangle3_weights[2124]), .feature_threshold(feature_thresholds[2124]), .feature_above(feature_aboves[2124]), .feature_below(feature_belows[2124]), .scan_win_std_dev(scan_win_std_dev[2124]), .feature_accum(feature_accums[2124]));
  accum_calculator ac2125(.scan_win(scan_win2125), .rectangle1_x(rectangle1_xs[2125]), .rectangle1_y(rectangle1_ys[2125]), .rectangle1_width(rectangle1_widths[2125]), .rectangle1_height(rectangle1_heights[2125]), .rectangle1_weight(rectangle1_weights[2125]), .rectangle2_x(rectangle2_xs[2125]), .rectangle2_y(rectangle2_ys[2125]), .rectangle2_width(rectangle2_widths[2125]), .rectangle2_height(rectangle2_heights[2125]), .rectangle2_weight(rectangle2_weights[2125]), .rectangle3_x(rectangle3_xs[2125]), .rectangle3_y(rectangle3_ys[2125]), .rectangle3_width(rectangle3_widths[2125]), .rectangle3_height(rectangle3_heights[2125]), .rectangle3_weight(rectangle3_weights[2125]), .feature_threshold(feature_thresholds[2125]), .feature_above(feature_aboves[2125]), .feature_below(feature_belows[2125]), .scan_win_std_dev(scan_win_std_dev[2125]), .feature_accum(feature_accums[2125]));
  accum_calculator ac2126(.scan_win(scan_win2126), .rectangle1_x(rectangle1_xs[2126]), .rectangle1_y(rectangle1_ys[2126]), .rectangle1_width(rectangle1_widths[2126]), .rectangle1_height(rectangle1_heights[2126]), .rectangle1_weight(rectangle1_weights[2126]), .rectangle2_x(rectangle2_xs[2126]), .rectangle2_y(rectangle2_ys[2126]), .rectangle2_width(rectangle2_widths[2126]), .rectangle2_height(rectangle2_heights[2126]), .rectangle2_weight(rectangle2_weights[2126]), .rectangle3_x(rectangle3_xs[2126]), .rectangle3_y(rectangle3_ys[2126]), .rectangle3_width(rectangle3_widths[2126]), .rectangle3_height(rectangle3_heights[2126]), .rectangle3_weight(rectangle3_weights[2126]), .feature_threshold(feature_thresholds[2126]), .feature_above(feature_aboves[2126]), .feature_below(feature_belows[2126]), .scan_win_std_dev(scan_win_std_dev[2126]), .feature_accum(feature_accums[2126]));
  accum_calculator ac2127(.scan_win(scan_win2127), .rectangle1_x(rectangle1_xs[2127]), .rectangle1_y(rectangle1_ys[2127]), .rectangle1_width(rectangle1_widths[2127]), .rectangle1_height(rectangle1_heights[2127]), .rectangle1_weight(rectangle1_weights[2127]), .rectangle2_x(rectangle2_xs[2127]), .rectangle2_y(rectangle2_ys[2127]), .rectangle2_width(rectangle2_widths[2127]), .rectangle2_height(rectangle2_heights[2127]), .rectangle2_weight(rectangle2_weights[2127]), .rectangle3_x(rectangle3_xs[2127]), .rectangle3_y(rectangle3_ys[2127]), .rectangle3_width(rectangle3_widths[2127]), .rectangle3_height(rectangle3_heights[2127]), .rectangle3_weight(rectangle3_weights[2127]), .feature_threshold(feature_thresholds[2127]), .feature_above(feature_aboves[2127]), .feature_below(feature_belows[2127]), .scan_win_std_dev(scan_win_std_dev[2127]), .feature_accum(feature_accums[2127]));
  accum_calculator ac2128(.scan_win(scan_win2128), .rectangle1_x(rectangle1_xs[2128]), .rectangle1_y(rectangle1_ys[2128]), .rectangle1_width(rectangle1_widths[2128]), .rectangle1_height(rectangle1_heights[2128]), .rectangle1_weight(rectangle1_weights[2128]), .rectangle2_x(rectangle2_xs[2128]), .rectangle2_y(rectangle2_ys[2128]), .rectangle2_width(rectangle2_widths[2128]), .rectangle2_height(rectangle2_heights[2128]), .rectangle2_weight(rectangle2_weights[2128]), .rectangle3_x(rectangle3_xs[2128]), .rectangle3_y(rectangle3_ys[2128]), .rectangle3_width(rectangle3_widths[2128]), .rectangle3_height(rectangle3_heights[2128]), .rectangle3_weight(rectangle3_weights[2128]), .feature_threshold(feature_thresholds[2128]), .feature_above(feature_aboves[2128]), .feature_below(feature_belows[2128]), .scan_win_std_dev(scan_win_std_dev[2128]), .feature_accum(feature_accums[2128]));
  accum_calculator ac2129(.scan_win(scan_win2129), .rectangle1_x(rectangle1_xs[2129]), .rectangle1_y(rectangle1_ys[2129]), .rectangle1_width(rectangle1_widths[2129]), .rectangle1_height(rectangle1_heights[2129]), .rectangle1_weight(rectangle1_weights[2129]), .rectangle2_x(rectangle2_xs[2129]), .rectangle2_y(rectangle2_ys[2129]), .rectangle2_width(rectangle2_widths[2129]), .rectangle2_height(rectangle2_heights[2129]), .rectangle2_weight(rectangle2_weights[2129]), .rectangle3_x(rectangle3_xs[2129]), .rectangle3_y(rectangle3_ys[2129]), .rectangle3_width(rectangle3_widths[2129]), .rectangle3_height(rectangle3_heights[2129]), .rectangle3_weight(rectangle3_weights[2129]), .feature_threshold(feature_thresholds[2129]), .feature_above(feature_aboves[2129]), .feature_below(feature_belows[2129]), .scan_win_std_dev(scan_win_std_dev[2129]), .feature_accum(feature_accums[2129]));
  accum_calculator ac2130(.scan_win(scan_win2130), .rectangle1_x(rectangle1_xs[2130]), .rectangle1_y(rectangle1_ys[2130]), .rectangle1_width(rectangle1_widths[2130]), .rectangle1_height(rectangle1_heights[2130]), .rectangle1_weight(rectangle1_weights[2130]), .rectangle2_x(rectangle2_xs[2130]), .rectangle2_y(rectangle2_ys[2130]), .rectangle2_width(rectangle2_widths[2130]), .rectangle2_height(rectangle2_heights[2130]), .rectangle2_weight(rectangle2_weights[2130]), .rectangle3_x(rectangle3_xs[2130]), .rectangle3_y(rectangle3_ys[2130]), .rectangle3_width(rectangle3_widths[2130]), .rectangle3_height(rectangle3_heights[2130]), .rectangle3_weight(rectangle3_weights[2130]), .feature_threshold(feature_thresholds[2130]), .feature_above(feature_aboves[2130]), .feature_below(feature_belows[2130]), .scan_win_std_dev(scan_win_std_dev[2130]), .feature_accum(feature_accums[2130]));
  accum_calculator ac2131(.scan_win(scan_win2131), .rectangle1_x(rectangle1_xs[2131]), .rectangle1_y(rectangle1_ys[2131]), .rectangle1_width(rectangle1_widths[2131]), .rectangle1_height(rectangle1_heights[2131]), .rectangle1_weight(rectangle1_weights[2131]), .rectangle2_x(rectangle2_xs[2131]), .rectangle2_y(rectangle2_ys[2131]), .rectangle2_width(rectangle2_widths[2131]), .rectangle2_height(rectangle2_heights[2131]), .rectangle2_weight(rectangle2_weights[2131]), .rectangle3_x(rectangle3_xs[2131]), .rectangle3_y(rectangle3_ys[2131]), .rectangle3_width(rectangle3_widths[2131]), .rectangle3_height(rectangle3_heights[2131]), .rectangle3_weight(rectangle3_weights[2131]), .feature_threshold(feature_thresholds[2131]), .feature_above(feature_aboves[2131]), .feature_below(feature_belows[2131]), .scan_win_std_dev(scan_win_std_dev[2131]), .feature_accum(feature_accums[2131]));
  accum_calculator ac2132(.scan_win(scan_win2132), .rectangle1_x(rectangle1_xs[2132]), .rectangle1_y(rectangle1_ys[2132]), .rectangle1_width(rectangle1_widths[2132]), .rectangle1_height(rectangle1_heights[2132]), .rectangle1_weight(rectangle1_weights[2132]), .rectangle2_x(rectangle2_xs[2132]), .rectangle2_y(rectangle2_ys[2132]), .rectangle2_width(rectangle2_widths[2132]), .rectangle2_height(rectangle2_heights[2132]), .rectangle2_weight(rectangle2_weights[2132]), .rectangle3_x(rectangle3_xs[2132]), .rectangle3_y(rectangle3_ys[2132]), .rectangle3_width(rectangle3_widths[2132]), .rectangle3_height(rectangle3_heights[2132]), .rectangle3_weight(rectangle3_weights[2132]), .feature_threshold(feature_thresholds[2132]), .feature_above(feature_aboves[2132]), .feature_below(feature_belows[2132]), .scan_win_std_dev(scan_win_std_dev[2132]), .feature_accum(feature_accums[2132]));
  accum_calculator ac2133(.scan_win(scan_win2133), .rectangle1_x(rectangle1_xs[2133]), .rectangle1_y(rectangle1_ys[2133]), .rectangle1_width(rectangle1_widths[2133]), .rectangle1_height(rectangle1_heights[2133]), .rectangle1_weight(rectangle1_weights[2133]), .rectangle2_x(rectangle2_xs[2133]), .rectangle2_y(rectangle2_ys[2133]), .rectangle2_width(rectangle2_widths[2133]), .rectangle2_height(rectangle2_heights[2133]), .rectangle2_weight(rectangle2_weights[2133]), .rectangle3_x(rectangle3_xs[2133]), .rectangle3_y(rectangle3_ys[2133]), .rectangle3_width(rectangle3_widths[2133]), .rectangle3_height(rectangle3_heights[2133]), .rectangle3_weight(rectangle3_weights[2133]), .feature_threshold(feature_thresholds[2133]), .feature_above(feature_aboves[2133]), .feature_below(feature_belows[2133]), .scan_win_std_dev(scan_win_std_dev[2133]), .feature_accum(feature_accums[2133]));
  accum_calculator ac2134(.scan_win(scan_win2134), .rectangle1_x(rectangle1_xs[2134]), .rectangle1_y(rectangle1_ys[2134]), .rectangle1_width(rectangle1_widths[2134]), .rectangle1_height(rectangle1_heights[2134]), .rectangle1_weight(rectangle1_weights[2134]), .rectangle2_x(rectangle2_xs[2134]), .rectangle2_y(rectangle2_ys[2134]), .rectangle2_width(rectangle2_widths[2134]), .rectangle2_height(rectangle2_heights[2134]), .rectangle2_weight(rectangle2_weights[2134]), .rectangle3_x(rectangle3_xs[2134]), .rectangle3_y(rectangle3_ys[2134]), .rectangle3_width(rectangle3_widths[2134]), .rectangle3_height(rectangle3_heights[2134]), .rectangle3_weight(rectangle3_weights[2134]), .feature_threshold(feature_thresholds[2134]), .feature_above(feature_aboves[2134]), .feature_below(feature_belows[2134]), .scan_win_std_dev(scan_win_std_dev[2134]), .feature_accum(feature_accums[2134]));
  accum_calculator ac2135(.scan_win(scan_win2135), .rectangle1_x(rectangle1_xs[2135]), .rectangle1_y(rectangle1_ys[2135]), .rectangle1_width(rectangle1_widths[2135]), .rectangle1_height(rectangle1_heights[2135]), .rectangle1_weight(rectangle1_weights[2135]), .rectangle2_x(rectangle2_xs[2135]), .rectangle2_y(rectangle2_ys[2135]), .rectangle2_width(rectangle2_widths[2135]), .rectangle2_height(rectangle2_heights[2135]), .rectangle2_weight(rectangle2_weights[2135]), .rectangle3_x(rectangle3_xs[2135]), .rectangle3_y(rectangle3_ys[2135]), .rectangle3_width(rectangle3_widths[2135]), .rectangle3_height(rectangle3_heights[2135]), .rectangle3_weight(rectangle3_weights[2135]), .feature_threshold(feature_thresholds[2135]), .feature_above(feature_aboves[2135]), .feature_below(feature_belows[2135]), .scan_win_std_dev(scan_win_std_dev[2135]), .feature_accum(feature_accums[2135]));
  accum_calculator ac2136(.scan_win(scan_win2136), .rectangle1_x(rectangle1_xs[2136]), .rectangle1_y(rectangle1_ys[2136]), .rectangle1_width(rectangle1_widths[2136]), .rectangle1_height(rectangle1_heights[2136]), .rectangle1_weight(rectangle1_weights[2136]), .rectangle2_x(rectangle2_xs[2136]), .rectangle2_y(rectangle2_ys[2136]), .rectangle2_width(rectangle2_widths[2136]), .rectangle2_height(rectangle2_heights[2136]), .rectangle2_weight(rectangle2_weights[2136]), .rectangle3_x(rectangle3_xs[2136]), .rectangle3_y(rectangle3_ys[2136]), .rectangle3_width(rectangle3_widths[2136]), .rectangle3_height(rectangle3_heights[2136]), .rectangle3_weight(rectangle3_weights[2136]), .feature_threshold(feature_thresholds[2136]), .feature_above(feature_aboves[2136]), .feature_below(feature_belows[2136]), .scan_win_std_dev(scan_win_std_dev[2136]), .feature_accum(feature_accums[2136]));
  accum_calculator ac2137(.scan_win(scan_win2137), .rectangle1_x(rectangle1_xs[2137]), .rectangle1_y(rectangle1_ys[2137]), .rectangle1_width(rectangle1_widths[2137]), .rectangle1_height(rectangle1_heights[2137]), .rectangle1_weight(rectangle1_weights[2137]), .rectangle2_x(rectangle2_xs[2137]), .rectangle2_y(rectangle2_ys[2137]), .rectangle2_width(rectangle2_widths[2137]), .rectangle2_height(rectangle2_heights[2137]), .rectangle2_weight(rectangle2_weights[2137]), .rectangle3_x(rectangle3_xs[2137]), .rectangle3_y(rectangle3_ys[2137]), .rectangle3_width(rectangle3_widths[2137]), .rectangle3_height(rectangle3_heights[2137]), .rectangle3_weight(rectangle3_weights[2137]), .feature_threshold(feature_thresholds[2137]), .feature_above(feature_aboves[2137]), .feature_below(feature_belows[2137]), .scan_win_std_dev(scan_win_std_dev[2137]), .feature_accum(feature_accums[2137]));
  accum_calculator ac2138(.scan_win(scan_win2138), .rectangle1_x(rectangle1_xs[2138]), .rectangle1_y(rectangle1_ys[2138]), .rectangle1_width(rectangle1_widths[2138]), .rectangle1_height(rectangle1_heights[2138]), .rectangle1_weight(rectangle1_weights[2138]), .rectangle2_x(rectangle2_xs[2138]), .rectangle2_y(rectangle2_ys[2138]), .rectangle2_width(rectangle2_widths[2138]), .rectangle2_height(rectangle2_heights[2138]), .rectangle2_weight(rectangle2_weights[2138]), .rectangle3_x(rectangle3_xs[2138]), .rectangle3_y(rectangle3_ys[2138]), .rectangle3_width(rectangle3_widths[2138]), .rectangle3_height(rectangle3_heights[2138]), .rectangle3_weight(rectangle3_weights[2138]), .feature_threshold(feature_thresholds[2138]), .feature_above(feature_aboves[2138]), .feature_below(feature_belows[2138]), .scan_win_std_dev(scan_win_std_dev[2138]), .feature_accum(feature_accums[2138]));
  accum_calculator ac2139(.scan_win(scan_win2139), .rectangle1_x(rectangle1_xs[2139]), .rectangle1_y(rectangle1_ys[2139]), .rectangle1_width(rectangle1_widths[2139]), .rectangle1_height(rectangle1_heights[2139]), .rectangle1_weight(rectangle1_weights[2139]), .rectangle2_x(rectangle2_xs[2139]), .rectangle2_y(rectangle2_ys[2139]), .rectangle2_width(rectangle2_widths[2139]), .rectangle2_height(rectangle2_heights[2139]), .rectangle2_weight(rectangle2_weights[2139]), .rectangle3_x(rectangle3_xs[2139]), .rectangle3_y(rectangle3_ys[2139]), .rectangle3_width(rectangle3_widths[2139]), .rectangle3_height(rectangle3_heights[2139]), .rectangle3_weight(rectangle3_weights[2139]), .feature_threshold(feature_thresholds[2139]), .feature_above(feature_aboves[2139]), .feature_below(feature_belows[2139]), .scan_win_std_dev(scan_win_std_dev[2139]), .feature_accum(feature_accums[2139]));
  accum_calculator ac2140(.scan_win(scan_win2140), .rectangle1_x(rectangle1_xs[2140]), .rectangle1_y(rectangle1_ys[2140]), .rectangle1_width(rectangle1_widths[2140]), .rectangle1_height(rectangle1_heights[2140]), .rectangle1_weight(rectangle1_weights[2140]), .rectangle2_x(rectangle2_xs[2140]), .rectangle2_y(rectangle2_ys[2140]), .rectangle2_width(rectangle2_widths[2140]), .rectangle2_height(rectangle2_heights[2140]), .rectangle2_weight(rectangle2_weights[2140]), .rectangle3_x(rectangle3_xs[2140]), .rectangle3_y(rectangle3_ys[2140]), .rectangle3_width(rectangle3_widths[2140]), .rectangle3_height(rectangle3_heights[2140]), .rectangle3_weight(rectangle3_weights[2140]), .feature_threshold(feature_thresholds[2140]), .feature_above(feature_aboves[2140]), .feature_below(feature_belows[2140]), .scan_win_std_dev(scan_win_std_dev[2140]), .feature_accum(feature_accums[2140]));
  accum_calculator ac2141(.scan_win(scan_win2141), .rectangle1_x(rectangle1_xs[2141]), .rectangle1_y(rectangle1_ys[2141]), .rectangle1_width(rectangle1_widths[2141]), .rectangle1_height(rectangle1_heights[2141]), .rectangle1_weight(rectangle1_weights[2141]), .rectangle2_x(rectangle2_xs[2141]), .rectangle2_y(rectangle2_ys[2141]), .rectangle2_width(rectangle2_widths[2141]), .rectangle2_height(rectangle2_heights[2141]), .rectangle2_weight(rectangle2_weights[2141]), .rectangle3_x(rectangle3_xs[2141]), .rectangle3_y(rectangle3_ys[2141]), .rectangle3_width(rectangle3_widths[2141]), .rectangle3_height(rectangle3_heights[2141]), .rectangle3_weight(rectangle3_weights[2141]), .feature_threshold(feature_thresholds[2141]), .feature_above(feature_aboves[2141]), .feature_below(feature_belows[2141]), .scan_win_std_dev(scan_win_std_dev[2141]), .feature_accum(feature_accums[2141]));
  accum_calculator ac2142(.scan_win(scan_win2142), .rectangle1_x(rectangle1_xs[2142]), .rectangle1_y(rectangle1_ys[2142]), .rectangle1_width(rectangle1_widths[2142]), .rectangle1_height(rectangle1_heights[2142]), .rectangle1_weight(rectangle1_weights[2142]), .rectangle2_x(rectangle2_xs[2142]), .rectangle2_y(rectangle2_ys[2142]), .rectangle2_width(rectangle2_widths[2142]), .rectangle2_height(rectangle2_heights[2142]), .rectangle2_weight(rectangle2_weights[2142]), .rectangle3_x(rectangle3_xs[2142]), .rectangle3_y(rectangle3_ys[2142]), .rectangle3_width(rectangle3_widths[2142]), .rectangle3_height(rectangle3_heights[2142]), .rectangle3_weight(rectangle3_weights[2142]), .feature_threshold(feature_thresholds[2142]), .feature_above(feature_aboves[2142]), .feature_below(feature_belows[2142]), .scan_win_std_dev(scan_win_std_dev[2142]), .feature_accum(feature_accums[2142]));
  accum_calculator ac2143(.scan_win(scan_win2143), .rectangle1_x(rectangle1_xs[2143]), .rectangle1_y(rectangle1_ys[2143]), .rectangle1_width(rectangle1_widths[2143]), .rectangle1_height(rectangle1_heights[2143]), .rectangle1_weight(rectangle1_weights[2143]), .rectangle2_x(rectangle2_xs[2143]), .rectangle2_y(rectangle2_ys[2143]), .rectangle2_width(rectangle2_widths[2143]), .rectangle2_height(rectangle2_heights[2143]), .rectangle2_weight(rectangle2_weights[2143]), .rectangle3_x(rectangle3_xs[2143]), .rectangle3_y(rectangle3_ys[2143]), .rectangle3_width(rectangle3_widths[2143]), .rectangle3_height(rectangle3_heights[2143]), .rectangle3_weight(rectangle3_weights[2143]), .feature_threshold(feature_thresholds[2143]), .feature_above(feature_aboves[2143]), .feature_below(feature_belows[2143]), .scan_win_std_dev(scan_win_std_dev[2143]), .feature_accum(feature_accums[2143]));
  accum_calculator ac2144(.scan_win(scan_win2144), .rectangle1_x(rectangle1_xs[2144]), .rectangle1_y(rectangle1_ys[2144]), .rectangle1_width(rectangle1_widths[2144]), .rectangle1_height(rectangle1_heights[2144]), .rectangle1_weight(rectangle1_weights[2144]), .rectangle2_x(rectangle2_xs[2144]), .rectangle2_y(rectangle2_ys[2144]), .rectangle2_width(rectangle2_widths[2144]), .rectangle2_height(rectangle2_heights[2144]), .rectangle2_weight(rectangle2_weights[2144]), .rectangle3_x(rectangle3_xs[2144]), .rectangle3_y(rectangle3_ys[2144]), .rectangle3_width(rectangle3_widths[2144]), .rectangle3_height(rectangle3_heights[2144]), .rectangle3_weight(rectangle3_weights[2144]), .feature_threshold(feature_thresholds[2144]), .feature_above(feature_aboves[2144]), .feature_below(feature_belows[2144]), .scan_win_std_dev(scan_win_std_dev[2144]), .feature_accum(feature_accums[2144]));
  accum_calculator ac2145(.scan_win(scan_win2145), .rectangle1_x(rectangle1_xs[2145]), .rectangle1_y(rectangle1_ys[2145]), .rectangle1_width(rectangle1_widths[2145]), .rectangle1_height(rectangle1_heights[2145]), .rectangle1_weight(rectangle1_weights[2145]), .rectangle2_x(rectangle2_xs[2145]), .rectangle2_y(rectangle2_ys[2145]), .rectangle2_width(rectangle2_widths[2145]), .rectangle2_height(rectangle2_heights[2145]), .rectangle2_weight(rectangle2_weights[2145]), .rectangle3_x(rectangle3_xs[2145]), .rectangle3_y(rectangle3_ys[2145]), .rectangle3_width(rectangle3_widths[2145]), .rectangle3_height(rectangle3_heights[2145]), .rectangle3_weight(rectangle3_weights[2145]), .feature_threshold(feature_thresholds[2145]), .feature_above(feature_aboves[2145]), .feature_below(feature_belows[2145]), .scan_win_std_dev(scan_win_std_dev[2145]), .feature_accum(feature_accums[2145]));
  accum_calculator ac2146(.scan_win(scan_win2146), .rectangle1_x(rectangle1_xs[2146]), .rectangle1_y(rectangle1_ys[2146]), .rectangle1_width(rectangle1_widths[2146]), .rectangle1_height(rectangle1_heights[2146]), .rectangle1_weight(rectangle1_weights[2146]), .rectangle2_x(rectangle2_xs[2146]), .rectangle2_y(rectangle2_ys[2146]), .rectangle2_width(rectangle2_widths[2146]), .rectangle2_height(rectangle2_heights[2146]), .rectangle2_weight(rectangle2_weights[2146]), .rectangle3_x(rectangle3_xs[2146]), .rectangle3_y(rectangle3_ys[2146]), .rectangle3_width(rectangle3_widths[2146]), .rectangle3_height(rectangle3_heights[2146]), .rectangle3_weight(rectangle3_weights[2146]), .feature_threshold(feature_thresholds[2146]), .feature_above(feature_aboves[2146]), .feature_below(feature_belows[2146]), .scan_win_std_dev(scan_win_std_dev[2146]), .feature_accum(feature_accums[2146]));
  accum_calculator ac2147(.scan_win(scan_win2147), .rectangle1_x(rectangle1_xs[2147]), .rectangle1_y(rectangle1_ys[2147]), .rectangle1_width(rectangle1_widths[2147]), .rectangle1_height(rectangle1_heights[2147]), .rectangle1_weight(rectangle1_weights[2147]), .rectangle2_x(rectangle2_xs[2147]), .rectangle2_y(rectangle2_ys[2147]), .rectangle2_width(rectangle2_widths[2147]), .rectangle2_height(rectangle2_heights[2147]), .rectangle2_weight(rectangle2_weights[2147]), .rectangle3_x(rectangle3_xs[2147]), .rectangle3_y(rectangle3_ys[2147]), .rectangle3_width(rectangle3_widths[2147]), .rectangle3_height(rectangle3_heights[2147]), .rectangle3_weight(rectangle3_weights[2147]), .feature_threshold(feature_thresholds[2147]), .feature_above(feature_aboves[2147]), .feature_below(feature_belows[2147]), .scan_win_std_dev(scan_win_std_dev[2147]), .feature_accum(feature_accums[2147]));
  accum_calculator ac2148(.scan_win(scan_win2148), .rectangle1_x(rectangle1_xs[2148]), .rectangle1_y(rectangle1_ys[2148]), .rectangle1_width(rectangle1_widths[2148]), .rectangle1_height(rectangle1_heights[2148]), .rectangle1_weight(rectangle1_weights[2148]), .rectangle2_x(rectangle2_xs[2148]), .rectangle2_y(rectangle2_ys[2148]), .rectangle2_width(rectangle2_widths[2148]), .rectangle2_height(rectangle2_heights[2148]), .rectangle2_weight(rectangle2_weights[2148]), .rectangle3_x(rectangle3_xs[2148]), .rectangle3_y(rectangle3_ys[2148]), .rectangle3_width(rectangle3_widths[2148]), .rectangle3_height(rectangle3_heights[2148]), .rectangle3_weight(rectangle3_weights[2148]), .feature_threshold(feature_thresholds[2148]), .feature_above(feature_aboves[2148]), .feature_below(feature_belows[2148]), .scan_win_std_dev(scan_win_std_dev[2148]), .feature_accum(feature_accums[2148]));
  accum_calculator ac2149(.scan_win(scan_win2149), .rectangle1_x(rectangle1_xs[2149]), .rectangle1_y(rectangle1_ys[2149]), .rectangle1_width(rectangle1_widths[2149]), .rectangle1_height(rectangle1_heights[2149]), .rectangle1_weight(rectangle1_weights[2149]), .rectangle2_x(rectangle2_xs[2149]), .rectangle2_y(rectangle2_ys[2149]), .rectangle2_width(rectangle2_widths[2149]), .rectangle2_height(rectangle2_heights[2149]), .rectangle2_weight(rectangle2_weights[2149]), .rectangle3_x(rectangle3_xs[2149]), .rectangle3_y(rectangle3_ys[2149]), .rectangle3_width(rectangle3_widths[2149]), .rectangle3_height(rectangle3_heights[2149]), .rectangle3_weight(rectangle3_weights[2149]), .feature_threshold(feature_thresholds[2149]), .feature_above(feature_aboves[2149]), .feature_below(feature_belows[2149]), .scan_win_std_dev(scan_win_std_dev[2149]), .feature_accum(feature_accums[2149]));
  accum_calculator ac2150(.scan_win(scan_win2150), .rectangle1_x(rectangle1_xs[2150]), .rectangle1_y(rectangle1_ys[2150]), .rectangle1_width(rectangle1_widths[2150]), .rectangle1_height(rectangle1_heights[2150]), .rectangle1_weight(rectangle1_weights[2150]), .rectangle2_x(rectangle2_xs[2150]), .rectangle2_y(rectangle2_ys[2150]), .rectangle2_width(rectangle2_widths[2150]), .rectangle2_height(rectangle2_heights[2150]), .rectangle2_weight(rectangle2_weights[2150]), .rectangle3_x(rectangle3_xs[2150]), .rectangle3_y(rectangle3_ys[2150]), .rectangle3_width(rectangle3_widths[2150]), .rectangle3_height(rectangle3_heights[2150]), .rectangle3_weight(rectangle3_weights[2150]), .feature_threshold(feature_thresholds[2150]), .feature_above(feature_aboves[2150]), .feature_below(feature_belows[2150]), .scan_win_std_dev(scan_win_std_dev[2150]), .feature_accum(feature_accums[2150]));
  accum_calculator ac2151(.scan_win(scan_win2151), .rectangle1_x(rectangle1_xs[2151]), .rectangle1_y(rectangle1_ys[2151]), .rectangle1_width(rectangle1_widths[2151]), .rectangle1_height(rectangle1_heights[2151]), .rectangle1_weight(rectangle1_weights[2151]), .rectangle2_x(rectangle2_xs[2151]), .rectangle2_y(rectangle2_ys[2151]), .rectangle2_width(rectangle2_widths[2151]), .rectangle2_height(rectangle2_heights[2151]), .rectangle2_weight(rectangle2_weights[2151]), .rectangle3_x(rectangle3_xs[2151]), .rectangle3_y(rectangle3_ys[2151]), .rectangle3_width(rectangle3_widths[2151]), .rectangle3_height(rectangle3_heights[2151]), .rectangle3_weight(rectangle3_weights[2151]), .feature_threshold(feature_thresholds[2151]), .feature_above(feature_aboves[2151]), .feature_below(feature_belows[2151]), .scan_win_std_dev(scan_win_std_dev[2151]), .feature_accum(feature_accums[2151]));
  accum_calculator ac2152(.scan_win(scan_win2152), .rectangle1_x(rectangle1_xs[2152]), .rectangle1_y(rectangle1_ys[2152]), .rectangle1_width(rectangle1_widths[2152]), .rectangle1_height(rectangle1_heights[2152]), .rectangle1_weight(rectangle1_weights[2152]), .rectangle2_x(rectangle2_xs[2152]), .rectangle2_y(rectangle2_ys[2152]), .rectangle2_width(rectangle2_widths[2152]), .rectangle2_height(rectangle2_heights[2152]), .rectangle2_weight(rectangle2_weights[2152]), .rectangle3_x(rectangle3_xs[2152]), .rectangle3_y(rectangle3_ys[2152]), .rectangle3_width(rectangle3_widths[2152]), .rectangle3_height(rectangle3_heights[2152]), .rectangle3_weight(rectangle3_weights[2152]), .feature_threshold(feature_thresholds[2152]), .feature_above(feature_aboves[2152]), .feature_below(feature_belows[2152]), .scan_win_std_dev(scan_win_std_dev[2152]), .feature_accum(feature_accums[2152]));
  accum_calculator ac2153(.scan_win(scan_win2153), .rectangle1_x(rectangle1_xs[2153]), .rectangle1_y(rectangle1_ys[2153]), .rectangle1_width(rectangle1_widths[2153]), .rectangle1_height(rectangle1_heights[2153]), .rectangle1_weight(rectangle1_weights[2153]), .rectangle2_x(rectangle2_xs[2153]), .rectangle2_y(rectangle2_ys[2153]), .rectangle2_width(rectangle2_widths[2153]), .rectangle2_height(rectangle2_heights[2153]), .rectangle2_weight(rectangle2_weights[2153]), .rectangle3_x(rectangle3_xs[2153]), .rectangle3_y(rectangle3_ys[2153]), .rectangle3_width(rectangle3_widths[2153]), .rectangle3_height(rectangle3_heights[2153]), .rectangle3_weight(rectangle3_weights[2153]), .feature_threshold(feature_thresholds[2153]), .feature_above(feature_aboves[2153]), .feature_below(feature_belows[2153]), .scan_win_std_dev(scan_win_std_dev[2153]), .feature_accum(feature_accums[2153]));
  accum_calculator ac2154(.scan_win(scan_win2154), .rectangle1_x(rectangle1_xs[2154]), .rectangle1_y(rectangle1_ys[2154]), .rectangle1_width(rectangle1_widths[2154]), .rectangle1_height(rectangle1_heights[2154]), .rectangle1_weight(rectangle1_weights[2154]), .rectangle2_x(rectangle2_xs[2154]), .rectangle2_y(rectangle2_ys[2154]), .rectangle2_width(rectangle2_widths[2154]), .rectangle2_height(rectangle2_heights[2154]), .rectangle2_weight(rectangle2_weights[2154]), .rectangle3_x(rectangle3_xs[2154]), .rectangle3_y(rectangle3_ys[2154]), .rectangle3_width(rectangle3_widths[2154]), .rectangle3_height(rectangle3_heights[2154]), .rectangle3_weight(rectangle3_weights[2154]), .feature_threshold(feature_thresholds[2154]), .feature_above(feature_aboves[2154]), .feature_below(feature_belows[2154]), .scan_win_std_dev(scan_win_std_dev[2154]), .feature_accum(feature_accums[2154]));
  accum_calculator ac2155(.scan_win(scan_win2155), .rectangle1_x(rectangle1_xs[2155]), .rectangle1_y(rectangle1_ys[2155]), .rectangle1_width(rectangle1_widths[2155]), .rectangle1_height(rectangle1_heights[2155]), .rectangle1_weight(rectangle1_weights[2155]), .rectangle2_x(rectangle2_xs[2155]), .rectangle2_y(rectangle2_ys[2155]), .rectangle2_width(rectangle2_widths[2155]), .rectangle2_height(rectangle2_heights[2155]), .rectangle2_weight(rectangle2_weights[2155]), .rectangle3_x(rectangle3_xs[2155]), .rectangle3_y(rectangle3_ys[2155]), .rectangle3_width(rectangle3_widths[2155]), .rectangle3_height(rectangle3_heights[2155]), .rectangle3_weight(rectangle3_weights[2155]), .feature_threshold(feature_thresholds[2155]), .feature_above(feature_aboves[2155]), .feature_below(feature_belows[2155]), .scan_win_std_dev(scan_win_std_dev[2155]), .feature_accum(feature_accums[2155]));
  accum_calculator ac2156(.scan_win(scan_win2156), .rectangle1_x(rectangle1_xs[2156]), .rectangle1_y(rectangle1_ys[2156]), .rectangle1_width(rectangle1_widths[2156]), .rectangle1_height(rectangle1_heights[2156]), .rectangle1_weight(rectangle1_weights[2156]), .rectangle2_x(rectangle2_xs[2156]), .rectangle2_y(rectangle2_ys[2156]), .rectangle2_width(rectangle2_widths[2156]), .rectangle2_height(rectangle2_heights[2156]), .rectangle2_weight(rectangle2_weights[2156]), .rectangle3_x(rectangle3_xs[2156]), .rectangle3_y(rectangle3_ys[2156]), .rectangle3_width(rectangle3_widths[2156]), .rectangle3_height(rectangle3_heights[2156]), .rectangle3_weight(rectangle3_weights[2156]), .feature_threshold(feature_thresholds[2156]), .feature_above(feature_aboves[2156]), .feature_below(feature_belows[2156]), .scan_win_std_dev(scan_win_std_dev[2156]), .feature_accum(feature_accums[2156]));
  accum_calculator ac2157(.scan_win(scan_win2157), .rectangle1_x(rectangle1_xs[2157]), .rectangle1_y(rectangle1_ys[2157]), .rectangle1_width(rectangle1_widths[2157]), .rectangle1_height(rectangle1_heights[2157]), .rectangle1_weight(rectangle1_weights[2157]), .rectangle2_x(rectangle2_xs[2157]), .rectangle2_y(rectangle2_ys[2157]), .rectangle2_width(rectangle2_widths[2157]), .rectangle2_height(rectangle2_heights[2157]), .rectangle2_weight(rectangle2_weights[2157]), .rectangle3_x(rectangle3_xs[2157]), .rectangle3_y(rectangle3_ys[2157]), .rectangle3_width(rectangle3_widths[2157]), .rectangle3_height(rectangle3_heights[2157]), .rectangle3_weight(rectangle3_weights[2157]), .feature_threshold(feature_thresholds[2157]), .feature_above(feature_aboves[2157]), .feature_below(feature_belows[2157]), .scan_win_std_dev(scan_win_std_dev[2157]), .feature_accum(feature_accums[2157]));
  accum_calculator ac2158(.scan_win(scan_win2158), .rectangle1_x(rectangle1_xs[2158]), .rectangle1_y(rectangle1_ys[2158]), .rectangle1_width(rectangle1_widths[2158]), .rectangle1_height(rectangle1_heights[2158]), .rectangle1_weight(rectangle1_weights[2158]), .rectangle2_x(rectangle2_xs[2158]), .rectangle2_y(rectangle2_ys[2158]), .rectangle2_width(rectangle2_widths[2158]), .rectangle2_height(rectangle2_heights[2158]), .rectangle2_weight(rectangle2_weights[2158]), .rectangle3_x(rectangle3_xs[2158]), .rectangle3_y(rectangle3_ys[2158]), .rectangle3_width(rectangle3_widths[2158]), .rectangle3_height(rectangle3_heights[2158]), .rectangle3_weight(rectangle3_weights[2158]), .feature_threshold(feature_thresholds[2158]), .feature_above(feature_aboves[2158]), .feature_below(feature_belows[2158]), .scan_win_std_dev(scan_win_std_dev[2158]), .feature_accum(feature_accums[2158]));
  accum_calculator ac2159(.scan_win(scan_win2159), .rectangle1_x(rectangle1_xs[2159]), .rectangle1_y(rectangle1_ys[2159]), .rectangle1_width(rectangle1_widths[2159]), .rectangle1_height(rectangle1_heights[2159]), .rectangle1_weight(rectangle1_weights[2159]), .rectangle2_x(rectangle2_xs[2159]), .rectangle2_y(rectangle2_ys[2159]), .rectangle2_width(rectangle2_widths[2159]), .rectangle2_height(rectangle2_heights[2159]), .rectangle2_weight(rectangle2_weights[2159]), .rectangle3_x(rectangle3_xs[2159]), .rectangle3_y(rectangle3_ys[2159]), .rectangle3_width(rectangle3_widths[2159]), .rectangle3_height(rectangle3_heights[2159]), .rectangle3_weight(rectangle3_weights[2159]), .feature_threshold(feature_thresholds[2159]), .feature_above(feature_aboves[2159]), .feature_below(feature_belows[2159]), .scan_win_std_dev(scan_win_std_dev[2159]), .feature_accum(feature_accums[2159]));
  accum_calculator ac2160(.scan_win(scan_win2160), .rectangle1_x(rectangle1_xs[2160]), .rectangle1_y(rectangle1_ys[2160]), .rectangle1_width(rectangle1_widths[2160]), .rectangle1_height(rectangle1_heights[2160]), .rectangle1_weight(rectangle1_weights[2160]), .rectangle2_x(rectangle2_xs[2160]), .rectangle2_y(rectangle2_ys[2160]), .rectangle2_width(rectangle2_widths[2160]), .rectangle2_height(rectangle2_heights[2160]), .rectangle2_weight(rectangle2_weights[2160]), .rectangle3_x(rectangle3_xs[2160]), .rectangle3_y(rectangle3_ys[2160]), .rectangle3_width(rectangle3_widths[2160]), .rectangle3_height(rectangle3_heights[2160]), .rectangle3_weight(rectangle3_weights[2160]), .feature_threshold(feature_thresholds[2160]), .feature_above(feature_aboves[2160]), .feature_below(feature_belows[2160]), .scan_win_std_dev(scan_win_std_dev[2160]), .feature_accum(feature_accums[2160]));
  accum_calculator ac2161(.scan_win(scan_win2161), .rectangle1_x(rectangle1_xs[2161]), .rectangle1_y(rectangle1_ys[2161]), .rectangle1_width(rectangle1_widths[2161]), .rectangle1_height(rectangle1_heights[2161]), .rectangle1_weight(rectangle1_weights[2161]), .rectangle2_x(rectangle2_xs[2161]), .rectangle2_y(rectangle2_ys[2161]), .rectangle2_width(rectangle2_widths[2161]), .rectangle2_height(rectangle2_heights[2161]), .rectangle2_weight(rectangle2_weights[2161]), .rectangle3_x(rectangle3_xs[2161]), .rectangle3_y(rectangle3_ys[2161]), .rectangle3_width(rectangle3_widths[2161]), .rectangle3_height(rectangle3_heights[2161]), .rectangle3_weight(rectangle3_weights[2161]), .feature_threshold(feature_thresholds[2161]), .feature_above(feature_aboves[2161]), .feature_below(feature_belows[2161]), .scan_win_std_dev(scan_win_std_dev[2161]), .feature_accum(feature_accums[2161]));
  accum_calculator ac2162(.scan_win(scan_win2162), .rectangle1_x(rectangle1_xs[2162]), .rectangle1_y(rectangle1_ys[2162]), .rectangle1_width(rectangle1_widths[2162]), .rectangle1_height(rectangle1_heights[2162]), .rectangle1_weight(rectangle1_weights[2162]), .rectangle2_x(rectangle2_xs[2162]), .rectangle2_y(rectangle2_ys[2162]), .rectangle2_width(rectangle2_widths[2162]), .rectangle2_height(rectangle2_heights[2162]), .rectangle2_weight(rectangle2_weights[2162]), .rectangle3_x(rectangle3_xs[2162]), .rectangle3_y(rectangle3_ys[2162]), .rectangle3_width(rectangle3_widths[2162]), .rectangle3_height(rectangle3_heights[2162]), .rectangle3_weight(rectangle3_weights[2162]), .feature_threshold(feature_thresholds[2162]), .feature_above(feature_aboves[2162]), .feature_below(feature_belows[2162]), .scan_win_std_dev(scan_win_std_dev[2162]), .feature_accum(feature_accums[2162]));
  accum_calculator ac2163(.scan_win(scan_win2163), .rectangle1_x(rectangle1_xs[2163]), .rectangle1_y(rectangle1_ys[2163]), .rectangle1_width(rectangle1_widths[2163]), .rectangle1_height(rectangle1_heights[2163]), .rectangle1_weight(rectangle1_weights[2163]), .rectangle2_x(rectangle2_xs[2163]), .rectangle2_y(rectangle2_ys[2163]), .rectangle2_width(rectangle2_widths[2163]), .rectangle2_height(rectangle2_heights[2163]), .rectangle2_weight(rectangle2_weights[2163]), .rectangle3_x(rectangle3_xs[2163]), .rectangle3_y(rectangle3_ys[2163]), .rectangle3_width(rectangle3_widths[2163]), .rectangle3_height(rectangle3_heights[2163]), .rectangle3_weight(rectangle3_weights[2163]), .feature_threshold(feature_thresholds[2163]), .feature_above(feature_aboves[2163]), .feature_below(feature_belows[2163]), .scan_win_std_dev(scan_win_std_dev[2163]), .feature_accum(feature_accums[2163]));
  accum_calculator ac2164(.scan_win(scan_win2164), .rectangle1_x(rectangle1_xs[2164]), .rectangle1_y(rectangle1_ys[2164]), .rectangle1_width(rectangle1_widths[2164]), .rectangle1_height(rectangle1_heights[2164]), .rectangle1_weight(rectangle1_weights[2164]), .rectangle2_x(rectangle2_xs[2164]), .rectangle2_y(rectangle2_ys[2164]), .rectangle2_width(rectangle2_widths[2164]), .rectangle2_height(rectangle2_heights[2164]), .rectangle2_weight(rectangle2_weights[2164]), .rectangle3_x(rectangle3_xs[2164]), .rectangle3_y(rectangle3_ys[2164]), .rectangle3_width(rectangle3_widths[2164]), .rectangle3_height(rectangle3_heights[2164]), .rectangle3_weight(rectangle3_weights[2164]), .feature_threshold(feature_thresholds[2164]), .feature_above(feature_aboves[2164]), .feature_below(feature_belows[2164]), .scan_win_std_dev(scan_win_std_dev[2164]), .feature_accum(feature_accums[2164]));
  accum_calculator ac2165(.scan_win(scan_win2165), .rectangle1_x(rectangle1_xs[2165]), .rectangle1_y(rectangle1_ys[2165]), .rectangle1_width(rectangle1_widths[2165]), .rectangle1_height(rectangle1_heights[2165]), .rectangle1_weight(rectangle1_weights[2165]), .rectangle2_x(rectangle2_xs[2165]), .rectangle2_y(rectangle2_ys[2165]), .rectangle2_width(rectangle2_widths[2165]), .rectangle2_height(rectangle2_heights[2165]), .rectangle2_weight(rectangle2_weights[2165]), .rectangle3_x(rectangle3_xs[2165]), .rectangle3_y(rectangle3_ys[2165]), .rectangle3_width(rectangle3_widths[2165]), .rectangle3_height(rectangle3_heights[2165]), .rectangle3_weight(rectangle3_weights[2165]), .feature_threshold(feature_thresholds[2165]), .feature_above(feature_aboves[2165]), .feature_below(feature_belows[2165]), .scan_win_std_dev(scan_win_std_dev[2165]), .feature_accum(feature_accums[2165]));
  accum_calculator ac2166(.scan_win(scan_win2166), .rectangle1_x(rectangle1_xs[2166]), .rectangle1_y(rectangle1_ys[2166]), .rectangle1_width(rectangle1_widths[2166]), .rectangle1_height(rectangle1_heights[2166]), .rectangle1_weight(rectangle1_weights[2166]), .rectangle2_x(rectangle2_xs[2166]), .rectangle2_y(rectangle2_ys[2166]), .rectangle2_width(rectangle2_widths[2166]), .rectangle2_height(rectangle2_heights[2166]), .rectangle2_weight(rectangle2_weights[2166]), .rectangle3_x(rectangle3_xs[2166]), .rectangle3_y(rectangle3_ys[2166]), .rectangle3_width(rectangle3_widths[2166]), .rectangle3_height(rectangle3_heights[2166]), .rectangle3_weight(rectangle3_weights[2166]), .feature_threshold(feature_thresholds[2166]), .feature_above(feature_aboves[2166]), .feature_below(feature_belows[2166]), .scan_win_std_dev(scan_win_std_dev[2166]), .feature_accum(feature_accums[2166]));
  accum_calculator ac2167(.scan_win(scan_win2167), .rectangle1_x(rectangle1_xs[2167]), .rectangle1_y(rectangle1_ys[2167]), .rectangle1_width(rectangle1_widths[2167]), .rectangle1_height(rectangle1_heights[2167]), .rectangle1_weight(rectangle1_weights[2167]), .rectangle2_x(rectangle2_xs[2167]), .rectangle2_y(rectangle2_ys[2167]), .rectangle2_width(rectangle2_widths[2167]), .rectangle2_height(rectangle2_heights[2167]), .rectangle2_weight(rectangle2_weights[2167]), .rectangle3_x(rectangle3_xs[2167]), .rectangle3_y(rectangle3_ys[2167]), .rectangle3_width(rectangle3_widths[2167]), .rectangle3_height(rectangle3_heights[2167]), .rectangle3_weight(rectangle3_weights[2167]), .feature_threshold(feature_thresholds[2167]), .feature_above(feature_aboves[2167]), .feature_below(feature_belows[2167]), .scan_win_std_dev(scan_win_std_dev[2167]), .feature_accum(feature_accums[2167]));
  accum_calculator ac2168(.scan_win(scan_win2168), .rectangle1_x(rectangle1_xs[2168]), .rectangle1_y(rectangle1_ys[2168]), .rectangle1_width(rectangle1_widths[2168]), .rectangle1_height(rectangle1_heights[2168]), .rectangle1_weight(rectangle1_weights[2168]), .rectangle2_x(rectangle2_xs[2168]), .rectangle2_y(rectangle2_ys[2168]), .rectangle2_width(rectangle2_widths[2168]), .rectangle2_height(rectangle2_heights[2168]), .rectangle2_weight(rectangle2_weights[2168]), .rectangle3_x(rectangle3_xs[2168]), .rectangle3_y(rectangle3_ys[2168]), .rectangle3_width(rectangle3_widths[2168]), .rectangle3_height(rectangle3_heights[2168]), .rectangle3_weight(rectangle3_weights[2168]), .feature_threshold(feature_thresholds[2168]), .feature_above(feature_aboves[2168]), .feature_below(feature_belows[2168]), .scan_win_std_dev(scan_win_std_dev[2168]), .feature_accum(feature_accums[2168]));
  accum_calculator ac2169(.scan_win(scan_win2169), .rectangle1_x(rectangle1_xs[2169]), .rectangle1_y(rectangle1_ys[2169]), .rectangle1_width(rectangle1_widths[2169]), .rectangle1_height(rectangle1_heights[2169]), .rectangle1_weight(rectangle1_weights[2169]), .rectangle2_x(rectangle2_xs[2169]), .rectangle2_y(rectangle2_ys[2169]), .rectangle2_width(rectangle2_widths[2169]), .rectangle2_height(rectangle2_heights[2169]), .rectangle2_weight(rectangle2_weights[2169]), .rectangle3_x(rectangle3_xs[2169]), .rectangle3_y(rectangle3_ys[2169]), .rectangle3_width(rectangle3_widths[2169]), .rectangle3_height(rectangle3_heights[2169]), .rectangle3_weight(rectangle3_weights[2169]), .feature_threshold(feature_thresholds[2169]), .feature_above(feature_aboves[2169]), .feature_below(feature_belows[2169]), .scan_win_std_dev(scan_win_std_dev[2169]), .feature_accum(feature_accums[2169]));
  accum_calculator ac2170(.scan_win(scan_win2170), .rectangle1_x(rectangle1_xs[2170]), .rectangle1_y(rectangle1_ys[2170]), .rectangle1_width(rectangle1_widths[2170]), .rectangle1_height(rectangle1_heights[2170]), .rectangle1_weight(rectangle1_weights[2170]), .rectangle2_x(rectangle2_xs[2170]), .rectangle2_y(rectangle2_ys[2170]), .rectangle2_width(rectangle2_widths[2170]), .rectangle2_height(rectangle2_heights[2170]), .rectangle2_weight(rectangle2_weights[2170]), .rectangle3_x(rectangle3_xs[2170]), .rectangle3_y(rectangle3_ys[2170]), .rectangle3_width(rectangle3_widths[2170]), .rectangle3_height(rectangle3_heights[2170]), .rectangle3_weight(rectangle3_weights[2170]), .feature_threshold(feature_thresholds[2170]), .feature_above(feature_aboves[2170]), .feature_below(feature_belows[2170]), .scan_win_std_dev(scan_win_std_dev[2170]), .feature_accum(feature_accums[2170]));
  accum_calculator ac2171(.scan_win(scan_win2171), .rectangle1_x(rectangle1_xs[2171]), .rectangle1_y(rectangle1_ys[2171]), .rectangle1_width(rectangle1_widths[2171]), .rectangle1_height(rectangle1_heights[2171]), .rectangle1_weight(rectangle1_weights[2171]), .rectangle2_x(rectangle2_xs[2171]), .rectangle2_y(rectangle2_ys[2171]), .rectangle2_width(rectangle2_widths[2171]), .rectangle2_height(rectangle2_heights[2171]), .rectangle2_weight(rectangle2_weights[2171]), .rectangle3_x(rectangle3_xs[2171]), .rectangle3_y(rectangle3_ys[2171]), .rectangle3_width(rectangle3_widths[2171]), .rectangle3_height(rectangle3_heights[2171]), .rectangle3_weight(rectangle3_weights[2171]), .feature_threshold(feature_thresholds[2171]), .feature_above(feature_aboves[2171]), .feature_below(feature_belows[2171]), .scan_win_std_dev(scan_win_std_dev[2171]), .feature_accum(feature_accums[2171]));
  accum_calculator ac2172(.scan_win(scan_win2172), .rectangle1_x(rectangle1_xs[2172]), .rectangle1_y(rectangle1_ys[2172]), .rectangle1_width(rectangle1_widths[2172]), .rectangle1_height(rectangle1_heights[2172]), .rectangle1_weight(rectangle1_weights[2172]), .rectangle2_x(rectangle2_xs[2172]), .rectangle2_y(rectangle2_ys[2172]), .rectangle2_width(rectangle2_widths[2172]), .rectangle2_height(rectangle2_heights[2172]), .rectangle2_weight(rectangle2_weights[2172]), .rectangle3_x(rectangle3_xs[2172]), .rectangle3_y(rectangle3_ys[2172]), .rectangle3_width(rectangle3_widths[2172]), .rectangle3_height(rectangle3_heights[2172]), .rectangle3_weight(rectangle3_weights[2172]), .feature_threshold(feature_thresholds[2172]), .feature_above(feature_aboves[2172]), .feature_below(feature_belows[2172]), .scan_win_std_dev(scan_win_std_dev[2172]), .feature_accum(feature_accums[2172]));
  accum_calculator ac2173(.scan_win(scan_win2173), .rectangle1_x(rectangle1_xs[2173]), .rectangle1_y(rectangle1_ys[2173]), .rectangle1_width(rectangle1_widths[2173]), .rectangle1_height(rectangle1_heights[2173]), .rectangle1_weight(rectangle1_weights[2173]), .rectangle2_x(rectangle2_xs[2173]), .rectangle2_y(rectangle2_ys[2173]), .rectangle2_width(rectangle2_widths[2173]), .rectangle2_height(rectangle2_heights[2173]), .rectangle2_weight(rectangle2_weights[2173]), .rectangle3_x(rectangle3_xs[2173]), .rectangle3_y(rectangle3_ys[2173]), .rectangle3_width(rectangle3_widths[2173]), .rectangle3_height(rectangle3_heights[2173]), .rectangle3_weight(rectangle3_weights[2173]), .feature_threshold(feature_thresholds[2173]), .feature_above(feature_aboves[2173]), .feature_below(feature_belows[2173]), .scan_win_std_dev(scan_win_std_dev[2173]), .feature_accum(feature_accums[2173]));
  accum_calculator ac2174(.scan_win(scan_win2174), .rectangle1_x(rectangle1_xs[2174]), .rectangle1_y(rectangle1_ys[2174]), .rectangle1_width(rectangle1_widths[2174]), .rectangle1_height(rectangle1_heights[2174]), .rectangle1_weight(rectangle1_weights[2174]), .rectangle2_x(rectangle2_xs[2174]), .rectangle2_y(rectangle2_ys[2174]), .rectangle2_width(rectangle2_widths[2174]), .rectangle2_height(rectangle2_heights[2174]), .rectangle2_weight(rectangle2_weights[2174]), .rectangle3_x(rectangle3_xs[2174]), .rectangle3_y(rectangle3_ys[2174]), .rectangle3_width(rectangle3_widths[2174]), .rectangle3_height(rectangle3_heights[2174]), .rectangle3_weight(rectangle3_weights[2174]), .feature_threshold(feature_thresholds[2174]), .feature_above(feature_aboves[2174]), .feature_below(feature_belows[2174]), .scan_win_std_dev(scan_win_std_dev[2174]), .feature_accum(feature_accums[2174]));
  accum_calculator ac2175(.scan_win(scan_win2175), .rectangle1_x(rectangle1_xs[2175]), .rectangle1_y(rectangle1_ys[2175]), .rectangle1_width(rectangle1_widths[2175]), .rectangle1_height(rectangle1_heights[2175]), .rectangle1_weight(rectangle1_weights[2175]), .rectangle2_x(rectangle2_xs[2175]), .rectangle2_y(rectangle2_ys[2175]), .rectangle2_width(rectangle2_widths[2175]), .rectangle2_height(rectangle2_heights[2175]), .rectangle2_weight(rectangle2_weights[2175]), .rectangle3_x(rectangle3_xs[2175]), .rectangle3_y(rectangle3_ys[2175]), .rectangle3_width(rectangle3_widths[2175]), .rectangle3_height(rectangle3_heights[2175]), .rectangle3_weight(rectangle3_weights[2175]), .feature_threshold(feature_thresholds[2175]), .feature_above(feature_aboves[2175]), .feature_below(feature_belows[2175]), .scan_win_std_dev(scan_win_std_dev[2175]), .feature_accum(feature_accums[2175]));
  accum_calculator ac2176(.scan_win(scan_win2176), .rectangle1_x(rectangle1_xs[2176]), .rectangle1_y(rectangle1_ys[2176]), .rectangle1_width(rectangle1_widths[2176]), .rectangle1_height(rectangle1_heights[2176]), .rectangle1_weight(rectangle1_weights[2176]), .rectangle2_x(rectangle2_xs[2176]), .rectangle2_y(rectangle2_ys[2176]), .rectangle2_width(rectangle2_widths[2176]), .rectangle2_height(rectangle2_heights[2176]), .rectangle2_weight(rectangle2_weights[2176]), .rectangle3_x(rectangle3_xs[2176]), .rectangle3_y(rectangle3_ys[2176]), .rectangle3_width(rectangle3_widths[2176]), .rectangle3_height(rectangle3_heights[2176]), .rectangle3_weight(rectangle3_weights[2176]), .feature_threshold(feature_thresholds[2176]), .feature_above(feature_aboves[2176]), .feature_below(feature_belows[2176]), .scan_win_std_dev(scan_win_std_dev[2176]), .feature_accum(feature_accums[2176]));
  accum_calculator ac2177(.scan_win(scan_win2177), .rectangle1_x(rectangle1_xs[2177]), .rectangle1_y(rectangle1_ys[2177]), .rectangle1_width(rectangle1_widths[2177]), .rectangle1_height(rectangle1_heights[2177]), .rectangle1_weight(rectangle1_weights[2177]), .rectangle2_x(rectangle2_xs[2177]), .rectangle2_y(rectangle2_ys[2177]), .rectangle2_width(rectangle2_widths[2177]), .rectangle2_height(rectangle2_heights[2177]), .rectangle2_weight(rectangle2_weights[2177]), .rectangle3_x(rectangle3_xs[2177]), .rectangle3_y(rectangle3_ys[2177]), .rectangle3_width(rectangle3_widths[2177]), .rectangle3_height(rectangle3_heights[2177]), .rectangle3_weight(rectangle3_weights[2177]), .feature_threshold(feature_thresholds[2177]), .feature_above(feature_aboves[2177]), .feature_below(feature_belows[2177]), .scan_win_std_dev(scan_win_std_dev[2177]), .feature_accum(feature_accums[2177]));
  accum_calculator ac2178(.scan_win(scan_win2178), .rectangle1_x(rectangle1_xs[2178]), .rectangle1_y(rectangle1_ys[2178]), .rectangle1_width(rectangle1_widths[2178]), .rectangle1_height(rectangle1_heights[2178]), .rectangle1_weight(rectangle1_weights[2178]), .rectangle2_x(rectangle2_xs[2178]), .rectangle2_y(rectangle2_ys[2178]), .rectangle2_width(rectangle2_widths[2178]), .rectangle2_height(rectangle2_heights[2178]), .rectangle2_weight(rectangle2_weights[2178]), .rectangle3_x(rectangle3_xs[2178]), .rectangle3_y(rectangle3_ys[2178]), .rectangle3_width(rectangle3_widths[2178]), .rectangle3_height(rectangle3_heights[2178]), .rectangle3_weight(rectangle3_weights[2178]), .feature_threshold(feature_thresholds[2178]), .feature_above(feature_aboves[2178]), .feature_below(feature_belows[2178]), .scan_win_std_dev(scan_win_std_dev[2178]), .feature_accum(feature_accums[2178]));
  accum_calculator ac2179(.scan_win(scan_win2179), .rectangle1_x(rectangle1_xs[2179]), .rectangle1_y(rectangle1_ys[2179]), .rectangle1_width(rectangle1_widths[2179]), .rectangle1_height(rectangle1_heights[2179]), .rectangle1_weight(rectangle1_weights[2179]), .rectangle2_x(rectangle2_xs[2179]), .rectangle2_y(rectangle2_ys[2179]), .rectangle2_width(rectangle2_widths[2179]), .rectangle2_height(rectangle2_heights[2179]), .rectangle2_weight(rectangle2_weights[2179]), .rectangle3_x(rectangle3_xs[2179]), .rectangle3_y(rectangle3_ys[2179]), .rectangle3_width(rectangle3_widths[2179]), .rectangle3_height(rectangle3_heights[2179]), .rectangle3_weight(rectangle3_weights[2179]), .feature_threshold(feature_thresholds[2179]), .feature_above(feature_aboves[2179]), .feature_below(feature_belows[2179]), .scan_win_std_dev(scan_win_std_dev[2179]), .feature_accum(feature_accums[2179]));
  accum_calculator ac2180(.scan_win(scan_win2180), .rectangle1_x(rectangle1_xs[2180]), .rectangle1_y(rectangle1_ys[2180]), .rectangle1_width(rectangle1_widths[2180]), .rectangle1_height(rectangle1_heights[2180]), .rectangle1_weight(rectangle1_weights[2180]), .rectangle2_x(rectangle2_xs[2180]), .rectangle2_y(rectangle2_ys[2180]), .rectangle2_width(rectangle2_widths[2180]), .rectangle2_height(rectangle2_heights[2180]), .rectangle2_weight(rectangle2_weights[2180]), .rectangle3_x(rectangle3_xs[2180]), .rectangle3_y(rectangle3_ys[2180]), .rectangle3_width(rectangle3_widths[2180]), .rectangle3_height(rectangle3_heights[2180]), .rectangle3_weight(rectangle3_weights[2180]), .feature_threshold(feature_thresholds[2180]), .feature_above(feature_aboves[2180]), .feature_below(feature_belows[2180]), .scan_win_std_dev(scan_win_std_dev[2180]), .feature_accum(feature_accums[2180]));
  accum_calculator ac2181(.scan_win(scan_win2181), .rectangle1_x(rectangle1_xs[2181]), .rectangle1_y(rectangle1_ys[2181]), .rectangle1_width(rectangle1_widths[2181]), .rectangle1_height(rectangle1_heights[2181]), .rectangle1_weight(rectangle1_weights[2181]), .rectangle2_x(rectangle2_xs[2181]), .rectangle2_y(rectangle2_ys[2181]), .rectangle2_width(rectangle2_widths[2181]), .rectangle2_height(rectangle2_heights[2181]), .rectangle2_weight(rectangle2_weights[2181]), .rectangle3_x(rectangle3_xs[2181]), .rectangle3_y(rectangle3_ys[2181]), .rectangle3_width(rectangle3_widths[2181]), .rectangle3_height(rectangle3_heights[2181]), .rectangle3_weight(rectangle3_weights[2181]), .feature_threshold(feature_thresholds[2181]), .feature_above(feature_aboves[2181]), .feature_below(feature_belows[2181]), .scan_win_std_dev(scan_win_std_dev[2181]), .feature_accum(feature_accums[2181]));
  accum_calculator ac2182(.scan_win(scan_win2182), .rectangle1_x(rectangle1_xs[2182]), .rectangle1_y(rectangle1_ys[2182]), .rectangle1_width(rectangle1_widths[2182]), .rectangle1_height(rectangle1_heights[2182]), .rectangle1_weight(rectangle1_weights[2182]), .rectangle2_x(rectangle2_xs[2182]), .rectangle2_y(rectangle2_ys[2182]), .rectangle2_width(rectangle2_widths[2182]), .rectangle2_height(rectangle2_heights[2182]), .rectangle2_weight(rectangle2_weights[2182]), .rectangle3_x(rectangle3_xs[2182]), .rectangle3_y(rectangle3_ys[2182]), .rectangle3_width(rectangle3_widths[2182]), .rectangle3_height(rectangle3_heights[2182]), .rectangle3_weight(rectangle3_weights[2182]), .feature_threshold(feature_thresholds[2182]), .feature_above(feature_aboves[2182]), .feature_below(feature_belows[2182]), .scan_win_std_dev(scan_win_std_dev[2182]), .feature_accum(feature_accums[2182]));
  accum_calculator ac2183(.scan_win(scan_win2183), .rectangle1_x(rectangle1_xs[2183]), .rectangle1_y(rectangle1_ys[2183]), .rectangle1_width(rectangle1_widths[2183]), .rectangle1_height(rectangle1_heights[2183]), .rectangle1_weight(rectangle1_weights[2183]), .rectangle2_x(rectangle2_xs[2183]), .rectangle2_y(rectangle2_ys[2183]), .rectangle2_width(rectangle2_widths[2183]), .rectangle2_height(rectangle2_heights[2183]), .rectangle2_weight(rectangle2_weights[2183]), .rectangle3_x(rectangle3_xs[2183]), .rectangle3_y(rectangle3_ys[2183]), .rectangle3_width(rectangle3_widths[2183]), .rectangle3_height(rectangle3_heights[2183]), .rectangle3_weight(rectangle3_weights[2183]), .feature_threshold(feature_thresholds[2183]), .feature_above(feature_aboves[2183]), .feature_below(feature_belows[2183]), .scan_win_std_dev(scan_win_std_dev[2183]), .feature_accum(feature_accums[2183]));
  accum_calculator ac2184(.scan_win(scan_win2184), .rectangle1_x(rectangle1_xs[2184]), .rectangle1_y(rectangle1_ys[2184]), .rectangle1_width(rectangle1_widths[2184]), .rectangle1_height(rectangle1_heights[2184]), .rectangle1_weight(rectangle1_weights[2184]), .rectangle2_x(rectangle2_xs[2184]), .rectangle2_y(rectangle2_ys[2184]), .rectangle2_width(rectangle2_widths[2184]), .rectangle2_height(rectangle2_heights[2184]), .rectangle2_weight(rectangle2_weights[2184]), .rectangle3_x(rectangle3_xs[2184]), .rectangle3_y(rectangle3_ys[2184]), .rectangle3_width(rectangle3_widths[2184]), .rectangle3_height(rectangle3_heights[2184]), .rectangle3_weight(rectangle3_weights[2184]), .feature_threshold(feature_thresholds[2184]), .feature_above(feature_aboves[2184]), .feature_below(feature_belows[2184]), .scan_win_std_dev(scan_win_std_dev[2184]), .feature_accum(feature_accums[2184]));
  accum_calculator ac2185(.scan_win(scan_win2185), .rectangle1_x(rectangle1_xs[2185]), .rectangle1_y(rectangle1_ys[2185]), .rectangle1_width(rectangle1_widths[2185]), .rectangle1_height(rectangle1_heights[2185]), .rectangle1_weight(rectangle1_weights[2185]), .rectangle2_x(rectangle2_xs[2185]), .rectangle2_y(rectangle2_ys[2185]), .rectangle2_width(rectangle2_widths[2185]), .rectangle2_height(rectangle2_heights[2185]), .rectangle2_weight(rectangle2_weights[2185]), .rectangle3_x(rectangle3_xs[2185]), .rectangle3_y(rectangle3_ys[2185]), .rectangle3_width(rectangle3_widths[2185]), .rectangle3_height(rectangle3_heights[2185]), .rectangle3_weight(rectangle3_weights[2185]), .feature_threshold(feature_thresholds[2185]), .feature_above(feature_aboves[2185]), .feature_below(feature_belows[2185]), .scan_win_std_dev(scan_win_std_dev[2185]), .feature_accum(feature_accums[2185]));
  accum_calculator ac2186(.scan_win(scan_win2186), .rectangle1_x(rectangle1_xs[2186]), .rectangle1_y(rectangle1_ys[2186]), .rectangle1_width(rectangle1_widths[2186]), .rectangle1_height(rectangle1_heights[2186]), .rectangle1_weight(rectangle1_weights[2186]), .rectangle2_x(rectangle2_xs[2186]), .rectangle2_y(rectangle2_ys[2186]), .rectangle2_width(rectangle2_widths[2186]), .rectangle2_height(rectangle2_heights[2186]), .rectangle2_weight(rectangle2_weights[2186]), .rectangle3_x(rectangle3_xs[2186]), .rectangle3_y(rectangle3_ys[2186]), .rectangle3_width(rectangle3_widths[2186]), .rectangle3_height(rectangle3_heights[2186]), .rectangle3_weight(rectangle3_weights[2186]), .feature_threshold(feature_thresholds[2186]), .feature_above(feature_aboves[2186]), .feature_below(feature_belows[2186]), .scan_win_std_dev(scan_win_std_dev[2186]), .feature_accum(feature_accums[2186]));
  accum_calculator ac2187(.scan_win(scan_win2187), .rectangle1_x(rectangle1_xs[2187]), .rectangle1_y(rectangle1_ys[2187]), .rectangle1_width(rectangle1_widths[2187]), .rectangle1_height(rectangle1_heights[2187]), .rectangle1_weight(rectangle1_weights[2187]), .rectangle2_x(rectangle2_xs[2187]), .rectangle2_y(rectangle2_ys[2187]), .rectangle2_width(rectangle2_widths[2187]), .rectangle2_height(rectangle2_heights[2187]), .rectangle2_weight(rectangle2_weights[2187]), .rectangle3_x(rectangle3_xs[2187]), .rectangle3_y(rectangle3_ys[2187]), .rectangle3_width(rectangle3_widths[2187]), .rectangle3_height(rectangle3_heights[2187]), .rectangle3_weight(rectangle3_weights[2187]), .feature_threshold(feature_thresholds[2187]), .feature_above(feature_aboves[2187]), .feature_below(feature_belows[2187]), .scan_win_std_dev(scan_win_std_dev[2187]), .feature_accum(feature_accums[2187]));
  accum_calculator ac2188(.scan_win(scan_win2188), .rectangle1_x(rectangle1_xs[2188]), .rectangle1_y(rectangle1_ys[2188]), .rectangle1_width(rectangle1_widths[2188]), .rectangle1_height(rectangle1_heights[2188]), .rectangle1_weight(rectangle1_weights[2188]), .rectangle2_x(rectangle2_xs[2188]), .rectangle2_y(rectangle2_ys[2188]), .rectangle2_width(rectangle2_widths[2188]), .rectangle2_height(rectangle2_heights[2188]), .rectangle2_weight(rectangle2_weights[2188]), .rectangle3_x(rectangle3_xs[2188]), .rectangle3_y(rectangle3_ys[2188]), .rectangle3_width(rectangle3_widths[2188]), .rectangle3_height(rectangle3_heights[2188]), .rectangle3_weight(rectangle3_weights[2188]), .feature_threshold(feature_thresholds[2188]), .feature_above(feature_aboves[2188]), .feature_below(feature_belows[2188]), .scan_win_std_dev(scan_win_std_dev[2188]), .feature_accum(feature_accums[2188]));
  accum_calculator ac2189(.scan_win(scan_win2189), .rectangle1_x(rectangle1_xs[2189]), .rectangle1_y(rectangle1_ys[2189]), .rectangle1_width(rectangle1_widths[2189]), .rectangle1_height(rectangle1_heights[2189]), .rectangle1_weight(rectangle1_weights[2189]), .rectangle2_x(rectangle2_xs[2189]), .rectangle2_y(rectangle2_ys[2189]), .rectangle2_width(rectangle2_widths[2189]), .rectangle2_height(rectangle2_heights[2189]), .rectangle2_weight(rectangle2_weights[2189]), .rectangle3_x(rectangle3_xs[2189]), .rectangle3_y(rectangle3_ys[2189]), .rectangle3_width(rectangle3_widths[2189]), .rectangle3_height(rectangle3_heights[2189]), .rectangle3_weight(rectangle3_weights[2189]), .feature_threshold(feature_thresholds[2189]), .feature_above(feature_aboves[2189]), .feature_below(feature_belows[2189]), .scan_win_std_dev(scan_win_std_dev[2189]), .feature_accum(feature_accums[2189]));
  accum_calculator ac2190(.scan_win(scan_win2190), .rectangle1_x(rectangle1_xs[2190]), .rectangle1_y(rectangle1_ys[2190]), .rectangle1_width(rectangle1_widths[2190]), .rectangle1_height(rectangle1_heights[2190]), .rectangle1_weight(rectangle1_weights[2190]), .rectangle2_x(rectangle2_xs[2190]), .rectangle2_y(rectangle2_ys[2190]), .rectangle2_width(rectangle2_widths[2190]), .rectangle2_height(rectangle2_heights[2190]), .rectangle2_weight(rectangle2_weights[2190]), .rectangle3_x(rectangle3_xs[2190]), .rectangle3_y(rectangle3_ys[2190]), .rectangle3_width(rectangle3_widths[2190]), .rectangle3_height(rectangle3_heights[2190]), .rectangle3_weight(rectangle3_weights[2190]), .feature_threshold(feature_thresholds[2190]), .feature_above(feature_aboves[2190]), .feature_below(feature_belows[2190]), .scan_win_std_dev(scan_win_std_dev[2190]), .feature_accum(feature_accums[2190]));
  accum_calculator ac2191(.scan_win(scan_win2191), .rectangle1_x(rectangle1_xs[2191]), .rectangle1_y(rectangle1_ys[2191]), .rectangle1_width(rectangle1_widths[2191]), .rectangle1_height(rectangle1_heights[2191]), .rectangle1_weight(rectangle1_weights[2191]), .rectangle2_x(rectangle2_xs[2191]), .rectangle2_y(rectangle2_ys[2191]), .rectangle2_width(rectangle2_widths[2191]), .rectangle2_height(rectangle2_heights[2191]), .rectangle2_weight(rectangle2_weights[2191]), .rectangle3_x(rectangle3_xs[2191]), .rectangle3_y(rectangle3_ys[2191]), .rectangle3_width(rectangle3_widths[2191]), .rectangle3_height(rectangle3_heights[2191]), .rectangle3_weight(rectangle3_weights[2191]), .feature_threshold(feature_thresholds[2191]), .feature_above(feature_aboves[2191]), .feature_below(feature_belows[2191]), .scan_win_std_dev(scan_win_std_dev[2191]), .feature_accum(feature_accums[2191]));
  accum_calculator ac2192(.scan_win(scan_win2192), .rectangle1_x(rectangle1_xs[2192]), .rectangle1_y(rectangle1_ys[2192]), .rectangle1_width(rectangle1_widths[2192]), .rectangle1_height(rectangle1_heights[2192]), .rectangle1_weight(rectangle1_weights[2192]), .rectangle2_x(rectangle2_xs[2192]), .rectangle2_y(rectangle2_ys[2192]), .rectangle2_width(rectangle2_widths[2192]), .rectangle2_height(rectangle2_heights[2192]), .rectangle2_weight(rectangle2_weights[2192]), .rectangle3_x(rectangle3_xs[2192]), .rectangle3_y(rectangle3_ys[2192]), .rectangle3_width(rectangle3_widths[2192]), .rectangle3_height(rectangle3_heights[2192]), .rectangle3_weight(rectangle3_weights[2192]), .feature_threshold(feature_thresholds[2192]), .feature_above(feature_aboves[2192]), .feature_below(feature_belows[2192]), .scan_win_std_dev(scan_win_std_dev[2192]), .feature_accum(feature_accums[2192]));
  accum_calculator ac2193(.scan_win(scan_win2193), .rectangle1_x(rectangle1_xs[2193]), .rectangle1_y(rectangle1_ys[2193]), .rectangle1_width(rectangle1_widths[2193]), .rectangle1_height(rectangle1_heights[2193]), .rectangle1_weight(rectangle1_weights[2193]), .rectangle2_x(rectangle2_xs[2193]), .rectangle2_y(rectangle2_ys[2193]), .rectangle2_width(rectangle2_widths[2193]), .rectangle2_height(rectangle2_heights[2193]), .rectangle2_weight(rectangle2_weights[2193]), .rectangle3_x(rectangle3_xs[2193]), .rectangle3_y(rectangle3_ys[2193]), .rectangle3_width(rectangle3_widths[2193]), .rectangle3_height(rectangle3_heights[2193]), .rectangle3_weight(rectangle3_weights[2193]), .feature_threshold(feature_thresholds[2193]), .feature_above(feature_aboves[2193]), .feature_below(feature_belows[2193]), .scan_win_std_dev(scan_win_std_dev[2193]), .feature_accum(feature_accums[2193]));
  accum_calculator ac2194(.scan_win(scan_win2194), .rectangle1_x(rectangle1_xs[2194]), .rectangle1_y(rectangle1_ys[2194]), .rectangle1_width(rectangle1_widths[2194]), .rectangle1_height(rectangle1_heights[2194]), .rectangle1_weight(rectangle1_weights[2194]), .rectangle2_x(rectangle2_xs[2194]), .rectangle2_y(rectangle2_ys[2194]), .rectangle2_width(rectangle2_widths[2194]), .rectangle2_height(rectangle2_heights[2194]), .rectangle2_weight(rectangle2_weights[2194]), .rectangle3_x(rectangle3_xs[2194]), .rectangle3_y(rectangle3_ys[2194]), .rectangle3_width(rectangle3_widths[2194]), .rectangle3_height(rectangle3_heights[2194]), .rectangle3_weight(rectangle3_weights[2194]), .feature_threshold(feature_thresholds[2194]), .feature_above(feature_aboves[2194]), .feature_below(feature_belows[2194]), .scan_win_std_dev(scan_win_std_dev[2194]), .feature_accum(feature_accums[2194]));
  accum_calculator ac2195(.scan_win(scan_win2195), .rectangle1_x(rectangle1_xs[2195]), .rectangle1_y(rectangle1_ys[2195]), .rectangle1_width(rectangle1_widths[2195]), .rectangle1_height(rectangle1_heights[2195]), .rectangle1_weight(rectangle1_weights[2195]), .rectangle2_x(rectangle2_xs[2195]), .rectangle2_y(rectangle2_ys[2195]), .rectangle2_width(rectangle2_widths[2195]), .rectangle2_height(rectangle2_heights[2195]), .rectangle2_weight(rectangle2_weights[2195]), .rectangle3_x(rectangle3_xs[2195]), .rectangle3_y(rectangle3_ys[2195]), .rectangle3_width(rectangle3_widths[2195]), .rectangle3_height(rectangle3_heights[2195]), .rectangle3_weight(rectangle3_weights[2195]), .feature_threshold(feature_thresholds[2195]), .feature_above(feature_aboves[2195]), .feature_below(feature_belows[2195]), .scan_win_std_dev(scan_win_std_dev[2195]), .feature_accum(feature_accums[2195]));
  accum_calculator ac2196(.scan_win(scan_win2196), .rectangle1_x(rectangle1_xs[2196]), .rectangle1_y(rectangle1_ys[2196]), .rectangle1_width(rectangle1_widths[2196]), .rectangle1_height(rectangle1_heights[2196]), .rectangle1_weight(rectangle1_weights[2196]), .rectangle2_x(rectangle2_xs[2196]), .rectangle2_y(rectangle2_ys[2196]), .rectangle2_width(rectangle2_widths[2196]), .rectangle2_height(rectangle2_heights[2196]), .rectangle2_weight(rectangle2_weights[2196]), .rectangle3_x(rectangle3_xs[2196]), .rectangle3_y(rectangle3_ys[2196]), .rectangle3_width(rectangle3_widths[2196]), .rectangle3_height(rectangle3_heights[2196]), .rectangle3_weight(rectangle3_weights[2196]), .feature_threshold(feature_thresholds[2196]), .feature_above(feature_aboves[2196]), .feature_below(feature_belows[2196]), .scan_win_std_dev(scan_win_std_dev[2196]), .feature_accum(feature_accums[2196]));
  accum_calculator ac2197(.scan_win(scan_win2197), .rectangle1_x(rectangle1_xs[2197]), .rectangle1_y(rectangle1_ys[2197]), .rectangle1_width(rectangle1_widths[2197]), .rectangle1_height(rectangle1_heights[2197]), .rectangle1_weight(rectangle1_weights[2197]), .rectangle2_x(rectangle2_xs[2197]), .rectangle2_y(rectangle2_ys[2197]), .rectangle2_width(rectangle2_widths[2197]), .rectangle2_height(rectangle2_heights[2197]), .rectangle2_weight(rectangle2_weights[2197]), .rectangle3_x(rectangle3_xs[2197]), .rectangle3_y(rectangle3_ys[2197]), .rectangle3_width(rectangle3_widths[2197]), .rectangle3_height(rectangle3_heights[2197]), .rectangle3_weight(rectangle3_weights[2197]), .feature_threshold(feature_thresholds[2197]), .feature_above(feature_aboves[2197]), .feature_below(feature_belows[2197]), .scan_win_std_dev(scan_win_std_dev[2197]), .feature_accum(feature_accums[2197]));
  accum_calculator ac2198(.scan_win(scan_win2198), .rectangle1_x(rectangle1_xs[2198]), .rectangle1_y(rectangle1_ys[2198]), .rectangle1_width(rectangle1_widths[2198]), .rectangle1_height(rectangle1_heights[2198]), .rectangle1_weight(rectangle1_weights[2198]), .rectangle2_x(rectangle2_xs[2198]), .rectangle2_y(rectangle2_ys[2198]), .rectangle2_width(rectangle2_widths[2198]), .rectangle2_height(rectangle2_heights[2198]), .rectangle2_weight(rectangle2_weights[2198]), .rectangle3_x(rectangle3_xs[2198]), .rectangle3_y(rectangle3_ys[2198]), .rectangle3_width(rectangle3_widths[2198]), .rectangle3_height(rectangle3_heights[2198]), .rectangle3_weight(rectangle3_weights[2198]), .feature_threshold(feature_thresholds[2198]), .feature_above(feature_aboves[2198]), .feature_below(feature_belows[2198]), .scan_win_std_dev(scan_win_std_dev[2198]), .feature_accum(feature_accums[2198]));
  accum_calculator ac2199(.scan_win(scan_win2199), .rectangle1_x(rectangle1_xs[2199]), .rectangle1_y(rectangle1_ys[2199]), .rectangle1_width(rectangle1_widths[2199]), .rectangle1_height(rectangle1_heights[2199]), .rectangle1_weight(rectangle1_weights[2199]), .rectangle2_x(rectangle2_xs[2199]), .rectangle2_y(rectangle2_ys[2199]), .rectangle2_width(rectangle2_widths[2199]), .rectangle2_height(rectangle2_heights[2199]), .rectangle2_weight(rectangle2_weights[2199]), .rectangle3_x(rectangle3_xs[2199]), .rectangle3_y(rectangle3_ys[2199]), .rectangle3_width(rectangle3_widths[2199]), .rectangle3_height(rectangle3_heights[2199]), .rectangle3_weight(rectangle3_weights[2199]), .feature_threshold(feature_thresholds[2199]), .feature_above(feature_aboves[2199]), .feature_below(feature_belows[2199]), .scan_win_std_dev(scan_win_std_dev[2199]), .feature_accum(feature_accums[2199]));
  accum_calculator ac2200(.scan_win(scan_win2200), .rectangle1_x(rectangle1_xs[2200]), .rectangle1_y(rectangle1_ys[2200]), .rectangle1_width(rectangle1_widths[2200]), .rectangle1_height(rectangle1_heights[2200]), .rectangle1_weight(rectangle1_weights[2200]), .rectangle2_x(rectangle2_xs[2200]), .rectangle2_y(rectangle2_ys[2200]), .rectangle2_width(rectangle2_widths[2200]), .rectangle2_height(rectangle2_heights[2200]), .rectangle2_weight(rectangle2_weights[2200]), .rectangle3_x(rectangle3_xs[2200]), .rectangle3_y(rectangle3_ys[2200]), .rectangle3_width(rectangle3_widths[2200]), .rectangle3_height(rectangle3_heights[2200]), .rectangle3_weight(rectangle3_weights[2200]), .feature_threshold(feature_thresholds[2200]), .feature_above(feature_aboves[2200]), .feature_below(feature_belows[2200]), .scan_win_std_dev(scan_win_std_dev[2200]), .feature_accum(feature_accums[2200]));
  accum_calculator ac2201(.scan_win(scan_win2201), .rectangle1_x(rectangle1_xs[2201]), .rectangle1_y(rectangle1_ys[2201]), .rectangle1_width(rectangle1_widths[2201]), .rectangle1_height(rectangle1_heights[2201]), .rectangle1_weight(rectangle1_weights[2201]), .rectangle2_x(rectangle2_xs[2201]), .rectangle2_y(rectangle2_ys[2201]), .rectangle2_width(rectangle2_widths[2201]), .rectangle2_height(rectangle2_heights[2201]), .rectangle2_weight(rectangle2_weights[2201]), .rectangle3_x(rectangle3_xs[2201]), .rectangle3_y(rectangle3_ys[2201]), .rectangle3_width(rectangle3_widths[2201]), .rectangle3_height(rectangle3_heights[2201]), .rectangle3_weight(rectangle3_weights[2201]), .feature_threshold(feature_thresholds[2201]), .feature_above(feature_aboves[2201]), .feature_below(feature_belows[2201]), .scan_win_std_dev(scan_win_std_dev[2201]), .feature_accum(feature_accums[2201]));
  accum_calculator ac2202(.scan_win(scan_win2202), .rectangle1_x(rectangle1_xs[2202]), .rectangle1_y(rectangle1_ys[2202]), .rectangle1_width(rectangle1_widths[2202]), .rectangle1_height(rectangle1_heights[2202]), .rectangle1_weight(rectangle1_weights[2202]), .rectangle2_x(rectangle2_xs[2202]), .rectangle2_y(rectangle2_ys[2202]), .rectangle2_width(rectangle2_widths[2202]), .rectangle2_height(rectangle2_heights[2202]), .rectangle2_weight(rectangle2_weights[2202]), .rectangle3_x(rectangle3_xs[2202]), .rectangle3_y(rectangle3_ys[2202]), .rectangle3_width(rectangle3_widths[2202]), .rectangle3_height(rectangle3_heights[2202]), .rectangle3_weight(rectangle3_weights[2202]), .feature_threshold(feature_thresholds[2202]), .feature_above(feature_aboves[2202]), .feature_below(feature_belows[2202]), .scan_win_std_dev(scan_win_std_dev[2202]), .feature_accum(feature_accums[2202]));
  accum_calculator ac2203(.scan_win(scan_win2203), .rectangle1_x(rectangle1_xs[2203]), .rectangle1_y(rectangle1_ys[2203]), .rectangle1_width(rectangle1_widths[2203]), .rectangle1_height(rectangle1_heights[2203]), .rectangle1_weight(rectangle1_weights[2203]), .rectangle2_x(rectangle2_xs[2203]), .rectangle2_y(rectangle2_ys[2203]), .rectangle2_width(rectangle2_widths[2203]), .rectangle2_height(rectangle2_heights[2203]), .rectangle2_weight(rectangle2_weights[2203]), .rectangle3_x(rectangle3_xs[2203]), .rectangle3_y(rectangle3_ys[2203]), .rectangle3_width(rectangle3_widths[2203]), .rectangle3_height(rectangle3_heights[2203]), .rectangle3_weight(rectangle3_weights[2203]), .feature_threshold(feature_thresholds[2203]), .feature_above(feature_aboves[2203]), .feature_below(feature_belows[2203]), .scan_win_std_dev(scan_win_std_dev[2203]), .feature_accum(feature_accums[2203]));
  accum_calculator ac2204(.scan_win(scan_win2204), .rectangle1_x(rectangle1_xs[2204]), .rectangle1_y(rectangle1_ys[2204]), .rectangle1_width(rectangle1_widths[2204]), .rectangle1_height(rectangle1_heights[2204]), .rectangle1_weight(rectangle1_weights[2204]), .rectangle2_x(rectangle2_xs[2204]), .rectangle2_y(rectangle2_ys[2204]), .rectangle2_width(rectangle2_widths[2204]), .rectangle2_height(rectangle2_heights[2204]), .rectangle2_weight(rectangle2_weights[2204]), .rectangle3_x(rectangle3_xs[2204]), .rectangle3_y(rectangle3_ys[2204]), .rectangle3_width(rectangle3_widths[2204]), .rectangle3_height(rectangle3_heights[2204]), .rectangle3_weight(rectangle3_weights[2204]), .feature_threshold(feature_thresholds[2204]), .feature_above(feature_aboves[2204]), .feature_below(feature_belows[2204]), .scan_win_std_dev(scan_win_std_dev[2204]), .feature_accum(feature_accums[2204]));
  accum_calculator ac2205(.scan_win(scan_win2205), .rectangle1_x(rectangle1_xs[2205]), .rectangle1_y(rectangle1_ys[2205]), .rectangle1_width(rectangle1_widths[2205]), .rectangle1_height(rectangle1_heights[2205]), .rectangle1_weight(rectangle1_weights[2205]), .rectangle2_x(rectangle2_xs[2205]), .rectangle2_y(rectangle2_ys[2205]), .rectangle2_width(rectangle2_widths[2205]), .rectangle2_height(rectangle2_heights[2205]), .rectangle2_weight(rectangle2_weights[2205]), .rectangle3_x(rectangle3_xs[2205]), .rectangle3_y(rectangle3_ys[2205]), .rectangle3_width(rectangle3_widths[2205]), .rectangle3_height(rectangle3_heights[2205]), .rectangle3_weight(rectangle3_weights[2205]), .feature_threshold(feature_thresholds[2205]), .feature_above(feature_aboves[2205]), .feature_below(feature_belows[2205]), .scan_win_std_dev(scan_win_std_dev[2205]), .feature_accum(feature_accums[2205]));
  accum_calculator ac2206(.scan_win(scan_win2206), .rectangle1_x(rectangle1_xs[2206]), .rectangle1_y(rectangle1_ys[2206]), .rectangle1_width(rectangle1_widths[2206]), .rectangle1_height(rectangle1_heights[2206]), .rectangle1_weight(rectangle1_weights[2206]), .rectangle2_x(rectangle2_xs[2206]), .rectangle2_y(rectangle2_ys[2206]), .rectangle2_width(rectangle2_widths[2206]), .rectangle2_height(rectangle2_heights[2206]), .rectangle2_weight(rectangle2_weights[2206]), .rectangle3_x(rectangle3_xs[2206]), .rectangle3_y(rectangle3_ys[2206]), .rectangle3_width(rectangle3_widths[2206]), .rectangle3_height(rectangle3_heights[2206]), .rectangle3_weight(rectangle3_weights[2206]), .feature_threshold(feature_thresholds[2206]), .feature_above(feature_aboves[2206]), .feature_below(feature_belows[2206]), .scan_win_std_dev(scan_win_std_dev[2206]), .feature_accum(feature_accums[2206]));
  accum_calculator ac2207(.scan_win(scan_win2207), .rectangle1_x(rectangle1_xs[2207]), .rectangle1_y(rectangle1_ys[2207]), .rectangle1_width(rectangle1_widths[2207]), .rectangle1_height(rectangle1_heights[2207]), .rectangle1_weight(rectangle1_weights[2207]), .rectangle2_x(rectangle2_xs[2207]), .rectangle2_y(rectangle2_ys[2207]), .rectangle2_width(rectangle2_widths[2207]), .rectangle2_height(rectangle2_heights[2207]), .rectangle2_weight(rectangle2_weights[2207]), .rectangle3_x(rectangle3_xs[2207]), .rectangle3_y(rectangle3_ys[2207]), .rectangle3_width(rectangle3_widths[2207]), .rectangle3_height(rectangle3_heights[2207]), .rectangle3_weight(rectangle3_weights[2207]), .feature_threshold(feature_thresholds[2207]), .feature_above(feature_aboves[2207]), .feature_below(feature_belows[2207]), .scan_win_std_dev(scan_win_std_dev[2207]), .feature_accum(feature_accums[2207]));
  accum_calculator ac2208(.scan_win(scan_win2208), .rectangle1_x(rectangle1_xs[2208]), .rectangle1_y(rectangle1_ys[2208]), .rectangle1_width(rectangle1_widths[2208]), .rectangle1_height(rectangle1_heights[2208]), .rectangle1_weight(rectangle1_weights[2208]), .rectangle2_x(rectangle2_xs[2208]), .rectangle2_y(rectangle2_ys[2208]), .rectangle2_width(rectangle2_widths[2208]), .rectangle2_height(rectangle2_heights[2208]), .rectangle2_weight(rectangle2_weights[2208]), .rectangle3_x(rectangle3_xs[2208]), .rectangle3_y(rectangle3_ys[2208]), .rectangle3_width(rectangle3_widths[2208]), .rectangle3_height(rectangle3_heights[2208]), .rectangle3_weight(rectangle3_weights[2208]), .feature_threshold(feature_thresholds[2208]), .feature_above(feature_aboves[2208]), .feature_below(feature_belows[2208]), .scan_win_std_dev(scan_win_std_dev[2208]), .feature_accum(feature_accums[2208]));
  accum_calculator ac2209(.scan_win(scan_win2209), .rectangle1_x(rectangle1_xs[2209]), .rectangle1_y(rectangle1_ys[2209]), .rectangle1_width(rectangle1_widths[2209]), .rectangle1_height(rectangle1_heights[2209]), .rectangle1_weight(rectangle1_weights[2209]), .rectangle2_x(rectangle2_xs[2209]), .rectangle2_y(rectangle2_ys[2209]), .rectangle2_width(rectangle2_widths[2209]), .rectangle2_height(rectangle2_heights[2209]), .rectangle2_weight(rectangle2_weights[2209]), .rectangle3_x(rectangle3_xs[2209]), .rectangle3_y(rectangle3_ys[2209]), .rectangle3_width(rectangle3_widths[2209]), .rectangle3_height(rectangle3_heights[2209]), .rectangle3_weight(rectangle3_weights[2209]), .feature_threshold(feature_thresholds[2209]), .feature_above(feature_aboves[2209]), .feature_below(feature_belows[2209]), .scan_win_std_dev(scan_win_std_dev[2209]), .feature_accum(feature_accums[2209]));
  accum_calculator ac2210(.scan_win(scan_win2210), .rectangle1_x(rectangle1_xs[2210]), .rectangle1_y(rectangle1_ys[2210]), .rectangle1_width(rectangle1_widths[2210]), .rectangle1_height(rectangle1_heights[2210]), .rectangle1_weight(rectangle1_weights[2210]), .rectangle2_x(rectangle2_xs[2210]), .rectangle2_y(rectangle2_ys[2210]), .rectangle2_width(rectangle2_widths[2210]), .rectangle2_height(rectangle2_heights[2210]), .rectangle2_weight(rectangle2_weights[2210]), .rectangle3_x(rectangle3_xs[2210]), .rectangle3_y(rectangle3_ys[2210]), .rectangle3_width(rectangle3_widths[2210]), .rectangle3_height(rectangle3_heights[2210]), .rectangle3_weight(rectangle3_weights[2210]), .feature_threshold(feature_thresholds[2210]), .feature_above(feature_aboves[2210]), .feature_below(feature_belows[2210]), .scan_win_std_dev(scan_win_std_dev[2210]), .feature_accum(feature_accums[2210]));
  accum_calculator ac2211(.scan_win(scan_win2211), .rectangle1_x(rectangle1_xs[2211]), .rectangle1_y(rectangle1_ys[2211]), .rectangle1_width(rectangle1_widths[2211]), .rectangle1_height(rectangle1_heights[2211]), .rectangle1_weight(rectangle1_weights[2211]), .rectangle2_x(rectangle2_xs[2211]), .rectangle2_y(rectangle2_ys[2211]), .rectangle2_width(rectangle2_widths[2211]), .rectangle2_height(rectangle2_heights[2211]), .rectangle2_weight(rectangle2_weights[2211]), .rectangle3_x(rectangle3_xs[2211]), .rectangle3_y(rectangle3_ys[2211]), .rectangle3_width(rectangle3_widths[2211]), .rectangle3_height(rectangle3_heights[2211]), .rectangle3_weight(rectangle3_weights[2211]), .feature_threshold(feature_thresholds[2211]), .feature_above(feature_aboves[2211]), .feature_below(feature_belows[2211]), .scan_win_std_dev(scan_win_std_dev[2211]), .feature_accum(feature_accums[2211]));
  accum_calculator ac2212(.scan_win(scan_win2212), .rectangle1_x(rectangle1_xs[2212]), .rectangle1_y(rectangle1_ys[2212]), .rectangle1_width(rectangle1_widths[2212]), .rectangle1_height(rectangle1_heights[2212]), .rectangle1_weight(rectangle1_weights[2212]), .rectangle2_x(rectangle2_xs[2212]), .rectangle2_y(rectangle2_ys[2212]), .rectangle2_width(rectangle2_widths[2212]), .rectangle2_height(rectangle2_heights[2212]), .rectangle2_weight(rectangle2_weights[2212]), .rectangle3_x(rectangle3_xs[2212]), .rectangle3_y(rectangle3_ys[2212]), .rectangle3_width(rectangle3_widths[2212]), .rectangle3_height(rectangle3_heights[2212]), .rectangle3_weight(rectangle3_weights[2212]), .feature_threshold(feature_thresholds[2212]), .feature_above(feature_aboves[2212]), .feature_below(feature_belows[2212]), .scan_win_std_dev(scan_win_std_dev[2212]), .feature_accum(feature_accums[2212]));
  accum_calculator ac2213(.scan_win(scan_win2213), .rectangle1_x(rectangle1_xs[2213]), .rectangle1_y(rectangle1_ys[2213]), .rectangle1_width(rectangle1_widths[2213]), .rectangle1_height(rectangle1_heights[2213]), .rectangle1_weight(rectangle1_weights[2213]), .rectangle2_x(rectangle2_xs[2213]), .rectangle2_y(rectangle2_ys[2213]), .rectangle2_width(rectangle2_widths[2213]), .rectangle2_height(rectangle2_heights[2213]), .rectangle2_weight(rectangle2_weights[2213]), .rectangle3_x(rectangle3_xs[2213]), .rectangle3_y(rectangle3_ys[2213]), .rectangle3_width(rectangle3_widths[2213]), .rectangle3_height(rectangle3_heights[2213]), .rectangle3_weight(rectangle3_weights[2213]), .feature_threshold(feature_thresholds[2213]), .feature_above(feature_aboves[2213]), .feature_below(feature_belows[2213]), .scan_win_std_dev(scan_win_std_dev[2213]), .feature_accum(feature_accums[2213]));
  accum_calculator ac2214(.scan_win(scan_win2214), .rectangle1_x(rectangle1_xs[2214]), .rectangle1_y(rectangle1_ys[2214]), .rectangle1_width(rectangle1_widths[2214]), .rectangle1_height(rectangle1_heights[2214]), .rectangle1_weight(rectangle1_weights[2214]), .rectangle2_x(rectangle2_xs[2214]), .rectangle2_y(rectangle2_ys[2214]), .rectangle2_width(rectangle2_widths[2214]), .rectangle2_height(rectangle2_heights[2214]), .rectangle2_weight(rectangle2_weights[2214]), .rectangle3_x(rectangle3_xs[2214]), .rectangle3_y(rectangle3_ys[2214]), .rectangle3_width(rectangle3_widths[2214]), .rectangle3_height(rectangle3_heights[2214]), .rectangle3_weight(rectangle3_weights[2214]), .feature_threshold(feature_thresholds[2214]), .feature_above(feature_aboves[2214]), .feature_below(feature_belows[2214]), .scan_win_std_dev(scan_win_std_dev[2214]), .feature_accum(feature_accums[2214]));
  accum_calculator ac2215(.scan_win(scan_win2215), .rectangle1_x(rectangle1_xs[2215]), .rectangle1_y(rectangle1_ys[2215]), .rectangle1_width(rectangle1_widths[2215]), .rectangle1_height(rectangle1_heights[2215]), .rectangle1_weight(rectangle1_weights[2215]), .rectangle2_x(rectangle2_xs[2215]), .rectangle2_y(rectangle2_ys[2215]), .rectangle2_width(rectangle2_widths[2215]), .rectangle2_height(rectangle2_heights[2215]), .rectangle2_weight(rectangle2_weights[2215]), .rectangle3_x(rectangle3_xs[2215]), .rectangle3_y(rectangle3_ys[2215]), .rectangle3_width(rectangle3_widths[2215]), .rectangle3_height(rectangle3_heights[2215]), .rectangle3_weight(rectangle3_weights[2215]), .feature_threshold(feature_thresholds[2215]), .feature_above(feature_aboves[2215]), .feature_below(feature_belows[2215]), .scan_win_std_dev(scan_win_std_dev[2215]), .feature_accum(feature_accums[2215]));
  accum_calculator ac2216(.scan_win(scan_win2216), .rectangle1_x(rectangle1_xs[2216]), .rectangle1_y(rectangle1_ys[2216]), .rectangle1_width(rectangle1_widths[2216]), .rectangle1_height(rectangle1_heights[2216]), .rectangle1_weight(rectangle1_weights[2216]), .rectangle2_x(rectangle2_xs[2216]), .rectangle2_y(rectangle2_ys[2216]), .rectangle2_width(rectangle2_widths[2216]), .rectangle2_height(rectangle2_heights[2216]), .rectangle2_weight(rectangle2_weights[2216]), .rectangle3_x(rectangle3_xs[2216]), .rectangle3_y(rectangle3_ys[2216]), .rectangle3_width(rectangle3_widths[2216]), .rectangle3_height(rectangle3_heights[2216]), .rectangle3_weight(rectangle3_weights[2216]), .feature_threshold(feature_thresholds[2216]), .feature_above(feature_aboves[2216]), .feature_below(feature_belows[2216]), .scan_win_std_dev(scan_win_std_dev[2216]), .feature_accum(feature_accums[2216]));
  accum_calculator ac2217(.scan_win(scan_win2217), .rectangle1_x(rectangle1_xs[2217]), .rectangle1_y(rectangle1_ys[2217]), .rectangle1_width(rectangle1_widths[2217]), .rectangle1_height(rectangle1_heights[2217]), .rectangle1_weight(rectangle1_weights[2217]), .rectangle2_x(rectangle2_xs[2217]), .rectangle2_y(rectangle2_ys[2217]), .rectangle2_width(rectangle2_widths[2217]), .rectangle2_height(rectangle2_heights[2217]), .rectangle2_weight(rectangle2_weights[2217]), .rectangle3_x(rectangle3_xs[2217]), .rectangle3_y(rectangle3_ys[2217]), .rectangle3_width(rectangle3_widths[2217]), .rectangle3_height(rectangle3_heights[2217]), .rectangle3_weight(rectangle3_weights[2217]), .feature_threshold(feature_thresholds[2217]), .feature_above(feature_aboves[2217]), .feature_below(feature_belows[2217]), .scan_win_std_dev(scan_win_std_dev[2217]), .feature_accum(feature_accums[2217]));
  accum_calculator ac2218(.scan_win(scan_win2218), .rectangle1_x(rectangle1_xs[2218]), .rectangle1_y(rectangle1_ys[2218]), .rectangle1_width(rectangle1_widths[2218]), .rectangle1_height(rectangle1_heights[2218]), .rectangle1_weight(rectangle1_weights[2218]), .rectangle2_x(rectangle2_xs[2218]), .rectangle2_y(rectangle2_ys[2218]), .rectangle2_width(rectangle2_widths[2218]), .rectangle2_height(rectangle2_heights[2218]), .rectangle2_weight(rectangle2_weights[2218]), .rectangle3_x(rectangle3_xs[2218]), .rectangle3_y(rectangle3_ys[2218]), .rectangle3_width(rectangle3_widths[2218]), .rectangle3_height(rectangle3_heights[2218]), .rectangle3_weight(rectangle3_weights[2218]), .feature_threshold(feature_thresholds[2218]), .feature_above(feature_aboves[2218]), .feature_below(feature_belows[2218]), .scan_win_std_dev(scan_win_std_dev[2218]), .feature_accum(feature_accums[2218]));
  accum_calculator ac2219(.scan_win(scan_win2219), .rectangle1_x(rectangle1_xs[2219]), .rectangle1_y(rectangle1_ys[2219]), .rectangle1_width(rectangle1_widths[2219]), .rectangle1_height(rectangle1_heights[2219]), .rectangle1_weight(rectangle1_weights[2219]), .rectangle2_x(rectangle2_xs[2219]), .rectangle2_y(rectangle2_ys[2219]), .rectangle2_width(rectangle2_widths[2219]), .rectangle2_height(rectangle2_heights[2219]), .rectangle2_weight(rectangle2_weights[2219]), .rectangle3_x(rectangle3_xs[2219]), .rectangle3_y(rectangle3_ys[2219]), .rectangle3_width(rectangle3_widths[2219]), .rectangle3_height(rectangle3_heights[2219]), .rectangle3_weight(rectangle3_weights[2219]), .feature_threshold(feature_thresholds[2219]), .feature_above(feature_aboves[2219]), .feature_below(feature_belows[2219]), .scan_win_std_dev(scan_win_std_dev[2219]), .feature_accum(feature_accums[2219]));
  accum_calculator ac2220(.scan_win(scan_win2220), .rectangle1_x(rectangle1_xs[2220]), .rectangle1_y(rectangle1_ys[2220]), .rectangle1_width(rectangle1_widths[2220]), .rectangle1_height(rectangle1_heights[2220]), .rectangle1_weight(rectangle1_weights[2220]), .rectangle2_x(rectangle2_xs[2220]), .rectangle2_y(rectangle2_ys[2220]), .rectangle2_width(rectangle2_widths[2220]), .rectangle2_height(rectangle2_heights[2220]), .rectangle2_weight(rectangle2_weights[2220]), .rectangle3_x(rectangle3_xs[2220]), .rectangle3_y(rectangle3_ys[2220]), .rectangle3_width(rectangle3_widths[2220]), .rectangle3_height(rectangle3_heights[2220]), .rectangle3_weight(rectangle3_weights[2220]), .feature_threshold(feature_thresholds[2220]), .feature_above(feature_aboves[2220]), .feature_below(feature_belows[2220]), .scan_win_std_dev(scan_win_std_dev[2220]), .feature_accum(feature_accums[2220]));
  accum_calculator ac2221(.scan_win(scan_win2221), .rectangle1_x(rectangle1_xs[2221]), .rectangle1_y(rectangle1_ys[2221]), .rectangle1_width(rectangle1_widths[2221]), .rectangle1_height(rectangle1_heights[2221]), .rectangle1_weight(rectangle1_weights[2221]), .rectangle2_x(rectangle2_xs[2221]), .rectangle2_y(rectangle2_ys[2221]), .rectangle2_width(rectangle2_widths[2221]), .rectangle2_height(rectangle2_heights[2221]), .rectangle2_weight(rectangle2_weights[2221]), .rectangle3_x(rectangle3_xs[2221]), .rectangle3_y(rectangle3_ys[2221]), .rectangle3_width(rectangle3_widths[2221]), .rectangle3_height(rectangle3_heights[2221]), .rectangle3_weight(rectangle3_weights[2221]), .feature_threshold(feature_thresholds[2221]), .feature_above(feature_aboves[2221]), .feature_below(feature_belows[2221]), .scan_win_std_dev(scan_win_std_dev[2221]), .feature_accum(feature_accums[2221]));
  accum_calculator ac2222(.scan_win(scan_win2222), .rectangle1_x(rectangle1_xs[2222]), .rectangle1_y(rectangle1_ys[2222]), .rectangle1_width(rectangle1_widths[2222]), .rectangle1_height(rectangle1_heights[2222]), .rectangle1_weight(rectangle1_weights[2222]), .rectangle2_x(rectangle2_xs[2222]), .rectangle2_y(rectangle2_ys[2222]), .rectangle2_width(rectangle2_widths[2222]), .rectangle2_height(rectangle2_heights[2222]), .rectangle2_weight(rectangle2_weights[2222]), .rectangle3_x(rectangle3_xs[2222]), .rectangle3_y(rectangle3_ys[2222]), .rectangle3_width(rectangle3_widths[2222]), .rectangle3_height(rectangle3_heights[2222]), .rectangle3_weight(rectangle3_weights[2222]), .feature_threshold(feature_thresholds[2222]), .feature_above(feature_aboves[2222]), .feature_below(feature_belows[2222]), .scan_win_std_dev(scan_win_std_dev[2222]), .feature_accum(feature_accums[2222]));
  accum_calculator ac2223(.scan_win(scan_win2223), .rectangle1_x(rectangle1_xs[2223]), .rectangle1_y(rectangle1_ys[2223]), .rectangle1_width(rectangle1_widths[2223]), .rectangle1_height(rectangle1_heights[2223]), .rectangle1_weight(rectangle1_weights[2223]), .rectangle2_x(rectangle2_xs[2223]), .rectangle2_y(rectangle2_ys[2223]), .rectangle2_width(rectangle2_widths[2223]), .rectangle2_height(rectangle2_heights[2223]), .rectangle2_weight(rectangle2_weights[2223]), .rectangle3_x(rectangle3_xs[2223]), .rectangle3_y(rectangle3_ys[2223]), .rectangle3_width(rectangle3_widths[2223]), .rectangle3_height(rectangle3_heights[2223]), .rectangle3_weight(rectangle3_weights[2223]), .feature_threshold(feature_thresholds[2223]), .feature_above(feature_aboves[2223]), .feature_below(feature_belows[2223]), .scan_win_std_dev(scan_win_std_dev[2223]), .feature_accum(feature_accums[2223]));
  accum_calculator ac2224(.scan_win(scan_win2224), .rectangle1_x(rectangle1_xs[2224]), .rectangle1_y(rectangle1_ys[2224]), .rectangle1_width(rectangle1_widths[2224]), .rectangle1_height(rectangle1_heights[2224]), .rectangle1_weight(rectangle1_weights[2224]), .rectangle2_x(rectangle2_xs[2224]), .rectangle2_y(rectangle2_ys[2224]), .rectangle2_width(rectangle2_widths[2224]), .rectangle2_height(rectangle2_heights[2224]), .rectangle2_weight(rectangle2_weights[2224]), .rectangle3_x(rectangle3_xs[2224]), .rectangle3_y(rectangle3_ys[2224]), .rectangle3_width(rectangle3_widths[2224]), .rectangle3_height(rectangle3_heights[2224]), .rectangle3_weight(rectangle3_weights[2224]), .feature_threshold(feature_thresholds[2224]), .feature_above(feature_aboves[2224]), .feature_below(feature_belows[2224]), .scan_win_std_dev(scan_win_std_dev[2224]), .feature_accum(feature_accums[2224]));
  accum_calculator ac2225(.scan_win(scan_win2225), .rectangle1_x(rectangle1_xs[2225]), .rectangle1_y(rectangle1_ys[2225]), .rectangle1_width(rectangle1_widths[2225]), .rectangle1_height(rectangle1_heights[2225]), .rectangle1_weight(rectangle1_weights[2225]), .rectangle2_x(rectangle2_xs[2225]), .rectangle2_y(rectangle2_ys[2225]), .rectangle2_width(rectangle2_widths[2225]), .rectangle2_height(rectangle2_heights[2225]), .rectangle2_weight(rectangle2_weights[2225]), .rectangle3_x(rectangle3_xs[2225]), .rectangle3_y(rectangle3_ys[2225]), .rectangle3_width(rectangle3_widths[2225]), .rectangle3_height(rectangle3_heights[2225]), .rectangle3_weight(rectangle3_weights[2225]), .feature_threshold(feature_thresholds[2225]), .feature_above(feature_aboves[2225]), .feature_below(feature_belows[2225]), .scan_win_std_dev(scan_win_std_dev[2225]), .feature_accum(feature_accums[2225]));
  accum_calculator ac2226(.scan_win(scan_win2226), .rectangle1_x(rectangle1_xs[2226]), .rectangle1_y(rectangle1_ys[2226]), .rectangle1_width(rectangle1_widths[2226]), .rectangle1_height(rectangle1_heights[2226]), .rectangle1_weight(rectangle1_weights[2226]), .rectangle2_x(rectangle2_xs[2226]), .rectangle2_y(rectangle2_ys[2226]), .rectangle2_width(rectangle2_widths[2226]), .rectangle2_height(rectangle2_heights[2226]), .rectangle2_weight(rectangle2_weights[2226]), .rectangle3_x(rectangle3_xs[2226]), .rectangle3_y(rectangle3_ys[2226]), .rectangle3_width(rectangle3_widths[2226]), .rectangle3_height(rectangle3_heights[2226]), .rectangle3_weight(rectangle3_weights[2226]), .feature_threshold(feature_thresholds[2226]), .feature_above(feature_aboves[2226]), .feature_below(feature_belows[2226]), .scan_win_std_dev(scan_win_std_dev[2226]), .feature_accum(feature_accums[2226]));
  accum_calculator ac2227(.scan_win(scan_win2227), .rectangle1_x(rectangle1_xs[2227]), .rectangle1_y(rectangle1_ys[2227]), .rectangle1_width(rectangle1_widths[2227]), .rectangle1_height(rectangle1_heights[2227]), .rectangle1_weight(rectangle1_weights[2227]), .rectangle2_x(rectangle2_xs[2227]), .rectangle2_y(rectangle2_ys[2227]), .rectangle2_width(rectangle2_widths[2227]), .rectangle2_height(rectangle2_heights[2227]), .rectangle2_weight(rectangle2_weights[2227]), .rectangle3_x(rectangle3_xs[2227]), .rectangle3_y(rectangle3_ys[2227]), .rectangle3_width(rectangle3_widths[2227]), .rectangle3_height(rectangle3_heights[2227]), .rectangle3_weight(rectangle3_weights[2227]), .feature_threshold(feature_thresholds[2227]), .feature_above(feature_aboves[2227]), .feature_below(feature_belows[2227]), .scan_win_std_dev(scan_win_std_dev[2227]), .feature_accum(feature_accums[2227]));
  accum_calculator ac2228(.scan_win(scan_win2228), .rectangle1_x(rectangle1_xs[2228]), .rectangle1_y(rectangle1_ys[2228]), .rectangle1_width(rectangle1_widths[2228]), .rectangle1_height(rectangle1_heights[2228]), .rectangle1_weight(rectangle1_weights[2228]), .rectangle2_x(rectangle2_xs[2228]), .rectangle2_y(rectangle2_ys[2228]), .rectangle2_width(rectangle2_widths[2228]), .rectangle2_height(rectangle2_heights[2228]), .rectangle2_weight(rectangle2_weights[2228]), .rectangle3_x(rectangle3_xs[2228]), .rectangle3_y(rectangle3_ys[2228]), .rectangle3_width(rectangle3_widths[2228]), .rectangle3_height(rectangle3_heights[2228]), .rectangle3_weight(rectangle3_weights[2228]), .feature_threshold(feature_thresholds[2228]), .feature_above(feature_aboves[2228]), .feature_below(feature_belows[2228]), .scan_win_std_dev(scan_win_std_dev[2228]), .feature_accum(feature_accums[2228]));
  accum_calculator ac2229(.scan_win(scan_win2229), .rectangle1_x(rectangle1_xs[2229]), .rectangle1_y(rectangle1_ys[2229]), .rectangle1_width(rectangle1_widths[2229]), .rectangle1_height(rectangle1_heights[2229]), .rectangle1_weight(rectangle1_weights[2229]), .rectangle2_x(rectangle2_xs[2229]), .rectangle2_y(rectangle2_ys[2229]), .rectangle2_width(rectangle2_widths[2229]), .rectangle2_height(rectangle2_heights[2229]), .rectangle2_weight(rectangle2_weights[2229]), .rectangle3_x(rectangle3_xs[2229]), .rectangle3_y(rectangle3_ys[2229]), .rectangle3_width(rectangle3_widths[2229]), .rectangle3_height(rectangle3_heights[2229]), .rectangle3_weight(rectangle3_weights[2229]), .feature_threshold(feature_thresholds[2229]), .feature_above(feature_aboves[2229]), .feature_below(feature_belows[2229]), .scan_win_std_dev(scan_win_std_dev[2229]), .feature_accum(feature_accums[2229]));
  accum_calculator ac2230(.scan_win(scan_win2230), .rectangle1_x(rectangle1_xs[2230]), .rectangle1_y(rectangle1_ys[2230]), .rectangle1_width(rectangle1_widths[2230]), .rectangle1_height(rectangle1_heights[2230]), .rectangle1_weight(rectangle1_weights[2230]), .rectangle2_x(rectangle2_xs[2230]), .rectangle2_y(rectangle2_ys[2230]), .rectangle2_width(rectangle2_widths[2230]), .rectangle2_height(rectangle2_heights[2230]), .rectangle2_weight(rectangle2_weights[2230]), .rectangle3_x(rectangle3_xs[2230]), .rectangle3_y(rectangle3_ys[2230]), .rectangle3_width(rectangle3_widths[2230]), .rectangle3_height(rectangle3_heights[2230]), .rectangle3_weight(rectangle3_weights[2230]), .feature_threshold(feature_thresholds[2230]), .feature_above(feature_aboves[2230]), .feature_below(feature_belows[2230]), .scan_win_std_dev(scan_win_std_dev[2230]), .feature_accum(feature_accums[2230]));
  accum_calculator ac2231(.scan_win(scan_win2231), .rectangle1_x(rectangle1_xs[2231]), .rectangle1_y(rectangle1_ys[2231]), .rectangle1_width(rectangle1_widths[2231]), .rectangle1_height(rectangle1_heights[2231]), .rectangle1_weight(rectangle1_weights[2231]), .rectangle2_x(rectangle2_xs[2231]), .rectangle2_y(rectangle2_ys[2231]), .rectangle2_width(rectangle2_widths[2231]), .rectangle2_height(rectangle2_heights[2231]), .rectangle2_weight(rectangle2_weights[2231]), .rectangle3_x(rectangle3_xs[2231]), .rectangle3_y(rectangle3_ys[2231]), .rectangle3_width(rectangle3_widths[2231]), .rectangle3_height(rectangle3_heights[2231]), .rectangle3_weight(rectangle3_weights[2231]), .feature_threshold(feature_thresholds[2231]), .feature_above(feature_aboves[2231]), .feature_below(feature_belows[2231]), .scan_win_std_dev(scan_win_std_dev[2231]), .feature_accum(feature_accums[2231]));
  accum_calculator ac2232(.scan_win(scan_win2232), .rectangle1_x(rectangle1_xs[2232]), .rectangle1_y(rectangle1_ys[2232]), .rectangle1_width(rectangle1_widths[2232]), .rectangle1_height(rectangle1_heights[2232]), .rectangle1_weight(rectangle1_weights[2232]), .rectangle2_x(rectangle2_xs[2232]), .rectangle2_y(rectangle2_ys[2232]), .rectangle2_width(rectangle2_widths[2232]), .rectangle2_height(rectangle2_heights[2232]), .rectangle2_weight(rectangle2_weights[2232]), .rectangle3_x(rectangle3_xs[2232]), .rectangle3_y(rectangle3_ys[2232]), .rectangle3_width(rectangle3_widths[2232]), .rectangle3_height(rectangle3_heights[2232]), .rectangle3_weight(rectangle3_weights[2232]), .feature_threshold(feature_thresholds[2232]), .feature_above(feature_aboves[2232]), .feature_below(feature_belows[2232]), .scan_win_std_dev(scan_win_std_dev[2232]), .feature_accum(feature_accums[2232]));
  accum_calculator ac2233(.scan_win(scan_win2233), .rectangle1_x(rectangle1_xs[2233]), .rectangle1_y(rectangle1_ys[2233]), .rectangle1_width(rectangle1_widths[2233]), .rectangle1_height(rectangle1_heights[2233]), .rectangle1_weight(rectangle1_weights[2233]), .rectangle2_x(rectangle2_xs[2233]), .rectangle2_y(rectangle2_ys[2233]), .rectangle2_width(rectangle2_widths[2233]), .rectangle2_height(rectangle2_heights[2233]), .rectangle2_weight(rectangle2_weights[2233]), .rectangle3_x(rectangle3_xs[2233]), .rectangle3_y(rectangle3_ys[2233]), .rectangle3_width(rectangle3_widths[2233]), .rectangle3_height(rectangle3_heights[2233]), .rectangle3_weight(rectangle3_weights[2233]), .feature_threshold(feature_thresholds[2233]), .feature_above(feature_aboves[2233]), .feature_below(feature_belows[2233]), .scan_win_std_dev(scan_win_std_dev[2233]), .feature_accum(feature_accums[2233]));
  accum_calculator ac2234(.scan_win(scan_win2234), .rectangle1_x(rectangle1_xs[2234]), .rectangle1_y(rectangle1_ys[2234]), .rectangle1_width(rectangle1_widths[2234]), .rectangle1_height(rectangle1_heights[2234]), .rectangle1_weight(rectangle1_weights[2234]), .rectangle2_x(rectangle2_xs[2234]), .rectangle2_y(rectangle2_ys[2234]), .rectangle2_width(rectangle2_widths[2234]), .rectangle2_height(rectangle2_heights[2234]), .rectangle2_weight(rectangle2_weights[2234]), .rectangle3_x(rectangle3_xs[2234]), .rectangle3_y(rectangle3_ys[2234]), .rectangle3_width(rectangle3_widths[2234]), .rectangle3_height(rectangle3_heights[2234]), .rectangle3_weight(rectangle3_weights[2234]), .feature_threshold(feature_thresholds[2234]), .feature_above(feature_aboves[2234]), .feature_below(feature_belows[2234]), .scan_win_std_dev(scan_win_std_dev[2234]), .feature_accum(feature_accums[2234]));
  accum_calculator ac2235(.scan_win(scan_win2235), .rectangle1_x(rectangle1_xs[2235]), .rectangle1_y(rectangle1_ys[2235]), .rectangle1_width(rectangle1_widths[2235]), .rectangle1_height(rectangle1_heights[2235]), .rectangle1_weight(rectangle1_weights[2235]), .rectangle2_x(rectangle2_xs[2235]), .rectangle2_y(rectangle2_ys[2235]), .rectangle2_width(rectangle2_widths[2235]), .rectangle2_height(rectangle2_heights[2235]), .rectangle2_weight(rectangle2_weights[2235]), .rectangle3_x(rectangle3_xs[2235]), .rectangle3_y(rectangle3_ys[2235]), .rectangle3_width(rectangle3_widths[2235]), .rectangle3_height(rectangle3_heights[2235]), .rectangle3_weight(rectangle3_weights[2235]), .feature_threshold(feature_thresholds[2235]), .feature_above(feature_aboves[2235]), .feature_below(feature_belows[2235]), .scan_win_std_dev(scan_win_std_dev[2235]), .feature_accum(feature_accums[2235]));
  accum_calculator ac2236(.scan_win(scan_win2236), .rectangle1_x(rectangle1_xs[2236]), .rectangle1_y(rectangle1_ys[2236]), .rectangle1_width(rectangle1_widths[2236]), .rectangle1_height(rectangle1_heights[2236]), .rectangle1_weight(rectangle1_weights[2236]), .rectangle2_x(rectangle2_xs[2236]), .rectangle2_y(rectangle2_ys[2236]), .rectangle2_width(rectangle2_widths[2236]), .rectangle2_height(rectangle2_heights[2236]), .rectangle2_weight(rectangle2_weights[2236]), .rectangle3_x(rectangle3_xs[2236]), .rectangle3_y(rectangle3_ys[2236]), .rectangle3_width(rectangle3_widths[2236]), .rectangle3_height(rectangle3_heights[2236]), .rectangle3_weight(rectangle3_weights[2236]), .feature_threshold(feature_thresholds[2236]), .feature_above(feature_aboves[2236]), .feature_below(feature_belows[2236]), .scan_win_std_dev(scan_win_std_dev[2236]), .feature_accum(feature_accums[2236]));
  accum_calculator ac2237(.scan_win(scan_win2237), .rectangle1_x(rectangle1_xs[2237]), .rectangle1_y(rectangle1_ys[2237]), .rectangle1_width(rectangle1_widths[2237]), .rectangle1_height(rectangle1_heights[2237]), .rectangle1_weight(rectangle1_weights[2237]), .rectangle2_x(rectangle2_xs[2237]), .rectangle2_y(rectangle2_ys[2237]), .rectangle2_width(rectangle2_widths[2237]), .rectangle2_height(rectangle2_heights[2237]), .rectangle2_weight(rectangle2_weights[2237]), .rectangle3_x(rectangle3_xs[2237]), .rectangle3_y(rectangle3_ys[2237]), .rectangle3_width(rectangle3_widths[2237]), .rectangle3_height(rectangle3_heights[2237]), .rectangle3_weight(rectangle3_weights[2237]), .feature_threshold(feature_thresholds[2237]), .feature_above(feature_aboves[2237]), .feature_below(feature_belows[2237]), .scan_win_std_dev(scan_win_std_dev[2237]), .feature_accum(feature_accums[2237]));
  accum_calculator ac2238(.scan_win(scan_win2238), .rectangle1_x(rectangle1_xs[2238]), .rectangle1_y(rectangle1_ys[2238]), .rectangle1_width(rectangle1_widths[2238]), .rectangle1_height(rectangle1_heights[2238]), .rectangle1_weight(rectangle1_weights[2238]), .rectangle2_x(rectangle2_xs[2238]), .rectangle2_y(rectangle2_ys[2238]), .rectangle2_width(rectangle2_widths[2238]), .rectangle2_height(rectangle2_heights[2238]), .rectangle2_weight(rectangle2_weights[2238]), .rectangle3_x(rectangle3_xs[2238]), .rectangle3_y(rectangle3_ys[2238]), .rectangle3_width(rectangle3_widths[2238]), .rectangle3_height(rectangle3_heights[2238]), .rectangle3_weight(rectangle3_weights[2238]), .feature_threshold(feature_thresholds[2238]), .feature_above(feature_aboves[2238]), .feature_below(feature_belows[2238]), .scan_win_std_dev(scan_win_std_dev[2238]), .feature_accum(feature_accums[2238]));
  accum_calculator ac2239(.scan_win(scan_win2239), .rectangle1_x(rectangle1_xs[2239]), .rectangle1_y(rectangle1_ys[2239]), .rectangle1_width(rectangle1_widths[2239]), .rectangle1_height(rectangle1_heights[2239]), .rectangle1_weight(rectangle1_weights[2239]), .rectangle2_x(rectangle2_xs[2239]), .rectangle2_y(rectangle2_ys[2239]), .rectangle2_width(rectangle2_widths[2239]), .rectangle2_height(rectangle2_heights[2239]), .rectangle2_weight(rectangle2_weights[2239]), .rectangle3_x(rectangle3_xs[2239]), .rectangle3_y(rectangle3_ys[2239]), .rectangle3_width(rectangle3_widths[2239]), .rectangle3_height(rectangle3_heights[2239]), .rectangle3_weight(rectangle3_weights[2239]), .feature_threshold(feature_thresholds[2239]), .feature_above(feature_aboves[2239]), .feature_below(feature_belows[2239]), .scan_win_std_dev(scan_win_std_dev[2239]), .feature_accum(feature_accums[2239]));
  accum_calculator ac2240(.scan_win(scan_win2240), .rectangle1_x(rectangle1_xs[2240]), .rectangle1_y(rectangle1_ys[2240]), .rectangle1_width(rectangle1_widths[2240]), .rectangle1_height(rectangle1_heights[2240]), .rectangle1_weight(rectangle1_weights[2240]), .rectangle2_x(rectangle2_xs[2240]), .rectangle2_y(rectangle2_ys[2240]), .rectangle2_width(rectangle2_widths[2240]), .rectangle2_height(rectangle2_heights[2240]), .rectangle2_weight(rectangle2_weights[2240]), .rectangle3_x(rectangle3_xs[2240]), .rectangle3_y(rectangle3_ys[2240]), .rectangle3_width(rectangle3_widths[2240]), .rectangle3_height(rectangle3_heights[2240]), .rectangle3_weight(rectangle3_weights[2240]), .feature_threshold(feature_thresholds[2240]), .feature_above(feature_aboves[2240]), .feature_below(feature_belows[2240]), .scan_win_std_dev(scan_win_std_dev[2240]), .feature_accum(feature_accums[2240]));
  accum_calculator ac2241(.scan_win(scan_win2241), .rectangle1_x(rectangle1_xs[2241]), .rectangle1_y(rectangle1_ys[2241]), .rectangle1_width(rectangle1_widths[2241]), .rectangle1_height(rectangle1_heights[2241]), .rectangle1_weight(rectangle1_weights[2241]), .rectangle2_x(rectangle2_xs[2241]), .rectangle2_y(rectangle2_ys[2241]), .rectangle2_width(rectangle2_widths[2241]), .rectangle2_height(rectangle2_heights[2241]), .rectangle2_weight(rectangle2_weights[2241]), .rectangle3_x(rectangle3_xs[2241]), .rectangle3_y(rectangle3_ys[2241]), .rectangle3_width(rectangle3_widths[2241]), .rectangle3_height(rectangle3_heights[2241]), .rectangle3_weight(rectangle3_weights[2241]), .feature_threshold(feature_thresholds[2241]), .feature_above(feature_aboves[2241]), .feature_below(feature_belows[2241]), .scan_win_std_dev(scan_win_std_dev[2241]), .feature_accum(feature_accums[2241]));
  accum_calculator ac2242(.scan_win(scan_win2242), .rectangle1_x(rectangle1_xs[2242]), .rectangle1_y(rectangle1_ys[2242]), .rectangle1_width(rectangle1_widths[2242]), .rectangle1_height(rectangle1_heights[2242]), .rectangle1_weight(rectangle1_weights[2242]), .rectangle2_x(rectangle2_xs[2242]), .rectangle2_y(rectangle2_ys[2242]), .rectangle2_width(rectangle2_widths[2242]), .rectangle2_height(rectangle2_heights[2242]), .rectangle2_weight(rectangle2_weights[2242]), .rectangle3_x(rectangle3_xs[2242]), .rectangle3_y(rectangle3_ys[2242]), .rectangle3_width(rectangle3_widths[2242]), .rectangle3_height(rectangle3_heights[2242]), .rectangle3_weight(rectangle3_weights[2242]), .feature_threshold(feature_thresholds[2242]), .feature_above(feature_aboves[2242]), .feature_below(feature_belows[2242]), .scan_win_std_dev(scan_win_std_dev[2242]), .feature_accum(feature_accums[2242]));
  accum_calculator ac2243(.scan_win(scan_win2243), .rectangle1_x(rectangle1_xs[2243]), .rectangle1_y(rectangle1_ys[2243]), .rectangle1_width(rectangle1_widths[2243]), .rectangle1_height(rectangle1_heights[2243]), .rectangle1_weight(rectangle1_weights[2243]), .rectangle2_x(rectangle2_xs[2243]), .rectangle2_y(rectangle2_ys[2243]), .rectangle2_width(rectangle2_widths[2243]), .rectangle2_height(rectangle2_heights[2243]), .rectangle2_weight(rectangle2_weights[2243]), .rectangle3_x(rectangle3_xs[2243]), .rectangle3_y(rectangle3_ys[2243]), .rectangle3_width(rectangle3_widths[2243]), .rectangle3_height(rectangle3_heights[2243]), .rectangle3_weight(rectangle3_weights[2243]), .feature_threshold(feature_thresholds[2243]), .feature_above(feature_aboves[2243]), .feature_below(feature_belows[2243]), .scan_win_std_dev(scan_win_std_dev[2243]), .feature_accum(feature_accums[2243]));
  accum_calculator ac2244(.scan_win(scan_win2244), .rectangle1_x(rectangle1_xs[2244]), .rectangle1_y(rectangle1_ys[2244]), .rectangle1_width(rectangle1_widths[2244]), .rectangle1_height(rectangle1_heights[2244]), .rectangle1_weight(rectangle1_weights[2244]), .rectangle2_x(rectangle2_xs[2244]), .rectangle2_y(rectangle2_ys[2244]), .rectangle2_width(rectangle2_widths[2244]), .rectangle2_height(rectangle2_heights[2244]), .rectangle2_weight(rectangle2_weights[2244]), .rectangle3_x(rectangle3_xs[2244]), .rectangle3_y(rectangle3_ys[2244]), .rectangle3_width(rectangle3_widths[2244]), .rectangle3_height(rectangle3_heights[2244]), .rectangle3_weight(rectangle3_weights[2244]), .feature_threshold(feature_thresholds[2244]), .feature_above(feature_aboves[2244]), .feature_below(feature_belows[2244]), .scan_win_std_dev(scan_win_std_dev[2244]), .feature_accum(feature_accums[2244]));
  accum_calculator ac2245(.scan_win(scan_win2245), .rectangle1_x(rectangle1_xs[2245]), .rectangle1_y(rectangle1_ys[2245]), .rectangle1_width(rectangle1_widths[2245]), .rectangle1_height(rectangle1_heights[2245]), .rectangle1_weight(rectangle1_weights[2245]), .rectangle2_x(rectangle2_xs[2245]), .rectangle2_y(rectangle2_ys[2245]), .rectangle2_width(rectangle2_widths[2245]), .rectangle2_height(rectangle2_heights[2245]), .rectangle2_weight(rectangle2_weights[2245]), .rectangle3_x(rectangle3_xs[2245]), .rectangle3_y(rectangle3_ys[2245]), .rectangle3_width(rectangle3_widths[2245]), .rectangle3_height(rectangle3_heights[2245]), .rectangle3_weight(rectangle3_weights[2245]), .feature_threshold(feature_thresholds[2245]), .feature_above(feature_aboves[2245]), .feature_below(feature_belows[2245]), .scan_win_std_dev(scan_win_std_dev[2245]), .feature_accum(feature_accums[2245]));
  accum_calculator ac2246(.scan_win(scan_win2246), .rectangle1_x(rectangle1_xs[2246]), .rectangle1_y(rectangle1_ys[2246]), .rectangle1_width(rectangle1_widths[2246]), .rectangle1_height(rectangle1_heights[2246]), .rectangle1_weight(rectangle1_weights[2246]), .rectangle2_x(rectangle2_xs[2246]), .rectangle2_y(rectangle2_ys[2246]), .rectangle2_width(rectangle2_widths[2246]), .rectangle2_height(rectangle2_heights[2246]), .rectangle2_weight(rectangle2_weights[2246]), .rectangle3_x(rectangle3_xs[2246]), .rectangle3_y(rectangle3_ys[2246]), .rectangle3_width(rectangle3_widths[2246]), .rectangle3_height(rectangle3_heights[2246]), .rectangle3_weight(rectangle3_weights[2246]), .feature_threshold(feature_thresholds[2246]), .feature_above(feature_aboves[2246]), .feature_below(feature_belows[2246]), .scan_win_std_dev(scan_win_std_dev[2246]), .feature_accum(feature_accums[2246]));
  accum_calculator ac2247(.scan_win(scan_win2247), .rectangle1_x(rectangle1_xs[2247]), .rectangle1_y(rectangle1_ys[2247]), .rectangle1_width(rectangle1_widths[2247]), .rectangle1_height(rectangle1_heights[2247]), .rectangle1_weight(rectangle1_weights[2247]), .rectangle2_x(rectangle2_xs[2247]), .rectangle2_y(rectangle2_ys[2247]), .rectangle2_width(rectangle2_widths[2247]), .rectangle2_height(rectangle2_heights[2247]), .rectangle2_weight(rectangle2_weights[2247]), .rectangle3_x(rectangle3_xs[2247]), .rectangle3_y(rectangle3_ys[2247]), .rectangle3_width(rectangle3_widths[2247]), .rectangle3_height(rectangle3_heights[2247]), .rectangle3_weight(rectangle3_weights[2247]), .feature_threshold(feature_thresholds[2247]), .feature_above(feature_aboves[2247]), .feature_below(feature_belows[2247]), .scan_win_std_dev(scan_win_std_dev[2247]), .feature_accum(feature_accums[2247]));
  accum_calculator ac2248(.scan_win(scan_win2248), .rectangle1_x(rectangle1_xs[2248]), .rectangle1_y(rectangle1_ys[2248]), .rectangle1_width(rectangle1_widths[2248]), .rectangle1_height(rectangle1_heights[2248]), .rectangle1_weight(rectangle1_weights[2248]), .rectangle2_x(rectangle2_xs[2248]), .rectangle2_y(rectangle2_ys[2248]), .rectangle2_width(rectangle2_widths[2248]), .rectangle2_height(rectangle2_heights[2248]), .rectangle2_weight(rectangle2_weights[2248]), .rectangle3_x(rectangle3_xs[2248]), .rectangle3_y(rectangle3_ys[2248]), .rectangle3_width(rectangle3_widths[2248]), .rectangle3_height(rectangle3_heights[2248]), .rectangle3_weight(rectangle3_weights[2248]), .feature_threshold(feature_thresholds[2248]), .feature_above(feature_aboves[2248]), .feature_below(feature_belows[2248]), .scan_win_std_dev(scan_win_std_dev[2248]), .feature_accum(feature_accums[2248]));
  accum_calculator ac2249(.scan_win(scan_win2249), .rectangle1_x(rectangle1_xs[2249]), .rectangle1_y(rectangle1_ys[2249]), .rectangle1_width(rectangle1_widths[2249]), .rectangle1_height(rectangle1_heights[2249]), .rectangle1_weight(rectangle1_weights[2249]), .rectangle2_x(rectangle2_xs[2249]), .rectangle2_y(rectangle2_ys[2249]), .rectangle2_width(rectangle2_widths[2249]), .rectangle2_height(rectangle2_heights[2249]), .rectangle2_weight(rectangle2_weights[2249]), .rectangle3_x(rectangle3_xs[2249]), .rectangle3_y(rectangle3_ys[2249]), .rectangle3_width(rectangle3_widths[2249]), .rectangle3_height(rectangle3_heights[2249]), .rectangle3_weight(rectangle3_weights[2249]), .feature_threshold(feature_thresholds[2249]), .feature_above(feature_aboves[2249]), .feature_below(feature_belows[2249]), .scan_win_std_dev(scan_win_std_dev[2249]), .feature_accum(feature_accums[2249]));
  accum_calculator ac2250(.scan_win(scan_win2250), .rectangle1_x(rectangle1_xs[2250]), .rectangle1_y(rectangle1_ys[2250]), .rectangle1_width(rectangle1_widths[2250]), .rectangle1_height(rectangle1_heights[2250]), .rectangle1_weight(rectangle1_weights[2250]), .rectangle2_x(rectangle2_xs[2250]), .rectangle2_y(rectangle2_ys[2250]), .rectangle2_width(rectangle2_widths[2250]), .rectangle2_height(rectangle2_heights[2250]), .rectangle2_weight(rectangle2_weights[2250]), .rectangle3_x(rectangle3_xs[2250]), .rectangle3_y(rectangle3_ys[2250]), .rectangle3_width(rectangle3_widths[2250]), .rectangle3_height(rectangle3_heights[2250]), .rectangle3_weight(rectangle3_weights[2250]), .feature_threshold(feature_thresholds[2250]), .feature_above(feature_aboves[2250]), .feature_below(feature_belows[2250]), .scan_win_std_dev(scan_win_std_dev[2250]), .feature_accum(feature_accums[2250]));
  accum_calculator ac2251(.scan_win(scan_win2251), .rectangle1_x(rectangle1_xs[2251]), .rectangle1_y(rectangle1_ys[2251]), .rectangle1_width(rectangle1_widths[2251]), .rectangle1_height(rectangle1_heights[2251]), .rectangle1_weight(rectangle1_weights[2251]), .rectangle2_x(rectangle2_xs[2251]), .rectangle2_y(rectangle2_ys[2251]), .rectangle2_width(rectangle2_widths[2251]), .rectangle2_height(rectangle2_heights[2251]), .rectangle2_weight(rectangle2_weights[2251]), .rectangle3_x(rectangle3_xs[2251]), .rectangle3_y(rectangle3_ys[2251]), .rectangle3_width(rectangle3_widths[2251]), .rectangle3_height(rectangle3_heights[2251]), .rectangle3_weight(rectangle3_weights[2251]), .feature_threshold(feature_thresholds[2251]), .feature_above(feature_aboves[2251]), .feature_below(feature_belows[2251]), .scan_win_std_dev(scan_win_std_dev[2251]), .feature_accum(feature_accums[2251]));
  accum_calculator ac2252(.scan_win(scan_win2252), .rectangle1_x(rectangle1_xs[2252]), .rectangle1_y(rectangle1_ys[2252]), .rectangle1_width(rectangle1_widths[2252]), .rectangle1_height(rectangle1_heights[2252]), .rectangle1_weight(rectangle1_weights[2252]), .rectangle2_x(rectangle2_xs[2252]), .rectangle2_y(rectangle2_ys[2252]), .rectangle2_width(rectangle2_widths[2252]), .rectangle2_height(rectangle2_heights[2252]), .rectangle2_weight(rectangle2_weights[2252]), .rectangle3_x(rectangle3_xs[2252]), .rectangle3_y(rectangle3_ys[2252]), .rectangle3_width(rectangle3_widths[2252]), .rectangle3_height(rectangle3_heights[2252]), .rectangle3_weight(rectangle3_weights[2252]), .feature_threshold(feature_thresholds[2252]), .feature_above(feature_aboves[2252]), .feature_below(feature_belows[2252]), .scan_win_std_dev(scan_win_std_dev[2252]), .feature_accum(feature_accums[2252]));
  accum_calculator ac2253(.scan_win(scan_win2253), .rectangle1_x(rectangle1_xs[2253]), .rectangle1_y(rectangle1_ys[2253]), .rectangle1_width(rectangle1_widths[2253]), .rectangle1_height(rectangle1_heights[2253]), .rectangle1_weight(rectangle1_weights[2253]), .rectangle2_x(rectangle2_xs[2253]), .rectangle2_y(rectangle2_ys[2253]), .rectangle2_width(rectangle2_widths[2253]), .rectangle2_height(rectangle2_heights[2253]), .rectangle2_weight(rectangle2_weights[2253]), .rectangle3_x(rectangle3_xs[2253]), .rectangle3_y(rectangle3_ys[2253]), .rectangle3_width(rectangle3_widths[2253]), .rectangle3_height(rectangle3_heights[2253]), .rectangle3_weight(rectangle3_weights[2253]), .feature_threshold(feature_thresholds[2253]), .feature_above(feature_aboves[2253]), .feature_below(feature_belows[2253]), .scan_win_std_dev(scan_win_std_dev[2253]), .feature_accum(feature_accums[2253]));
  accum_calculator ac2254(.scan_win(scan_win2254), .rectangle1_x(rectangle1_xs[2254]), .rectangle1_y(rectangle1_ys[2254]), .rectangle1_width(rectangle1_widths[2254]), .rectangle1_height(rectangle1_heights[2254]), .rectangle1_weight(rectangle1_weights[2254]), .rectangle2_x(rectangle2_xs[2254]), .rectangle2_y(rectangle2_ys[2254]), .rectangle2_width(rectangle2_widths[2254]), .rectangle2_height(rectangle2_heights[2254]), .rectangle2_weight(rectangle2_weights[2254]), .rectangle3_x(rectangle3_xs[2254]), .rectangle3_y(rectangle3_ys[2254]), .rectangle3_width(rectangle3_widths[2254]), .rectangle3_height(rectangle3_heights[2254]), .rectangle3_weight(rectangle3_weights[2254]), .feature_threshold(feature_thresholds[2254]), .feature_above(feature_aboves[2254]), .feature_below(feature_belows[2254]), .scan_win_std_dev(scan_win_std_dev[2254]), .feature_accum(feature_accums[2254]));
  accum_calculator ac2255(.scan_win(scan_win2255), .rectangle1_x(rectangle1_xs[2255]), .rectangle1_y(rectangle1_ys[2255]), .rectangle1_width(rectangle1_widths[2255]), .rectangle1_height(rectangle1_heights[2255]), .rectangle1_weight(rectangle1_weights[2255]), .rectangle2_x(rectangle2_xs[2255]), .rectangle2_y(rectangle2_ys[2255]), .rectangle2_width(rectangle2_widths[2255]), .rectangle2_height(rectangle2_heights[2255]), .rectangle2_weight(rectangle2_weights[2255]), .rectangle3_x(rectangle3_xs[2255]), .rectangle3_y(rectangle3_ys[2255]), .rectangle3_width(rectangle3_widths[2255]), .rectangle3_height(rectangle3_heights[2255]), .rectangle3_weight(rectangle3_weights[2255]), .feature_threshold(feature_thresholds[2255]), .feature_above(feature_aboves[2255]), .feature_below(feature_belows[2255]), .scan_win_std_dev(scan_win_std_dev[2255]), .feature_accum(feature_accums[2255]));
  accum_calculator ac2256(.scan_win(scan_win2256), .rectangle1_x(rectangle1_xs[2256]), .rectangle1_y(rectangle1_ys[2256]), .rectangle1_width(rectangle1_widths[2256]), .rectangle1_height(rectangle1_heights[2256]), .rectangle1_weight(rectangle1_weights[2256]), .rectangle2_x(rectangle2_xs[2256]), .rectangle2_y(rectangle2_ys[2256]), .rectangle2_width(rectangle2_widths[2256]), .rectangle2_height(rectangle2_heights[2256]), .rectangle2_weight(rectangle2_weights[2256]), .rectangle3_x(rectangle3_xs[2256]), .rectangle3_y(rectangle3_ys[2256]), .rectangle3_width(rectangle3_widths[2256]), .rectangle3_height(rectangle3_heights[2256]), .rectangle3_weight(rectangle3_weights[2256]), .feature_threshold(feature_thresholds[2256]), .feature_above(feature_aboves[2256]), .feature_below(feature_belows[2256]), .scan_win_std_dev(scan_win_std_dev[2256]), .feature_accum(feature_accums[2256]));
  accum_calculator ac2257(.scan_win(scan_win2257), .rectangle1_x(rectangle1_xs[2257]), .rectangle1_y(rectangle1_ys[2257]), .rectangle1_width(rectangle1_widths[2257]), .rectangle1_height(rectangle1_heights[2257]), .rectangle1_weight(rectangle1_weights[2257]), .rectangle2_x(rectangle2_xs[2257]), .rectangle2_y(rectangle2_ys[2257]), .rectangle2_width(rectangle2_widths[2257]), .rectangle2_height(rectangle2_heights[2257]), .rectangle2_weight(rectangle2_weights[2257]), .rectangle3_x(rectangle3_xs[2257]), .rectangle3_y(rectangle3_ys[2257]), .rectangle3_width(rectangle3_widths[2257]), .rectangle3_height(rectangle3_heights[2257]), .rectangle3_weight(rectangle3_weights[2257]), .feature_threshold(feature_thresholds[2257]), .feature_above(feature_aboves[2257]), .feature_below(feature_belows[2257]), .scan_win_std_dev(scan_win_std_dev[2257]), .feature_accum(feature_accums[2257]));
  accum_calculator ac2258(.scan_win(scan_win2258), .rectangle1_x(rectangle1_xs[2258]), .rectangle1_y(rectangle1_ys[2258]), .rectangle1_width(rectangle1_widths[2258]), .rectangle1_height(rectangle1_heights[2258]), .rectangle1_weight(rectangle1_weights[2258]), .rectangle2_x(rectangle2_xs[2258]), .rectangle2_y(rectangle2_ys[2258]), .rectangle2_width(rectangle2_widths[2258]), .rectangle2_height(rectangle2_heights[2258]), .rectangle2_weight(rectangle2_weights[2258]), .rectangle3_x(rectangle3_xs[2258]), .rectangle3_y(rectangle3_ys[2258]), .rectangle3_width(rectangle3_widths[2258]), .rectangle3_height(rectangle3_heights[2258]), .rectangle3_weight(rectangle3_weights[2258]), .feature_threshold(feature_thresholds[2258]), .feature_above(feature_aboves[2258]), .feature_below(feature_belows[2258]), .scan_win_std_dev(scan_win_std_dev[2258]), .feature_accum(feature_accums[2258]));
  accum_calculator ac2259(.scan_win(scan_win2259), .rectangle1_x(rectangle1_xs[2259]), .rectangle1_y(rectangle1_ys[2259]), .rectangle1_width(rectangle1_widths[2259]), .rectangle1_height(rectangle1_heights[2259]), .rectangle1_weight(rectangle1_weights[2259]), .rectangle2_x(rectangle2_xs[2259]), .rectangle2_y(rectangle2_ys[2259]), .rectangle2_width(rectangle2_widths[2259]), .rectangle2_height(rectangle2_heights[2259]), .rectangle2_weight(rectangle2_weights[2259]), .rectangle3_x(rectangle3_xs[2259]), .rectangle3_y(rectangle3_ys[2259]), .rectangle3_width(rectangle3_widths[2259]), .rectangle3_height(rectangle3_heights[2259]), .rectangle3_weight(rectangle3_weights[2259]), .feature_threshold(feature_thresholds[2259]), .feature_above(feature_aboves[2259]), .feature_below(feature_belows[2259]), .scan_win_std_dev(scan_win_std_dev[2259]), .feature_accum(feature_accums[2259]));
  accum_calculator ac2260(.scan_win(scan_win2260), .rectangle1_x(rectangle1_xs[2260]), .rectangle1_y(rectangle1_ys[2260]), .rectangle1_width(rectangle1_widths[2260]), .rectangle1_height(rectangle1_heights[2260]), .rectangle1_weight(rectangle1_weights[2260]), .rectangle2_x(rectangle2_xs[2260]), .rectangle2_y(rectangle2_ys[2260]), .rectangle2_width(rectangle2_widths[2260]), .rectangle2_height(rectangle2_heights[2260]), .rectangle2_weight(rectangle2_weights[2260]), .rectangle3_x(rectangle3_xs[2260]), .rectangle3_y(rectangle3_ys[2260]), .rectangle3_width(rectangle3_widths[2260]), .rectangle3_height(rectangle3_heights[2260]), .rectangle3_weight(rectangle3_weights[2260]), .feature_threshold(feature_thresholds[2260]), .feature_above(feature_aboves[2260]), .feature_below(feature_belows[2260]), .scan_win_std_dev(scan_win_std_dev[2260]), .feature_accum(feature_accums[2260]));
  accum_calculator ac2261(.scan_win(scan_win2261), .rectangle1_x(rectangle1_xs[2261]), .rectangle1_y(rectangle1_ys[2261]), .rectangle1_width(rectangle1_widths[2261]), .rectangle1_height(rectangle1_heights[2261]), .rectangle1_weight(rectangle1_weights[2261]), .rectangle2_x(rectangle2_xs[2261]), .rectangle2_y(rectangle2_ys[2261]), .rectangle2_width(rectangle2_widths[2261]), .rectangle2_height(rectangle2_heights[2261]), .rectangle2_weight(rectangle2_weights[2261]), .rectangle3_x(rectangle3_xs[2261]), .rectangle3_y(rectangle3_ys[2261]), .rectangle3_width(rectangle3_widths[2261]), .rectangle3_height(rectangle3_heights[2261]), .rectangle3_weight(rectangle3_weights[2261]), .feature_threshold(feature_thresholds[2261]), .feature_above(feature_aboves[2261]), .feature_below(feature_belows[2261]), .scan_win_std_dev(scan_win_std_dev[2261]), .feature_accum(feature_accums[2261]));
  accum_calculator ac2262(.scan_win(scan_win2262), .rectangle1_x(rectangle1_xs[2262]), .rectangle1_y(rectangle1_ys[2262]), .rectangle1_width(rectangle1_widths[2262]), .rectangle1_height(rectangle1_heights[2262]), .rectangle1_weight(rectangle1_weights[2262]), .rectangle2_x(rectangle2_xs[2262]), .rectangle2_y(rectangle2_ys[2262]), .rectangle2_width(rectangle2_widths[2262]), .rectangle2_height(rectangle2_heights[2262]), .rectangle2_weight(rectangle2_weights[2262]), .rectangle3_x(rectangle3_xs[2262]), .rectangle3_y(rectangle3_ys[2262]), .rectangle3_width(rectangle3_widths[2262]), .rectangle3_height(rectangle3_heights[2262]), .rectangle3_weight(rectangle3_weights[2262]), .feature_threshold(feature_thresholds[2262]), .feature_above(feature_aboves[2262]), .feature_below(feature_belows[2262]), .scan_win_std_dev(scan_win_std_dev[2262]), .feature_accum(feature_accums[2262]));
  accum_calculator ac2263(.scan_win(scan_win2263), .rectangle1_x(rectangle1_xs[2263]), .rectangle1_y(rectangle1_ys[2263]), .rectangle1_width(rectangle1_widths[2263]), .rectangle1_height(rectangle1_heights[2263]), .rectangle1_weight(rectangle1_weights[2263]), .rectangle2_x(rectangle2_xs[2263]), .rectangle2_y(rectangle2_ys[2263]), .rectangle2_width(rectangle2_widths[2263]), .rectangle2_height(rectangle2_heights[2263]), .rectangle2_weight(rectangle2_weights[2263]), .rectangle3_x(rectangle3_xs[2263]), .rectangle3_y(rectangle3_ys[2263]), .rectangle3_width(rectangle3_widths[2263]), .rectangle3_height(rectangle3_heights[2263]), .rectangle3_weight(rectangle3_weights[2263]), .feature_threshold(feature_thresholds[2263]), .feature_above(feature_aboves[2263]), .feature_below(feature_belows[2263]), .scan_win_std_dev(scan_win_std_dev[2263]), .feature_accum(feature_accums[2263]));
  accum_calculator ac2264(.scan_win(scan_win2264), .rectangle1_x(rectangle1_xs[2264]), .rectangle1_y(rectangle1_ys[2264]), .rectangle1_width(rectangle1_widths[2264]), .rectangle1_height(rectangle1_heights[2264]), .rectangle1_weight(rectangle1_weights[2264]), .rectangle2_x(rectangle2_xs[2264]), .rectangle2_y(rectangle2_ys[2264]), .rectangle2_width(rectangle2_widths[2264]), .rectangle2_height(rectangle2_heights[2264]), .rectangle2_weight(rectangle2_weights[2264]), .rectangle3_x(rectangle3_xs[2264]), .rectangle3_y(rectangle3_ys[2264]), .rectangle3_width(rectangle3_widths[2264]), .rectangle3_height(rectangle3_heights[2264]), .rectangle3_weight(rectangle3_weights[2264]), .feature_threshold(feature_thresholds[2264]), .feature_above(feature_aboves[2264]), .feature_below(feature_belows[2264]), .scan_win_std_dev(scan_win_std_dev[2264]), .feature_accum(feature_accums[2264]));
  accum_calculator ac2265(.scan_win(scan_win2265), .rectangle1_x(rectangle1_xs[2265]), .rectangle1_y(rectangle1_ys[2265]), .rectangle1_width(rectangle1_widths[2265]), .rectangle1_height(rectangle1_heights[2265]), .rectangle1_weight(rectangle1_weights[2265]), .rectangle2_x(rectangle2_xs[2265]), .rectangle2_y(rectangle2_ys[2265]), .rectangle2_width(rectangle2_widths[2265]), .rectangle2_height(rectangle2_heights[2265]), .rectangle2_weight(rectangle2_weights[2265]), .rectangle3_x(rectangle3_xs[2265]), .rectangle3_y(rectangle3_ys[2265]), .rectangle3_width(rectangle3_widths[2265]), .rectangle3_height(rectangle3_heights[2265]), .rectangle3_weight(rectangle3_weights[2265]), .feature_threshold(feature_thresholds[2265]), .feature_above(feature_aboves[2265]), .feature_below(feature_belows[2265]), .scan_win_std_dev(scan_win_std_dev[2265]), .feature_accum(feature_accums[2265]));
  accum_calculator ac2266(.scan_win(scan_win2266), .rectangle1_x(rectangle1_xs[2266]), .rectangle1_y(rectangle1_ys[2266]), .rectangle1_width(rectangle1_widths[2266]), .rectangle1_height(rectangle1_heights[2266]), .rectangle1_weight(rectangle1_weights[2266]), .rectangle2_x(rectangle2_xs[2266]), .rectangle2_y(rectangle2_ys[2266]), .rectangle2_width(rectangle2_widths[2266]), .rectangle2_height(rectangle2_heights[2266]), .rectangle2_weight(rectangle2_weights[2266]), .rectangle3_x(rectangle3_xs[2266]), .rectangle3_y(rectangle3_ys[2266]), .rectangle3_width(rectangle3_widths[2266]), .rectangle3_height(rectangle3_heights[2266]), .rectangle3_weight(rectangle3_weights[2266]), .feature_threshold(feature_thresholds[2266]), .feature_above(feature_aboves[2266]), .feature_below(feature_belows[2266]), .scan_win_std_dev(scan_win_std_dev[2266]), .feature_accum(feature_accums[2266]));
  accum_calculator ac2267(.scan_win(scan_win2267), .rectangle1_x(rectangle1_xs[2267]), .rectangle1_y(rectangle1_ys[2267]), .rectangle1_width(rectangle1_widths[2267]), .rectangle1_height(rectangle1_heights[2267]), .rectangle1_weight(rectangle1_weights[2267]), .rectangle2_x(rectangle2_xs[2267]), .rectangle2_y(rectangle2_ys[2267]), .rectangle2_width(rectangle2_widths[2267]), .rectangle2_height(rectangle2_heights[2267]), .rectangle2_weight(rectangle2_weights[2267]), .rectangle3_x(rectangle3_xs[2267]), .rectangle3_y(rectangle3_ys[2267]), .rectangle3_width(rectangle3_widths[2267]), .rectangle3_height(rectangle3_heights[2267]), .rectangle3_weight(rectangle3_weights[2267]), .feature_threshold(feature_thresholds[2267]), .feature_above(feature_aboves[2267]), .feature_below(feature_belows[2267]), .scan_win_std_dev(scan_win_std_dev[2267]), .feature_accum(feature_accums[2267]));
  accum_calculator ac2268(.scan_win(scan_win2268), .rectangle1_x(rectangle1_xs[2268]), .rectangle1_y(rectangle1_ys[2268]), .rectangle1_width(rectangle1_widths[2268]), .rectangle1_height(rectangle1_heights[2268]), .rectangle1_weight(rectangle1_weights[2268]), .rectangle2_x(rectangle2_xs[2268]), .rectangle2_y(rectangle2_ys[2268]), .rectangle2_width(rectangle2_widths[2268]), .rectangle2_height(rectangle2_heights[2268]), .rectangle2_weight(rectangle2_weights[2268]), .rectangle3_x(rectangle3_xs[2268]), .rectangle3_y(rectangle3_ys[2268]), .rectangle3_width(rectangle3_widths[2268]), .rectangle3_height(rectangle3_heights[2268]), .rectangle3_weight(rectangle3_weights[2268]), .feature_threshold(feature_thresholds[2268]), .feature_above(feature_aboves[2268]), .feature_below(feature_belows[2268]), .scan_win_std_dev(scan_win_std_dev[2268]), .feature_accum(feature_accums[2268]));
  accum_calculator ac2269(.scan_win(scan_win2269), .rectangle1_x(rectangle1_xs[2269]), .rectangle1_y(rectangle1_ys[2269]), .rectangle1_width(rectangle1_widths[2269]), .rectangle1_height(rectangle1_heights[2269]), .rectangle1_weight(rectangle1_weights[2269]), .rectangle2_x(rectangle2_xs[2269]), .rectangle2_y(rectangle2_ys[2269]), .rectangle2_width(rectangle2_widths[2269]), .rectangle2_height(rectangle2_heights[2269]), .rectangle2_weight(rectangle2_weights[2269]), .rectangle3_x(rectangle3_xs[2269]), .rectangle3_y(rectangle3_ys[2269]), .rectangle3_width(rectangle3_widths[2269]), .rectangle3_height(rectangle3_heights[2269]), .rectangle3_weight(rectangle3_weights[2269]), .feature_threshold(feature_thresholds[2269]), .feature_above(feature_aboves[2269]), .feature_below(feature_belows[2269]), .scan_win_std_dev(scan_win_std_dev[2269]), .feature_accum(feature_accums[2269]));
  accum_calculator ac2270(.scan_win(scan_win2270), .rectangle1_x(rectangle1_xs[2270]), .rectangle1_y(rectangle1_ys[2270]), .rectangle1_width(rectangle1_widths[2270]), .rectangle1_height(rectangle1_heights[2270]), .rectangle1_weight(rectangle1_weights[2270]), .rectangle2_x(rectangle2_xs[2270]), .rectangle2_y(rectangle2_ys[2270]), .rectangle2_width(rectangle2_widths[2270]), .rectangle2_height(rectangle2_heights[2270]), .rectangle2_weight(rectangle2_weights[2270]), .rectangle3_x(rectangle3_xs[2270]), .rectangle3_y(rectangle3_ys[2270]), .rectangle3_width(rectangle3_widths[2270]), .rectangle3_height(rectangle3_heights[2270]), .rectangle3_weight(rectangle3_weights[2270]), .feature_threshold(feature_thresholds[2270]), .feature_above(feature_aboves[2270]), .feature_below(feature_belows[2270]), .scan_win_std_dev(scan_win_std_dev[2270]), .feature_accum(feature_accums[2270]));
  accum_calculator ac2271(.scan_win(scan_win2271), .rectangle1_x(rectangle1_xs[2271]), .rectangle1_y(rectangle1_ys[2271]), .rectangle1_width(rectangle1_widths[2271]), .rectangle1_height(rectangle1_heights[2271]), .rectangle1_weight(rectangle1_weights[2271]), .rectangle2_x(rectangle2_xs[2271]), .rectangle2_y(rectangle2_ys[2271]), .rectangle2_width(rectangle2_widths[2271]), .rectangle2_height(rectangle2_heights[2271]), .rectangle2_weight(rectangle2_weights[2271]), .rectangle3_x(rectangle3_xs[2271]), .rectangle3_y(rectangle3_ys[2271]), .rectangle3_width(rectangle3_widths[2271]), .rectangle3_height(rectangle3_heights[2271]), .rectangle3_weight(rectangle3_weights[2271]), .feature_threshold(feature_thresholds[2271]), .feature_above(feature_aboves[2271]), .feature_below(feature_belows[2271]), .scan_win_std_dev(scan_win_std_dev[2271]), .feature_accum(feature_accums[2271]));
  accum_calculator ac2272(.scan_win(scan_win2272), .rectangle1_x(rectangle1_xs[2272]), .rectangle1_y(rectangle1_ys[2272]), .rectangle1_width(rectangle1_widths[2272]), .rectangle1_height(rectangle1_heights[2272]), .rectangle1_weight(rectangle1_weights[2272]), .rectangle2_x(rectangle2_xs[2272]), .rectangle2_y(rectangle2_ys[2272]), .rectangle2_width(rectangle2_widths[2272]), .rectangle2_height(rectangle2_heights[2272]), .rectangle2_weight(rectangle2_weights[2272]), .rectangle3_x(rectangle3_xs[2272]), .rectangle3_y(rectangle3_ys[2272]), .rectangle3_width(rectangle3_widths[2272]), .rectangle3_height(rectangle3_heights[2272]), .rectangle3_weight(rectangle3_weights[2272]), .feature_threshold(feature_thresholds[2272]), .feature_above(feature_aboves[2272]), .feature_below(feature_belows[2272]), .scan_win_std_dev(scan_win_std_dev[2272]), .feature_accum(feature_accums[2272]));
  accum_calculator ac2273(.scan_win(scan_win2273), .rectangle1_x(rectangle1_xs[2273]), .rectangle1_y(rectangle1_ys[2273]), .rectangle1_width(rectangle1_widths[2273]), .rectangle1_height(rectangle1_heights[2273]), .rectangle1_weight(rectangle1_weights[2273]), .rectangle2_x(rectangle2_xs[2273]), .rectangle2_y(rectangle2_ys[2273]), .rectangle2_width(rectangle2_widths[2273]), .rectangle2_height(rectangle2_heights[2273]), .rectangle2_weight(rectangle2_weights[2273]), .rectangle3_x(rectangle3_xs[2273]), .rectangle3_y(rectangle3_ys[2273]), .rectangle3_width(rectangle3_widths[2273]), .rectangle3_height(rectangle3_heights[2273]), .rectangle3_weight(rectangle3_weights[2273]), .feature_threshold(feature_thresholds[2273]), .feature_above(feature_aboves[2273]), .feature_below(feature_belows[2273]), .scan_win_std_dev(scan_win_std_dev[2273]), .feature_accum(feature_accums[2273]));
  accum_calculator ac2274(.scan_win(scan_win2274), .rectangle1_x(rectangle1_xs[2274]), .rectangle1_y(rectangle1_ys[2274]), .rectangle1_width(rectangle1_widths[2274]), .rectangle1_height(rectangle1_heights[2274]), .rectangle1_weight(rectangle1_weights[2274]), .rectangle2_x(rectangle2_xs[2274]), .rectangle2_y(rectangle2_ys[2274]), .rectangle2_width(rectangle2_widths[2274]), .rectangle2_height(rectangle2_heights[2274]), .rectangle2_weight(rectangle2_weights[2274]), .rectangle3_x(rectangle3_xs[2274]), .rectangle3_y(rectangle3_ys[2274]), .rectangle3_width(rectangle3_widths[2274]), .rectangle3_height(rectangle3_heights[2274]), .rectangle3_weight(rectangle3_weights[2274]), .feature_threshold(feature_thresholds[2274]), .feature_above(feature_aboves[2274]), .feature_below(feature_belows[2274]), .scan_win_std_dev(scan_win_std_dev[2274]), .feature_accum(feature_accums[2274]));
  accum_calculator ac2275(.scan_win(scan_win2275), .rectangle1_x(rectangle1_xs[2275]), .rectangle1_y(rectangle1_ys[2275]), .rectangle1_width(rectangle1_widths[2275]), .rectangle1_height(rectangle1_heights[2275]), .rectangle1_weight(rectangle1_weights[2275]), .rectangle2_x(rectangle2_xs[2275]), .rectangle2_y(rectangle2_ys[2275]), .rectangle2_width(rectangle2_widths[2275]), .rectangle2_height(rectangle2_heights[2275]), .rectangle2_weight(rectangle2_weights[2275]), .rectangle3_x(rectangle3_xs[2275]), .rectangle3_y(rectangle3_ys[2275]), .rectangle3_width(rectangle3_widths[2275]), .rectangle3_height(rectangle3_heights[2275]), .rectangle3_weight(rectangle3_weights[2275]), .feature_threshold(feature_thresholds[2275]), .feature_above(feature_aboves[2275]), .feature_below(feature_belows[2275]), .scan_win_std_dev(scan_win_std_dev[2275]), .feature_accum(feature_accums[2275]));
  accum_calculator ac2276(.scan_win(scan_win2276), .rectangle1_x(rectangle1_xs[2276]), .rectangle1_y(rectangle1_ys[2276]), .rectangle1_width(rectangle1_widths[2276]), .rectangle1_height(rectangle1_heights[2276]), .rectangle1_weight(rectangle1_weights[2276]), .rectangle2_x(rectangle2_xs[2276]), .rectangle2_y(rectangle2_ys[2276]), .rectangle2_width(rectangle2_widths[2276]), .rectangle2_height(rectangle2_heights[2276]), .rectangle2_weight(rectangle2_weights[2276]), .rectangle3_x(rectangle3_xs[2276]), .rectangle3_y(rectangle3_ys[2276]), .rectangle3_width(rectangle3_widths[2276]), .rectangle3_height(rectangle3_heights[2276]), .rectangle3_weight(rectangle3_weights[2276]), .feature_threshold(feature_thresholds[2276]), .feature_above(feature_aboves[2276]), .feature_below(feature_belows[2276]), .scan_win_std_dev(scan_win_std_dev[2276]), .feature_accum(feature_accums[2276]));
  accum_calculator ac2277(.scan_win(scan_win2277), .rectangle1_x(rectangle1_xs[2277]), .rectangle1_y(rectangle1_ys[2277]), .rectangle1_width(rectangle1_widths[2277]), .rectangle1_height(rectangle1_heights[2277]), .rectangle1_weight(rectangle1_weights[2277]), .rectangle2_x(rectangle2_xs[2277]), .rectangle2_y(rectangle2_ys[2277]), .rectangle2_width(rectangle2_widths[2277]), .rectangle2_height(rectangle2_heights[2277]), .rectangle2_weight(rectangle2_weights[2277]), .rectangle3_x(rectangle3_xs[2277]), .rectangle3_y(rectangle3_ys[2277]), .rectangle3_width(rectangle3_widths[2277]), .rectangle3_height(rectangle3_heights[2277]), .rectangle3_weight(rectangle3_weights[2277]), .feature_threshold(feature_thresholds[2277]), .feature_above(feature_aboves[2277]), .feature_below(feature_belows[2277]), .scan_win_std_dev(scan_win_std_dev[2277]), .feature_accum(feature_accums[2277]));
  accum_calculator ac2278(.scan_win(scan_win2278), .rectangle1_x(rectangle1_xs[2278]), .rectangle1_y(rectangle1_ys[2278]), .rectangle1_width(rectangle1_widths[2278]), .rectangle1_height(rectangle1_heights[2278]), .rectangle1_weight(rectangle1_weights[2278]), .rectangle2_x(rectangle2_xs[2278]), .rectangle2_y(rectangle2_ys[2278]), .rectangle2_width(rectangle2_widths[2278]), .rectangle2_height(rectangle2_heights[2278]), .rectangle2_weight(rectangle2_weights[2278]), .rectangle3_x(rectangle3_xs[2278]), .rectangle3_y(rectangle3_ys[2278]), .rectangle3_width(rectangle3_widths[2278]), .rectangle3_height(rectangle3_heights[2278]), .rectangle3_weight(rectangle3_weights[2278]), .feature_threshold(feature_thresholds[2278]), .feature_above(feature_aboves[2278]), .feature_below(feature_belows[2278]), .scan_win_std_dev(scan_win_std_dev[2278]), .feature_accum(feature_accums[2278]));
  accum_calculator ac2279(.scan_win(scan_win2279), .rectangle1_x(rectangle1_xs[2279]), .rectangle1_y(rectangle1_ys[2279]), .rectangle1_width(rectangle1_widths[2279]), .rectangle1_height(rectangle1_heights[2279]), .rectangle1_weight(rectangle1_weights[2279]), .rectangle2_x(rectangle2_xs[2279]), .rectangle2_y(rectangle2_ys[2279]), .rectangle2_width(rectangle2_widths[2279]), .rectangle2_height(rectangle2_heights[2279]), .rectangle2_weight(rectangle2_weights[2279]), .rectangle3_x(rectangle3_xs[2279]), .rectangle3_y(rectangle3_ys[2279]), .rectangle3_width(rectangle3_widths[2279]), .rectangle3_height(rectangle3_heights[2279]), .rectangle3_weight(rectangle3_weights[2279]), .feature_threshold(feature_thresholds[2279]), .feature_above(feature_aboves[2279]), .feature_below(feature_belows[2279]), .scan_win_std_dev(scan_win_std_dev[2279]), .feature_accum(feature_accums[2279]));
  accum_calculator ac2280(.scan_win(scan_win2280), .rectangle1_x(rectangle1_xs[2280]), .rectangle1_y(rectangle1_ys[2280]), .rectangle1_width(rectangle1_widths[2280]), .rectangle1_height(rectangle1_heights[2280]), .rectangle1_weight(rectangle1_weights[2280]), .rectangle2_x(rectangle2_xs[2280]), .rectangle2_y(rectangle2_ys[2280]), .rectangle2_width(rectangle2_widths[2280]), .rectangle2_height(rectangle2_heights[2280]), .rectangle2_weight(rectangle2_weights[2280]), .rectangle3_x(rectangle3_xs[2280]), .rectangle3_y(rectangle3_ys[2280]), .rectangle3_width(rectangle3_widths[2280]), .rectangle3_height(rectangle3_heights[2280]), .rectangle3_weight(rectangle3_weights[2280]), .feature_threshold(feature_thresholds[2280]), .feature_above(feature_aboves[2280]), .feature_below(feature_belows[2280]), .scan_win_std_dev(scan_win_std_dev[2280]), .feature_accum(feature_accums[2280]));
  accum_calculator ac2281(.scan_win(scan_win2281), .rectangle1_x(rectangle1_xs[2281]), .rectangle1_y(rectangle1_ys[2281]), .rectangle1_width(rectangle1_widths[2281]), .rectangle1_height(rectangle1_heights[2281]), .rectangle1_weight(rectangle1_weights[2281]), .rectangle2_x(rectangle2_xs[2281]), .rectangle2_y(rectangle2_ys[2281]), .rectangle2_width(rectangle2_widths[2281]), .rectangle2_height(rectangle2_heights[2281]), .rectangle2_weight(rectangle2_weights[2281]), .rectangle3_x(rectangle3_xs[2281]), .rectangle3_y(rectangle3_ys[2281]), .rectangle3_width(rectangle3_widths[2281]), .rectangle3_height(rectangle3_heights[2281]), .rectangle3_weight(rectangle3_weights[2281]), .feature_threshold(feature_thresholds[2281]), .feature_above(feature_aboves[2281]), .feature_below(feature_belows[2281]), .scan_win_std_dev(scan_win_std_dev[2281]), .feature_accum(feature_accums[2281]));
  accum_calculator ac2282(.scan_win(scan_win2282), .rectangle1_x(rectangle1_xs[2282]), .rectangle1_y(rectangle1_ys[2282]), .rectangle1_width(rectangle1_widths[2282]), .rectangle1_height(rectangle1_heights[2282]), .rectangle1_weight(rectangle1_weights[2282]), .rectangle2_x(rectangle2_xs[2282]), .rectangle2_y(rectangle2_ys[2282]), .rectangle2_width(rectangle2_widths[2282]), .rectangle2_height(rectangle2_heights[2282]), .rectangle2_weight(rectangle2_weights[2282]), .rectangle3_x(rectangle3_xs[2282]), .rectangle3_y(rectangle3_ys[2282]), .rectangle3_width(rectangle3_widths[2282]), .rectangle3_height(rectangle3_heights[2282]), .rectangle3_weight(rectangle3_weights[2282]), .feature_threshold(feature_thresholds[2282]), .feature_above(feature_aboves[2282]), .feature_below(feature_belows[2282]), .scan_win_std_dev(scan_win_std_dev[2282]), .feature_accum(feature_accums[2282]));
  accum_calculator ac2283(.scan_win(scan_win2283), .rectangle1_x(rectangle1_xs[2283]), .rectangle1_y(rectangle1_ys[2283]), .rectangle1_width(rectangle1_widths[2283]), .rectangle1_height(rectangle1_heights[2283]), .rectangle1_weight(rectangle1_weights[2283]), .rectangle2_x(rectangle2_xs[2283]), .rectangle2_y(rectangle2_ys[2283]), .rectangle2_width(rectangle2_widths[2283]), .rectangle2_height(rectangle2_heights[2283]), .rectangle2_weight(rectangle2_weights[2283]), .rectangle3_x(rectangle3_xs[2283]), .rectangle3_y(rectangle3_ys[2283]), .rectangle3_width(rectangle3_widths[2283]), .rectangle3_height(rectangle3_heights[2283]), .rectangle3_weight(rectangle3_weights[2283]), .feature_threshold(feature_thresholds[2283]), .feature_above(feature_aboves[2283]), .feature_below(feature_belows[2283]), .scan_win_std_dev(scan_win_std_dev[2283]), .feature_accum(feature_accums[2283]));
  accum_calculator ac2284(.scan_win(scan_win2284), .rectangle1_x(rectangle1_xs[2284]), .rectangle1_y(rectangle1_ys[2284]), .rectangle1_width(rectangle1_widths[2284]), .rectangle1_height(rectangle1_heights[2284]), .rectangle1_weight(rectangle1_weights[2284]), .rectangle2_x(rectangle2_xs[2284]), .rectangle2_y(rectangle2_ys[2284]), .rectangle2_width(rectangle2_widths[2284]), .rectangle2_height(rectangle2_heights[2284]), .rectangle2_weight(rectangle2_weights[2284]), .rectangle3_x(rectangle3_xs[2284]), .rectangle3_y(rectangle3_ys[2284]), .rectangle3_width(rectangle3_widths[2284]), .rectangle3_height(rectangle3_heights[2284]), .rectangle3_weight(rectangle3_weights[2284]), .feature_threshold(feature_thresholds[2284]), .feature_above(feature_aboves[2284]), .feature_below(feature_belows[2284]), .scan_win_std_dev(scan_win_std_dev[2284]), .feature_accum(feature_accums[2284]));
  accum_calculator ac2285(.scan_win(scan_win2285), .rectangle1_x(rectangle1_xs[2285]), .rectangle1_y(rectangle1_ys[2285]), .rectangle1_width(rectangle1_widths[2285]), .rectangle1_height(rectangle1_heights[2285]), .rectangle1_weight(rectangle1_weights[2285]), .rectangle2_x(rectangle2_xs[2285]), .rectangle2_y(rectangle2_ys[2285]), .rectangle2_width(rectangle2_widths[2285]), .rectangle2_height(rectangle2_heights[2285]), .rectangle2_weight(rectangle2_weights[2285]), .rectangle3_x(rectangle3_xs[2285]), .rectangle3_y(rectangle3_ys[2285]), .rectangle3_width(rectangle3_widths[2285]), .rectangle3_height(rectangle3_heights[2285]), .rectangle3_weight(rectangle3_weights[2285]), .feature_threshold(feature_thresholds[2285]), .feature_above(feature_aboves[2285]), .feature_below(feature_belows[2285]), .scan_win_std_dev(scan_win_std_dev[2285]), .feature_accum(feature_accums[2285]));
  accum_calculator ac2286(.scan_win(scan_win2286), .rectangle1_x(rectangle1_xs[2286]), .rectangle1_y(rectangle1_ys[2286]), .rectangle1_width(rectangle1_widths[2286]), .rectangle1_height(rectangle1_heights[2286]), .rectangle1_weight(rectangle1_weights[2286]), .rectangle2_x(rectangle2_xs[2286]), .rectangle2_y(rectangle2_ys[2286]), .rectangle2_width(rectangle2_widths[2286]), .rectangle2_height(rectangle2_heights[2286]), .rectangle2_weight(rectangle2_weights[2286]), .rectangle3_x(rectangle3_xs[2286]), .rectangle3_y(rectangle3_ys[2286]), .rectangle3_width(rectangle3_widths[2286]), .rectangle3_height(rectangle3_heights[2286]), .rectangle3_weight(rectangle3_weights[2286]), .feature_threshold(feature_thresholds[2286]), .feature_above(feature_aboves[2286]), .feature_below(feature_belows[2286]), .scan_win_std_dev(scan_win_std_dev[2286]), .feature_accum(feature_accums[2286]));
  accum_calculator ac2287(.scan_win(scan_win2287), .rectangle1_x(rectangle1_xs[2287]), .rectangle1_y(rectangle1_ys[2287]), .rectangle1_width(rectangle1_widths[2287]), .rectangle1_height(rectangle1_heights[2287]), .rectangle1_weight(rectangle1_weights[2287]), .rectangle2_x(rectangle2_xs[2287]), .rectangle2_y(rectangle2_ys[2287]), .rectangle2_width(rectangle2_widths[2287]), .rectangle2_height(rectangle2_heights[2287]), .rectangle2_weight(rectangle2_weights[2287]), .rectangle3_x(rectangle3_xs[2287]), .rectangle3_y(rectangle3_ys[2287]), .rectangle3_width(rectangle3_widths[2287]), .rectangle3_height(rectangle3_heights[2287]), .rectangle3_weight(rectangle3_weights[2287]), .feature_threshold(feature_thresholds[2287]), .feature_above(feature_aboves[2287]), .feature_below(feature_belows[2287]), .scan_win_std_dev(scan_win_std_dev[2287]), .feature_accum(feature_accums[2287]));
  accum_calculator ac2288(.scan_win(scan_win2288), .rectangle1_x(rectangle1_xs[2288]), .rectangle1_y(rectangle1_ys[2288]), .rectangle1_width(rectangle1_widths[2288]), .rectangle1_height(rectangle1_heights[2288]), .rectangle1_weight(rectangle1_weights[2288]), .rectangle2_x(rectangle2_xs[2288]), .rectangle2_y(rectangle2_ys[2288]), .rectangle2_width(rectangle2_widths[2288]), .rectangle2_height(rectangle2_heights[2288]), .rectangle2_weight(rectangle2_weights[2288]), .rectangle3_x(rectangle3_xs[2288]), .rectangle3_y(rectangle3_ys[2288]), .rectangle3_width(rectangle3_widths[2288]), .rectangle3_height(rectangle3_heights[2288]), .rectangle3_weight(rectangle3_weights[2288]), .feature_threshold(feature_thresholds[2288]), .feature_above(feature_aboves[2288]), .feature_below(feature_belows[2288]), .scan_win_std_dev(scan_win_std_dev[2288]), .feature_accum(feature_accums[2288]));
  accum_calculator ac2289(.scan_win(scan_win2289), .rectangle1_x(rectangle1_xs[2289]), .rectangle1_y(rectangle1_ys[2289]), .rectangle1_width(rectangle1_widths[2289]), .rectangle1_height(rectangle1_heights[2289]), .rectangle1_weight(rectangle1_weights[2289]), .rectangle2_x(rectangle2_xs[2289]), .rectangle2_y(rectangle2_ys[2289]), .rectangle2_width(rectangle2_widths[2289]), .rectangle2_height(rectangle2_heights[2289]), .rectangle2_weight(rectangle2_weights[2289]), .rectangle3_x(rectangle3_xs[2289]), .rectangle3_y(rectangle3_ys[2289]), .rectangle3_width(rectangle3_widths[2289]), .rectangle3_height(rectangle3_heights[2289]), .rectangle3_weight(rectangle3_weights[2289]), .feature_threshold(feature_thresholds[2289]), .feature_above(feature_aboves[2289]), .feature_below(feature_belows[2289]), .scan_win_std_dev(scan_win_std_dev[2289]), .feature_accum(feature_accums[2289]));
  accum_calculator ac2290(.scan_win(scan_win2290), .rectangle1_x(rectangle1_xs[2290]), .rectangle1_y(rectangle1_ys[2290]), .rectangle1_width(rectangle1_widths[2290]), .rectangle1_height(rectangle1_heights[2290]), .rectangle1_weight(rectangle1_weights[2290]), .rectangle2_x(rectangle2_xs[2290]), .rectangle2_y(rectangle2_ys[2290]), .rectangle2_width(rectangle2_widths[2290]), .rectangle2_height(rectangle2_heights[2290]), .rectangle2_weight(rectangle2_weights[2290]), .rectangle3_x(rectangle3_xs[2290]), .rectangle3_y(rectangle3_ys[2290]), .rectangle3_width(rectangle3_widths[2290]), .rectangle3_height(rectangle3_heights[2290]), .rectangle3_weight(rectangle3_weights[2290]), .feature_threshold(feature_thresholds[2290]), .feature_above(feature_aboves[2290]), .feature_below(feature_belows[2290]), .scan_win_std_dev(scan_win_std_dev[2290]), .feature_accum(feature_accums[2290]));
  accum_calculator ac2291(.scan_win(scan_win2291), .rectangle1_x(rectangle1_xs[2291]), .rectangle1_y(rectangle1_ys[2291]), .rectangle1_width(rectangle1_widths[2291]), .rectangle1_height(rectangle1_heights[2291]), .rectangle1_weight(rectangle1_weights[2291]), .rectangle2_x(rectangle2_xs[2291]), .rectangle2_y(rectangle2_ys[2291]), .rectangle2_width(rectangle2_widths[2291]), .rectangle2_height(rectangle2_heights[2291]), .rectangle2_weight(rectangle2_weights[2291]), .rectangle3_x(rectangle3_xs[2291]), .rectangle3_y(rectangle3_ys[2291]), .rectangle3_width(rectangle3_widths[2291]), .rectangle3_height(rectangle3_heights[2291]), .rectangle3_weight(rectangle3_weights[2291]), .feature_threshold(feature_thresholds[2291]), .feature_above(feature_aboves[2291]), .feature_below(feature_belows[2291]), .scan_win_std_dev(scan_win_std_dev[2291]), .feature_accum(feature_accums[2291]));
  accum_calculator ac2292(.scan_win(scan_win2292), .rectangle1_x(rectangle1_xs[2292]), .rectangle1_y(rectangle1_ys[2292]), .rectangle1_width(rectangle1_widths[2292]), .rectangle1_height(rectangle1_heights[2292]), .rectangle1_weight(rectangle1_weights[2292]), .rectangle2_x(rectangle2_xs[2292]), .rectangle2_y(rectangle2_ys[2292]), .rectangle2_width(rectangle2_widths[2292]), .rectangle2_height(rectangle2_heights[2292]), .rectangle2_weight(rectangle2_weights[2292]), .rectangle3_x(rectangle3_xs[2292]), .rectangle3_y(rectangle3_ys[2292]), .rectangle3_width(rectangle3_widths[2292]), .rectangle3_height(rectangle3_heights[2292]), .rectangle3_weight(rectangle3_weights[2292]), .feature_threshold(feature_thresholds[2292]), .feature_above(feature_aboves[2292]), .feature_below(feature_belows[2292]), .scan_win_std_dev(scan_win_std_dev[2292]), .feature_accum(feature_accums[2292]));
  accum_calculator ac2293(.scan_win(scan_win2293), .rectangle1_x(rectangle1_xs[2293]), .rectangle1_y(rectangle1_ys[2293]), .rectangle1_width(rectangle1_widths[2293]), .rectangle1_height(rectangle1_heights[2293]), .rectangle1_weight(rectangle1_weights[2293]), .rectangle2_x(rectangle2_xs[2293]), .rectangle2_y(rectangle2_ys[2293]), .rectangle2_width(rectangle2_widths[2293]), .rectangle2_height(rectangle2_heights[2293]), .rectangle2_weight(rectangle2_weights[2293]), .rectangle3_x(rectangle3_xs[2293]), .rectangle3_y(rectangle3_ys[2293]), .rectangle3_width(rectangle3_widths[2293]), .rectangle3_height(rectangle3_heights[2293]), .rectangle3_weight(rectangle3_weights[2293]), .feature_threshold(feature_thresholds[2293]), .feature_above(feature_aboves[2293]), .feature_below(feature_belows[2293]), .scan_win_std_dev(scan_win_std_dev[2293]), .feature_accum(feature_accums[2293]));
  accum_calculator ac2294(.scan_win(scan_win2294), .rectangle1_x(rectangle1_xs[2294]), .rectangle1_y(rectangle1_ys[2294]), .rectangle1_width(rectangle1_widths[2294]), .rectangle1_height(rectangle1_heights[2294]), .rectangle1_weight(rectangle1_weights[2294]), .rectangle2_x(rectangle2_xs[2294]), .rectangle2_y(rectangle2_ys[2294]), .rectangle2_width(rectangle2_widths[2294]), .rectangle2_height(rectangle2_heights[2294]), .rectangle2_weight(rectangle2_weights[2294]), .rectangle3_x(rectangle3_xs[2294]), .rectangle3_y(rectangle3_ys[2294]), .rectangle3_width(rectangle3_widths[2294]), .rectangle3_height(rectangle3_heights[2294]), .rectangle3_weight(rectangle3_weights[2294]), .feature_threshold(feature_thresholds[2294]), .feature_above(feature_aboves[2294]), .feature_below(feature_belows[2294]), .scan_win_std_dev(scan_win_std_dev[2294]), .feature_accum(feature_accums[2294]));
  accum_calculator ac2295(.scan_win(scan_win2295), .rectangle1_x(rectangle1_xs[2295]), .rectangle1_y(rectangle1_ys[2295]), .rectangle1_width(rectangle1_widths[2295]), .rectangle1_height(rectangle1_heights[2295]), .rectangle1_weight(rectangle1_weights[2295]), .rectangle2_x(rectangle2_xs[2295]), .rectangle2_y(rectangle2_ys[2295]), .rectangle2_width(rectangle2_widths[2295]), .rectangle2_height(rectangle2_heights[2295]), .rectangle2_weight(rectangle2_weights[2295]), .rectangle3_x(rectangle3_xs[2295]), .rectangle3_y(rectangle3_ys[2295]), .rectangle3_width(rectangle3_widths[2295]), .rectangle3_height(rectangle3_heights[2295]), .rectangle3_weight(rectangle3_weights[2295]), .feature_threshold(feature_thresholds[2295]), .feature_above(feature_aboves[2295]), .feature_below(feature_belows[2295]), .scan_win_std_dev(scan_win_std_dev[2295]), .feature_accum(feature_accums[2295]));
  accum_calculator ac2296(.scan_win(scan_win2296), .rectangle1_x(rectangle1_xs[2296]), .rectangle1_y(rectangle1_ys[2296]), .rectangle1_width(rectangle1_widths[2296]), .rectangle1_height(rectangle1_heights[2296]), .rectangle1_weight(rectangle1_weights[2296]), .rectangle2_x(rectangle2_xs[2296]), .rectangle2_y(rectangle2_ys[2296]), .rectangle2_width(rectangle2_widths[2296]), .rectangle2_height(rectangle2_heights[2296]), .rectangle2_weight(rectangle2_weights[2296]), .rectangle3_x(rectangle3_xs[2296]), .rectangle3_y(rectangle3_ys[2296]), .rectangle3_width(rectangle3_widths[2296]), .rectangle3_height(rectangle3_heights[2296]), .rectangle3_weight(rectangle3_weights[2296]), .feature_threshold(feature_thresholds[2296]), .feature_above(feature_aboves[2296]), .feature_below(feature_belows[2296]), .scan_win_std_dev(scan_win_std_dev[2296]), .feature_accum(feature_accums[2296]));
  accum_calculator ac2297(.scan_win(scan_win2297), .rectangle1_x(rectangle1_xs[2297]), .rectangle1_y(rectangle1_ys[2297]), .rectangle1_width(rectangle1_widths[2297]), .rectangle1_height(rectangle1_heights[2297]), .rectangle1_weight(rectangle1_weights[2297]), .rectangle2_x(rectangle2_xs[2297]), .rectangle2_y(rectangle2_ys[2297]), .rectangle2_width(rectangle2_widths[2297]), .rectangle2_height(rectangle2_heights[2297]), .rectangle2_weight(rectangle2_weights[2297]), .rectangle3_x(rectangle3_xs[2297]), .rectangle3_y(rectangle3_ys[2297]), .rectangle3_width(rectangle3_widths[2297]), .rectangle3_height(rectangle3_heights[2297]), .rectangle3_weight(rectangle3_weights[2297]), .feature_threshold(feature_thresholds[2297]), .feature_above(feature_aboves[2297]), .feature_below(feature_belows[2297]), .scan_win_std_dev(scan_win_std_dev[2297]), .feature_accum(feature_accums[2297]));
  accum_calculator ac2298(.scan_win(scan_win2298), .rectangle1_x(rectangle1_xs[2298]), .rectangle1_y(rectangle1_ys[2298]), .rectangle1_width(rectangle1_widths[2298]), .rectangle1_height(rectangle1_heights[2298]), .rectangle1_weight(rectangle1_weights[2298]), .rectangle2_x(rectangle2_xs[2298]), .rectangle2_y(rectangle2_ys[2298]), .rectangle2_width(rectangle2_widths[2298]), .rectangle2_height(rectangle2_heights[2298]), .rectangle2_weight(rectangle2_weights[2298]), .rectangle3_x(rectangle3_xs[2298]), .rectangle3_y(rectangle3_ys[2298]), .rectangle3_width(rectangle3_widths[2298]), .rectangle3_height(rectangle3_heights[2298]), .rectangle3_weight(rectangle3_weights[2298]), .feature_threshold(feature_thresholds[2298]), .feature_above(feature_aboves[2298]), .feature_below(feature_belows[2298]), .scan_win_std_dev(scan_win_std_dev[2298]), .feature_accum(feature_accums[2298]));
  accum_calculator ac2299(.scan_win(scan_win2299), .rectangle1_x(rectangle1_xs[2299]), .rectangle1_y(rectangle1_ys[2299]), .rectangle1_width(rectangle1_widths[2299]), .rectangle1_height(rectangle1_heights[2299]), .rectangle1_weight(rectangle1_weights[2299]), .rectangle2_x(rectangle2_xs[2299]), .rectangle2_y(rectangle2_ys[2299]), .rectangle2_width(rectangle2_widths[2299]), .rectangle2_height(rectangle2_heights[2299]), .rectangle2_weight(rectangle2_weights[2299]), .rectangle3_x(rectangle3_xs[2299]), .rectangle3_y(rectangle3_ys[2299]), .rectangle3_width(rectangle3_widths[2299]), .rectangle3_height(rectangle3_heights[2299]), .rectangle3_weight(rectangle3_weights[2299]), .feature_threshold(feature_thresholds[2299]), .feature_above(feature_aboves[2299]), .feature_below(feature_belows[2299]), .scan_win_std_dev(scan_win_std_dev[2299]), .feature_accum(feature_accums[2299]));
  accum_calculator ac2300(.scan_win(scan_win2300), .rectangle1_x(rectangle1_xs[2300]), .rectangle1_y(rectangle1_ys[2300]), .rectangle1_width(rectangle1_widths[2300]), .rectangle1_height(rectangle1_heights[2300]), .rectangle1_weight(rectangle1_weights[2300]), .rectangle2_x(rectangle2_xs[2300]), .rectangle2_y(rectangle2_ys[2300]), .rectangle2_width(rectangle2_widths[2300]), .rectangle2_height(rectangle2_heights[2300]), .rectangle2_weight(rectangle2_weights[2300]), .rectangle3_x(rectangle3_xs[2300]), .rectangle3_y(rectangle3_ys[2300]), .rectangle3_width(rectangle3_widths[2300]), .rectangle3_height(rectangle3_heights[2300]), .rectangle3_weight(rectangle3_weights[2300]), .feature_threshold(feature_thresholds[2300]), .feature_above(feature_aboves[2300]), .feature_below(feature_belows[2300]), .scan_win_std_dev(scan_win_std_dev[2300]), .feature_accum(feature_accums[2300]));
  accum_calculator ac2301(.scan_win(scan_win2301), .rectangle1_x(rectangle1_xs[2301]), .rectangle1_y(rectangle1_ys[2301]), .rectangle1_width(rectangle1_widths[2301]), .rectangle1_height(rectangle1_heights[2301]), .rectangle1_weight(rectangle1_weights[2301]), .rectangle2_x(rectangle2_xs[2301]), .rectangle2_y(rectangle2_ys[2301]), .rectangle2_width(rectangle2_widths[2301]), .rectangle2_height(rectangle2_heights[2301]), .rectangle2_weight(rectangle2_weights[2301]), .rectangle3_x(rectangle3_xs[2301]), .rectangle3_y(rectangle3_ys[2301]), .rectangle3_width(rectangle3_widths[2301]), .rectangle3_height(rectangle3_heights[2301]), .rectangle3_weight(rectangle3_weights[2301]), .feature_threshold(feature_thresholds[2301]), .feature_above(feature_aboves[2301]), .feature_below(feature_belows[2301]), .scan_win_std_dev(scan_win_std_dev[2301]), .feature_accum(feature_accums[2301]));
  accum_calculator ac2302(.scan_win(scan_win2302), .rectangle1_x(rectangle1_xs[2302]), .rectangle1_y(rectangle1_ys[2302]), .rectangle1_width(rectangle1_widths[2302]), .rectangle1_height(rectangle1_heights[2302]), .rectangle1_weight(rectangle1_weights[2302]), .rectangle2_x(rectangle2_xs[2302]), .rectangle2_y(rectangle2_ys[2302]), .rectangle2_width(rectangle2_widths[2302]), .rectangle2_height(rectangle2_heights[2302]), .rectangle2_weight(rectangle2_weights[2302]), .rectangle3_x(rectangle3_xs[2302]), .rectangle3_y(rectangle3_ys[2302]), .rectangle3_width(rectangle3_widths[2302]), .rectangle3_height(rectangle3_heights[2302]), .rectangle3_weight(rectangle3_weights[2302]), .feature_threshold(feature_thresholds[2302]), .feature_above(feature_aboves[2302]), .feature_below(feature_belows[2302]), .scan_win_std_dev(scan_win_std_dev[2302]), .feature_accum(feature_accums[2302]));
  accum_calculator ac2303(.scan_win(scan_win2303), .rectangle1_x(rectangle1_xs[2303]), .rectangle1_y(rectangle1_ys[2303]), .rectangle1_width(rectangle1_widths[2303]), .rectangle1_height(rectangle1_heights[2303]), .rectangle1_weight(rectangle1_weights[2303]), .rectangle2_x(rectangle2_xs[2303]), .rectangle2_y(rectangle2_ys[2303]), .rectangle2_width(rectangle2_widths[2303]), .rectangle2_height(rectangle2_heights[2303]), .rectangle2_weight(rectangle2_weights[2303]), .rectangle3_x(rectangle3_xs[2303]), .rectangle3_y(rectangle3_ys[2303]), .rectangle3_width(rectangle3_widths[2303]), .rectangle3_height(rectangle3_heights[2303]), .rectangle3_weight(rectangle3_weights[2303]), .feature_threshold(feature_thresholds[2303]), .feature_above(feature_aboves[2303]), .feature_below(feature_belows[2303]), .scan_win_std_dev(scan_win_std_dev[2303]), .feature_accum(feature_accums[2303]));
  accum_calculator ac2304(.scan_win(scan_win2304), .rectangle1_x(rectangle1_xs[2304]), .rectangle1_y(rectangle1_ys[2304]), .rectangle1_width(rectangle1_widths[2304]), .rectangle1_height(rectangle1_heights[2304]), .rectangle1_weight(rectangle1_weights[2304]), .rectangle2_x(rectangle2_xs[2304]), .rectangle2_y(rectangle2_ys[2304]), .rectangle2_width(rectangle2_widths[2304]), .rectangle2_height(rectangle2_heights[2304]), .rectangle2_weight(rectangle2_weights[2304]), .rectangle3_x(rectangle3_xs[2304]), .rectangle3_y(rectangle3_ys[2304]), .rectangle3_width(rectangle3_widths[2304]), .rectangle3_height(rectangle3_heights[2304]), .rectangle3_weight(rectangle3_weights[2304]), .feature_threshold(feature_thresholds[2304]), .feature_above(feature_aboves[2304]), .feature_below(feature_belows[2304]), .scan_win_std_dev(scan_win_std_dev[2304]), .feature_accum(feature_accums[2304]));
  accum_calculator ac2305(.scan_win(scan_win2305), .rectangle1_x(rectangle1_xs[2305]), .rectangle1_y(rectangle1_ys[2305]), .rectangle1_width(rectangle1_widths[2305]), .rectangle1_height(rectangle1_heights[2305]), .rectangle1_weight(rectangle1_weights[2305]), .rectangle2_x(rectangle2_xs[2305]), .rectangle2_y(rectangle2_ys[2305]), .rectangle2_width(rectangle2_widths[2305]), .rectangle2_height(rectangle2_heights[2305]), .rectangle2_weight(rectangle2_weights[2305]), .rectangle3_x(rectangle3_xs[2305]), .rectangle3_y(rectangle3_ys[2305]), .rectangle3_width(rectangle3_widths[2305]), .rectangle3_height(rectangle3_heights[2305]), .rectangle3_weight(rectangle3_weights[2305]), .feature_threshold(feature_thresholds[2305]), .feature_above(feature_aboves[2305]), .feature_below(feature_belows[2305]), .scan_win_std_dev(scan_win_std_dev[2305]), .feature_accum(feature_accums[2305]));
  accum_calculator ac2306(.scan_win(scan_win2306), .rectangle1_x(rectangle1_xs[2306]), .rectangle1_y(rectangle1_ys[2306]), .rectangle1_width(rectangle1_widths[2306]), .rectangle1_height(rectangle1_heights[2306]), .rectangle1_weight(rectangle1_weights[2306]), .rectangle2_x(rectangle2_xs[2306]), .rectangle2_y(rectangle2_ys[2306]), .rectangle2_width(rectangle2_widths[2306]), .rectangle2_height(rectangle2_heights[2306]), .rectangle2_weight(rectangle2_weights[2306]), .rectangle3_x(rectangle3_xs[2306]), .rectangle3_y(rectangle3_ys[2306]), .rectangle3_width(rectangle3_widths[2306]), .rectangle3_height(rectangle3_heights[2306]), .rectangle3_weight(rectangle3_weights[2306]), .feature_threshold(feature_thresholds[2306]), .feature_above(feature_aboves[2306]), .feature_below(feature_belows[2306]), .scan_win_std_dev(scan_win_std_dev[2306]), .feature_accum(feature_accums[2306]));
  accum_calculator ac2307(.scan_win(scan_win2307), .rectangle1_x(rectangle1_xs[2307]), .rectangle1_y(rectangle1_ys[2307]), .rectangle1_width(rectangle1_widths[2307]), .rectangle1_height(rectangle1_heights[2307]), .rectangle1_weight(rectangle1_weights[2307]), .rectangle2_x(rectangle2_xs[2307]), .rectangle2_y(rectangle2_ys[2307]), .rectangle2_width(rectangle2_widths[2307]), .rectangle2_height(rectangle2_heights[2307]), .rectangle2_weight(rectangle2_weights[2307]), .rectangle3_x(rectangle3_xs[2307]), .rectangle3_y(rectangle3_ys[2307]), .rectangle3_width(rectangle3_widths[2307]), .rectangle3_height(rectangle3_heights[2307]), .rectangle3_weight(rectangle3_weights[2307]), .feature_threshold(feature_thresholds[2307]), .feature_above(feature_aboves[2307]), .feature_below(feature_belows[2307]), .scan_win_std_dev(scan_win_std_dev[2307]), .feature_accum(feature_accums[2307]));
  accum_calculator ac2308(.scan_win(scan_win2308), .rectangle1_x(rectangle1_xs[2308]), .rectangle1_y(rectangle1_ys[2308]), .rectangle1_width(rectangle1_widths[2308]), .rectangle1_height(rectangle1_heights[2308]), .rectangle1_weight(rectangle1_weights[2308]), .rectangle2_x(rectangle2_xs[2308]), .rectangle2_y(rectangle2_ys[2308]), .rectangle2_width(rectangle2_widths[2308]), .rectangle2_height(rectangle2_heights[2308]), .rectangle2_weight(rectangle2_weights[2308]), .rectangle3_x(rectangle3_xs[2308]), .rectangle3_y(rectangle3_ys[2308]), .rectangle3_width(rectangle3_widths[2308]), .rectangle3_height(rectangle3_heights[2308]), .rectangle3_weight(rectangle3_weights[2308]), .feature_threshold(feature_thresholds[2308]), .feature_above(feature_aboves[2308]), .feature_below(feature_belows[2308]), .scan_win_std_dev(scan_win_std_dev[2308]), .feature_accum(feature_accums[2308]));
  accum_calculator ac2309(.scan_win(scan_win2309), .rectangle1_x(rectangle1_xs[2309]), .rectangle1_y(rectangle1_ys[2309]), .rectangle1_width(rectangle1_widths[2309]), .rectangle1_height(rectangle1_heights[2309]), .rectangle1_weight(rectangle1_weights[2309]), .rectangle2_x(rectangle2_xs[2309]), .rectangle2_y(rectangle2_ys[2309]), .rectangle2_width(rectangle2_widths[2309]), .rectangle2_height(rectangle2_heights[2309]), .rectangle2_weight(rectangle2_weights[2309]), .rectangle3_x(rectangle3_xs[2309]), .rectangle3_y(rectangle3_ys[2309]), .rectangle3_width(rectangle3_widths[2309]), .rectangle3_height(rectangle3_heights[2309]), .rectangle3_weight(rectangle3_weights[2309]), .feature_threshold(feature_thresholds[2309]), .feature_above(feature_aboves[2309]), .feature_below(feature_belows[2309]), .scan_win_std_dev(scan_win_std_dev[2309]), .feature_accum(feature_accums[2309]));
  accum_calculator ac2310(.scan_win(scan_win2310), .rectangle1_x(rectangle1_xs[2310]), .rectangle1_y(rectangle1_ys[2310]), .rectangle1_width(rectangle1_widths[2310]), .rectangle1_height(rectangle1_heights[2310]), .rectangle1_weight(rectangle1_weights[2310]), .rectangle2_x(rectangle2_xs[2310]), .rectangle2_y(rectangle2_ys[2310]), .rectangle2_width(rectangle2_widths[2310]), .rectangle2_height(rectangle2_heights[2310]), .rectangle2_weight(rectangle2_weights[2310]), .rectangle3_x(rectangle3_xs[2310]), .rectangle3_y(rectangle3_ys[2310]), .rectangle3_width(rectangle3_widths[2310]), .rectangle3_height(rectangle3_heights[2310]), .rectangle3_weight(rectangle3_weights[2310]), .feature_threshold(feature_thresholds[2310]), .feature_above(feature_aboves[2310]), .feature_below(feature_belows[2310]), .scan_win_std_dev(scan_win_std_dev[2310]), .feature_accum(feature_accums[2310]));
  accum_calculator ac2311(.scan_win(scan_win2311), .rectangle1_x(rectangle1_xs[2311]), .rectangle1_y(rectangle1_ys[2311]), .rectangle1_width(rectangle1_widths[2311]), .rectangle1_height(rectangle1_heights[2311]), .rectangle1_weight(rectangle1_weights[2311]), .rectangle2_x(rectangle2_xs[2311]), .rectangle2_y(rectangle2_ys[2311]), .rectangle2_width(rectangle2_widths[2311]), .rectangle2_height(rectangle2_heights[2311]), .rectangle2_weight(rectangle2_weights[2311]), .rectangle3_x(rectangle3_xs[2311]), .rectangle3_y(rectangle3_ys[2311]), .rectangle3_width(rectangle3_widths[2311]), .rectangle3_height(rectangle3_heights[2311]), .rectangle3_weight(rectangle3_weights[2311]), .feature_threshold(feature_thresholds[2311]), .feature_above(feature_aboves[2311]), .feature_below(feature_belows[2311]), .scan_win_std_dev(scan_win_std_dev[2311]), .feature_accum(feature_accums[2311]));
  accum_calculator ac2312(.scan_win(scan_win2312), .rectangle1_x(rectangle1_xs[2312]), .rectangle1_y(rectangle1_ys[2312]), .rectangle1_width(rectangle1_widths[2312]), .rectangle1_height(rectangle1_heights[2312]), .rectangle1_weight(rectangle1_weights[2312]), .rectangle2_x(rectangle2_xs[2312]), .rectangle2_y(rectangle2_ys[2312]), .rectangle2_width(rectangle2_widths[2312]), .rectangle2_height(rectangle2_heights[2312]), .rectangle2_weight(rectangle2_weights[2312]), .rectangle3_x(rectangle3_xs[2312]), .rectangle3_y(rectangle3_ys[2312]), .rectangle3_width(rectangle3_widths[2312]), .rectangle3_height(rectangle3_heights[2312]), .rectangle3_weight(rectangle3_weights[2312]), .feature_threshold(feature_thresholds[2312]), .feature_above(feature_aboves[2312]), .feature_below(feature_belows[2312]), .scan_win_std_dev(scan_win_std_dev[2312]), .feature_accum(feature_accums[2312]));
  accum_calculator ac2313(.scan_win(scan_win2313), .rectangle1_x(rectangle1_xs[2313]), .rectangle1_y(rectangle1_ys[2313]), .rectangle1_width(rectangle1_widths[2313]), .rectangle1_height(rectangle1_heights[2313]), .rectangle1_weight(rectangle1_weights[2313]), .rectangle2_x(rectangle2_xs[2313]), .rectangle2_y(rectangle2_ys[2313]), .rectangle2_width(rectangle2_widths[2313]), .rectangle2_height(rectangle2_heights[2313]), .rectangle2_weight(rectangle2_weights[2313]), .rectangle3_x(rectangle3_xs[2313]), .rectangle3_y(rectangle3_ys[2313]), .rectangle3_width(rectangle3_widths[2313]), .rectangle3_height(rectangle3_heights[2313]), .rectangle3_weight(rectangle3_weights[2313]), .feature_threshold(feature_thresholds[2313]), .feature_above(feature_aboves[2313]), .feature_below(feature_belows[2313]), .scan_win_std_dev(scan_win_std_dev[2313]), .feature_accum(feature_accums[2313]));
  accum_calculator ac2314(.scan_win(scan_win2314), .rectangle1_x(rectangle1_xs[2314]), .rectangle1_y(rectangle1_ys[2314]), .rectangle1_width(rectangle1_widths[2314]), .rectangle1_height(rectangle1_heights[2314]), .rectangle1_weight(rectangle1_weights[2314]), .rectangle2_x(rectangle2_xs[2314]), .rectangle2_y(rectangle2_ys[2314]), .rectangle2_width(rectangle2_widths[2314]), .rectangle2_height(rectangle2_heights[2314]), .rectangle2_weight(rectangle2_weights[2314]), .rectangle3_x(rectangle3_xs[2314]), .rectangle3_y(rectangle3_ys[2314]), .rectangle3_width(rectangle3_widths[2314]), .rectangle3_height(rectangle3_heights[2314]), .rectangle3_weight(rectangle3_weights[2314]), .feature_threshold(feature_thresholds[2314]), .feature_above(feature_aboves[2314]), .feature_below(feature_belows[2314]), .scan_win_std_dev(scan_win_std_dev[2314]), .feature_accum(feature_accums[2314]));
  accum_calculator ac2315(.scan_win(scan_win2315), .rectangle1_x(rectangle1_xs[2315]), .rectangle1_y(rectangle1_ys[2315]), .rectangle1_width(rectangle1_widths[2315]), .rectangle1_height(rectangle1_heights[2315]), .rectangle1_weight(rectangle1_weights[2315]), .rectangle2_x(rectangle2_xs[2315]), .rectangle2_y(rectangle2_ys[2315]), .rectangle2_width(rectangle2_widths[2315]), .rectangle2_height(rectangle2_heights[2315]), .rectangle2_weight(rectangle2_weights[2315]), .rectangle3_x(rectangle3_xs[2315]), .rectangle3_y(rectangle3_ys[2315]), .rectangle3_width(rectangle3_widths[2315]), .rectangle3_height(rectangle3_heights[2315]), .rectangle3_weight(rectangle3_weights[2315]), .feature_threshold(feature_thresholds[2315]), .feature_above(feature_aboves[2315]), .feature_below(feature_belows[2315]), .scan_win_std_dev(scan_win_std_dev[2315]), .feature_accum(feature_accums[2315]));
  accum_calculator ac2316(.scan_win(scan_win2316), .rectangle1_x(rectangle1_xs[2316]), .rectangle1_y(rectangle1_ys[2316]), .rectangle1_width(rectangle1_widths[2316]), .rectangle1_height(rectangle1_heights[2316]), .rectangle1_weight(rectangle1_weights[2316]), .rectangle2_x(rectangle2_xs[2316]), .rectangle2_y(rectangle2_ys[2316]), .rectangle2_width(rectangle2_widths[2316]), .rectangle2_height(rectangle2_heights[2316]), .rectangle2_weight(rectangle2_weights[2316]), .rectangle3_x(rectangle3_xs[2316]), .rectangle3_y(rectangle3_ys[2316]), .rectangle3_width(rectangle3_widths[2316]), .rectangle3_height(rectangle3_heights[2316]), .rectangle3_weight(rectangle3_weights[2316]), .feature_threshold(feature_thresholds[2316]), .feature_above(feature_aboves[2316]), .feature_below(feature_belows[2316]), .scan_win_std_dev(scan_win_std_dev[2316]), .feature_accum(feature_accums[2316]));
  accum_calculator ac2317(.scan_win(scan_win2317), .rectangle1_x(rectangle1_xs[2317]), .rectangle1_y(rectangle1_ys[2317]), .rectangle1_width(rectangle1_widths[2317]), .rectangle1_height(rectangle1_heights[2317]), .rectangle1_weight(rectangle1_weights[2317]), .rectangle2_x(rectangle2_xs[2317]), .rectangle2_y(rectangle2_ys[2317]), .rectangle2_width(rectangle2_widths[2317]), .rectangle2_height(rectangle2_heights[2317]), .rectangle2_weight(rectangle2_weights[2317]), .rectangle3_x(rectangle3_xs[2317]), .rectangle3_y(rectangle3_ys[2317]), .rectangle3_width(rectangle3_widths[2317]), .rectangle3_height(rectangle3_heights[2317]), .rectangle3_weight(rectangle3_weights[2317]), .feature_threshold(feature_thresholds[2317]), .feature_above(feature_aboves[2317]), .feature_below(feature_belows[2317]), .scan_win_std_dev(scan_win_std_dev[2317]), .feature_accum(feature_accums[2317]));
  accum_calculator ac2318(.scan_win(scan_win2318), .rectangle1_x(rectangle1_xs[2318]), .rectangle1_y(rectangle1_ys[2318]), .rectangle1_width(rectangle1_widths[2318]), .rectangle1_height(rectangle1_heights[2318]), .rectangle1_weight(rectangle1_weights[2318]), .rectangle2_x(rectangle2_xs[2318]), .rectangle2_y(rectangle2_ys[2318]), .rectangle2_width(rectangle2_widths[2318]), .rectangle2_height(rectangle2_heights[2318]), .rectangle2_weight(rectangle2_weights[2318]), .rectangle3_x(rectangle3_xs[2318]), .rectangle3_y(rectangle3_ys[2318]), .rectangle3_width(rectangle3_widths[2318]), .rectangle3_height(rectangle3_heights[2318]), .rectangle3_weight(rectangle3_weights[2318]), .feature_threshold(feature_thresholds[2318]), .feature_above(feature_aboves[2318]), .feature_below(feature_belows[2318]), .scan_win_std_dev(scan_win_std_dev[2318]), .feature_accum(feature_accums[2318]));
  accum_calculator ac2319(.scan_win(scan_win2319), .rectangle1_x(rectangle1_xs[2319]), .rectangle1_y(rectangle1_ys[2319]), .rectangle1_width(rectangle1_widths[2319]), .rectangle1_height(rectangle1_heights[2319]), .rectangle1_weight(rectangle1_weights[2319]), .rectangle2_x(rectangle2_xs[2319]), .rectangle2_y(rectangle2_ys[2319]), .rectangle2_width(rectangle2_widths[2319]), .rectangle2_height(rectangle2_heights[2319]), .rectangle2_weight(rectangle2_weights[2319]), .rectangle3_x(rectangle3_xs[2319]), .rectangle3_y(rectangle3_ys[2319]), .rectangle3_width(rectangle3_widths[2319]), .rectangle3_height(rectangle3_heights[2319]), .rectangle3_weight(rectangle3_weights[2319]), .feature_threshold(feature_thresholds[2319]), .feature_above(feature_aboves[2319]), .feature_below(feature_belows[2319]), .scan_win_std_dev(scan_win_std_dev[2319]), .feature_accum(feature_accums[2319]));
  accum_calculator ac2320(.scan_win(scan_win2320), .rectangle1_x(rectangle1_xs[2320]), .rectangle1_y(rectangle1_ys[2320]), .rectangle1_width(rectangle1_widths[2320]), .rectangle1_height(rectangle1_heights[2320]), .rectangle1_weight(rectangle1_weights[2320]), .rectangle2_x(rectangle2_xs[2320]), .rectangle2_y(rectangle2_ys[2320]), .rectangle2_width(rectangle2_widths[2320]), .rectangle2_height(rectangle2_heights[2320]), .rectangle2_weight(rectangle2_weights[2320]), .rectangle3_x(rectangle3_xs[2320]), .rectangle3_y(rectangle3_ys[2320]), .rectangle3_width(rectangle3_widths[2320]), .rectangle3_height(rectangle3_heights[2320]), .rectangle3_weight(rectangle3_weights[2320]), .feature_threshold(feature_thresholds[2320]), .feature_above(feature_aboves[2320]), .feature_below(feature_belows[2320]), .scan_win_std_dev(scan_win_std_dev[2320]), .feature_accum(feature_accums[2320]));
  accum_calculator ac2321(.scan_win(scan_win2321), .rectangle1_x(rectangle1_xs[2321]), .rectangle1_y(rectangle1_ys[2321]), .rectangle1_width(rectangle1_widths[2321]), .rectangle1_height(rectangle1_heights[2321]), .rectangle1_weight(rectangle1_weights[2321]), .rectangle2_x(rectangle2_xs[2321]), .rectangle2_y(rectangle2_ys[2321]), .rectangle2_width(rectangle2_widths[2321]), .rectangle2_height(rectangle2_heights[2321]), .rectangle2_weight(rectangle2_weights[2321]), .rectangle3_x(rectangle3_xs[2321]), .rectangle3_y(rectangle3_ys[2321]), .rectangle3_width(rectangle3_widths[2321]), .rectangle3_height(rectangle3_heights[2321]), .rectangle3_weight(rectangle3_weights[2321]), .feature_threshold(feature_thresholds[2321]), .feature_above(feature_aboves[2321]), .feature_below(feature_belows[2321]), .scan_win_std_dev(scan_win_std_dev[2321]), .feature_accum(feature_accums[2321]));
  accum_calculator ac2322(.scan_win(scan_win2322), .rectangle1_x(rectangle1_xs[2322]), .rectangle1_y(rectangle1_ys[2322]), .rectangle1_width(rectangle1_widths[2322]), .rectangle1_height(rectangle1_heights[2322]), .rectangle1_weight(rectangle1_weights[2322]), .rectangle2_x(rectangle2_xs[2322]), .rectangle2_y(rectangle2_ys[2322]), .rectangle2_width(rectangle2_widths[2322]), .rectangle2_height(rectangle2_heights[2322]), .rectangle2_weight(rectangle2_weights[2322]), .rectangle3_x(rectangle3_xs[2322]), .rectangle3_y(rectangle3_ys[2322]), .rectangle3_width(rectangle3_widths[2322]), .rectangle3_height(rectangle3_heights[2322]), .rectangle3_weight(rectangle3_weights[2322]), .feature_threshold(feature_thresholds[2322]), .feature_above(feature_aboves[2322]), .feature_below(feature_belows[2322]), .scan_win_std_dev(scan_win_std_dev[2322]), .feature_accum(feature_accums[2322]));
  accum_calculator ac2323(.scan_win(scan_win2323), .rectangle1_x(rectangle1_xs[2323]), .rectangle1_y(rectangle1_ys[2323]), .rectangle1_width(rectangle1_widths[2323]), .rectangle1_height(rectangle1_heights[2323]), .rectangle1_weight(rectangle1_weights[2323]), .rectangle2_x(rectangle2_xs[2323]), .rectangle2_y(rectangle2_ys[2323]), .rectangle2_width(rectangle2_widths[2323]), .rectangle2_height(rectangle2_heights[2323]), .rectangle2_weight(rectangle2_weights[2323]), .rectangle3_x(rectangle3_xs[2323]), .rectangle3_y(rectangle3_ys[2323]), .rectangle3_width(rectangle3_widths[2323]), .rectangle3_height(rectangle3_heights[2323]), .rectangle3_weight(rectangle3_weights[2323]), .feature_threshold(feature_thresholds[2323]), .feature_above(feature_aboves[2323]), .feature_below(feature_belows[2323]), .scan_win_std_dev(scan_win_std_dev[2323]), .feature_accum(feature_accums[2323]));
  accum_calculator ac2324(.scan_win(scan_win2324), .rectangle1_x(rectangle1_xs[2324]), .rectangle1_y(rectangle1_ys[2324]), .rectangle1_width(rectangle1_widths[2324]), .rectangle1_height(rectangle1_heights[2324]), .rectangle1_weight(rectangle1_weights[2324]), .rectangle2_x(rectangle2_xs[2324]), .rectangle2_y(rectangle2_ys[2324]), .rectangle2_width(rectangle2_widths[2324]), .rectangle2_height(rectangle2_heights[2324]), .rectangle2_weight(rectangle2_weights[2324]), .rectangle3_x(rectangle3_xs[2324]), .rectangle3_y(rectangle3_ys[2324]), .rectangle3_width(rectangle3_widths[2324]), .rectangle3_height(rectangle3_heights[2324]), .rectangle3_weight(rectangle3_weights[2324]), .feature_threshold(feature_thresholds[2324]), .feature_above(feature_aboves[2324]), .feature_below(feature_belows[2324]), .scan_win_std_dev(scan_win_std_dev[2324]), .feature_accum(feature_accums[2324]));
  accum_calculator ac2325(.scan_win(scan_win2325), .rectangle1_x(rectangle1_xs[2325]), .rectangle1_y(rectangle1_ys[2325]), .rectangle1_width(rectangle1_widths[2325]), .rectangle1_height(rectangle1_heights[2325]), .rectangle1_weight(rectangle1_weights[2325]), .rectangle2_x(rectangle2_xs[2325]), .rectangle2_y(rectangle2_ys[2325]), .rectangle2_width(rectangle2_widths[2325]), .rectangle2_height(rectangle2_heights[2325]), .rectangle2_weight(rectangle2_weights[2325]), .rectangle3_x(rectangle3_xs[2325]), .rectangle3_y(rectangle3_ys[2325]), .rectangle3_width(rectangle3_widths[2325]), .rectangle3_height(rectangle3_heights[2325]), .rectangle3_weight(rectangle3_weights[2325]), .feature_threshold(feature_thresholds[2325]), .feature_above(feature_aboves[2325]), .feature_below(feature_belows[2325]), .scan_win_std_dev(scan_win_std_dev[2325]), .feature_accum(feature_accums[2325]));
  accum_calculator ac2326(.scan_win(scan_win2326), .rectangle1_x(rectangle1_xs[2326]), .rectangle1_y(rectangle1_ys[2326]), .rectangle1_width(rectangle1_widths[2326]), .rectangle1_height(rectangle1_heights[2326]), .rectangle1_weight(rectangle1_weights[2326]), .rectangle2_x(rectangle2_xs[2326]), .rectangle2_y(rectangle2_ys[2326]), .rectangle2_width(rectangle2_widths[2326]), .rectangle2_height(rectangle2_heights[2326]), .rectangle2_weight(rectangle2_weights[2326]), .rectangle3_x(rectangle3_xs[2326]), .rectangle3_y(rectangle3_ys[2326]), .rectangle3_width(rectangle3_widths[2326]), .rectangle3_height(rectangle3_heights[2326]), .rectangle3_weight(rectangle3_weights[2326]), .feature_threshold(feature_thresholds[2326]), .feature_above(feature_aboves[2326]), .feature_below(feature_belows[2326]), .scan_win_std_dev(scan_win_std_dev[2326]), .feature_accum(feature_accums[2326]));
  accum_calculator ac2327(.scan_win(scan_win2327), .rectangle1_x(rectangle1_xs[2327]), .rectangle1_y(rectangle1_ys[2327]), .rectangle1_width(rectangle1_widths[2327]), .rectangle1_height(rectangle1_heights[2327]), .rectangle1_weight(rectangle1_weights[2327]), .rectangle2_x(rectangle2_xs[2327]), .rectangle2_y(rectangle2_ys[2327]), .rectangle2_width(rectangle2_widths[2327]), .rectangle2_height(rectangle2_heights[2327]), .rectangle2_weight(rectangle2_weights[2327]), .rectangle3_x(rectangle3_xs[2327]), .rectangle3_y(rectangle3_ys[2327]), .rectangle3_width(rectangle3_widths[2327]), .rectangle3_height(rectangle3_heights[2327]), .rectangle3_weight(rectangle3_weights[2327]), .feature_threshold(feature_thresholds[2327]), .feature_above(feature_aboves[2327]), .feature_below(feature_belows[2327]), .scan_win_std_dev(scan_win_std_dev[2327]), .feature_accum(feature_accums[2327]));
  accum_calculator ac2328(.scan_win(scan_win2328), .rectangle1_x(rectangle1_xs[2328]), .rectangle1_y(rectangle1_ys[2328]), .rectangle1_width(rectangle1_widths[2328]), .rectangle1_height(rectangle1_heights[2328]), .rectangle1_weight(rectangle1_weights[2328]), .rectangle2_x(rectangle2_xs[2328]), .rectangle2_y(rectangle2_ys[2328]), .rectangle2_width(rectangle2_widths[2328]), .rectangle2_height(rectangle2_heights[2328]), .rectangle2_weight(rectangle2_weights[2328]), .rectangle3_x(rectangle3_xs[2328]), .rectangle3_y(rectangle3_ys[2328]), .rectangle3_width(rectangle3_widths[2328]), .rectangle3_height(rectangle3_heights[2328]), .rectangle3_weight(rectangle3_weights[2328]), .feature_threshold(feature_thresholds[2328]), .feature_above(feature_aboves[2328]), .feature_below(feature_belows[2328]), .scan_win_std_dev(scan_win_std_dev[2328]), .feature_accum(feature_accums[2328]));
  accum_calculator ac2329(.scan_win(scan_win2329), .rectangle1_x(rectangle1_xs[2329]), .rectangle1_y(rectangle1_ys[2329]), .rectangle1_width(rectangle1_widths[2329]), .rectangle1_height(rectangle1_heights[2329]), .rectangle1_weight(rectangle1_weights[2329]), .rectangle2_x(rectangle2_xs[2329]), .rectangle2_y(rectangle2_ys[2329]), .rectangle2_width(rectangle2_widths[2329]), .rectangle2_height(rectangle2_heights[2329]), .rectangle2_weight(rectangle2_weights[2329]), .rectangle3_x(rectangle3_xs[2329]), .rectangle3_y(rectangle3_ys[2329]), .rectangle3_width(rectangle3_widths[2329]), .rectangle3_height(rectangle3_heights[2329]), .rectangle3_weight(rectangle3_weights[2329]), .feature_threshold(feature_thresholds[2329]), .feature_above(feature_aboves[2329]), .feature_below(feature_belows[2329]), .scan_win_std_dev(scan_win_std_dev[2329]), .feature_accum(feature_accums[2329]));
  accum_calculator ac2330(.scan_win(scan_win2330), .rectangle1_x(rectangle1_xs[2330]), .rectangle1_y(rectangle1_ys[2330]), .rectangle1_width(rectangle1_widths[2330]), .rectangle1_height(rectangle1_heights[2330]), .rectangle1_weight(rectangle1_weights[2330]), .rectangle2_x(rectangle2_xs[2330]), .rectangle2_y(rectangle2_ys[2330]), .rectangle2_width(rectangle2_widths[2330]), .rectangle2_height(rectangle2_heights[2330]), .rectangle2_weight(rectangle2_weights[2330]), .rectangle3_x(rectangle3_xs[2330]), .rectangle3_y(rectangle3_ys[2330]), .rectangle3_width(rectangle3_widths[2330]), .rectangle3_height(rectangle3_heights[2330]), .rectangle3_weight(rectangle3_weights[2330]), .feature_threshold(feature_thresholds[2330]), .feature_above(feature_aboves[2330]), .feature_below(feature_belows[2330]), .scan_win_std_dev(scan_win_std_dev[2330]), .feature_accum(feature_accums[2330]));
  accum_calculator ac2331(.scan_win(scan_win2331), .rectangle1_x(rectangle1_xs[2331]), .rectangle1_y(rectangle1_ys[2331]), .rectangle1_width(rectangle1_widths[2331]), .rectangle1_height(rectangle1_heights[2331]), .rectangle1_weight(rectangle1_weights[2331]), .rectangle2_x(rectangle2_xs[2331]), .rectangle2_y(rectangle2_ys[2331]), .rectangle2_width(rectangle2_widths[2331]), .rectangle2_height(rectangle2_heights[2331]), .rectangle2_weight(rectangle2_weights[2331]), .rectangle3_x(rectangle3_xs[2331]), .rectangle3_y(rectangle3_ys[2331]), .rectangle3_width(rectangle3_widths[2331]), .rectangle3_height(rectangle3_heights[2331]), .rectangle3_weight(rectangle3_weights[2331]), .feature_threshold(feature_thresholds[2331]), .feature_above(feature_aboves[2331]), .feature_below(feature_belows[2331]), .scan_win_std_dev(scan_win_std_dev[2331]), .feature_accum(feature_accums[2331]));
  accum_calculator ac2332(.scan_win(scan_win2332), .rectangle1_x(rectangle1_xs[2332]), .rectangle1_y(rectangle1_ys[2332]), .rectangle1_width(rectangle1_widths[2332]), .rectangle1_height(rectangle1_heights[2332]), .rectangle1_weight(rectangle1_weights[2332]), .rectangle2_x(rectangle2_xs[2332]), .rectangle2_y(rectangle2_ys[2332]), .rectangle2_width(rectangle2_widths[2332]), .rectangle2_height(rectangle2_heights[2332]), .rectangle2_weight(rectangle2_weights[2332]), .rectangle3_x(rectangle3_xs[2332]), .rectangle3_y(rectangle3_ys[2332]), .rectangle3_width(rectangle3_widths[2332]), .rectangle3_height(rectangle3_heights[2332]), .rectangle3_weight(rectangle3_weights[2332]), .feature_threshold(feature_thresholds[2332]), .feature_above(feature_aboves[2332]), .feature_below(feature_belows[2332]), .scan_win_std_dev(scan_win_std_dev[2332]), .feature_accum(feature_accums[2332]));
  accum_calculator ac2333(.scan_win(scan_win2333), .rectangle1_x(rectangle1_xs[2333]), .rectangle1_y(rectangle1_ys[2333]), .rectangle1_width(rectangle1_widths[2333]), .rectangle1_height(rectangle1_heights[2333]), .rectangle1_weight(rectangle1_weights[2333]), .rectangle2_x(rectangle2_xs[2333]), .rectangle2_y(rectangle2_ys[2333]), .rectangle2_width(rectangle2_widths[2333]), .rectangle2_height(rectangle2_heights[2333]), .rectangle2_weight(rectangle2_weights[2333]), .rectangle3_x(rectangle3_xs[2333]), .rectangle3_y(rectangle3_ys[2333]), .rectangle3_width(rectangle3_widths[2333]), .rectangle3_height(rectangle3_heights[2333]), .rectangle3_weight(rectangle3_weights[2333]), .feature_threshold(feature_thresholds[2333]), .feature_above(feature_aboves[2333]), .feature_below(feature_belows[2333]), .scan_win_std_dev(scan_win_std_dev[2333]), .feature_accum(feature_accums[2333]));
  accum_calculator ac2334(.scan_win(scan_win2334), .rectangle1_x(rectangle1_xs[2334]), .rectangle1_y(rectangle1_ys[2334]), .rectangle1_width(rectangle1_widths[2334]), .rectangle1_height(rectangle1_heights[2334]), .rectangle1_weight(rectangle1_weights[2334]), .rectangle2_x(rectangle2_xs[2334]), .rectangle2_y(rectangle2_ys[2334]), .rectangle2_width(rectangle2_widths[2334]), .rectangle2_height(rectangle2_heights[2334]), .rectangle2_weight(rectangle2_weights[2334]), .rectangle3_x(rectangle3_xs[2334]), .rectangle3_y(rectangle3_ys[2334]), .rectangle3_width(rectangle3_widths[2334]), .rectangle3_height(rectangle3_heights[2334]), .rectangle3_weight(rectangle3_weights[2334]), .feature_threshold(feature_thresholds[2334]), .feature_above(feature_aboves[2334]), .feature_below(feature_belows[2334]), .scan_win_std_dev(scan_win_std_dev[2334]), .feature_accum(feature_accums[2334]));
  accum_calculator ac2335(.scan_win(scan_win2335), .rectangle1_x(rectangle1_xs[2335]), .rectangle1_y(rectangle1_ys[2335]), .rectangle1_width(rectangle1_widths[2335]), .rectangle1_height(rectangle1_heights[2335]), .rectangle1_weight(rectangle1_weights[2335]), .rectangle2_x(rectangle2_xs[2335]), .rectangle2_y(rectangle2_ys[2335]), .rectangle2_width(rectangle2_widths[2335]), .rectangle2_height(rectangle2_heights[2335]), .rectangle2_weight(rectangle2_weights[2335]), .rectangle3_x(rectangle3_xs[2335]), .rectangle3_y(rectangle3_ys[2335]), .rectangle3_width(rectangle3_widths[2335]), .rectangle3_height(rectangle3_heights[2335]), .rectangle3_weight(rectangle3_weights[2335]), .feature_threshold(feature_thresholds[2335]), .feature_above(feature_aboves[2335]), .feature_below(feature_belows[2335]), .scan_win_std_dev(scan_win_std_dev[2335]), .feature_accum(feature_accums[2335]));
  accum_calculator ac2336(.scan_win(scan_win2336), .rectangle1_x(rectangle1_xs[2336]), .rectangle1_y(rectangle1_ys[2336]), .rectangle1_width(rectangle1_widths[2336]), .rectangle1_height(rectangle1_heights[2336]), .rectangle1_weight(rectangle1_weights[2336]), .rectangle2_x(rectangle2_xs[2336]), .rectangle2_y(rectangle2_ys[2336]), .rectangle2_width(rectangle2_widths[2336]), .rectangle2_height(rectangle2_heights[2336]), .rectangle2_weight(rectangle2_weights[2336]), .rectangle3_x(rectangle3_xs[2336]), .rectangle3_y(rectangle3_ys[2336]), .rectangle3_width(rectangle3_widths[2336]), .rectangle3_height(rectangle3_heights[2336]), .rectangle3_weight(rectangle3_weights[2336]), .feature_threshold(feature_thresholds[2336]), .feature_above(feature_aboves[2336]), .feature_below(feature_belows[2336]), .scan_win_std_dev(scan_win_std_dev[2336]), .feature_accum(feature_accums[2336]));
  accum_calculator ac2337(.scan_win(scan_win2337), .rectangle1_x(rectangle1_xs[2337]), .rectangle1_y(rectangle1_ys[2337]), .rectangle1_width(rectangle1_widths[2337]), .rectangle1_height(rectangle1_heights[2337]), .rectangle1_weight(rectangle1_weights[2337]), .rectangle2_x(rectangle2_xs[2337]), .rectangle2_y(rectangle2_ys[2337]), .rectangle2_width(rectangle2_widths[2337]), .rectangle2_height(rectangle2_heights[2337]), .rectangle2_weight(rectangle2_weights[2337]), .rectangle3_x(rectangle3_xs[2337]), .rectangle3_y(rectangle3_ys[2337]), .rectangle3_width(rectangle3_widths[2337]), .rectangle3_height(rectangle3_heights[2337]), .rectangle3_weight(rectangle3_weights[2337]), .feature_threshold(feature_thresholds[2337]), .feature_above(feature_aboves[2337]), .feature_below(feature_belows[2337]), .scan_win_std_dev(scan_win_std_dev[2337]), .feature_accum(feature_accums[2337]));
  accum_calculator ac2338(.scan_win(scan_win2338), .rectangle1_x(rectangle1_xs[2338]), .rectangle1_y(rectangle1_ys[2338]), .rectangle1_width(rectangle1_widths[2338]), .rectangle1_height(rectangle1_heights[2338]), .rectangle1_weight(rectangle1_weights[2338]), .rectangle2_x(rectangle2_xs[2338]), .rectangle2_y(rectangle2_ys[2338]), .rectangle2_width(rectangle2_widths[2338]), .rectangle2_height(rectangle2_heights[2338]), .rectangle2_weight(rectangle2_weights[2338]), .rectangle3_x(rectangle3_xs[2338]), .rectangle3_y(rectangle3_ys[2338]), .rectangle3_width(rectangle3_widths[2338]), .rectangle3_height(rectangle3_heights[2338]), .rectangle3_weight(rectangle3_weights[2338]), .feature_threshold(feature_thresholds[2338]), .feature_above(feature_aboves[2338]), .feature_below(feature_belows[2338]), .scan_win_std_dev(scan_win_std_dev[2338]), .feature_accum(feature_accums[2338]));
  accum_calculator ac2339(.scan_win(scan_win2339), .rectangle1_x(rectangle1_xs[2339]), .rectangle1_y(rectangle1_ys[2339]), .rectangle1_width(rectangle1_widths[2339]), .rectangle1_height(rectangle1_heights[2339]), .rectangle1_weight(rectangle1_weights[2339]), .rectangle2_x(rectangle2_xs[2339]), .rectangle2_y(rectangle2_ys[2339]), .rectangle2_width(rectangle2_widths[2339]), .rectangle2_height(rectangle2_heights[2339]), .rectangle2_weight(rectangle2_weights[2339]), .rectangle3_x(rectangle3_xs[2339]), .rectangle3_y(rectangle3_ys[2339]), .rectangle3_width(rectangle3_widths[2339]), .rectangle3_height(rectangle3_heights[2339]), .rectangle3_weight(rectangle3_weights[2339]), .feature_threshold(feature_thresholds[2339]), .feature_above(feature_aboves[2339]), .feature_below(feature_belows[2339]), .scan_win_std_dev(scan_win_std_dev[2339]), .feature_accum(feature_accums[2339]));
  accum_calculator ac2340(.scan_win(scan_win2340), .rectangle1_x(rectangle1_xs[2340]), .rectangle1_y(rectangle1_ys[2340]), .rectangle1_width(rectangle1_widths[2340]), .rectangle1_height(rectangle1_heights[2340]), .rectangle1_weight(rectangle1_weights[2340]), .rectangle2_x(rectangle2_xs[2340]), .rectangle2_y(rectangle2_ys[2340]), .rectangle2_width(rectangle2_widths[2340]), .rectangle2_height(rectangle2_heights[2340]), .rectangle2_weight(rectangle2_weights[2340]), .rectangle3_x(rectangle3_xs[2340]), .rectangle3_y(rectangle3_ys[2340]), .rectangle3_width(rectangle3_widths[2340]), .rectangle3_height(rectangle3_heights[2340]), .rectangle3_weight(rectangle3_weights[2340]), .feature_threshold(feature_thresholds[2340]), .feature_above(feature_aboves[2340]), .feature_below(feature_belows[2340]), .scan_win_std_dev(scan_win_std_dev[2340]), .feature_accum(feature_accums[2340]));
  accum_calculator ac2341(.scan_win(scan_win2341), .rectangle1_x(rectangle1_xs[2341]), .rectangle1_y(rectangle1_ys[2341]), .rectangle1_width(rectangle1_widths[2341]), .rectangle1_height(rectangle1_heights[2341]), .rectangle1_weight(rectangle1_weights[2341]), .rectangle2_x(rectangle2_xs[2341]), .rectangle2_y(rectangle2_ys[2341]), .rectangle2_width(rectangle2_widths[2341]), .rectangle2_height(rectangle2_heights[2341]), .rectangle2_weight(rectangle2_weights[2341]), .rectangle3_x(rectangle3_xs[2341]), .rectangle3_y(rectangle3_ys[2341]), .rectangle3_width(rectangle3_widths[2341]), .rectangle3_height(rectangle3_heights[2341]), .rectangle3_weight(rectangle3_weights[2341]), .feature_threshold(feature_thresholds[2341]), .feature_above(feature_aboves[2341]), .feature_below(feature_belows[2341]), .scan_win_std_dev(scan_win_std_dev[2341]), .feature_accum(feature_accums[2341]));
  accum_calculator ac2342(.scan_win(scan_win2342), .rectangle1_x(rectangle1_xs[2342]), .rectangle1_y(rectangle1_ys[2342]), .rectangle1_width(rectangle1_widths[2342]), .rectangle1_height(rectangle1_heights[2342]), .rectangle1_weight(rectangle1_weights[2342]), .rectangle2_x(rectangle2_xs[2342]), .rectangle2_y(rectangle2_ys[2342]), .rectangle2_width(rectangle2_widths[2342]), .rectangle2_height(rectangle2_heights[2342]), .rectangle2_weight(rectangle2_weights[2342]), .rectangle3_x(rectangle3_xs[2342]), .rectangle3_y(rectangle3_ys[2342]), .rectangle3_width(rectangle3_widths[2342]), .rectangle3_height(rectangle3_heights[2342]), .rectangle3_weight(rectangle3_weights[2342]), .feature_threshold(feature_thresholds[2342]), .feature_above(feature_aboves[2342]), .feature_below(feature_belows[2342]), .scan_win_std_dev(scan_win_std_dev[2342]), .feature_accum(feature_accums[2342]));
  accum_calculator ac2343(.scan_win(scan_win2343), .rectangle1_x(rectangle1_xs[2343]), .rectangle1_y(rectangle1_ys[2343]), .rectangle1_width(rectangle1_widths[2343]), .rectangle1_height(rectangle1_heights[2343]), .rectangle1_weight(rectangle1_weights[2343]), .rectangle2_x(rectangle2_xs[2343]), .rectangle2_y(rectangle2_ys[2343]), .rectangle2_width(rectangle2_widths[2343]), .rectangle2_height(rectangle2_heights[2343]), .rectangle2_weight(rectangle2_weights[2343]), .rectangle3_x(rectangle3_xs[2343]), .rectangle3_y(rectangle3_ys[2343]), .rectangle3_width(rectangle3_widths[2343]), .rectangle3_height(rectangle3_heights[2343]), .rectangle3_weight(rectangle3_weights[2343]), .feature_threshold(feature_thresholds[2343]), .feature_above(feature_aboves[2343]), .feature_below(feature_belows[2343]), .scan_win_std_dev(scan_win_std_dev[2343]), .feature_accum(feature_accums[2343]));
  accum_calculator ac2344(.scan_win(scan_win2344), .rectangle1_x(rectangle1_xs[2344]), .rectangle1_y(rectangle1_ys[2344]), .rectangle1_width(rectangle1_widths[2344]), .rectangle1_height(rectangle1_heights[2344]), .rectangle1_weight(rectangle1_weights[2344]), .rectangle2_x(rectangle2_xs[2344]), .rectangle2_y(rectangle2_ys[2344]), .rectangle2_width(rectangle2_widths[2344]), .rectangle2_height(rectangle2_heights[2344]), .rectangle2_weight(rectangle2_weights[2344]), .rectangle3_x(rectangle3_xs[2344]), .rectangle3_y(rectangle3_ys[2344]), .rectangle3_width(rectangle3_widths[2344]), .rectangle3_height(rectangle3_heights[2344]), .rectangle3_weight(rectangle3_weights[2344]), .feature_threshold(feature_thresholds[2344]), .feature_above(feature_aboves[2344]), .feature_below(feature_belows[2344]), .scan_win_std_dev(scan_win_std_dev[2344]), .feature_accum(feature_accums[2344]));
  accum_calculator ac2345(.scan_win(scan_win2345), .rectangle1_x(rectangle1_xs[2345]), .rectangle1_y(rectangle1_ys[2345]), .rectangle1_width(rectangle1_widths[2345]), .rectangle1_height(rectangle1_heights[2345]), .rectangle1_weight(rectangle1_weights[2345]), .rectangle2_x(rectangle2_xs[2345]), .rectangle2_y(rectangle2_ys[2345]), .rectangle2_width(rectangle2_widths[2345]), .rectangle2_height(rectangle2_heights[2345]), .rectangle2_weight(rectangle2_weights[2345]), .rectangle3_x(rectangle3_xs[2345]), .rectangle3_y(rectangle3_ys[2345]), .rectangle3_width(rectangle3_widths[2345]), .rectangle3_height(rectangle3_heights[2345]), .rectangle3_weight(rectangle3_weights[2345]), .feature_threshold(feature_thresholds[2345]), .feature_above(feature_aboves[2345]), .feature_below(feature_belows[2345]), .scan_win_std_dev(scan_win_std_dev[2345]), .feature_accum(feature_accums[2345]));
  accum_calculator ac2346(.scan_win(scan_win2346), .rectangle1_x(rectangle1_xs[2346]), .rectangle1_y(rectangle1_ys[2346]), .rectangle1_width(rectangle1_widths[2346]), .rectangle1_height(rectangle1_heights[2346]), .rectangle1_weight(rectangle1_weights[2346]), .rectangle2_x(rectangle2_xs[2346]), .rectangle2_y(rectangle2_ys[2346]), .rectangle2_width(rectangle2_widths[2346]), .rectangle2_height(rectangle2_heights[2346]), .rectangle2_weight(rectangle2_weights[2346]), .rectangle3_x(rectangle3_xs[2346]), .rectangle3_y(rectangle3_ys[2346]), .rectangle3_width(rectangle3_widths[2346]), .rectangle3_height(rectangle3_heights[2346]), .rectangle3_weight(rectangle3_weights[2346]), .feature_threshold(feature_thresholds[2346]), .feature_above(feature_aboves[2346]), .feature_below(feature_belows[2346]), .scan_win_std_dev(scan_win_std_dev[2346]), .feature_accum(feature_accums[2346]));
  accum_calculator ac2347(.scan_win(scan_win2347), .rectangle1_x(rectangle1_xs[2347]), .rectangle1_y(rectangle1_ys[2347]), .rectangle1_width(rectangle1_widths[2347]), .rectangle1_height(rectangle1_heights[2347]), .rectangle1_weight(rectangle1_weights[2347]), .rectangle2_x(rectangle2_xs[2347]), .rectangle2_y(rectangle2_ys[2347]), .rectangle2_width(rectangle2_widths[2347]), .rectangle2_height(rectangle2_heights[2347]), .rectangle2_weight(rectangle2_weights[2347]), .rectangle3_x(rectangle3_xs[2347]), .rectangle3_y(rectangle3_ys[2347]), .rectangle3_width(rectangle3_widths[2347]), .rectangle3_height(rectangle3_heights[2347]), .rectangle3_weight(rectangle3_weights[2347]), .feature_threshold(feature_thresholds[2347]), .feature_above(feature_aboves[2347]), .feature_below(feature_belows[2347]), .scan_win_std_dev(scan_win_std_dev[2347]), .feature_accum(feature_accums[2347]));
  accum_calculator ac2348(.scan_win(scan_win2348), .rectangle1_x(rectangle1_xs[2348]), .rectangle1_y(rectangle1_ys[2348]), .rectangle1_width(rectangle1_widths[2348]), .rectangle1_height(rectangle1_heights[2348]), .rectangle1_weight(rectangle1_weights[2348]), .rectangle2_x(rectangle2_xs[2348]), .rectangle2_y(rectangle2_ys[2348]), .rectangle2_width(rectangle2_widths[2348]), .rectangle2_height(rectangle2_heights[2348]), .rectangle2_weight(rectangle2_weights[2348]), .rectangle3_x(rectangle3_xs[2348]), .rectangle3_y(rectangle3_ys[2348]), .rectangle3_width(rectangle3_widths[2348]), .rectangle3_height(rectangle3_heights[2348]), .rectangle3_weight(rectangle3_weights[2348]), .feature_threshold(feature_thresholds[2348]), .feature_above(feature_aboves[2348]), .feature_below(feature_belows[2348]), .scan_win_std_dev(scan_win_std_dev[2348]), .feature_accum(feature_accums[2348]));
  accum_calculator ac2349(.scan_win(scan_win2349), .rectangle1_x(rectangle1_xs[2349]), .rectangle1_y(rectangle1_ys[2349]), .rectangle1_width(rectangle1_widths[2349]), .rectangle1_height(rectangle1_heights[2349]), .rectangle1_weight(rectangle1_weights[2349]), .rectangle2_x(rectangle2_xs[2349]), .rectangle2_y(rectangle2_ys[2349]), .rectangle2_width(rectangle2_widths[2349]), .rectangle2_height(rectangle2_heights[2349]), .rectangle2_weight(rectangle2_weights[2349]), .rectangle3_x(rectangle3_xs[2349]), .rectangle3_y(rectangle3_ys[2349]), .rectangle3_width(rectangle3_widths[2349]), .rectangle3_height(rectangle3_heights[2349]), .rectangle3_weight(rectangle3_weights[2349]), .feature_threshold(feature_thresholds[2349]), .feature_above(feature_aboves[2349]), .feature_below(feature_belows[2349]), .scan_win_std_dev(scan_win_std_dev[2349]), .feature_accum(feature_accums[2349]));
  accum_calculator ac2350(.scan_win(scan_win2350), .rectangle1_x(rectangle1_xs[2350]), .rectangle1_y(rectangle1_ys[2350]), .rectangle1_width(rectangle1_widths[2350]), .rectangle1_height(rectangle1_heights[2350]), .rectangle1_weight(rectangle1_weights[2350]), .rectangle2_x(rectangle2_xs[2350]), .rectangle2_y(rectangle2_ys[2350]), .rectangle2_width(rectangle2_widths[2350]), .rectangle2_height(rectangle2_heights[2350]), .rectangle2_weight(rectangle2_weights[2350]), .rectangle3_x(rectangle3_xs[2350]), .rectangle3_y(rectangle3_ys[2350]), .rectangle3_width(rectangle3_widths[2350]), .rectangle3_height(rectangle3_heights[2350]), .rectangle3_weight(rectangle3_weights[2350]), .feature_threshold(feature_thresholds[2350]), .feature_above(feature_aboves[2350]), .feature_below(feature_belows[2350]), .scan_win_std_dev(scan_win_std_dev[2350]), .feature_accum(feature_accums[2350]));
  accum_calculator ac2351(.scan_win(scan_win2351), .rectangle1_x(rectangle1_xs[2351]), .rectangle1_y(rectangle1_ys[2351]), .rectangle1_width(rectangle1_widths[2351]), .rectangle1_height(rectangle1_heights[2351]), .rectangle1_weight(rectangle1_weights[2351]), .rectangle2_x(rectangle2_xs[2351]), .rectangle2_y(rectangle2_ys[2351]), .rectangle2_width(rectangle2_widths[2351]), .rectangle2_height(rectangle2_heights[2351]), .rectangle2_weight(rectangle2_weights[2351]), .rectangle3_x(rectangle3_xs[2351]), .rectangle3_y(rectangle3_ys[2351]), .rectangle3_width(rectangle3_widths[2351]), .rectangle3_height(rectangle3_heights[2351]), .rectangle3_weight(rectangle3_weights[2351]), .feature_threshold(feature_thresholds[2351]), .feature_above(feature_aboves[2351]), .feature_below(feature_belows[2351]), .scan_win_std_dev(scan_win_std_dev[2351]), .feature_accum(feature_accums[2351]));
  accum_calculator ac2352(.scan_win(scan_win2352), .rectangle1_x(rectangle1_xs[2352]), .rectangle1_y(rectangle1_ys[2352]), .rectangle1_width(rectangle1_widths[2352]), .rectangle1_height(rectangle1_heights[2352]), .rectangle1_weight(rectangle1_weights[2352]), .rectangle2_x(rectangle2_xs[2352]), .rectangle2_y(rectangle2_ys[2352]), .rectangle2_width(rectangle2_widths[2352]), .rectangle2_height(rectangle2_heights[2352]), .rectangle2_weight(rectangle2_weights[2352]), .rectangle3_x(rectangle3_xs[2352]), .rectangle3_y(rectangle3_ys[2352]), .rectangle3_width(rectangle3_widths[2352]), .rectangle3_height(rectangle3_heights[2352]), .rectangle3_weight(rectangle3_weights[2352]), .feature_threshold(feature_thresholds[2352]), .feature_above(feature_aboves[2352]), .feature_below(feature_belows[2352]), .scan_win_std_dev(scan_win_std_dev[2352]), .feature_accum(feature_accums[2352]));
  accum_calculator ac2353(.scan_win(scan_win2353), .rectangle1_x(rectangle1_xs[2353]), .rectangle1_y(rectangle1_ys[2353]), .rectangle1_width(rectangle1_widths[2353]), .rectangle1_height(rectangle1_heights[2353]), .rectangle1_weight(rectangle1_weights[2353]), .rectangle2_x(rectangle2_xs[2353]), .rectangle2_y(rectangle2_ys[2353]), .rectangle2_width(rectangle2_widths[2353]), .rectangle2_height(rectangle2_heights[2353]), .rectangle2_weight(rectangle2_weights[2353]), .rectangle3_x(rectangle3_xs[2353]), .rectangle3_y(rectangle3_ys[2353]), .rectangle3_width(rectangle3_widths[2353]), .rectangle3_height(rectangle3_heights[2353]), .rectangle3_weight(rectangle3_weights[2353]), .feature_threshold(feature_thresholds[2353]), .feature_above(feature_aboves[2353]), .feature_below(feature_belows[2353]), .scan_win_std_dev(scan_win_std_dev[2353]), .feature_accum(feature_accums[2353]));
  accum_calculator ac2354(.scan_win(scan_win2354), .rectangle1_x(rectangle1_xs[2354]), .rectangle1_y(rectangle1_ys[2354]), .rectangle1_width(rectangle1_widths[2354]), .rectangle1_height(rectangle1_heights[2354]), .rectangle1_weight(rectangle1_weights[2354]), .rectangle2_x(rectangle2_xs[2354]), .rectangle2_y(rectangle2_ys[2354]), .rectangle2_width(rectangle2_widths[2354]), .rectangle2_height(rectangle2_heights[2354]), .rectangle2_weight(rectangle2_weights[2354]), .rectangle3_x(rectangle3_xs[2354]), .rectangle3_y(rectangle3_ys[2354]), .rectangle3_width(rectangle3_widths[2354]), .rectangle3_height(rectangle3_heights[2354]), .rectangle3_weight(rectangle3_weights[2354]), .feature_threshold(feature_thresholds[2354]), .feature_above(feature_aboves[2354]), .feature_below(feature_belows[2354]), .scan_win_std_dev(scan_win_std_dev[2354]), .feature_accum(feature_accums[2354]));
  accum_calculator ac2355(.scan_win(scan_win2355), .rectangle1_x(rectangle1_xs[2355]), .rectangle1_y(rectangle1_ys[2355]), .rectangle1_width(rectangle1_widths[2355]), .rectangle1_height(rectangle1_heights[2355]), .rectangle1_weight(rectangle1_weights[2355]), .rectangle2_x(rectangle2_xs[2355]), .rectangle2_y(rectangle2_ys[2355]), .rectangle2_width(rectangle2_widths[2355]), .rectangle2_height(rectangle2_heights[2355]), .rectangle2_weight(rectangle2_weights[2355]), .rectangle3_x(rectangle3_xs[2355]), .rectangle3_y(rectangle3_ys[2355]), .rectangle3_width(rectangle3_widths[2355]), .rectangle3_height(rectangle3_heights[2355]), .rectangle3_weight(rectangle3_weights[2355]), .feature_threshold(feature_thresholds[2355]), .feature_above(feature_aboves[2355]), .feature_below(feature_belows[2355]), .scan_win_std_dev(scan_win_std_dev[2355]), .feature_accum(feature_accums[2355]));
  accum_calculator ac2356(.scan_win(scan_win2356), .rectangle1_x(rectangle1_xs[2356]), .rectangle1_y(rectangle1_ys[2356]), .rectangle1_width(rectangle1_widths[2356]), .rectangle1_height(rectangle1_heights[2356]), .rectangle1_weight(rectangle1_weights[2356]), .rectangle2_x(rectangle2_xs[2356]), .rectangle2_y(rectangle2_ys[2356]), .rectangle2_width(rectangle2_widths[2356]), .rectangle2_height(rectangle2_heights[2356]), .rectangle2_weight(rectangle2_weights[2356]), .rectangle3_x(rectangle3_xs[2356]), .rectangle3_y(rectangle3_ys[2356]), .rectangle3_width(rectangle3_widths[2356]), .rectangle3_height(rectangle3_heights[2356]), .rectangle3_weight(rectangle3_weights[2356]), .feature_threshold(feature_thresholds[2356]), .feature_above(feature_aboves[2356]), .feature_below(feature_belows[2356]), .scan_win_std_dev(scan_win_std_dev[2356]), .feature_accum(feature_accums[2356]));
  accum_calculator ac2357(.scan_win(scan_win2357), .rectangle1_x(rectangle1_xs[2357]), .rectangle1_y(rectangle1_ys[2357]), .rectangle1_width(rectangle1_widths[2357]), .rectangle1_height(rectangle1_heights[2357]), .rectangle1_weight(rectangle1_weights[2357]), .rectangle2_x(rectangle2_xs[2357]), .rectangle2_y(rectangle2_ys[2357]), .rectangle2_width(rectangle2_widths[2357]), .rectangle2_height(rectangle2_heights[2357]), .rectangle2_weight(rectangle2_weights[2357]), .rectangle3_x(rectangle3_xs[2357]), .rectangle3_y(rectangle3_ys[2357]), .rectangle3_width(rectangle3_widths[2357]), .rectangle3_height(rectangle3_heights[2357]), .rectangle3_weight(rectangle3_weights[2357]), .feature_threshold(feature_thresholds[2357]), .feature_above(feature_aboves[2357]), .feature_below(feature_belows[2357]), .scan_win_std_dev(scan_win_std_dev[2357]), .feature_accum(feature_accums[2357]));
  accum_calculator ac2358(.scan_win(scan_win2358), .rectangle1_x(rectangle1_xs[2358]), .rectangle1_y(rectangle1_ys[2358]), .rectangle1_width(rectangle1_widths[2358]), .rectangle1_height(rectangle1_heights[2358]), .rectangle1_weight(rectangle1_weights[2358]), .rectangle2_x(rectangle2_xs[2358]), .rectangle2_y(rectangle2_ys[2358]), .rectangle2_width(rectangle2_widths[2358]), .rectangle2_height(rectangle2_heights[2358]), .rectangle2_weight(rectangle2_weights[2358]), .rectangle3_x(rectangle3_xs[2358]), .rectangle3_y(rectangle3_ys[2358]), .rectangle3_width(rectangle3_widths[2358]), .rectangle3_height(rectangle3_heights[2358]), .rectangle3_weight(rectangle3_weights[2358]), .feature_threshold(feature_thresholds[2358]), .feature_above(feature_aboves[2358]), .feature_below(feature_belows[2358]), .scan_win_std_dev(scan_win_std_dev[2358]), .feature_accum(feature_accums[2358]));
  accum_calculator ac2359(.scan_win(scan_win2359), .rectangle1_x(rectangle1_xs[2359]), .rectangle1_y(rectangle1_ys[2359]), .rectangle1_width(rectangle1_widths[2359]), .rectangle1_height(rectangle1_heights[2359]), .rectangle1_weight(rectangle1_weights[2359]), .rectangle2_x(rectangle2_xs[2359]), .rectangle2_y(rectangle2_ys[2359]), .rectangle2_width(rectangle2_widths[2359]), .rectangle2_height(rectangle2_heights[2359]), .rectangle2_weight(rectangle2_weights[2359]), .rectangle3_x(rectangle3_xs[2359]), .rectangle3_y(rectangle3_ys[2359]), .rectangle3_width(rectangle3_widths[2359]), .rectangle3_height(rectangle3_heights[2359]), .rectangle3_weight(rectangle3_weights[2359]), .feature_threshold(feature_thresholds[2359]), .feature_above(feature_aboves[2359]), .feature_below(feature_belows[2359]), .scan_win_std_dev(scan_win_std_dev[2359]), .feature_accum(feature_accums[2359]));
  accum_calculator ac2360(.scan_win(scan_win2360), .rectangle1_x(rectangle1_xs[2360]), .rectangle1_y(rectangle1_ys[2360]), .rectangle1_width(rectangle1_widths[2360]), .rectangle1_height(rectangle1_heights[2360]), .rectangle1_weight(rectangle1_weights[2360]), .rectangle2_x(rectangle2_xs[2360]), .rectangle2_y(rectangle2_ys[2360]), .rectangle2_width(rectangle2_widths[2360]), .rectangle2_height(rectangle2_heights[2360]), .rectangle2_weight(rectangle2_weights[2360]), .rectangle3_x(rectangle3_xs[2360]), .rectangle3_y(rectangle3_ys[2360]), .rectangle3_width(rectangle3_widths[2360]), .rectangle3_height(rectangle3_heights[2360]), .rectangle3_weight(rectangle3_weights[2360]), .feature_threshold(feature_thresholds[2360]), .feature_above(feature_aboves[2360]), .feature_below(feature_belows[2360]), .scan_win_std_dev(scan_win_std_dev[2360]), .feature_accum(feature_accums[2360]));
  accum_calculator ac2361(.scan_win(scan_win2361), .rectangle1_x(rectangle1_xs[2361]), .rectangle1_y(rectangle1_ys[2361]), .rectangle1_width(rectangle1_widths[2361]), .rectangle1_height(rectangle1_heights[2361]), .rectangle1_weight(rectangle1_weights[2361]), .rectangle2_x(rectangle2_xs[2361]), .rectangle2_y(rectangle2_ys[2361]), .rectangle2_width(rectangle2_widths[2361]), .rectangle2_height(rectangle2_heights[2361]), .rectangle2_weight(rectangle2_weights[2361]), .rectangle3_x(rectangle3_xs[2361]), .rectangle3_y(rectangle3_ys[2361]), .rectangle3_width(rectangle3_widths[2361]), .rectangle3_height(rectangle3_heights[2361]), .rectangle3_weight(rectangle3_weights[2361]), .feature_threshold(feature_thresholds[2361]), .feature_above(feature_aboves[2361]), .feature_below(feature_belows[2361]), .scan_win_std_dev(scan_win_std_dev[2361]), .feature_accum(feature_accums[2361]));
  accum_calculator ac2362(.scan_win(scan_win2362), .rectangle1_x(rectangle1_xs[2362]), .rectangle1_y(rectangle1_ys[2362]), .rectangle1_width(rectangle1_widths[2362]), .rectangle1_height(rectangle1_heights[2362]), .rectangle1_weight(rectangle1_weights[2362]), .rectangle2_x(rectangle2_xs[2362]), .rectangle2_y(rectangle2_ys[2362]), .rectangle2_width(rectangle2_widths[2362]), .rectangle2_height(rectangle2_heights[2362]), .rectangle2_weight(rectangle2_weights[2362]), .rectangle3_x(rectangle3_xs[2362]), .rectangle3_y(rectangle3_ys[2362]), .rectangle3_width(rectangle3_widths[2362]), .rectangle3_height(rectangle3_heights[2362]), .rectangle3_weight(rectangle3_weights[2362]), .feature_threshold(feature_thresholds[2362]), .feature_above(feature_aboves[2362]), .feature_below(feature_belows[2362]), .scan_win_std_dev(scan_win_std_dev[2362]), .feature_accum(feature_accums[2362]));
  accum_calculator ac2363(.scan_win(scan_win2363), .rectangle1_x(rectangle1_xs[2363]), .rectangle1_y(rectangle1_ys[2363]), .rectangle1_width(rectangle1_widths[2363]), .rectangle1_height(rectangle1_heights[2363]), .rectangle1_weight(rectangle1_weights[2363]), .rectangle2_x(rectangle2_xs[2363]), .rectangle2_y(rectangle2_ys[2363]), .rectangle2_width(rectangle2_widths[2363]), .rectangle2_height(rectangle2_heights[2363]), .rectangle2_weight(rectangle2_weights[2363]), .rectangle3_x(rectangle3_xs[2363]), .rectangle3_y(rectangle3_ys[2363]), .rectangle3_width(rectangle3_widths[2363]), .rectangle3_height(rectangle3_heights[2363]), .rectangle3_weight(rectangle3_weights[2363]), .feature_threshold(feature_thresholds[2363]), .feature_above(feature_aboves[2363]), .feature_below(feature_belows[2363]), .scan_win_std_dev(scan_win_std_dev[2363]), .feature_accum(feature_accums[2363]));
  accum_calculator ac2364(.scan_win(scan_win2364), .rectangle1_x(rectangle1_xs[2364]), .rectangle1_y(rectangle1_ys[2364]), .rectangle1_width(rectangle1_widths[2364]), .rectangle1_height(rectangle1_heights[2364]), .rectangle1_weight(rectangle1_weights[2364]), .rectangle2_x(rectangle2_xs[2364]), .rectangle2_y(rectangle2_ys[2364]), .rectangle2_width(rectangle2_widths[2364]), .rectangle2_height(rectangle2_heights[2364]), .rectangle2_weight(rectangle2_weights[2364]), .rectangle3_x(rectangle3_xs[2364]), .rectangle3_y(rectangle3_ys[2364]), .rectangle3_width(rectangle3_widths[2364]), .rectangle3_height(rectangle3_heights[2364]), .rectangle3_weight(rectangle3_weights[2364]), .feature_threshold(feature_thresholds[2364]), .feature_above(feature_aboves[2364]), .feature_below(feature_belows[2364]), .scan_win_std_dev(scan_win_std_dev[2364]), .feature_accum(feature_accums[2364]));
  accum_calculator ac2365(.scan_win(scan_win2365), .rectangle1_x(rectangle1_xs[2365]), .rectangle1_y(rectangle1_ys[2365]), .rectangle1_width(rectangle1_widths[2365]), .rectangle1_height(rectangle1_heights[2365]), .rectangle1_weight(rectangle1_weights[2365]), .rectangle2_x(rectangle2_xs[2365]), .rectangle2_y(rectangle2_ys[2365]), .rectangle2_width(rectangle2_widths[2365]), .rectangle2_height(rectangle2_heights[2365]), .rectangle2_weight(rectangle2_weights[2365]), .rectangle3_x(rectangle3_xs[2365]), .rectangle3_y(rectangle3_ys[2365]), .rectangle3_width(rectangle3_widths[2365]), .rectangle3_height(rectangle3_heights[2365]), .rectangle3_weight(rectangle3_weights[2365]), .feature_threshold(feature_thresholds[2365]), .feature_above(feature_aboves[2365]), .feature_below(feature_belows[2365]), .scan_win_std_dev(scan_win_std_dev[2365]), .feature_accum(feature_accums[2365]));
  accum_calculator ac2366(.scan_win(scan_win2366), .rectangle1_x(rectangle1_xs[2366]), .rectangle1_y(rectangle1_ys[2366]), .rectangle1_width(rectangle1_widths[2366]), .rectangle1_height(rectangle1_heights[2366]), .rectangle1_weight(rectangle1_weights[2366]), .rectangle2_x(rectangle2_xs[2366]), .rectangle2_y(rectangle2_ys[2366]), .rectangle2_width(rectangle2_widths[2366]), .rectangle2_height(rectangle2_heights[2366]), .rectangle2_weight(rectangle2_weights[2366]), .rectangle3_x(rectangle3_xs[2366]), .rectangle3_y(rectangle3_ys[2366]), .rectangle3_width(rectangle3_widths[2366]), .rectangle3_height(rectangle3_heights[2366]), .rectangle3_weight(rectangle3_weights[2366]), .feature_threshold(feature_thresholds[2366]), .feature_above(feature_aboves[2366]), .feature_below(feature_belows[2366]), .scan_win_std_dev(scan_win_std_dev[2366]), .feature_accum(feature_accums[2366]));
  accum_calculator ac2367(.scan_win(scan_win2367), .rectangle1_x(rectangle1_xs[2367]), .rectangle1_y(rectangle1_ys[2367]), .rectangle1_width(rectangle1_widths[2367]), .rectangle1_height(rectangle1_heights[2367]), .rectangle1_weight(rectangle1_weights[2367]), .rectangle2_x(rectangle2_xs[2367]), .rectangle2_y(rectangle2_ys[2367]), .rectangle2_width(rectangle2_widths[2367]), .rectangle2_height(rectangle2_heights[2367]), .rectangle2_weight(rectangle2_weights[2367]), .rectangle3_x(rectangle3_xs[2367]), .rectangle3_y(rectangle3_ys[2367]), .rectangle3_width(rectangle3_widths[2367]), .rectangle3_height(rectangle3_heights[2367]), .rectangle3_weight(rectangle3_weights[2367]), .feature_threshold(feature_thresholds[2367]), .feature_above(feature_aboves[2367]), .feature_below(feature_belows[2367]), .scan_win_std_dev(scan_win_std_dev[2367]), .feature_accum(feature_accums[2367]));
  accum_calculator ac2368(.scan_win(scan_win2368), .rectangle1_x(rectangle1_xs[2368]), .rectangle1_y(rectangle1_ys[2368]), .rectangle1_width(rectangle1_widths[2368]), .rectangle1_height(rectangle1_heights[2368]), .rectangle1_weight(rectangle1_weights[2368]), .rectangle2_x(rectangle2_xs[2368]), .rectangle2_y(rectangle2_ys[2368]), .rectangle2_width(rectangle2_widths[2368]), .rectangle2_height(rectangle2_heights[2368]), .rectangle2_weight(rectangle2_weights[2368]), .rectangle3_x(rectangle3_xs[2368]), .rectangle3_y(rectangle3_ys[2368]), .rectangle3_width(rectangle3_widths[2368]), .rectangle3_height(rectangle3_heights[2368]), .rectangle3_weight(rectangle3_weights[2368]), .feature_threshold(feature_thresholds[2368]), .feature_above(feature_aboves[2368]), .feature_below(feature_belows[2368]), .scan_win_std_dev(scan_win_std_dev[2368]), .feature_accum(feature_accums[2368]));
  accum_calculator ac2369(.scan_win(scan_win2369), .rectangle1_x(rectangle1_xs[2369]), .rectangle1_y(rectangle1_ys[2369]), .rectangle1_width(rectangle1_widths[2369]), .rectangle1_height(rectangle1_heights[2369]), .rectangle1_weight(rectangle1_weights[2369]), .rectangle2_x(rectangle2_xs[2369]), .rectangle2_y(rectangle2_ys[2369]), .rectangle2_width(rectangle2_widths[2369]), .rectangle2_height(rectangle2_heights[2369]), .rectangle2_weight(rectangle2_weights[2369]), .rectangle3_x(rectangle3_xs[2369]), .rectangle3_y(rectangle3_ys[2369]), .rectangle3_width(rectangle3_widths[2369]), .rectangle3_height(rectangle3_heights[2369]), .rectangle3_weight(rectangle3_weights[2369]), .feature_threshold(feature_thresholds[2369]), .feature_above(feature_aboves[2369]), .feature_below(feature_belows[2369]), .scan_win_std_dev(scan_win_std_dev[2369]), .feature_accum(feature_accums[2369]));
  accum_calculator ac2370(.scan_win(scan_win2370), .rectangle1_x(rectangle1_xs[2370]), .rectangle1_y(rectangle1_ys[2370]), .rectangle1_width(rectangle1_widths[2370]), .rectangle1_height(rectangle1_heights[2370]), .rectangle1_weight(rectangle1_weights[2370]), .rectangle2_x(rectangle2_xs[2370]), .rectangle2_y(rectangle2_ys[2370]), .rectangle2_width(rectangle2_widths[2370]), .rectangle2_height(rectangle2_heights[2370]), .rectangle2_weight(rectangle2_weights[2370]), .rectangle3_x(rectangle3_xs[2370]), .rectangle3_y(rectangle3_ys[2370]), .rectangle3_width(rectangle3_widths[2370]), .rectangle3_height(rectangle3_heights[2370]), .rectangle3_weight(rectangle3_weights[2370]), .feature_threshold(feature_thresholds[2370]), .feature_above(feature_aboves[2370]), .feature_below(feature_belows[2370]), .scan_win_std_dev(scan_win_std_dev[2370]), .feature_accum(feature_accums[2370]));
  accum_calculator ac2371(.scan_win(scan_win2371), .rectangle1_x(rectangle1_xs[2371]), .rectangle1_y(rectangle1_ys[2371]), .rectangle1_width(rectangle1_widths[2371]), .rectangle1_height(rectangle1_heights[2371]), .rectangle1_weight(rectangle1_weights[2371]), .rectangle2_x(rectangle2_xs[2371]), .rectangle2_y(rectangle2_ys[2371]), .rectangle2_width(rectangle2_widths[2371]), .rectangle2_height(rectangle2_heights[2371]), .rectangle2_weight(rectangle2_weights[2371]), .rectangle3_x(rectangle3_xs[2371]), .rectangle3_y(rectangle3_ys[2371]), .rectangle3_width(rectangle3_widths[2371]), .rectangle3_height(rectangle3_heights[2371]), .rectangle3_weight(rectangle3_weights[2371]), .feature_threshold(feature_thresholds[2371]), .feature_above(feature_aboves[2371]), .feature_below(feature_belows[2371]), .scan_win_std_dev(scan_win_std_dev[2371]), .feature_accum(feature_accums[2371]));
  accum_calculator ac2372(.scan_win(scan_win2372), .rectangle1_x(rectangle1_xs[2372]), .rectangle1_y(rectangle1_ys[2372]), .rectangle1_width(rectangle1_widths[2372]), .rectangle1_height(rectangle1_heights[2372]), .rectangle1_weight(rectangle1_weights[2372]), .rectangle2_x(rectangle2_xs[2372]), .rectangle2_y(rectangle2_ys[2372]), .rectangle2_width(rectangle2_widths[2372]), .rectangle2_height(rectangle2_heights[2372]), .rectangle2_weight(rectangle2_weights[2372]), .rectangle3_x(rectangle3_xs[2372]), .rectangle3_y(rectangle3_ys[2372]), .rectangle3_width(rectangle3_widths[2372]), .rectangle3_height(rectangle3_heights[2372]), .rectangle3_weight(rectangle3_weights[2372]), .feature_threshold(feature_thresholds[2372]), .feature_above(feature_aboves[2372]), .feature_below(feature_belows[2372]), .scan_win_std_dev(scan_win_std_dev[2372]), .feature_accum(feature_accums[2372]));
  accum_calculator ac2373(.scan_win(scan_win2373), .rectangle1_x(rectangle1_xs[2373]), .rectangle1_y(rectangle1_ys[2373]), .rectangle1_width(rectangle1_widths[2373]), .rectangle1_height(rectangle1_heights[2373]), .rectangle1_weight(rectangle1_weights[2373]), .rectangle2_x(rectangle2_xs[2373]), .rectangle2_y(rectangle2_ys[2373]), .rectangle2_width(rectangle2_widths[2373]), .rectangle2_height(rectangle2_heights[2373]), .rectangle2_weight(rectangle2_weights[2373]), .rectangle3_x(rectangle3_xs[2373]), .rectangle3_y(rectangle3_ys[2373]), .rectangle3_width(rectangle3_widths[2373]), .rectangle3_height(rectangle3_heights[2373]), .rectangle3_weight(rectangle3_weights[2373]), .feature_threshold(feature_thresholds[2373]), .feature_above(feature_aboves[2373]), .feature_below(feature_belows[2373]), .scan_win_std_dev(scan_win_std_dev[2373]), .feature_accum(feature_accums[2373]));
  accum_calculator ac2374(.scan_win(scan_win2374), .rectangle1_x(rectangle1_xs[2374]), .rectangle1_y(rectangle1_ys[2374]), .rectangle1_width(rectangle1_widths[2374]), .rectangle1_height(rectangle1_heights[2374]), .rectangle1_weight(rectangle1_weights[2374]), .rectangle2_x(rectangle2_xs[2374]), .rectangle2_y(rectangle2_ys[2374]), .rectangle2_width(rectangle2_widths[2374]), .rectangle2_height(rectangle2_heights[2374]), .rectangle2_weight(rectangle2_weights[2374]), .rectangle3_x(rectangle3_xs[2374]), .rectangle3_y(rectangle3_ys[2374]), .rectangle3_width(rectangle3_widths[2374]), .rectangle3_height(rectangle3_heights[2374]), .rectangle3_weight(rectangle3_weights[2374]), .feature_threshold(feature_thresholds[2374]), .feature_above(feature_aboves[2374]), .feature_below(feature_belows[2374]), .scan_win_std_dev(scan_win_std_dev[2374]), .feature_accum(feature_accums[2374]));
  accum_calculator ac2375(.scan_win(scan_win2375), .rectangle1_x(rectangle1_xs[2375]), .rectangle1_y(rectangle1_ys[2375]), .rectangle1_width(rectangle1_widths[2375]), .rectangle1_height(rectangle1_heights[2375]), .rectangle1_weight(rectangle1_weights[2375]), .rectangle2_x(rectangle2_xs[2375]), .rectangle2_y(rectangle2_ys[2375]), .rectangle2_width(rectangle2_widths[2375]), .rectangle2_height(rectangle2_heights[2375]), .rectangle2_weight(rectangle2_weights[2375]), .rectangle3_x(rectangle3_xs[2375]), .rectangle3_y(rectangle3_ys[2375]), .rectangle3_width(rectangle3_widths[2375]), .rectangle3_height(rectangle3_heights[2375]), .rectangle3_weight(rectangle3_weights[2375]), .feature_threshold(feature_thresholds[2375]), .feature_above(feature_aboves[2375]), .feature_below(feature_belows[2375]), .scan_win_std_dev(scan_win_std_dev[2375]), .feature_accum(feature_accums[2375]));
  accum_calculator ac2376(.scan_win(scan_win2376), .rectangle1_x(rectangle1_xs[2376]), .rectangle1_y(rectangle1_ys[2376]), .rectangle1_width(rectangle1_widths[2376]), .rectangle1_height(rectangle1_heights[2376]), .rectangle1_weight(rectangle1_weights[2376]), .rectangle2_x(rectangle2_xs[2376]), .rectangle2_y(rectangle2_ys[2376]), .rectangle2_width(rectangle2_widths[2376]), .rectangle2_height(rectangle2_heights[2376]), .rectangle2_weight(rectangle2_weights[2376]), .rectangle3_x(rectangle3_xs[2376]), .rectangle3_y(rectangle3_ys[2376]), .rectangle3_width(rectangle3_widths[2376]), .rectangle3_height(rectangle3_heights[2376]), .rectangle3_weight(rectangle3_weights[2376]), .feature_threshold(feature_thresholds[2376]), .feature_above(feature_aboves[2376]), .feature_below(feature_belows[2376]), .scan_win_std_dev(scan_win_std_dev[2376]), .feature_accum(feature_accums[2376]));
  accum_calculator ac2377(.scan_win(scan_win2377), .rectangle1_x(rectangle1_xs[2377]), .rectangle1_y(rectangle1_ys[2377]), .rectangle1_width(rectangle1_widths[2377]), .rectangle1_height(rectangle1_heights[2377]), .rectangle1_weight(rectangle1_weights[2377]), .rectangle2_x(rectangle2_xs[2377]), .rectangle2_y(rectangle2_ys[2377]), .rectangle2_width(rectangle2_widths[2377]), .rectangle2_height(rectangle2_heights[2377]), .rectangle2_weight(rectangle2_weights[2377]), .rectangle3_x(rectangle3_xs[2377]), .rectangle3_y(rectangle3_ys[2377]), .rectangle3_width(rectangle3_widths[2377]), .rectangle3_height(rectangle3_heights[2377]), .rectangle3_weight(rectangle3_weights[2377]), .feature_threshold(feature_thresholds[2377]), .feature_above(feature_aboves[2377]), .feature_below(feature_belows[2377]), .scan_win_std_dev(scan_win_std_dev[2377]), .feature_accum(feature_accums[2377]));
  accum_calculator ac2378(.scan_win(scan_win2378), .rectangle1_x(rectangle1_xs[2378]), .rectangle1_y(rectangle1_ys[2378]), .rectangle1_width(rectangle1_widths[2378]), .rectangle1_height(rectangle1_heights[2378]), .rectangle1_weight(rectangle1_weights[2378]), .rectangle2_x(rectangle2_xs[2378]), .rectangle2_y(rectangle2_ys[2378]), .rectangle2_width(rectangle2_widths[2378]), .rectangle2_height(rectangle2_heights[2378]), .rectangle2_weight(rectangle2_weights[2378]), .rectangle3_x(rectangle3_xs[2378]), .rectangle3_y(rectangle3_ys[2378]), .rectangle3_width(rectangle3_widths[2378]), .rectangle3_height(rectangle3_heights[2378]), .rectangle3_weight(rectangle3_weights[2378]), .feature_threshold(feature_thresholds[2378]), .feature_above(feature_aboves[2378]), .feature_below(feature_belows[2378]), .scan_win_std_dev(scan_win_std_dev[2378]), .feature_accum(feature_accums[2378]));
  accum_calculator ac2379(.scan_win(scan_win2379), .rectangle1_x(rectangle1_xs[2379]), .rectangle1_y(rectangle1_ys[2379]), .rectangle1_width(rectangle1_widths[2379]), .rectangle1_height(rectangle1_heights[2379]), .rectangle1_weight(rectangle1_weights[2379]), .rectangle2_x(rectangle2_xs[2379]), .rectangle2_y(rectangle2_ys[2379]), .rectangle2_width(rectangle2_widths[2379]), .rectangle2_height(rectangle2_heights[2379]), .rectangle2_weight(rectangle2_weights[2379]), .rectangle3_x(rectangle3_xs[2379]), .rectangle3_y(rectangle3_ys[2379]), .rectangle3_width(rectangle3_widths[2379]), .rectangle3_height(rectangle3_heights[2379]), .rectangle3_weight(rectangle3_weights[2379]), .feature_threshold(feature_thresholds[2379]), .feature_above(feature_aboves[2379]), .feature_below(feature_belows[2379]), .scan_win_std_dev(scan_win_std_dev[2379]), .feature_accum(feature_accums[2379]));
  accum_calculator ac2380(.scan_win(scan_win2380), .rectangle1_x(rectangle1_xs[2380]), .rectangle1_y(rectangle1_ys[2380]), .rectangle1_width(rectangle1_widths[2380]), .rectangle1_height(rectangle1_heights[2380]), .rectangle1_weight(rectangle1_weights[2380]), .rectangle2_x(rectangle2_xs[2380]), .rectangle2_y(rectangle2_ys[2380]), .rectangle2_width(rectangle2_widths[2380]), .rectangle2_height(rectangle2_heights[2380]), .rectangle2_weight(rectangle2_weights[2380]), .rectangle3_x(rectangle3_xs[2380]), .rectangle3_y(rectangle3_ys[2380]), .rectangle3_width(rectangle3_widths[2380]), .rectangle3_height(rectangle3_heights[2380]), .rectangle3_weight(rectangle3_weights[2380]), .feature_threshold(feature_thresholds[2380]), .feature_above(feature_aboves[2380]), .feature_below(feature_belows[2380]), .scan_win_std_dev(scan_win_std_dev[2380]), .feature_accum(feature_accums[2380]));
  accum_calculator ac2381(.scan_win(scan_win2381), .rectangle1_x(rectangle1_xs[2381]), .rectangle1_y(rectangle1_ys[2381]), .rectangle1_width(rectangle1_widths[2381]), .rectangle1_height(rectangle1_heights[2381]), .rectangle1_weight(rectangle1_weights[2381]), .rectangle2_x(rectangle2_xs[2381]), .rectangle2_y(rectangle2_ys[2381]), .rectangle2_width(rectangle2_widths[2381]), .rectangle2_height(rectangle2_heights[2381]), .rectangle2_weight(rectangle2_weights[2381]), .rectangle3_x(rectangle3_xs[2381]), .rectangle3_y(rectangle3_ys[2381]), .rectangle3_width(rectangle3_widths[2381]), .rectangle3_height(rectangle3_heights[2381]), .rectangle3_weight(rectangle3_weights[2381]), .feature_threshold(feature_thresholds[2381]), .feature_above(feature_aboves[2381]), .feature_below(feature_belows[2381]), .scan_win_std_dev(scan_win_std_dev[2381]), .feature_accum(feature_accums[2381]));
  accum_calculator ac2382(.scan_win(scan_win2382), .rectangle1_x(rectangle1_xs[2382]), .rectangle1_y(rectangle1_ys[2382]), .rectangle1_width(rectangle1_widths[2382]), .rectangle1_height(rectangle1_heights[2382]), .rectangle1_weight(rectangle1_weights[2382]), .rectangle2_x(rectangle2_xs[2382]), .rectangle2_y(rectangle2_ys[2382]), .rectangle2_width(rectangle2_widths[2382]), .rectangle2_height(rectangle2_heights[2382]), .rectangle2_weight(rectangle2_weights[2382]), .rectangle3_x(rectangle3_xs[2382]), .rectangle3_y(rectangle3_ys[2382]), .rectangle3_width(rectangle3_widths[2382]), .rectangle3_height(rectangle3_heights[2382]), .rectangle3_weight(rectangle3_weights[2382]), .feature_threshold(feature_thresholds[2382]), .feature_above(feature_aboves[2382]), .feature_below(feature_belows[2382]), .scan_win_std_dev(scan_win_std_dev[2382]), .feature_accum(feature_accums[2382]));
  accum_calculator ac2383(.scan_win(scan_win2383), .rectangle1_x(rectangle1_xs[2383]), .rectangle1_y(rectangle1_ys[2383]), .rectangle1_width(rectangle1_widths[2383]), .rectangle1_height(rectangle1_heights[2383]), .rectangle1_weight(rectangle1_weights[2383]), .rectangle2_x(rectangle2_xs[2383]), .rectangle2_y(rectangle2_ys[2383]), .rectangle2_width(rectangle2_widths[2383]), .rectangle2_height(rectangle2_heights[2383]), .rectangle2_weight(rectangle2_weights[2383]), .rectangle3_x(rectangle3_xs[2383]), .rectangle3_y(rectangle3_ys[2383]), .rectangle3_width(rectangle3_widths[2383]), .rectangle3_height(rectangle3_heights[2383]), .rectangle3_weight(rectangle3_weights[2383]), .feature_threshold(feature_thresholds[2383]), .feature_above(feature_aboves[2383]), .feature_below(feature_belows[2383]), .scan_win_std_dev(scan_win_std_dev[2383]), .feature_accum(feature_accums[2383]));
  accum_calculator ac2384(.scan_win(scan_win2384), .rectangle1_x(rectangle1_xs[2384]), .rectangle1_y(rectangle1_ys[2384]), .rectangle1_width(rectangle1_widths[2384]), .rectangle1_height(rectangle1_heights[2384]), .rectangle1_weight(rectangle1_weights[2384]), .rectangle2_x(rectangle2_xs[2384]), .rectangle2_y(rectangle2_ys[2384]), .rectangle2_width(rectangle2_widths[2384]), .rectangle2_height(rectangle2_heights[2384]), .rectangle2_weight(rectangle2_weights[2384]), .rectangle3_x(rectangle3_xs[2384]), .rectangle3_y(rectangle3_ys[2384]), .rectangle3_width(rectangle3_widths[2384]), .rectangle3_height(rectangle3_heights[2384]), .rectangle3_weight(rectangle3_weights[2384]), .feature_threshold(feature_thresholds[2384]), .feature_above(feature_aboves[2384]), .feature_below(feature_belows[2384]), .scan_win_std_dev(scan_win_std_dev[2384]), .feature_accum(feature_accums[2384]));
  accum_calculator ac2385(.scan_win(scan_win2385), .rectangle1_x(rectangle1_xs[2385]), .rectangle1_y(rectangle1_ys[2385]), .rectangle1_width(rectangle1_widths[2385]), .rectangle1_height(rectangle1_heights[2385]), .rectangle1_weight(rectangle1_weights[2385]), .rectangle2_x(rectangle2_xs[2385]), .rectangle2_y(rectangle2_ys[2385]), .rectangle2_width(rectangle2_widths[2385]), .rectangle2_height(rectangle2_heights[2385]), .rectangle2_weight(rectangle2_weights[2385]), .rectangle3_x(rectangle3_xs[2385]), .rectangle3_y(rectangle3_ys[2385]), .rectangle3_width(rectangle3_widths[2385]), .rectangle3_height(rectangle3_heights[2385]), .rectangle3_weight(rectangle3_weights[2385]), .feature_threshold(feature_thresholds[2385]), .feature_above(feature_aboves[2385]), .feature_below(feature_belows[2385]), .scan_win_std_dev(scan_win_std_dev[2385]), .feature_accum(feature_accums[2385]));
  accum_calculator ac2386(.scan_win(scan_win2386), .rectangle1_x(rectangle1_xs[2386]), .rectangle1_y(rectangle1_ys[2386]), .rectangle1_width(rectangle1_widths[2386]), .rectangle1_height(rectangle1_heights[2386]), .rectangle1_weight(rectangle1_weights[2386]), .rectangle2_x(rectangle2_xs[2386]), .rectangle2_y(rectangle2_ys[2386]), .rectangle2_width(rectangle2_widths[2386]), .rectangle2_height(rectangle2_heights[2386]), .rectangle2_weight(rectangle2_weights[2386]), .rectangle3_x(rectangle3_xs[2386]), .rectangle3_y(rectangle3_ys[2386]), .rectangle3_width(rectangle3_widths[2386]), .rectangle3_height(rectangle3_heights[2386]), .rectangle3_weight(rectangle3_weights[2386]), .feature_threshold(feature_thresholds[2386]), .feature_above(feature_aboves[2386]), .feature_below(feature_belows[2386]), .scan_win_std_dev(scan_win_std_dev[2386]), .feature_accum(feature_accums[2386]));
  accum_calculator ac2387(.scan_win(scan_win2387), .rectangle1_x(rectangle1_xs[2387]), .rectangle1_y(rectangle1_ys[2387]), .rectangle1_width(rectangle1_widths[2387]), .rectangle1_height(rectangle1_heights[2387]), .rectangle1_weight(rectangle1_weights[2387]), .rectangle2_x(rectangle2_xs[2387]), .rectangle2_y(rectangle2_ys[2387]), .rectangle2_width(rectangle2_widths[2387]), .rectangle2_height(rectangle2_heights[2387]), .rectangle2_weight(rectangle2_weights[2387]), .rectangle3_x(rectangle3_xs[2387]), .rectangle3_y(rectangle3_ys[2387]), .rectangle3_width(rectangle3_widths[2387]), .rectangle3_height(rectangle3_heights[2387]), .rectangle3_weight(rectangle3_weights[2387]), .feature_threshold(feature_thresholds[2387]), .feature_above(feature_aboves[2387]), .feature_below(feature_belows[2387]), .scan_win_std_dev(scan_win_std_dev[2387]), .feature_accum(feature_accums[2387]));
  accum_calculator ac2388(.scan_win(scan_win2388), .rectangle1_x(rectangle1_xs[2388]), .rectangle1_y(rectangle1_ys[2388]), .rectangle1_width(rectangle1_widths[2388]), .rectangle1_height(rectangle1_heights[2388]), .rectangle1_weight(rectangle1_weights[2388]), .rectangle2_x(rectangle2_xs[2388]), .rectangle2_y(rectangle2_ys[2388]), .rectangle2_width(rectangle2_widths[2388]), .rectangle2_height(rectangle2_heights[2388]), .rectangle2_weight(rectangle2_weights[2388]), .rectangle3_x(rectangle3_xs[2388]), .rectangle3_y(rectangle3_ys[2388]), .rectangle3_width(rectangle3_widths[2388]), .rectangle3_height(rectangle3_heights[2388]), .rectangle3_weight(rectangle3_weights[2388]), .feature_threshold(feature_thresholds[2388]), .feature_above(feature_aboves[2388]), .feature_below(feature_belows[2388]), .scan_win_std_dev(scan_win_std_dev[2388]), .feature_accum(feature_accums[2388]));
  accum_calculator ac2389(.scan_win(scan_win2389), .rectangle1_x(rectangle1_xs[2389]), .rectangle1_y(rectangle1_ys[2389]), .rectangle1_width(rectangle1_widths[2389]), .rectangle1_height(rectangle1_heights[2389]), .rectangle1_weight(rectangle1_weights[2389]), .rectangle2_x(rectangle2_xs[2389]), .rectangle2_y(rectangle2_ys[2389]), .rectangle2_width(rectangle2_widths[2389]), .rectangle2_height(rectangle2_heights[2389]), .rectangle2_weight(rectangle2_weights[2389]), .rectangle3_x(rectangle3_xs[2389]), .rectangle3_y(rectangle3_ys[2389]), .rectangle3_width(rectangle3_widths[2389]), .rectangle3_height(rectangle3_heights[2389]), .rectangle3_weight(rectangle3_weights[2389]), .feature_threshold(feature_thresholds[2389]), .feature_above(feature_aboves[2389]), .feature_below(feature_belows[2389]), .scan_win_std_dev(scan_win_std_dev[2389]), .feature_accum(feature_accums[2389]));
  accum_calculator ac2390(.scan_win(scan_win2390), .rectangle1_x(rectangle1_xs[2390]), .rectangle1_y(rectangle1_ys[2390]), .rectangle1_width(rectangle1_widths[2390]), .rectangle1_height(rectangle1_heights[2390]), .rectangle1_weight(rectangle1_weights[2390]), .rectangle2_x(rectangle2_xs[2390]), .rectangle2_y(rectangle2_ys[2390]), .rectangle2_width(rectangle2_widths[2390]), .rectangle2_height(rectangle2_heights[2390]), .rectangle2_weight(rectangle2_weights[2390]), .rectangle3_x(rectangle3_xs[2390]), .rectangle3_y(rectangle3_ys[2390]), .rectangle3_width(rectangle3_widths[2390]), .rectangle3_height(rectangle3_heights[2390]), .rectangle3_weight(rectangle3_weights[2390]), .feature_threshold(feature_thresholds[2390]), .feature_above(feature_aboves[2390]), .feature_below(feature_belows[2390]), .scan_win_std_dev(scan_win_std_dev[2390]), .feature_accum(feature_accums[2390]));
  accum_calculator ac2391(.scan_win(scan_win2391), .rectangle1_x(rectangle1_xs[2391]), .rectangle1_y(rectangle1_ys[2391]), .rectangle1_width(rectangle1_widths[2391]), .rectangle1_height(rectangle1_heights[2391]), .rectangle1_weight(rectangle1_weights[2391]), .rectangle2_x(rectangle2_xs[2391]), .rectangle2_y(rectangle2_ys[2391]), .rectangle2_width(rectangle2_widths[2391]), .rectangle2_height(rectangle2_heights[2391]), .rectangle2_weight(rectangle2_weights[2391]), .rectangle3_x(rectangle3_xs[2391]), .rectangle3_y(rectangle3_ys[2391]), .rectangle3_width(rectangle3_widths[2391]), .rectangle3_height(rectangle3_heights[2391]), .rectangle3_weight(rectangle3_weights[2391]), .feature_threshold(feature_thresholds[2391]), .feature_above(feature_aboves[2391]), .feature_below(feature_belows[2391]), .scan_win_std_dev(scan_win_std_dev[2391]), .feature_accum(feature_accums[2391]));
  accum_calculator ac2392(.scan_win(scan_win2392), .rectangle1_x(rectangle1_xs[2392]), .rectangle1_y(rectangle1_ys[2392]), .rectangle1_width(rectangle1_widths[2392]), .rectangle1_height(rectangle1_heights[2392]), .rectangle1_weight(rectangle1_weights[2392]), .rectangle2_x(rectangle2_xs[2392]), .rectangle2_y(rectangle2_ys[2392]), .rectangle2_width(rectangle2_widths[2392]), .rectangle2_height(rectangle2_heights[2392]), .rectangle2_weight(rectangle2_weights[2392]), .rectangle3_x(rectangle3_xs[2392]), .rectangle3_y(rectangle3_ys[2392]), .rectangle3_width(rectangle3_widths[2392]), .rectangle3_height(rectangle3_heights[2392]), .rectangle3_weight(rectangle3_weights[2392]), .feature_threshold(feature_thresholds[2392]), .feature_above(feature_aboves[2392]), .feature_below(feature_belows[2392]), .scan_win_std_dev(scan_win_std_dev[2392]), .feature_accum(feature_accums[2392]));
  accum_calculator ac2393(.scan_win(scan_win2393), .rectangle1_x(rectangle1_xs[2393]), .rectangle1_y(rectangle1_ys[2393]), .rectangle1_width(rectangle1_widths[2393]), .rectangle1_height(rectangle1_heights[2393]), .rectangle1_weight(rectangle1_weights[2393]), .rectangle2_x(rectangle2_xs[2393]), .rectangle2_y(rectangle2_ys[2393]), .rectangle2_width(rectangle2_widths[2393]), .rectangle2_height(rectangle2_heights[2393]), .rectangle2_weight(rectangle2_weights[2393]), .rectangle3_x(rectangle3_xs[2393]), .rectangle3_y(rectangle3_ys[2393]), .rectangle3_width(rectangle3_widths[2393]), .rectangle3_height(rectangle3_heights[2393]), .rectangle3_weight(rectangle3_weights[2393]), .feature_threshold(feature_thresholds[2393]), .feature_above(feature_aboves[2393]), .feature_below(feature_belows[2393]), .scan_win_std_dev(scan_win_std_dev[2393]), .feature_accum(feature_accums[2393]));
  accum_calculator ac2394(.scan_win(scan_win2394), .rectangle1_x(rectangle1_xs[2394]), .rectangle1_y(rectangle1_ys[2394]), .rectangle1_width(rectangle1_widths[2394]), .rectangle1_height(rectangle1_heights[2394]), .rectangle1_weight(rectangle1_weights[2394]), .rectangle2_x(rectangle2_xs[2394]), .rectangle2_y(rectangle2_ys[2394]), .rectangle2_width(rectangle2_widths[2394]), .rectangle2_height(rectangle2_heights[2394]), .rectangle2_weight(rectangle2_weights[2394]), .rectangle3_x(rectangle3_xs[2394]), .rectangle3_y(rectangle3_ys[2394]), .rectangle3_width(rectangle3_widths[2394]), .rectangle3_height(rectangle3_heights[2394]), .rectangle3_weight(rectangle3_weights[2394]), .feature_threshold(feature_thresholds[2394]), .feature_above(feature_aboves[2394]), .feature_below(feature_belows[2394]), .scan_win_std_dev(scan_win_std_dev[2394]), .feature_accum(feature_accums[2394]));
  accum_calculator ac2395(.scan_win(scan_win2395), .rectangle1_x(rectangle1_xs[2395]), .rectangle1_y(rectangle1_ys[2395]), .rectangle1_width(rectangle1_widths[2395]), .rectangle1_height(rectangle1_heights[2395]), .rectangle1_weight(rectangle1_weights[2395]), .rectangle2_x(rectangle2_xs[2395]), .rectangle2_y(rectangle2_ys[2395]), .rectangle2_width(rectangle2_widths[2395]), .rectangle2_height(rectangle2_heights[2395]), .rectangle2_weight(rectangle2_weights[2395]), .rectangle3_x(rectangle3_xs[2395]), .rectangle3_y(rectangle3_ys[2395]), .rectangle3_width(rectangle3_widths[2395]), .rectangle3_height(rectangle3_heights[2395]), .rectangle3_weight(rectangle3_weights[2395]), .feature_threshold(feature_thresholds[2395]), .feature_above(feature_aboves[2395]), .feature_below(feature_belows[2395]), .scan_win_std_dev(scan_win_std_dev[2395]), .feature_accum(feature_accums[2395]));
  accum_calculator ac2396(.scan_win(scan_win2396), .rectangle1_x(rectangle1_xs[2396]), .rectangle1_y(rectangle1_ys[2396]), .rectangle1_width(rectangle1_widths[2396]), .rectangle1_height(rectangle1_heights[2396]), .rectangle1_weight(rectangle1_weights[2396]), .rectangle2_x(rectangle2_xs[2396]), .rectangle2_y(rectangle2_ys[2396]), .rectangle2_width(rectangle2_widths[2396]), .rectangle2_height(rectangle2_heights[2396]), .rectangle2_weight(rectangle2_weights[2396]), .rectangle3_x(rectangle3_xs[2396]), .rectangle3_y(rectangle3_ys[2396]), .rectangle3_width(rectangle3_widths[2396]), .rectangle3_height(rectangle3_heights[2396]), .rectangle3_weight(rectangle3_weights[2396]), .feature_threshold(feature_thresholds[2396]), .feature_above(feature_aboves[2396]), .feature_below(feature_belows[2396]), .scan_win_std_dev(scan_win_std_dev[2396]), .feature_accum(feature_accums[2396]));
  accum_calculator ac2397(.scan_win(scan_win2397), .rectangle1_x(rectangle1_xs[2397]), .rectangle1_y(rectangle1_ys[2397]), .rectangle1_width(rectangle1_widths[2397]), .rectangle1_height(rectangle1_heights[2397]), .rectangle1_weight(rectangle1_weights[2397]), .rectangle2_x(rectangle2_xs[2397]), .rectangle2_y(rectangle2_ys[2397]), .rectangle2_width(rectangle2_widths[2397]), .rectangle2_height(rectangle2_heights[2397]), .rectangle2_weight(rectangle2_weights[2397]), .rectangle3_x(rectangle3_xs[2397]), .rectangle3_y(rectangle3_ys[2397]), .rectangle3_width(rectangle3_widths[2397]), .rectangle3_height(rectangle3_heights[2397]), .rectangle3_weight(rectangle3_weights[2397]), .feature_threshold(feature_thresholds[2397]), .feature_above(feature_aboves[2397]), .feature_below(feature_belows[2397]), .scan_win_std_dev(scan_win_std_dev[2397]), .feature_accum(feature_accums[2397]));
  accum_calculator ac2398(.scan_win(scan_win2398), .rectangle1_x(rectangle1_xs[2398]), .rectangle1_y(rectangle1_ys[2398]), .rectangle1_width(rectangle1_widths[2398]), .rectangle1_height(rectangle1_heights[2398]), .rectangle1_weight(rectangle1_weights[2398]), .rectangle2_x(rectangle2_xs[2398]), .rectangle2_y(rectangle2_ys[2398]), .rectangle2_width(rectangle2_widths[2398]), .rectangle2_height(rectangle2_heights[2398]), .rectangle2_weight(rectangle2_weights[2398]), .rectangle3_x(rectangle3_xs[2398]), .rectangle3_y(rectangle3_ys[2398]), .rectangle3_width(rectangle3_widths[2398]), .rectangle3_height(rectangle3_heights[2398]), .rectangle3_weight(rectangle3_weights[2398]), .feature_threshold(feature_thresholds[2398]), .feature_above(feature_aboves[2398]), .feature_below(feature_belows[2398]), .scan_win_std_dev(scan_win_std_dev[2398]), .feature_accum(feature_accums[2398]));
  accum_calculator ac2399(.scan_win(scan_win2399), .rectangle1_x(rectangle1_xs[2399]), .rectangle1_y(rectangle1_ys[2399]), .rectangle1_width(rectangle1_widths[2399]), .rectangle1_height(rectangle1_heights[2399]), .rectangle1_weight(rectangle1_weights[2399]), .rectangle2_x(rectangle2_xs[2399]), .rectangle2_y(rectangle2_ys[2399]), .rectangle2_width(rectangle2_widths[2399]), .rectangle2_height(rectangle2_heights[2399]), .rectangle2_weight(rectangle2_weights[2399]), .rectangle3_x(rectangle3_xs[2399]), .rectangle3_y(rectangle3_ys[2399]), .rectangle3_width(rectangle3_widths[2399]), .rectangle3_height(rectangle3_heights[2399]), .rectangle3_weight(rectangle3_weights[2399]), .feature_threshold(feature_thresholds[2399]), .feature_above(feature_aboves[2399]), .feature_below(feature_belows[2399]), .scan_win_std_dev(scan_win_std_dev[2399]), .feature_accum(feature_accums[2399]));
  accum_calculator ac2400(.scan_win(scan_win2400), .rectangle1_x(rectangle1_xs[2400]), .rectangle1_y(rectangle1_ys[2400]), .rectangle1_width(rectangle1_widths[2400]), .rectangle1_height(rectangle1_heights[2400]), .rectangle1_weight(rectangle1_weights[2400]), .rectangle2_x(rectangle2_xs[2400]), .rectangle2_y(rectangle2_ys[2400]), .rectangle2_width(rectangle2_widths[2400]), .rectangle2_height(rectangle2_heights[2400]), .rectangle2_weight(rectangle2_weights[2400]), .rectangle3_x(rectangle3_xs[2400]), .rectangle3_y(rectangle3_ys[2400]), .rectangle3_width(rectangle3_widths[2400]), .rectangle3_height(rectangle3_heights[2400]), .rectangle3_weight(rectangle3_weights[2400]), .feature_threshold(feature_thresholds[2400]), .feature_above(feature_aboves[2400]), .feature_below(feature_belows[2400]), .scan_win_std_dev(scan_win_std_dev[2400]), .feature_accum(feature_accums[2400]));
  accum_calculator ac2401(.scan_win(scan_win2401), .rectangle1_x(rectangle1_xs[2401]), .rectangle1_y(rectangle1_ys[2401]), .rectangle1_width(rectangle1_widths[2401]), .rectangle1_height(rectangle1_heights[2401]), .rectangle1_weight(rectangle1_weights[2401]), .rectangle2_x(rectangle2_xs[2401]), .rectangle2_y(rectangle2_ys[2401]), .rectangle2_width(rectangle2_widths[2401]), .rectangle2_height(rectangle2_heights[2401]), .rectangle2_weight(rectangle2_weights[2401]), .rectangle3_x(rectangle3_xs[2401]), .rectangle3_y(rectangle3_ys[2401]), .rectangle3_width(rectangle3_widths[2401]), .rectangle3_height(rectangle3_heights[2401]), .rectangle3_weight(rectangle3_weights[2401]), .feature_threshold(feature_thresholds[2401]), .feature_above(feature_aboves[2401]), .feature_below(feature_belows[2401]), .scan_win_std_dev(scan_win_std_dev[2401]), .feature_accum(feature_accums[2401]));
  accum_calculator ac2402(.scan_win(scan_win2402), .rectangle1_x(rectangle1_xs[2402]), .rectangle1_y(rectangle1_ys[2402]), .rectangle1_width(rectangle1_widths[2402]), .rectangle1_height(rectangle1_heights[2402]), .rectangle1_weight(rectangle1_weights[2402]), .rectangle2_x(rectangle2_xs[2402]), .rectangle2_y(rectangle2_ys[2402]), .rectangle2_width(rectangle2_widths[2402]), .rectangle2_height(rectangle2_heights[2402]), .rectangle2_weight(rectangle2_weights[2402]), .rectangle3_x(rectangle3_xs[2402]), .rectangle3_y(rectangle3_ys[2402]), .rectangle3_width(rectangle3_widths[2402]), .rectangle3_height(rectangle3_heights[2402]), .rectangle3_weight(rectangle3_weights[2402]), .feature_threshold(feature_thresholds[2402]), .feature_above(feature_aboves[2402]), .feature_below(feature_belows[2402]), .scan_win_std_dev(scan_win_std_dev[2402]), .feature_accum(feature_accums[2402]));
  accum_calculator ac2403(.scan_win(scan_win2403), .rectangle1_x(rectangle1_xs[2403]), .rectangle1_y(rectangle1_ys[2403]), .rectangle1_width(rectangle1_widths[2403]), .rectangle1_height(rectangle1_heights[2403]), .rectangle1_weight(rectangle1_weights[2403]), .rectangle2_x(rectangle2_xs[2403]), .rectangle2_y(rectangle2_ys[2403]), .rectangle2_width(rectangle2_widths[2403]), .rectangle2_height(rectangle2_heights[2403]), .rectangle2_weight(rectangle2_weights[2403]), .rectangle3_x(rectangle3_xs[2403]), .rectangle3_y(rectangle3_ys[2403]), .rectangle3_width(rectangle3_widths[2403]), .rectangle3_height(rectangle3_heights[2403]), .rectangle3_weight(rectangle3_weights[2403]), .feature_threshold(feature_thresholds[2403]), .feature_above(feature_aboves[2403]), .feature_below(feature_belows[2403]), .scan_win_std_dev(scan_win_std_dev[2403]), .feature_accum(feature_accums[2403]));
  accum_calculator ac2404(.scan_win(scan_win2404), .rectangle1_x(rectangle1_xs[2404]), .rectangle1_y(rectangle1_ys[2404]), .rectangle1_width(rectangle1_widths[2404]), .rectangle1_height(rectangle1_heights[2404]), .rectangle1_weight(rectangle1_weights[2404]), .rectangle2_x(rectangle2_xs[2404]), .rectangle2_y(rectangle2_ys[2404]), .rectangle2_width(rectangle2_widths[2404]), .rectangle2_height(rectangle2_heights[2404]), .rectangle2_weight(rectangle2_weights[2404]), .rectangle3_x(rectangle3_xs[2404]), .rectangle3_y(rectangle3_ys[2404]), .rectangle3_width(rectangle3_widths[2404]), .rectangle3_height(rectangle3_heights[2404]), .rectangle3_weight(rectangle3_weights[2404]), .feature_threshold(feature_thresholds[2404]), .feature_above(feature_aboves[2404]), .feature_below(feature_belows[2404]), .scan_win_std_dev(scan_win_std_dev[2404]), .feature_accum(feature_accums[2404]));
  accum_calculator ac2405(.scan_win(scan_win2405), .rectangle1_x(rectangle1_xs[2405]), .rectangle1_y(rectangle1_ys[2405]), .rectangle1_width(rectangle1_widths[2405]), .rectangle1_height(rectangle1_heights[2405]), .rectangle1_weight(rectangle1_weights[2405]), .rectangle2_x(rectangle2_xs[2405]), .rectangle2_y(rectangle2_ys[2405]), .rectangle2_width(rectangle2_widths[2405]), .rectangle2_height(rectangle2_heights[2405]), .rectangle2_weight(rectangle2_weights[2405]), .rectangle3_x(rectangle3_xs[2405]), .rectangle3_y(rectangle3_ys[2405]), .rectangle3_width(rectangle3_widths[2405]), .rectangle3_height(rectangle3_heights[2405]), .rectangle3_weight(rectangle3_weights[2405]), .feature_threshold(feature_thresholds[2405]), .feature_above(feature_aboves[2405]), .feature_below(feature_belows[2405]), .scan_win_std_dev(scan_win_std_dev[2405]), .feature_accum(feature_accums[2405]));
  accum_calculator ac2406(.scan_win(scan_win2406), .rectangle1_x(rectangle1_xs[2406]), .rectangle1_y(rectangle1_ys[2406]), .rectangle1_width(rectangle1_widths[2406]), .rectangle1_height(rectangle1_heights[2406]), .rectangle1_weight(rectangle1_weights[2406]), .rectangle2_x(rectangle2_xs[2406]), .rectangle2_y(rectangle2_ys[2406]), .rectangle2_width(rectangle2_widths[2406]), .rectangle2_height(rectangle2_heights[2406]), .rectangle2_weight(rectangle2_weights[2406]), .rectangle3_x(rectangle3_xs[2406]), .rectangle3_y(rectangle3_ys[2406]), .rectangle3_width(rectangle3_widths[2406]), .rectangle3_height(rectangle3_heights[2406]), .rectangle3_weight(rectangle3_weights[2406]), .feature_threshold(feature_thresholds[2406]), .feature_above(feature_aboves[2406]), .feature_below(feature_belows[2406]), .scan_win_std_dev(scan_win_std_dev[2406]), .feature_accum(feature_accums[2406]));
  accum_calculator ac2407(.scan_win(scan_win2407), .rectangle1_x(rectangle1_xs[2407]), .rectangle1_y(rectangle1_ys[2407]), .rectangle1_width(rectangle1_widths[2407]), .rectangle1_height(rectangle1_heights[2407]), .rectangle1_weight(rectangle1_weights[2407]), .rectangle2_x(rectangle2_xs[2407]), .rectangle2_y(rectangle2_ys[2407]), .rectangle2_width(rectangle2_widths[2407]), .rectangle2_height(rectangle2_heights[2407]), .rectangle2_weight(rectangle2_weights[2407]), .rectangle3_x(rectangle3_xs[2407]), .rectangle3_y(rectangle3_ys[2407]), .rectangle3_width(rectangle3_widths[2407]), .rectangle3_height(rectangle3_heights[2407]), .rectangle3_weight(rectangle3_weights[2407]), .feature_threshold(feature_thresholds[2407]), .feature_above(feature_aboves[2407]), .feature_below(feature_belows[2407]), .scan_win_std_dev(scan_win_std_dev[2407]), .feature_accum(feature_accums[2407]));
  accum_calculator ac2408(.scan_win(scan_win2408), .rectangle1_x(rectangle1_xs[2408]), .rectangle1_y(rectangle1_ys[2408]), .rectangle1_width(rectangle1_widths[2408]), .rectangle1_height(rectangle1_heights[2408]), .rectangle1_weight(rectangle1_weights[2408]), .rectangle2_x(rectangle2_xs[2408]), .rectangle2_y(rectangle2_ys[2408]), .rectangle2_width(rectangle2_widths[2408]), .rectangle2_height(rectangle2_heights[2408]), .rectangle2_weight(rectangle2_weights[2408]), .rectangle3_x(rectangle3_xs[2408]), .rectangle3_y(rectangle3_ys[2408]), .rectangle3_width(rectangle3_widths[2408]), .rectangle3_height(rectangle3_heights[2408]), .rectangle3_weight(rectangle3_weights[2408]), .feature_threshold(feature_thresholds[2408]), .feature_above(feature_aboves[2408]), .feature_below(feature_belows[2408]), .scan_win_std_dev(scan_win_std_dev[2408]), .feature_accum(feature_accums[2408]));
  accum_calculator ac2409(.scan_win(scan_win2409), .rectangle1_x(rectangle1_xs[2409]), .rectangle1_y(rectangle1_ys[2409]), .rectangle1_width(rectangle1_widths[2409]), .rectangle1_height(rectangle1_heights[2409]), .rectangle1_weight(rectangle1_weights[2409]), .rectangle2_x(rectangle2_xs[2409]), .rectangle2_y(rectangle2_ys[2409]), .rectangle2_width(rectangle2_widths[2409]), .rectangle2_height(rectangle2_heights[2409]), .rectangle2_weight(rectangle2_weights[2409]), .rectangle3_x(rectangle3_xs[2409]), .rectangle3_y(rectangle3_ys[2409]), .rectangle3_width(rectangle3_widths[2409]), .rectangle3_height(rectangle3_heights[2409]), .rectangle3_weight(rectangle3_weights[2409]), .feature_threshold(feature_thresholds[2409]), .feature_above(feature_aboves[2409]), .feature_below(feature_belows[2409]), .scan_win_std_dev(scan_win_std_dev[2409]), .feature_accum(feature_accums[2409]));
  accum_calculator ac2410(.scan_win(scan_win2410), .rectangle1_x(rectangle1_xs[2410]), .rectangle1_y(rectangle1_ys[2410]), .rectangle1_width(rectangle1_widths[2410]), .rectangle1_height(rectangle1_heights[2410]), .rectangle1_weight(rectangle1_weights[2410]), .rectangle2_x(rectangle2_xs[2410]), .rectangle2_y(rectangle2_ys[2410]), .rectangle2_width(rectangle2_widths[2410]), .rectangle2_height(rectangle2_heights[2410]), .rectangle2_weight(rectangle2_weights[2410]), .rectangle3_x(rectangle3_xs[2410]), .rectangle3_y(rectangle3_ys[2410]), .rectangle3_width(rectangle3_widths[2410]), .rectangle3_height(rectangle3_heights[2410]), .rectangle3_weight(rectangle3_weights[2410]), .feature_threshold(feature_thresholds[2410]), .feature_above(feature_aboves[2410]), .feature_below(feature_belows[2410]), .scan_win_std_dev(scan_win_std_dev[2410]), .feature_accum(feature_accums[2410]));
  accum_calculator ac2411(.scan_win(scan_win2411), .rectangle1_x(rectangle1_xs[2411]), .rectangle1_y(rectangle1_ys[2411]), .rectangle1_width(rectangle1_widths[2411]), .rectangle1_height(rectangle1_heights[2411]), .rectangle1_weight(rectangle1_weights[2411]), .rectangle2_x(rectangle2_xs[2411]), .rectangle2_y(rectangle2_ys[2411]), .rectangle2_width(rectangle2_widths[2411]), .rectangle2_height(rectangle2_heights[2411]), .rectangle2_weight(rectangle2_weights[2411]), .rectangle3_x(rectangle3_xs[2411]), .rectangle3_y(rectangle3_ys[2411]), .rectangle3_width(rectangle3_widths[2411]), .rectangle3_height(rectangle3_heights[2411]), .rectangle3_weight(rectangle3_weights[2411]), .feature_threshold(feature_thresholds[2411]), .feature_above(feature_aboves[2411]), .feature_below(feature_belows[2411]), .scan_win_std_dev(scan_win_std_dev[2411]), .feature_accum(feature_accums[2411]));
  accum_calculator ac2412(.scan_win(scan_win2412), .rectangle1_x(rectangle1_xs[2412]), .rectangle1_y(rectangle1_ys[2412]), .rectangle1_width(rectangle1_widths[2412]), .rectangle1_height(rectangle1_heights[2412]), .rectangle1_weight(rectangle1_weights[2412]), .rectangle2_x(rectangle2_xs[2412]), .rectangle2_y(rectangle2_ys[2412]), .rectangle2_width(rectangle2_widths[2412]), .rectangle2_height(rectangle2_heights[2412]), .rectangle2_weight(rectangle2_weights[2412]), .rectangle3_x(rectangle3_xs[2412]), .rectangle3_y(rectangle3_ys[2412]), .rectangle3_width(rectangle3_widths[2412]), .rectangle3_height(rectangle3_heights[2412]), .rectangle3_weight(rectangle3_weights[2412]), .feature_threshold(feature_thresholds[2412]), .feature_above(feature_aboves[2412]), .feature_below(feature_belows[2412]), .scan_win_std_dev(scan_win_std_dev[2412]), .feature_accum(feature_accums[2412]));
  accum_calculator ac2413(.scan_win(scan_win2413), .rectangle1_x(rectangle1_xs[2413]), .rectangle1_y(rectangle1_ys[2413]), .rectangle1_width(rectangle1_widths[2413]), .rectangle1_height(rectangle1_heights[2413]), .rectangle1_weight(rectangle1_weights[2413]), .rectangle2_x(rectangle2_xs[2413]), .rectangle2_y(rectangle2_ys[2413]), .rectangle2_width(rectangle2_widths[2413]), .rectangle2_height(rectangle2_heights[2413]), .rectangle2_weight(rectangle2_weights[2413]), .rectangle3_x(rectangle3_xs[2413]), .rectangle3_y(rectangle3_ys[2413]), .rectangle3_width(rectangle3_widths[2413]), .rectangle3_height(rectangle3_heights[2413]), .rectangle3_weight(rectangle3_weights[2413]), .feature_threshold(feature_thresholds[2413]), .feature_above(feature_aboves[2413]), .feature_below(feature_belows[2413]), .scan_win_std_dev(scan_win_std_dev[2413]), .feature_accum(feature_accums[2413]));
  accum_calculator ac2414(.scan_win(scan_win2414), .rectangle1_x(rectangle1_xs[2414]), .rectangle1_y(rectangle1_ys[2414]), .rectangle1_width(rectangle1_widths[2414]), .rectangle1_height(rectangle1_heights[2414]), .rectangle1_weight(rectangle1_weights[2414]), .rectangle2_x(rectangle2_xs[2414]), .rectangle2_y(rectangle2_ys[2414]), .rectangle2_width(rectangle2_widths[2414]), .rectangle2_height(rectangle2_heights[2414]), .rectangle2_weight(rectangle2_weights[2414]), .rectangle3_x(rectangle3_xs[2414]), .rectangle3_y(rectangle3_ys[2414]), .rectangle3_width(rectangle3_widths[2414]), .rectangle3_height(rectangle3_heights[2414]), .rectangle3_weight(rectangle3_weights[2414]), .feature_threshold(feature_thresholds[2414]), .feature_above(feature_aboves[2414]), .feature_below(feature_belows[2414]), .scan_win_std_dev(scan_win_std_dev[2414]), .feature_accum(feature_accums[2414]));
  accum_calculator ac2415(.scan_win(scan_win2415), .rectangle1_x(rectangle1_xs[2415]), .rectangle1_y(rectangle1_ys[2415]), .rectangle1_width(rectangle1_widths[2415]), .rectangle1_height(rectangle1_heights[2415]), .rectangle1_weight(rectangle1_weights[2415]), .rectangle2_x(rectangle2_xs[2415]), .rectangle2_y(rectangle2_ys[2415]), .rectangle2_width(rectangle2_widths[2415]), .rectangle2_height(rectangle2_heights[2415]), .rectangle2_weight(rectangle2_weights[2415]), .rectangle3_x(rectangle3_xs[2415]), .rectangle3_y(rectangle3_ys[2415]), .rectangle3_width(rectangle3_widths[2415]), .rectangle3_height(rectangle3_heights[2415]), .rectangle3_weight(rectangle3_weights[2415]), .feature_threshold(feature_thresholds[2415]), .feature_above(feature_aboves[2415]), .feature_below(feature_belows[2415]), .scan_win_std_dev(scan_win_std_dev[2415]), .feature_accum(feature_accums[2415]));
  accum_calculator ac2416(.scan_win(scan_win2416), .rectangle1_x(rectangle1_xs[2416]), .rectangle1_y(rectangle1_ys[2416]), .rectangle1_width(rectangle1_widths[2416]), .rectangle1_height(rectangle1_heights[2416]), .rectangle1_weight(rectangle1_weights[2416]), .rectangle2_x(rectangle2_xs[2416]), .rectangle2_y(rectangle2_ys[2416]), .rectangle2_width(rectangle2_widths[2416]), .rectangle2_height(rectangle2_heights[2416]), .rectangle2_weight(rectangle2_weights[2416]), .rectangle3_x(rectangle3_xs[2416]), .rectangle3_y(rectangle3_ys[2416]), .rectangle3_width(rectangle3_widths[2416]), .rectangle3_height(rectangle3_heights[2416]), .rectangle3_weight(rectangle3_weights[2416]), .feature_threshold(feature_thresholds[2416]), .feature_above(feature_aboves[2416]), .feature_below(feature_belows[2416]), .scan_win_std_dev(scan_win_std_dev[2416]), .feature_accum(feature_accums[2416]));
  accum_calculator ac2417(.scan_win(scan_win2417), .rectangle1_x(rectangle1_xs[2417]), .rectangle1_y(rectangle1_ys[2417]), .rectangle1_width(rectangle1_widths[2417]), .rectangle1_height(rectangle1_heights[2417]), .rectangle1_weight(rectangle1_weights[2417]), .rectangle2_x(rectangle2_xs[2417]), .rectangle2_y(rectangle2_ys[2417]), .rectangle2_width(rectangle2_widths[2417]), .rectangle2_height(rectangle2_heights[2417]), .rectangle2_weight(rectangle2_weights[2417]), .rectangle3_x(rectangle3_xs[2417]), .rectangle3_y(rectangle3_ys[2417]), .rectangle3_width(rectangle3_widths[2417]), .rectangle3_height(rectangle3_heights[2417]), .rectangle3_weight(rectangle3_weights[2417]), .feature_threshold(feature_thresholds[2417]), .feature_above(feature_aboves[2417]), .feature_below(feature_belows[2417]), .scan_win_std_dev(scan_win_std_dev[2417]), .feature_accum(feature_accums[2417]));
  accum_calculator ac2418(.scan_win(scan_win2418), .rectangle1_x(rectangle1_xs[2418]), .rectangle1_y(rectangle1_ys[2418]), .rectangle1_width(rectangle1_widths[2418]), .rectangle1_height(rectangle1_heights[2418]), .rectangle1_weight(rectangle1_weights[2418]), .rectangle2_x(rectangle2_xs[2418]), .rectangle2_y(rectangle2_ys[2418]), .rectangle2_width(rectangle2_widths[2418]), .rectangle2_height(rectangle2_heights[2418]), .rectangle2_weight(rectangle2_weights[2418]), .rectangle3_x(rectangle3_xs[2418]), .rectangle3_y(rectangle3_ys[2418]), .rectangle3_width(rectangle3_widths[2418]), .rectangle3_height(rectangle3_heights[2418]), .rectangle3_weight(rectangle3_weights[2418]), .feature_threshold(feature_thresholds[2418]), .feature_above(feature_aboves[2418]), .feature_below(feature_belows[2418]), .scan_win_std_dev(scan_win_std_dev[2418]), .feature_accum(feature_accums[2418]));
  accum_calculator ac2419(.scan_win(scan_win2419), .rectangle1_x(rectangle1_xs[2419]), .rectangle1_y(rectangle1_ys[2419]), .rectangle1_width(rectangle1_widths[2419]), .rectangle1_height(rectangle1_heights[2419]), .rectangle1_weight(rectangle1_weights[2419]), .rectangle2_x(rectangle2_xs[2419]), .rectangle2_y(rectangle2_ys[2419]), .rectangle2_width(rectangle2_widths[2419]), .rectangle2_height(rectangle2_heights[2419]), .rectangle2_weight(rectangle2_weights[2419]), .rectangle3_x(rectangle3_xs[2419]), .rectangle3_y(rectangle3_ys[2419]), .rectangle3_width(rectangle3_widths[2419]), .rectangle3_height(rectangle3_heights[2419]), .rectangle3_weight(rectangle3_weights[2419]), .feature_threshold(feature_thresholds[2419]), .feature_above(feature_aboves[2419]), .feature_below(feature_belows[2419]), .scan_win_std_dev(scan_win_std_dev[2419]), .feature_accum(feature_accums[2419]));
  accum_calculator ac2420(.scan_win(scan_win2420), .rectangle1_x(rectangle1_xs[2420]), .rectangle1_y(rectangle1_ys[2420]), .rectangle1_width(rectangle1_widths[2420]), .rectangle1_height(rectangle1_heights[2420]), .rectangle1_weight(rectangle1_weights[2420]), .rectangle2_x(rectangle2_xs[2420]), .rectangle2_y(rectangle2_ys[2420]), .rectangle2_width(rectangle2_widths[2420]), .rectangle2_height(rectangle2_heights[2420]), .rectangle2_weight(rectangle2_weights[2420]), .rectangle3_x(rectangle3_xs[2420]), .rectangle3_y(rectangle3_ys[2420]), .rectangle3_width(rectangle3_widths[2420]), .rectangle3_height(rectangle3_heights[2420]), .rectangle3_weight(rectangle3_weights[2420]), .feature_threshold(feature_thresholds[2420]), .feature_above(feature_aboves[2420]), .feature_below(feature_belows[2420]), .scan_win_std_dev(scan_win_std_dev[2420]), .feature_accum(feature_accums[2420]));
  accum_calculator ac2421(.scan_win(scan_win2421), .rectangle1_x(rectangle1_xs[2421]), .rectangle1_y(rectangle1_ys[2421]), .rectangle1_width(rectangle1_widths[2421]), .rectangle1_height(rectangle1_heights[2421]), .rectangle1_weight(rectangle1_weights[2421]), .rectangle2_x(rectangle2_xs[2421]), .rectangle2_y(rectangle2_ys[2421]), .rectangle2_width(rectangle2_widths[2421]), .rectangle2_height(rectangle2_heights[2421]), .rectangle2_weight(rectangle2_weights[2421]), .rectangle3_x(rectangle3_xs[2421]), .rectangle3_y(rectangle3_ys[2421]), .rectangle3_width(rectangle3_widths[2421]), .rectangle3_height(rectangle3_heights[2421]), .rectangle3_weight(rectangle3_weights[2421]), .feature_threshold(feature_thresholds[2421]), .feature_above(feature_aboves[2421]), .feature_below(feature_belows[2421]), .scan_win_std_dev(scan_win_std_dev[2421]), .feature_accum(feature_accums[2421]));
  accum_calculator ac2422(.scan_win(scan_win2422), .rectangle1_x(rectangle1_xs[2422]), .rectangle1_y(rectangle1_ys[2422]), .rectangle1_width(rectangle1_widths[2422]), .rectangle1_height(rectangle1_heights[2422]), .rectangle1_weight(rectangle1_weights[2422]), .rectangle2_x(rectangle2_xs[2422]), .rectangle2_y(rectangle2_ys[2422]), .rectangle2_width(rectangle2_widths[2422]), .rectangle2_height(rectangle2_heights[2422]), .rectangle2_weight(rectangle2_weights[2422]), .rectangle3_x(rectangle3_xs[2422]), .rectangle3_y(rectangle3_ys[2422]), .rectangle3_width(rectangle3_widths[2422]), .rectangle3_height(rectangle3_heights[2422]), .rectangle3_weight(rectangle3_weights[2422]), .feature_threshold(feature_thresholds[2422]), .feature_above(feature_aboves[2422]), .feature_below(feature_belows[2422]), .scan_win_std_dev(scan_win_std_dev[2422]), .feature_accum(feature_accums[2422]));
  accum_calculator ac2423(.scan_win(scan_win2423), .rectangle1_x(rectangle1_xs[2423]), .rectangle1_y(rectangle1_ys[2423]), .rectangle1_width(rectangle1_widths[2423]), .rectangle1_height(rectangle1_heights[2423]), .rectangle1_weight(rectangle1_weights[2423]), .rectangle2_x(rectangle2_xs[2423]), .rectangle2_y(rectangle2_ys[2423]), .rectangle2_width(rectangle2_widths[2423]), .rectangle2_height(rectangle2_heights[2423]), .rectangle2_weight(rectangle2_weights[2423]), .rectangle3_x(rectangle3_xs[2423]), .rectangle3_y(rectangle3_ys[2423]), .rectangle3_width(rectangle3_widths[2423]), .rectangle3_height(rectangle3_heights[2423]), .rectangle3_weight(rectangle3_weights[2423]), .feature_threshold(feature_thresholds[2423]), .feature_above(feature_aboves[2423]), .feature_below(feature_belows[2423]), .scan_win_std_dev(scan_win_std_dev[2423]), .feature_accum(feature_accums[2423]));
  accum_calculator ac2424(.scan_win(scan_win2424), .rectangle1_x(rectangle1_xs[2424]), .rectangle1_y(rectangle1_ys[2424]), .rectangle1_width(rectangle1_widths[2424]), .rectangle1_height(rectangle1_heights[2424]), .rectangle1_weight(rectangle1_weights[2424]), .rectangle2_x(rectangle2_xs[2424]), .rectangle2_y(rectangle2_ys[2424]), .rectangle2_width(rectangle2_widths[2424]), .rectangle2_height(rectangle2_heights[2424]), .rectangle2_weight(rectangle2_weights[2424]), .rectangle3_x(rectangle3_xs[2424]), .rectangle3_y(rectangle3_ys[2424]), .rectangle3_width(rectangle3_widths[2424]), .rectangle3_height(rectangle3_heights[2424]), .rectangle3_weight(rectangle3_weights[2424]), .feature_threshold(feature_thresholds[2424]), .feature_above(feature_aboves[2424]), .feature_below(feature_belows[2424]), .scan_win_std_dev(scan_win_std_dev[2424]), .feature_accum(feature_accums[2424]));
  accum_calculator ac2425(.scan_win(scan_win2425), .rectangle1_x(rectangle1_xs[2425]), .rectangle1_y(rectangle1_ys[2425]), .rectangle1_width(rectangle1_widths[2425]), .rectangle1_height(rectangle1_heights[2425]), .rectangle1_weight(rectangle1_weights[2425]), .rectangle2_x(rectangle2_xs[2425]), .rectangle2_y(rectangle2_ys[2425]), .rectangle2_width(rectangle2_widths[2425]), .rectangle2_height(rectangle2_heights[2425]), .rectangle2_weight(rectangle2_weights[2425]), .rectangle3_x(rectangle3_xs[2425]), .rectangle3_y(rectangle3_ys[2425]), .rectangle3_width(rectangle3_widths[2425]), .rectangle3_height(rectangle3_heights[2425]), .rectangle3_weight(rectangle3_weights[2425]), .feature_threshold(feature_thresholds[2425]), .feature_above(feature_aboves[2425]), .feature_below(feature_belows[2425]), .scan_win_std_dev(scan_win_std_dev[2425]), .feature_accum(feature_accums[2425]));
  accum_calculator ac2426(.scan_win(scan_win2426), .rectangle1_x(rectangle1_xs[2426]), .rectangle1_y(rectangle1_ys[2426]), .rectangle1_width(rectangle1_widths[2426]), .rectangle1_height(rectangle1_heights[2426]), .rectangle1_weight(rectangle1_weights[2426]), .rectangle2_x(rectangle2_xs[2426]), .rectangle2_y(rectangle2_ys[2426]), .rectangle2_width(rectangle2_widths[2426]), .rectangle2_height(rectangle2_heights[2426]), .rectangle2_weight(rectangle2_weights[2426]), .rectangle3_x(rectangle3_xs[2426]), .rectangle3_y(rectangle3_ys[2426]), .rectangle3_width(rectangle3_widths[2426]), .rectangle3_height(rectangle3_heights[2426]), .rectangle3_weight(rectangle3_weights[2426]), .feature_threshold(feature_thresholds[2426]), .feature_above(feature_aboves[2426]), .feature_below(feature_belows[2426]), .scan_win_std_dev(scan_win_std_dev[2426]), .feature_accum(feature_accums[2426]));
  accum_calculator ac2427(.scan_win(scan_win2427), .rectangle1_x(rectangle1_xs[2427]), .rectangle1_y(rectangle1_ys[2427]), .rectangle1_width(rectangle1_widths[2427]), .rectangle1_height(rectangle1_heights[2427]), .rectangle1_weight(rectangle1_weights[2427]), .rectangle2_x(rectangle2_xs[2427]), .rectangle2_y(rectangle2_ys[2427]), .rectangle2_width(rectangle2_widths[2427]), .rectangle2_height(rectangle2_heights[2427]), .rectangle2_weight(rectangle2_weights[2427]), .rectangle3_x(rectangle3_xs[2427]), .rectangle3_y(rectangle3_ys[2427]), .rectangle3_width(rectangle3_widths[2427]), .rectangle3_height(rectangle3_heights[2427]), .rectangle3_weight(rectangle3_weights[2427]), .feature_threshold(feature_thresholds[2427]), .feature_above(feature_aboves[2427]), .feature_below(feature_belows[2427]), .scan_win_std_dev(scan_win_std_dev[2427]), .feature_accum(feature_accums[2427]));
  accum_calculator ac2428(.scan_win(scan_win2428), .rectangle1_x(rectangle1_xs[2428]), .rectangle1_y(rectangle1_ys[2428]), .rectangle1_width(rectangle1_widths[2428]), .rectangle1_height(rectangle1_heights[2428]), .rectangle1_weight(rectangle1_weights[2428]), .rectangle2_x(rectangle2_xs[2428]), .rectangle2_y(rectangle2_ys[2428]), .rectangle2_width(rectangle2_widths[2428]), .rectangle2_height(rectangle2_heights[2428]), .rectangle2_weight(rectangle2_weights[2428]), .rectangle3_x(rectangle3_xs[2428]), .rectangle3_y(rectangle3_ys[2428]), .rectangle3_width(rectangle3_widths[2428]), .rectangle3_height(rectangle3_heights[2428]), .rectangle3_weight(rectangle3_weights[2428]), .feature_threshold(feature_thresholds[2428]), .feature_above(feature_aboves[2428]), .feature_below(feature_belows[2428]), .scan_win_std_dev(scan_win_std_dev[2428]), .feature_accum(feature_accums[2428]));
  accum_calculator ac2429(.scan_win(scan_win2429), .rectangle1_x(rectangle1_xs[2429]), .rectangle1_y(rectangle1_ys[2429]), .rectangle1_width(rectangle1_widths[2429]), .rectangle1_height(rectangle1_heights[2429]), .rectangle1_weight(rectangle1_weights[2429]), .rectangle2_x(rectangle2_xs[2429]), .rectangle2_y(rectangle2_ys[2429]), .rectangle2_width(rectangle2_widths[2429]), .rectangle2_height(rectangle2_heights[2429]), .rectangle2_weight(rectangle2_weights[2429]), .rectangle3_x(rectangle3_xs[2429]), .rectangle3_y(rectangle3_ys[2429]), .rectangle3_width(rectangle3_widths[2429]), .rectangle3_height(rectangle3_heights[2429]), .rectangle3_weight(rectangle3_weights[2429]), .feature_threshold(feature_thresholds[2429]), .feature_above(feature_aboves[2429]), .feature_below(feature_belows[2429]), .scan_win_std_dev(scan_win_std_dev[2429]), .feature_accum(feature_accums[2429]));
  accum_calculator ac2430(.scan_win(scan_win2430), .rectangle1_x(rectangle1_xs[2430]), .rectangle1_y(rectangle1_ys[2430]), .rectangle1_width(rectangle1_widths[2430]), .rectangle1_height(rectangle1_heights[2430]), .rectangle1_weight(rectangle1_weights[2430]), .rectangle2_x(rectangle2_xs[2430]), .rectangle2_y(rectangle2_ys[2430]), .rectangle2_width(rectangle2_widths[2430]), .rectangle2_height(rectangle2_heights[2430]), .rectangle2_weight(rectangle2_weights[2430]), .rectangle3_x(rectangle3_xs[2430]), .rectangle3_y(rectangle3_ys[2430]), .rectangle3_width(rectangle3_widths[2430]), .rectangle3_height(rectangle3_heights[2430]), .rectangle3_weight(rectangle3_weights[2430]), .feature_threshold(feature_thresholds[2430]), .feature_above(feature_aboves[2430]), .feature_below(feature_belows[2430]), .scan_win_std_dev(scan_win_std_dev[2430]), .feature_accum(feature_accums[2430]));
  accum_calculator ac2431(.scan_win(scan_win2431), .rectangle1_x(rectangle1_xs[2431]), .rectangle1_y(rectangle1_ys[2431]), .rectangle1_width(rectangle1_widths[2431]), .rectangle1_height(rectangle1_heights[2431]), .rectangle1_weight(rectangle1_weights[2431]), .rectangle2_x(rectangle2_xs[2431]), .rectangle2_y(rectangle2_ys[2431]), .rectangle2_width(rectangle2_widths[2431]), .rectangle2_height(rectangle2_heights[2431]), .rectangle2_weight(rectangle2_weights[2431]), .rectangle3_x(rectangle3_xs[2431]), .rectangle3_y(rectangle3_ys[2431]), .rectangle3_width(rectangle3_widths[2431]), .rectangle3_height(rectangle3_heights[2431]), .rectangle3_weight(rectangle3_weights[2431]), .feature_threshold(feature_thresholds[2431]), .feature_above(feature_aboves[2431]), .feature_below(feature_belows[2431]), .scan_win_std_dev(scan_win_std_dev[2431]), .feature_accum(feature_accums[2431]));
  accum_calculator ac2432(.scan_win(scan_win2432), .rectangle1_x(rectangle1_xs[2432]), .rectangle1_y(rectangle1_ys[2432]), .rectangle1_width(rectangle1_widths[2432]), .rectangle1_height(rectangle1_heights[2432]), .rectangle1_weight(rectangle1_weights[2432]), .rectangle2_x(rectangle2_xs[2432]), .rectangle2_y(rectangle2_ys[2432]), .rectangle2_width(rectangle2_widths[2432]), .rectangle2_height(rectangle2_heights[2432]), .rectangle2_weight(rectangle2_weights[2432]), .rectangle3_x(rectangle3_xs[2432]), .rectangle3_y(rectangle3_ys[2432]), .rectangle3_width(rectangle3_widths[2432]), .rectangle3_height(rectangle3_heights[2432]), .rectangle3_weight(rectangle3_weights[2432]), .feature_threshold(feature_thresholds[2432]), .feature_above(feature_aboves[2432]), .feature_below(feature_belows[2432]), .scan_win_std_dev(scan_win_std_dev[2432]), .feature_accum(feature_accums[2432]));
  accum_calculator ac2433(.scan_win(scan_win2433), .rectangle1_x(rectangle1_xs[2433]), .rectangle1_y(rectangle1_ys[2433]), .rectangle1_width(rectangle1_widths[2433]), .rectangle1_height(rectangle1_heights[2433]), .rectangle1_weight(rectangle1_weights[2433]), .rectangle2_x(rectangle2_xs[2433]), .rectangle2_y(rectangle2_ys[2433]), .rectangle2_width(rectangle2_widths[2433]), .rectangle2_height(rectangle2_heights[2433]), .rectangle2_weight(rectangle2_weights[2433]), .rectangle3_x(rectangle3_xs[2433]), .rectangle3_y(rectangle3_ys[2433]), .rectangle3_width(rectangle3_widths[2433]), .rectangle3_height(rectangle3_heights[2433]), .rectangle3_weight(rectangle3_weights[2433]), .feature_threshold(feature_thresholds[2433]), .feature_above(feature_aboves[2433]), .feature_below(feature_belows[2433]), .scan_win_std_dev(scan_win_std_dev[2433]), .feature_accum(feature_accums[2433]));
  accum_calculator ac2434(.scan_win(scan_win2434), .rectangle1_x(rectangle1_xs[2434]), .rectangle1_y(rectangle1_ys[2434]), .rectangle1_width(rectangle1_widths[2434]), .rectangle1_height(rectangle1_heights[2434]), .rectangle1_weight(rectangle1_weights[2434]), .rectangle2_x(rectangle2_xs[2434]), .rectangle2_y(rectangle2_ys[2434]), .rectangle2_width(rectangle2_widths[2434]), .rectangle2_height(rectangle2_heights[2434]), .rectangle2_weight(rectangle2_weights[2434]), .rectangle3_x(rectangle3_xs[2434]), .rectangle3_y(rectangle3_ys[2434]), .rectangle3_width(rectangle3_widths[2434]), .rectangle3_height(rectangle3_heights[2434]), .rectangle3_weight(rectangle3_weights[2434]), .feature_threshold(feature_thresholds[2434]), .feature_above(feature_aboves[2434]), .feature_below(feature_belows[2434]), .scan_win_std_dev(scan_win_std_dev[2434]), .feature_accum(feature_accums[2434]));
  accum_calculator ac2435(.scan_win(scan_win2435), .rectangle1_x(rectangle1_xs[2435]), .rectangle1_y(rectangle1_ys[2435]), .rectangle1_width(rectangle1_widths[2435]), .rectangle1_height(rectangle1_heights[2435]), .rectangle1_weight(rectangle1_weights[2435]), .rectangle2_x(rectangle2_xs[2435]), .rectangle2_y(rectangle2_ys[2435]), .rectangle2_width(rectangle2_widths[2435]), .rectangle2_height(rectangle2_heights[2435]), .rectangle2_weight(rectangle2_weights[2435]), .rectangle3_x(rectangle3_xs[2435]), .rectangle3_y(rectangle3_ys[2435]), .rectangle3_width(rectangle3_widths[2435]), .rectangle3_height(rectangle3_heights[2435]), .rectangle3_weight(rectangle3_weights[2435]), .feature_threshold(feature_thresholds[2435]), .feature_above(feature_aboves[2435]), .feature_below(feature_belows[2435]), .scan_win_std_dev(scan_win_std_dev[2435]), .feature_accum(feature_accums[2435]));
  accum_calculator ac2436(.scan_win(scan_win2436), .rectangle1_x(rectangle1_xs[2436]), .rectangle1_y(rectangle1_ys[2436]), .rectangle1_width(rectangle1_widths[2436]), .rectangle1_height(rectangle1_heights[2436]), .rectangle1_weight(rectangle1_weights[2436]), .rectangle2_x(rectangle2_xs[2436]), .rectangle2_y(rectangle2_ys[2436]), .rectangle2_width(rectangle2_widths[2436]), .rectangle2_height(rectangle2_heights[2436]), .rectangle2_weight(rectangle2_weights[2436]), .rectangle3_x(rectangle3_xs[2436]), .rectangle3_y(rectangle3_ys[2436]), .rectangle3_width(rectangle3_widths[2436]), .rectangle3_height(rectangle3_heights[2436]), .rectangle3_weight(rectangle3_weights[2436]), .feature_threshold(feature_thresholds[2436]), .feature_above(feature_aboves[2436]), .feature_below(feature_belows[2436]), .scan_win_std_dev(scan_win_std_dev[2436]), .feature_accum(feature_accums[2436]));
  accum_calculator ac2437(.scan_win(scan_win2437), .rectangle1_x(rectangle1_xs[2437]), .rectangle1_y(rectangle1_ys[2437]), .rectangle1_width(rectangle1_widths[2437]), .rectangle1_height(rectangle1_heights[2437]), .rectangle1_weight(rectangle1_weights[2437]), .rectangle2_x(rectangle2_xs[2437]), .rectangle2_y(rectangle2_ys[2437]), .rectangle2_width(rectangle2_widths[2437]), .rectangle2_height(rectangle2_heights[2437]), .rectangle2_weight(rectangle2_weights[2437]), .rectangle3_x(rectangle3_xs[2437]), .rectangle3_y(rectangle3_ys[2437]), .rectangle3_width(rectangle3_widths[2437]), .rectangle3_height(rectangle3_heights[2437]), .rectangle3_weight(rectangle3_weights[2437]), .feature_threshold(feature_thresholds[2437]), .feature_above(feature_aboves[2437]), .feature_below(feature_belows[2437]), .scan_win_std_dev(scan_win_std_dev[2437]), .feature_accum(feature_accums[2437]));
  accum_calculator ac2438(.scan_win(scan_win2438), .rectangle1_x(rectangle1_xs[2438]), .rectangle1_y(rectangle1_ys[2438]), .rectangle1_width(rectangle1_widths[2438]), .rectangle1_height(rectangle1_heights[2438]), .rectangle1_weight(rectangle1_weights[2438]), .rectangle2_x(rectangle2_xs[2438]), .rectangle2_y(rectangle2_ys[2438]), .rectangle2_width(rectangle2_widths[2438]), .rectangle2_height(rectangle2_heights[2438]), .rectangle2_weight(rectangle2_weights[2438]), .rectangle3_x(rectangle3_xs[2438]), .rectangle3_y(rectangle3_ys[2438]), .rectangle3_width(rectangle3_widths[2438]), .rectangle3_height(rectangle3_heights[2438]), .rectangle3_weight(rectangle3_weights[2438]), .feature_threshold(feature_thresholds[2438]), .feature_above(feature_aboves[2438]), .feature_below(feature_belows[2438]), .scan_win_std_dev(scan_win_std_dev[2438]), .feature_accum(feature_accums[2438]));
  accum_calculator ac2439(.scan_win(scan_win2439), .rectangle1_x(rectangle1_xs[2439]), .rectangle1_y(rectangle1_ys[2439]), .rectangle1_width(rectangle1_widths[2439]), .rectangle1_height(rectangle1_heights[2439]), .rectangle1_weight(rectangle1_weights[2439]), .rectangle2_x(rectangle2_xs[2439]), .rectangle2_y(rectangle2_ys[2439]), .rectangle2_width(rectangle2_widths[2439]), .rectangle2_height(rectangle2_heights[2439]), .rectangle2_weight(rectangle2_weights[2439]), .rectangle3_x(rectangle3_xs[2439]), .rectangle3_y(rectangle3_ys[2439]), .rectangle3_width(rectangle3_widths[2439]), .rectangle3_height(rectangle3_heights[2439]), .rectangle3_weight(rectangle3_weights[2439]), .feature_threshold(feature_thresholds[2439]), .feature_above(feature_aboves[2439]), .feature_below(feature_belows[2439]), .scan_win_std_dev(scan_win_std_dev[2439]), .feature_accum(feature_accums[2439]));
  accum_calculator ac2440(.scan_win(scan_win2440), .rectangle1_x(rectangle1_xs[2440]), .rectangle1_y(rectangle1_ys[2440]), .rectangle1_width(rectangle1_widths[2440]), .rectangle1_height(rectangle1_heights[2440]), .rectangle1_weight(rectangle1_weights[2440]), .rectangle2_x(rectangle2_xs[2440]), .rectangle2_y(rectangle2_ys[2440]), .rectangle2_width(rectangle2_widths[2440]), .rectangle2_height(rectangle2_heights[2440]), .rectangle2_weight(rectangle2_weights[2440]), .rectangle3_x(rectangle3_xs[2440]), .rectangle3_y(rectangle3_ys[2440]), .rectangle3_width(rectangle3_widths[2440]), .rectangle3_height(rectangle3_heights[2440]), .rectangle3_weight(rectangle3_weights[2440]), .feature_threshold(feature_thresholds[2440]), .feature_above(feature_aboves[2440]), .feature_below(feature_belows[2440]), .scan_win_std_dev(scan_win_std_dev[2440]), .feature_accum(feature_accums[2440]));
  accum_calculator ac2441(.scan_win(scan_win2441), .rectangle1_x(rectangle1_xs[2441]), .rectangle1_y(rectangle1_ys[2441]), .rectangle1_width(rectangle1_widths[2441]), .rectangle1_height(rectangle1_heights[2441]), .rectangle1_weight(rectangle1_weights[2441]), .rectangle2_x(rectangle2_xs[2441]), .rectangle2_y(rectangle2_ys[2441]), .rectangle2_width(rectangle2_widths[2441]), .rectangle2_height(rectangle2_heights[2441]), .rectangle2_weight(rectangle2_weights[2441]), .rectangle3_x(rectangle3_xs[2441]), .rectangle3_y(rectangle3_ys[2441]), .rectangle3_width(rectangle3_widths[2441]), .rectangle3_height(rectangle3_heights[2441]), .rectangle3_weight(rectangle3_weights[2441]), .feature_threshold(feature_thresholds[2441]), .feature_above(feature_aboves[2441]), .feature_below(feature_belows[2441]), .scan_win_std_dev(scan_win_std_dev[2441]), .feature_accum(feature_accums[2441]));
  accum_calculator ac2442(.scan_win(scan_win2442), .rectangle1_x(rectangle1_xs[2442]), .rectangle1_y(rectangle1_ys[2442]), .rectangle1_width(rectangle1_widths[2442]), .rectangle1_height(rectangle1_heights[2442]), .rectangle1_weight(rectangle1_weights[2442]), .rectangle2_x(rectangle2_xs[2442]), .rectangle2_y(rectangle2_ys[2442]), .rectangle2_width(rectangle2_widths[2442]), .rectangle2_height(rectangle2_heights[2442]), .rectangle2_weight(rectangle2_weights[2442]), .rectangle3_x(rectangle3_xs[2442]), .rectangle3_y(rectangle3_ys[2442]), .rectangle3_width(rectangle3_widths[2442]), .rectangle3_height(rectangle3_heights[2442]), .rectangle3_weight(rectangle3_weights[2442]), .feature_threshold(feature_thresholds[2442]), .feature_above(feature_aboves[2442]), .feature_below(feature_belows[2442]), .scan_win_std_dev(scan_win_std_dev[2442]), .feature_accum(feature_accums[2442]));
  accum_calculator ac2443(.scan_win(scan_win2443), .rectangle1_x(rectangle1_xs[2443]), .rectangle1_y(rectangle1_ys[2443]), .rectangle1_width(rectangle1_widths[2443]), .rectangle1_height(rectangle1_heights[2443]), .rectangle1_weight(rectangle1_weights[2443]), .rectangle2_x(rectangle2_xs[2443]), .rectangle2_y(rectangle2_ys[2443]), .rectangle2_width(rectangle2_widths[2443]), .rectangle2_height(rectangle2_heights[2443]), .rectangle2_weight(rectangle2_weights[2443]), .rectangle3_x(rectangle3_xs[2443]), .rectangle3_y(rectangle3_ys[2443]), .rectangle3_width(rectangle3_widths[2443]), .rectangle3_height(rectangle3_heights[2443]), .rectangle3_weight(rectangle3_weights[2443]), .feature_threshold(feature_thresholds[2443]), .feature_above(feature_aboves[2443]), .feature_below(feature_belows[2443]), .scan_win_std_dev(scan_win_std_dev[2443]), .feature_accum(feature_accums[2443]));
  accum_calculator ac2444(.scan_win(scan_win2444), .rectangle1_x(rectangle1_xs[2444]), .rectangle1_y(rectangle1_ys[2444]), .rectangle1_width(rectangle1_widths[2444]), .rectangle1_height(rectangle1_heights[2444]), .rectangle1_weight(rectangle1_weights[2444]), .rectangle2_x(rectangle2_xs[2444]), .rectangle2_y(rectangle2_ys[2444]), .rectangle2_width(rectangle2_widths[2444]), .rectangle2_height(rectangle2_heights[2444]), .rectangle2_weight(rectangle2_weights[2444]), .rectangle3_x(rectangle3_xs[2444]), .rectangle3_y(rectangle3_ys[2444]), .rectangle3_width(rectangle3_widths[2444]), .rectangle3_height(rectangle3_heights[2444]), .rectangle3_weight(rectangle3_weights[2444]), .feature_threshold(feature_thresholds[2444]), .feature_above(feature_aboves[2444]), .feature_below(feature_belows[2444]), .scan_win_std_dev(scan_win_std_dev[2444]), .feature_accum(feature_accums[2444]));
  accum_calculator ac2445(.scan_win(scan_win2445), .rectangle1_x(rectangle1_xs[2445]), .rectangle1_y(rectangle1_ys[2445]), .rectangle1_width(rectangle1_widths[2445]), .rectangle1_height(rectangle1_heights[2445]), .rectangle1_weight(rectangle1_weights[2445]), .rectangle2_x(rectangle2_xs[2445]), .rectangle2_y(rectangle2_ys[2445]), .rectangle2_width(rectangle2_widths[2445]), .rectangle2_height(rectangle2_heights[2445]), .rectangle2_weight(rectangle2_weights[2445]), .rectangle3_x(rectangle3_xs[2445]), .rectangle3_y(rectangle3_ys[2445]), .rectangle3_width(rectangle3_widths[2445]), .rectangle3_height(rectangle3_heights[2445]), .rectangle3_weight(rectangle3_weights[2445]), .feature_threshold(feature_thresholds[2445]), .feature_above(feature_aboves[2445]), .feature_below(feature_belows[2445]), .scan_win_std_dev(scan_win_std_dev[2445]), .feature_accum(feature_accums[2445]));
  accum_calculator ac2446(.scan_win(scan_win2446), .rectangle1_x(rectangle1_xs[2446]), .rectangle1_y(rectangle1_ys[2446]), .rectangle1_width(rectangle1_widths[2446]), .rectangle1_height(rectangle1_heights[2446]), .rectangle1_weight(rectangle1_weights[2446]), .rectangle2_x(rectangle2_xs[2446]), .rectangle2_y(rectangle2_ys[2446]), .rectangle2_width(rectangle2_widths[2446]), .rectangle2_height(rectangle2_heights[2446]), .rectangle2_weight(rectangle2_weights[2446]), .rectangle3_x(rectangle3_xs[2446]), .rectangle3_y(rectangle3_ys[2446]), .rectangle3_width(rectangle3_widths[2446]), .rectangle3_height(rectangle3_heights[2446]), .rectangle3_weight(rectangle3_weights[2446]), .feature_threshold(feature_thresholds[2446]), .feature_above(feature_aboves[2446]), .feature_below(feature_belows[2446]), .scan_win_std_dev(scan_win_std_dev[2446]), .feature_accum(feature_accums[2446]));
  accum_calculator ac2447(.scan_win(scan_win2447), .rectangle1_x(rectangle1_xs[2447]), .rectangle1_y(rectangle1_ys[2447]), .rectangle1_width(rectangle1_widths[2447]), .rectangle1_height(rectangle1_heights[2447]), .rectangle1_weight(rectangle1_weights[2447]), .rectangle2_x(rectangle2_xs[2447]), .rectangle2_y(rectangle2_ys[2447]), .rectangle2_width(rectangle2_widths[2447]), .rectangle2_height(rectangle2_heights[2447]), .rectangle2_weight(rectangle2_weights[2447]), .rectangle3_x(rectangle3_xs[2447]), .rectangle3_y(rectangle3_ys[2447]), .rectangle3_width(rectangle3_widths[2447]), .rectangle3_height(rectangle3_heights[2447]), .rectangle3_weight(rectangle3_weights[2447]), .feature_threshold(feature_thresholds[2447]), .feature_above(feature_aboves[2447]), .feature_below(feature_belows[2447]), .scan_win_std_dev(scan_win_std_dev[2447]), .feature_accum(feature_accums[2447]));
  accum_calculator ac2448(.scan_win(scan_win2448), .rectangle1_x(rectangle1_xs[2448]), .rectangle1_y(rectangle1_ys[2448]), .rectangle1_width(rectangle1_widths[2448]), .rectangle1_height(rectangle1_heights[2448]), .rectangle1_weight(rectangle1_weights[2448]), .rectangle2_x(rectangle2_xs[2448]), .rectangle2_y(rectangle2_ys[2448]), .rectangle2_width(rectangle2_widths[2448]), .rectangle2_height(rectangle2_heights[2448]), .rectangle2_weight(rectangle2_weights[2448]), .rectangle3_x(rectangle3_xs[2448]), .rectangle3_y(rectangle3_ys[2448]), .rectangle3_width(rectangle3_widths[2448]), .rectangle3_height(rectangle3_heights[2448]), .rectangle3_weight(rectangle3_weights[2448]), .feature_threshold(feature_thresholds[2448]), .feature_above(feature_aboves[2448]), .feature_below(feature_belows[2448]), .scan_win_std_dev(scan_win_std_dev[2448]), .feature_accum(feature_accums[2448]));
  accum_calculator ac2449(.scan_win(scan_win2449), .rectangle1_x(rectangle1_xs[2449]), .rectangle1_y(rectangle1_ys[2449]), .rectangle1_width(rectangle1_widths[2449]), .rectangle1_height(rectangle1_heights[2449]), .rectangle1_weight(rectangle1_weights[2449]), .rectangle2_x(rectangle2_xs[2449]), .rectangle2_y(rectangle2_ys[2449]), .rectangle2_width(rectangle2_widths[2449]), .rectangle2_height(rectangle2_heights[2449]), .rectangle2_weight(rectangle2_weights[2449]), .rectangle3_x(rectangle3_xs[2449]), .rectangle3_y(rectangle3_ys[2449]), .rectangle3_width(rectangle3_widths[2449]), .rectangle3_height(rectangle3_heights[2449]), .rectangle3_weight(rectangle3_weights[2449]), .feature_threshold(feature_thresholds[2449]), .feature_above(feature_aboves[2449]), .feature_below(feature_belows[2449]), .scan_win_std_dev(scan_win_std_dev[2449]), .feature_accum(feature_accums[2449]));
  accum_calculator ac2450(.scan_win(scan_win2450), .rectangle1_x(rectangle1_xs[2450]), .rectangle1_y(rectangle1_ys[2450]), .rectangle1_width(rectangle1_widths[2450]), .rectangle1_height(rectangle1_heights[2450]), .rectangle1_weight(rectangle1_weights[2450]), .rectangle2_x(rectangle2_xs[2450]), .rectangle2_y(rectangle2_ys[2450]), .rectangle2_width(rectangle2_widths[2450]), .rectangle2_height(rectangle2_heights[2450]), .rectangle2_weight(rectangle2_weights[2450]), .rectangle3_x(rectangle3_xs[2450]), .rectangle3_y(rectangle3_ys[2450]), .rectangle3_width(rectangle3_widths[2450]), .rectangle3_height(rectangle3_heights[2450]), .rectangle3_weight(rectangle3_weights[2450]), .feature_threshold(feature_thresholds[2450]), .feature_above(feature_aboves[2450]), .feature_below(feature_belows[2450]), .scan_win_std_dev(scan_win_std_dev[2450]), .feature_accum(feature_accums[2450]));
  accum_calculator ac2451(.scan_win(scan_win2451), .rectangle1_x(rectangle1_xs[2451]), .rectangle1_y(rectangle1_ys[2451]), .rectangle1_width(rectangle1_widths[2451]), .rectangle1_height(rectangle1_heights[2451]), .rectangle1_weight(rectangle1_weights[2451]), .rectangle2_x(rectangle2_xs[2451]), .rectangle2_y(rectangle2_ys[2451]), .rectangle2_width(rectangle2_widths[2451]), .rectangle2_height(rectangle2_heights[2451]), .rectangle2_weight(rectangle2_weights[2451]), .rectangle3_x(rectangle3_xs[2451]), .rectangle3_y(rectangle3_ys[2451]), .rectangle3_width(rectangle3_widths[2451]), .rectangle3_height(rectangle3_heights[2451]), .rectangle3_weight(rectangle3_weights[2451]), .feature_threshold(feature_thresholds[2451]), .feature_above(feature_aboves[2451]), .feature_below(feature_belows[2451]), .scan_win_std_dev(scan_win_std_dev[2451]), .feature_accum(feature_accums[2451]));
  accum_calculator ac2452(.scan_win(scan_win2452), .rectangle1_x(rectangle1_xs[2452]), .rectangle1_y(rectangle1_ys[2452]), .rectangle1_width(rectangle1_widths[2452]), .rectangle1_height(rectangle1_heights[2452]), .rectangle1_weight(rectangle1_weights[2452]), .rectangle2_x(rectangle2_xs[2452]), .rectangle2_y(rectangle2_ys[2452]), .rectangle2_width(rectangle2_widths[2452]), .rectangle2_height(rectangle2_heights[2452]), .rectangle2_weight(rectangle2_weights[2452]), .rectangle3_x(rectangle3_xs[2452]), .rectangle3_y(rectangle3_ys[2452]), .rectangle3_width(rectangle3_widths[2452]), .rectangle3_height(rectangle3_heights[2452]), .rectangle3_weight(rectangle3_weights[2452]), .feature_threshold(feature_thresholds[2452]), .feature_above(feature_aboves[2452]), .feature_below(feature_belows[2452]), .scan_win_std_dev(scan_win_std_dev[2452]), .feature_accum(feature_accums[2452]));
  accum_calculator ac2453(.scan_win(scan_win2453), .rectangle1_x(rectangle1_xs[2453]), .rectangle1_y(rectangle1_ys[2453]), .rectangle1_width(rectangle1_widths[2453]), .rectangle1_height(rectangle1_heights[2453]), .rectangle1_weight(rectangle1_weights[2453]), .rectangle2_x(rectangle2_xs[2453]), .rectangle2_y(rectangle2_ys[2453]), .rectangle2_width(rectangle2_widths[2453]), .rectangle2_height(rectangle2_heights[2453]), .rectangle2_weight(rectangle2_weights[2453]), .rectangle3_x(rectangle3_xs[2453]), .rectangle3_y(rectangle3_ys[2453]), .rectangle3_width(rectangle3_widths[2453]), .rectangle3_height(rectangle3_heights[2453]), .rectangle3_weight(rectangle3_weights[2453]), .feature_threshold(feature_thresholds[2453]), .feature_above(feature_aboves[2453]), .feature_below(feature_belows[2453]), .scan_win_std_dev(scan_win_std_dev[2453]), .feature_accum(feature_accums[2453]));
  accum_calculator ac2454(.scan_win(scan_win2454), .rectangle1_x(rectangle1_xs[2454]), .rectangle1_y(rectangle1_ys[2454]), .rectangle1_width(rectangle1_widths[2454]), .rectangle1_height(rectangle1_heights[2454]), .rectangle1_weight(rectangle1_weights[2454]), .rectangle2_x(rectangle2_xs[2454]), .rectangle2_y(rectangle2_ys[2454]), .rectangle2_width(rectangle2_widths[2454]), .rectangle2_height(rectangle2_heights[2454]), .rectangle2_weight(rectangle2_weights[2454]), .rectangle3_x(rectangle3_xs[2454]), .rectangle3_y(rectangle3_ys[2454]), .rectangle3_width(rectangle3_widths[2454]), .rectangle3_height(rectangle3_heights[2454]), .rectangle3_weight(rectangle3_weights[2454]), .feature_threshold(feature_thresholds[2454]), .feature_above(feature_aboves[2454]), .feature_below(feature_belows[2454]), .scan_win_std_dev(scan_win_std_dev[2454]), .feature_accum(feature_accums[2454]));
  accum_calculator ac2455(.scan_win(scan_win2455), .rectangle1_x(rectangle1_xs[2455]), .rectangle1_y(rectangle1_ys[2455]), .rectangle1_width(rectangle1_widths[2455]), .rectangle1_height(rectangle1_heights[2455]), .rectangle1_weight(rectangle1_weights[2455]), .rectangle2_x(rectangle2_xs[2455]), .rectangle2_y(rectangle2_ys[2455]), .rectangle2_width(rectangle2_widths[2455]), .rectangle2_height(rectangle2_heights[2455]), .rectangle2_weight(rectangle2_weights[2455]), .rectangle3_x(rectangle3_xs[2455]), .rectangle3_y(rectangle3_ys[2455]), .rectangle3_width(rectangle3_widths[2455]), .rectangle3_height(rectangle3_heights[2455]), .rectangle3_weight(rectangle3_weights[2455]), .feature_threshold(feature_thresholds[2455]), .feature_above(feature_aboves[2455]), .feature_below(feature_belows[2455]), .scan_win_std_dev(scan_win_std_dev[2455]), .feature_accum(feature_accums[2455]));
  accum_calculator ac2456(.scan_win(scan_win2456), .rectangle1_x(rectangle1_xs[2456]), .rectangle1_y(rectangle1_ys[2456]), .rectangle1_width(rectangle1_widths[2456]), .rectangle1_height(rectangle1_heights[2456]), .rectangle1_weight(rectangle1_weights[2456]), .rectangle2_x(rectangle2_xs[2456]), .rectangle2_y(rectangle2_ys[2456]), .rectangle2_width(rectangle2_widths[2456]), .rectangle2_height(rectangle2_heights[2456]), .rectangle2_weight(rectangle2_weights[2456]), .rectangle3_x(rectangle3_xs[2456]), .rectangle3_y(rectangle3_ys[2456]), .rectangle3_width(rectangle3_widths[2456]), .rectangle3_height(rectangle3_heights[2456]), .rectangle3_weight(rectangle3_weights[2456]), .feature_threshold(feature_thresholds[2456]), .feature_above(feature_aboves[2456]), .feature_below(feature_belows[2456]), .scan_win_std_dev(scan_win_std_dev[2456]), .feature_accum(feature_accums[2456]));
  accum_calculator ac2457(.scan_win(scan_win2457), .rectangle1_x(rectangle1_xs[2457]), .rectangle1_y(rectangle1_ys[2457]), .rectangle1_width(rectangle1_widths[2457]), .rectangle1_height(rectangle1_heights[2457]), .rectangle1_weight(rectangle1_weights[2457]), .rectangle2_x(rectangle2_xs[2457]), .rectangle2_y(rectangle2_ys[2457]), .rectangle2_width(rectangle2_widths[2457]), .rectangle2_height(rectangle2_heights[2457]), .rectangle2_weight(rectangle2_weights[2457]), .rectangle3_x(rectangle3_xs[2457]), .rectangle3_y(rectangle3_ys[2457]), .rectangle3_width(rectangle3_widths[2457]), .rectangle3_height(rectangle3_heights[2457]), .rectangle3_weight(rectangle3_weights[2457]), .feature_threshold(feature_thresholds[2457]), .feature_above(feature_aboves[2457]), .feature_below(feature_belows[2457]), .scan_win_std_dev(scan_win_std_dev[2457]), .feature_accum(feature_accums[2457]));
  accum_calculator ac2458(.scan_win(scan_win2458), .rectangle1_x(rectangle1_xs[2458]), .rectangle1_y(rectangle1_ys[2458]), .rectangle1_width(rectangle1_widths[2458]), .rectangle1_height(rectangle1_heights[2458]), .rectangle1_weight(rectangle1_weights[2458]), .rectangle2_x(rectangle2_xs[2458]), .rectangle2_y(rectangle2_ys[2458]), .rectangle2_width(rectangle2_widths[2458]), .rectangle2_height(rectangle2_heights[2458]), .rectangle2_weight(rectangle2_weights[2458]), .rectangle3_x(rectangle3_xs[2458]), .rectangle3_y(rectangle3_ys[2458]), .rectangle3_width(rectangle3_widths[2458]), .rectangle3_height(rectangle3_heights[2458]), .rectangle3_weight(rectangle3_weights[2458]), .feature_threshold(feature_thresholds[2458]), .feature_above(feature_aboves[2458]), .feature_below(feature_belows[2458]), .scan_win_std_dev(scan_win_std_dev[2458]), .feature_accum(feature_accums[2458]));
  accum_calculator ac2459(.scan_win(scan_win2459), .rectangle1_x(rectangle1_xs[2459]), .rectangle1_y(rectangle1_ys[2459]), .rectangle1_width(rectangle1_widths[2459]), .rectangle1_height(rectangle1_heights[2459]), .rectangle1_weight(rectangle1_weights[2459]), .rectangle2_x(rectangle2_xs[2459]), .rectangle2_y(rectangle2_ys[2459]), .rectangle2_width(rectangle2_widths[2459]), .rectangle2_height(rectangle2_heights[2459]), .rectangle2_weight(rectangle2_weights[2459]), .rectangle3_x(rectangle3_xs[2459]), .rectangle3_y(rectangle3_ys[2459]), .rectangle3_width(rectangle3_widths[2459]), .rectangle3_height(rectangle3_heights[2459]), .rectangle3_weight(rectangle3_weights[2459]), .feature_threshold(feature_thresholds[2459]), .feature_above(feature_aboves[2459]), .feature_below(feature_belows[2459]), .scan_win_std_dev(scan_win_std_dev[2459]), .feature_accum(feature_accums[2459]));
  accum_calculator ac2460(.scan_win(scan_win2460), .rectangle1_x(rectangle1_xs[2460]), .rectangle1_y(rectangle1_ys[2460]), .rectangle1_width(rectangle1_widths[2460]), .rectangle1_height(rectangle1_heights[2460]), .rectangle1_weight(rectangle1_weights[2460]), .rectangle2_x(rectangle2_xs[2460]), .rectangle2_y(rectangle2_ys[2460]), .rectangle2_width(rectangle2_widths[2460]), .rectangle2_height(rectangle2_heights[2460]), .rectangle2_weight(rectangle2_weights[2460]), .rectangle3_x(rectangle3_xs[2460]), .rectangle3_y(rectangle3_ys[2460]), .rectangle3_width(rectangle3_widths[2460]), .rectangle3_height(rectangle3_heights[2460]), .rectangle3_weight(rectangle3_weights[2460]), .feature_threshold(feature_thresholds[2460]), .feature_above(feature_aboves[2460]), .feature_below(feature_belows[2460]), .scan_win_std_dev(scan_win_std_dev[2460]), .feature_accum(feature_accums[2460]));
  accum_calculator ac2461(.scan_win(scan_win2461), .rectangle1_x(rectangle1_xs[2461]), .rectangle1_y(rectangle1_ys[2461]), .rectangle1_width(rectangle1_widths[2461]), .rectangle1_height(rectangle1_heights[2461]), .rectangle1_weight(rectangle1_weights[2461]), .rectangle2_x(rectangle2_xs[2461]), .rectangle2_y(rectangle2_ys[2461]), .rectangle2_width(rectangle2_widths[2461]), .rectangle2_height(rectangle2_heights[2461]), .rectangle2_weight(rectangle2_weights[2461]), .rectangle3_x(rectangle3_xs[2461]), .rectangle3_y(rectangle3_ys[2461]), .rectangle3_width(rectangle3_widths[2461]), .rectangle3_height(rectangle3_heights[2461]), .rectangle3_weight(rectangle3_weights[2461]), .feature_threshold(feature_thresholds[2461]), .feature_above(feature_aboves[2461]), .feature_below(feature_belows[2461]), .scan_win_std_dev(scan_win_std_dev[2461]), .feature_accum(feature_accums[2461]));
  accum_calculator ac2462(.scan_win(scan_win2462), .rectangle1_x(rectangle1_xs[2462]), .rectangle1_y(rectangle1_ys[2462]), .rectangle1_width(rectangle1_widths[2462]), .rectangle1_height(rectangle1_heights[2462]), .rectangle1_weight(rectangle1_weights[2462]), .rectangle2_x(rectangle2_xs[2462]), .rectangle2_y(rectangle2_ys[2462]), .rectangle2_width(rectangle2_widths[2462]), .rectangle2_height(rectangle2_heights[2462]), .rectangle2_weight(rectangle2_weights[2462]), .rectangle3_x(rectangle3_xs[2462]), .rectangle3_y(rectangle3_ys[2462]), .rectangle3_width(rectangle3_widths[2462]), .rectangle3_height(rectangle3_heights[2462]), .rectangle3_weight(rectangle3_weights[2462]), .feature_threshold(feature_thresholds[2462]), .feature_above(feature_aboves[2462]), .feature_below(feature_belows[2462]), .scan_win_std_dev(scan_win_std_dev[2462]), .feature_accum(feature_accums[2462]));
  accum_calculator ac2463(.scan_win(scan_win2463), .rectangle1_x(rectangle1_xs[2463]), .rectangle1_y(rectangle1_ys[2463]), .rectangle1_width(rectangle1_widths[2463]), .rectangle1_height(rectangle1_heights[2463]), .rectangle1_weight(rectangle1_weights[2463]), .rectangle2_x(rectangle2_xs[2463]), .rectangle2_y(rectangle2_ys[2463]), .rectangle2_width(rectangle2_widths[2463]), .rectangle2_height(rectangle2_heights[2463]), .rectangle2_weight(rectangle2_weights[2463]), .rectangle3_x(rectangle3_xs[2463]), .rectangle3_y(rectangle3_ys[2463]), .rectangle3_width(rectangle3_widths[2463]), .rectangle3_height(rectangle3_heights[2463]), .rectangle3_weight(rectangle3_weights[2463]), .feature_threshold(feature_thresholds[2463]), .feature_above(feature_aboves[2463]), .feature_below(feature_belows[2463]), .scan_win_std_dev(scan_win_std_dev[2463]), .feature_accum(feature_accums[2463]));
  accum_calculator ac2464(.scan_win(scan_win2464), .rectangle1_x(rectangle1_xs[2464]), .rectangle1_y(rectangle1_ys[2464]), .rectangle1_width(rectangle1_widths[2464]), .rectangle1_height(rectangle1_heights[2464]), .rectangle1_weight(rectangle1_weights[2464]), .rectangle2_x(rectangle2_xs[2464]), .rectangle2_y(rectangle2_ys[2464]), .rectangle2_width(rectangle2_widths[2464]), .rectangle2_height(rectangle2_heights[2464]), .rectangle2_weight(rectangle2_weights[2464]), .rectangle3_x(rectangle3_xs[2464]), .rectangle3_y(rectangle3_ys[2464]), .rectangle3_width(rectangle3_widths[2464]), .rectangle3_height(rectangle3_heights[2464]), .rectangle3_weight(rectangle3_weights[2464]), .feature_threshold(feature_thresholds[2464]), .feature_above(feature_aboves[2464]), .feature_below(feature_belows[2464]), .scan_win_std_dev(scan_win_std_dev[2464]), .feature_accum(feature_accums[2464]));
  accum_calculator ac2465(.scan_win(scan_win2465), .rectangle1_x(rectangle1_xs[2465]), .rectangle1_y(rectangle1_ys[2465]), .rectangle1_width(rectangle1_widths[2465]), .rectangle1_height(rectangle1_heights[2465]), .rectangle1_weight(rectangle1_weights[2465]), .rectangle2_x(rectangle2_xs[2465]), .rectangle2_y(rectangle2_ys[2465]), .rectangle2_width(rectangle2_widths[2465]), .rectangle2_height(rectangle2_heights[2465]), .rectangle2_weight(rectangle2_weights[2465]), .rectangle3_x(rectangle3_xs[2465]), .rectangle3_y(rectangle3_ys[2465]), .rectangle3_width(rectangle3_widths[2465]), .rectangle3_height(rectangle3_heights[2465]), .rectangle3_weight(rectangle3_weights[2465]), .feature_threshold(feature_thresholds[2465]), .feature_above(feature_aboves[2465]), .feature_below(feature_belows[2465]), .scan_win_std_dev(scan_win_std_dev[2465]), .feature_accum(feature_accums[2465]));
  accum_calculator ac2466(.scan_win(scan_win2466), .rectangle1_x(rectangle1_xs[2466]), .rectangle1_y(rectangle1_ys[2466]), .rectangle1_width(rectangle1_widths[2466]), .rectangle1_height(rectangle1_heights[2466]), .rectangle1_weight(rectangle1_weights[2466]), .rectangle2_x(rectangle2_xs[2466]), .rectangle2_y(rectangle2_ys[2466]), .rectangle2_width(rectangle2_widths[2466]), .rectangle2_height(rectangle2_heights[2466]), .rectangle2_weight(rectangle2_weights[2466]), .rectangle3_x(rectangle3_xs[2466]), .rectangle3_y(rectangle3_ys[2466]), .rectangle3_width(rectangle3_widths[2466]), .rectangle3_height(rectangle3_heights[2466]), .rectangle3_weight(rectangle3_weights[2466]), .feature_threshold(feature_thresholds[2466]), .feature_above(feature_aboves[2466]), .feature_below(feature_belows[2466]), .scan_win_std_dev(scan_win_std_dev[2466]), .feature_accum(feature_accums[2466]));
  accum_calculator ac2467(.scan_win(scan_win2467), .rectangle1_x(rectangle1_xs[2467]), .rectangle1_y(rectangle1_ys[2467]), .rectangle1_width(rectangle1_widths[2467]), .rectangle1_height(rectangle1_heights[2467]), .rectangle1_weight(rectangle1_weights[2467]), .rectangle2_x(rectangle2_xs[2467]), .rectangle2_y(rectangle2_ys[2467]), .rectangle2_width(rectangle2_widths[2467]), .rectangle2_height(rectangle2_heights[2467]), .rectangle2_weight(rectangle2_weights[2467]), .rectangle3_x(rectangle3_xs[2467]), .rectangle3_y(rectangle3_ys[2467]), .rectangle3_width(rectangle3_widths[2467]), .rectangle3_height(rectangle3_heights[2467]), .rectangle3_weight(rectangle3_weights[2467]), .feature_threshold(feature_thresholds[2467]), .feature_above(feature_aboves[2467]), .feature_below(feature_belows[2467]), .scan_win_std_dev(scan_win_std_dev[2467]), .feature_accum(feature_accums[2467]));
  accum_calculator ac2468(.scan_win(scan_win2468), .rectangle1_x(rectangle1_xs[2468]), .rectangle1_y(rectangle1_ys[2468]), .rectangle1_width(rectangle1_widths[2468]), .rectangle1_height(rectangle1_heights[2468]), .rectangle1_weight(rectangle1_weights[2468]), .rectangle2_x(rectangle2_xs[2468]), .rectangle2_y(rectangle2_ys[2468]), .rectangle2_width(rectangle2_widths[2468]), .rectangle2_height(rectangle2_heights[2468]), .rectangle2_weight(rectangle2_weights[2468]), .rectangle3_x(rectangle3_xs[2468]), .rectangle3_y(rectangle3_ys[2468]), .rectangle3_width(rectangle3_widths[2468]), .rectangle3_height(rectangle3_heights[2468]), .rectangle3_weight(rectangle3_weights[2468]), .feature_threshold(feature_thresholds[2468]), .feature_above(feature_aboves[2468]), .feature_below(feature_belows[2468]), .scan_win_std_dev(scan_win_std_dev[2468]), .feature_accum(feature_accums[2468]));
  accum_calculator ac2469(.scan_win(scan_win2469), .rectangle1_x(rectangle1_xs[2469]), .rectangle1_y(rectangle1_ys[2469]), .rectangle1_width(rectangle1_widths[2469]), .rectangle1_height(rectangle1_heights[2469]), .rectangle1_weight(rectangle1_weights[2469]), .rectangle2_x(rectangle2_xs[2469]), .rectangle2_y(rectangle2_ys[2469]), .rectangle2_width(rectangle2_widths[2469]), .rectangle2_height(rectangle2_heights[2469]), .rectangle2_weight(rectangle2_weights[2469]), .rectangle3_x(rectangle3_xs[2469]), .rectangle3_y(rectangle3_ys[2469]), .rectangle3_width(rectangle3_widths[2469]), .rectangle3_height(rectangle3_heights[2469]), .rectangle3_weight(rectangle3_weights[2469]), .feature_threshold(feature_thresholds[2469]), .feature_above(feature_aboves[2469]), .feature_below(feature_belows[2469]), .scan_win_std_dev(scan_win_std_dev[2469]), .feature_accum(feature_accums[2469]));
  accum_calculator ac2470(.scan_win(scan_win2470), .rectangle1_x(rectangle1_xs[2470]), .rectangle1_y(rectangle1_ys[2470]), .rectangle1_width(rectangle1_widths[2470]), .rectangle1_height(rectangle1_heights[2470]), .rectangle1_weight(rectangle1_weights[2470]), .rectangle2_x(rectangle2_xs[2470]), .rectangle2_y(rectangle2_ys[2470]), .rectangle2_width(rectangle2_widths[2470]), .rectangle2_height(rectangle2_heights[2470]), .rectangle2_weight(rectangle2_weights[2470]), .rectangle3_x(rectangle3_xs[2470]), .rectangle3_y(rectangle3_ys[2470]), .rectangle3_width(rectangle3_widths[2470]), .rectangle3_height(rectangle3_heights[2470]), .rectangle3_weight(rectangle3_weights[2470]), .feature_threshold(feature_thresholds[2470]), .feature_above(feature_aboves[2470]), .feature_below(feature_belows[2470]), .scan_win_std_dev(scan_win_std_dev[2470]), .feature_accum(feature_accums[2470]));
  accum_calculator ac2471(.scan_win(scan_win2471), .rectangle1_x(rectangle1_xs[2471]), .rectangle1_y(rectangle1_ys[2471]), .rectangle1_width(rectangle1_widths[2471]), .rectangle1_height(rectangle1_heights[2471]), .rectangle1_weight(rectangle1_weights[2471]), .rectangle2_x(rectangle2_xs[2471]), .rectangle2_y(rectangle2_ys[2471]), .rectangle2_width(rectangle2_widths[2471]), .rectangle2_height(rectangle2_heights[2471]), .rectangle2_weight(rectangle2_weights[2471]), .rectangle3_x(rectangle3_xs[2471]), .rectangle3_y(rectangle3_ys[2471]), .rectangle3_width(rectangle3_widths[2471]), .rectangle3_height(rectangle3_heights[2471]), .rectangle3_weight(rectangle3_weights[2471]), .feature_threshold(feature_thresholds[2471]), .feature_above(feature_aboves[2471]), .feature_below(feature_belows[2471]), .scan_win_std_dev(scan_win_std_dev[2471]), .feature_accum(feature_accums[2471]));
  accum_calculator ac2472(.scan_win(scan_win2472), .rectangle1_x(rectangle1_xs[2472]), .rectangle1_y(rectangle1_ys[2472]), .rectangle1_width(rectangle1_widths[2472]), .rectangle1_height(rectangle1_heights[2472]), .rectangle1_weight(rectangle1_weights[2472]), .rectangle2_x(rectangle2_xs[2472]), .rectangle2_y(rectangle2_ys[2472]), .rectangle2_width(rectangle2_widths[2472]), .rectangle2_height(rectangle2_heights[2472]), .rectangle2_weight(rectangle2_weights[2472]), .rectangle3_x(rectangle3_xs[2472]), .rectangle3_y(rectangle3_ys[2472]), .rectangle3_width(rectangle3_widths[2472]), .rectangle3_height(rectangle3_heights[2472]), .rectangle3_weight(rectangle3_weights[2472]), .feature_threshold(feature_thresholds[2472]), .feature_above(feature_aboves[2472]), .feature_below(feature_belows[2472]), .scan_win_std_dev(scan_win_std_dev[2472]), .feature_accum(feature_accums[2472]));
  accum_calculator ac2473(.scan_win(scan_win2473), .rectangle1_x(rectangle1_xs[2473]), .rectangle1_y(rectangle1_ys[2473]), .rectangle1_width(rectangle1_widths[2473]), .rectangle1_height(rectangle1_heights[2473]), .rectangle1_weight(rectangle1_weights[2473]), .rectangle2_x(rectangle2_xs[2473]), .rectangle2_y(rectangle2_ys[2473]), .rectangle2_width(rectangle2_widths[2473]), .rectangle2_height(rectangle2_heights[2473]), .rectangle2_weight(rectangle2_weights[2473]), .rectangle3_x(rectangle3_xs[2473]), .rectangle3_y(rectangle3_ys[2473]), .rectangle3_width(rectangle3_widths[2473]), .rectangle3_height(rectangle3_heights[2473]), .rectangle3_weight(rectangle3_weights[2473]), .feature_threshold(feature_thresholds[2473]), .feature_above(feature_aboves[2473]), .feature_below(feature_belows[2473]), .scan_win_std_dev(scan_win_std_dev[2473]), .feature_accum(feature_accums[2473]));
  accum_calculator ac2474(.scan_win(scan_win2474), .rectangle1_x(rectangle1_xs[2474]), .rectangle1_y(rectangle1_ys[2474]), .rectangle1_width(rectangle1_widths[2474]), .rectangle1_height(rectangle1_heights[2474]), .rectangle1_weight(rectangle1_weights[2474]), .rectangle2_x(rectangle2_xs[2474]), .rectangle2_y(rectangle2_ys[2474]), .rectangle2_width(rectangle2_widths[2474]), .rectangle2_height(rectangle2_heights[2474]), .rectangle2_weight(rectangle2_weights[2474]), .rectangle3_x(rectangle3_xs[2474]), .rectangle3_y(rectangle3_ys[2474]), .rectangle3_width(rectangle3_widths[2474]), .rectangle3_height(rectangle3_heights[2474]), .rectangle3_weight(rectangle3_weights[2474]), .feature_threshold(feature_thresholds[2474]), .feature_above(feature_aboves[2474]), .feature_below(feature_belows[2474]), .scan_win_std_dev(scan_win_std_dev[2474]), .feature_accum(feature_accums[2474]));
  accum_calculator ac2475(.scan_win(scan_win2475), .rectangle1_x(rectangle1_xs[2475]), .rectangle1_y(rectangle1_ys[2475]), .rectangle1_width(rectangle1_widths[2475]), .rectangle1_height(rectangle1_heights[2475]), .rectangle1_weight(rectangle1_weights[2475]), .rectangle2_x(rectangle2_xs[2475]), .rectangle2_y(rectangle2_ys[2475]), .rectangle2_width(rectangle2_widths[2475]), .rectangle2_height(rectangle2_heights[2475]), .rectangle2_weight(rectangle2_weights[2475]), .rectangle3_x(rectangle3_xs[2475]), .rectangle3_y(rectangle3_ys[2475]), .rectangle3_width(rectangle3_widths[2475]), .rectangle3_height(rectangle3_heights[2475]), .rectangle3_weight(rectangle3_weights[2475]), .feature_threshold(feature_thresholds[2475]), .feature_above(feature_aboves[2475]), .feature_below(feature_belows[2475]), .scan_win_std_dev(scan_win_std_dev[2475]), .feature_accum(feature_accums[2475]));
  accum_calculator ac2476(.scan_win(scan_win2476), .rectangle1_x(rectangle1_xs[2476]), .rectangle1_y(rectangle1_ys[2476]), .rectangle1_width(rectangle1_widths[2476]), .rectangle1_height(rectangle1_heights[2476]), .rectangle1_weight(rectangle1_weights[2476]), .rectangle2_x(rectangle2_xs[2476]), .rectangle2_y(rectangle2_ys[2476]), .rectangle2_width(rectangle2_widths[2476]), .rectangle2_height(rectangle2_heights[2476]), .rectangle2_weight(rectangle2_weights[2476]), .rectangle3_x(rectangle3_xs[2476]), .rectangle3_y(rectangle3_ys[2476]), .rectangle3_width(rectangle3_widths[2476]), .rectangle3_height(rectangle3_heights[2476]), .rectangle3_weight(rectangle3_weights[2476]), .feature_threshold(feature_thresholds[2476]), .feature_above(feature_aboves[2476]), .feature_below(feature_belows[2476]), .scan_win_std_dev(scan_win_std_dev[2476]), .feature_accum(feature_accums[2476]));
  accum_calculator ac2477(.scan_win(scan_win2477), .rectangle1_x(rectangle1_xs[2477]), .rectangle1_y(rectangle1_ys[2477]), .rectangle1_width(rectangle1_widths[2477]), .rectangle1_height(rectangle1_heights[2477]), .rectangle1_weight(rectangle1_weights[2477]), .rectangle2_x(rectangle2_xs[2477]), .rectangle2_y(rectangle2_ys[2477]), .rectangle2_width(rectangle2_widths[2477]), .rectangle2_height(rectangle2_heights[2477]), .rectangle2_weight(rectangle2_weights[2477]), .rectangle3_x(rectangle3_xs[2477]), .rectangle3_y(rectangle3_ys[2477]), .rectangle3_width(rectangle3_widths[2477]), .rectangle3_height(rectangle3_heights[2477]), .rectangle3_weight(rectangle3_weights[2477]), .feature_threshold(feature_thresholds[2477]), .feature_above(feature_aboves[2477]), .feature_below(feature_belows[2477]), .scan_win_std_dev(scan_win_std_dev[2477]), .feature_accum(feature_accums[2477]));
  accum_calculator ac2478(.scan_win(scan_win2478), .rectangle1_x(rectangle1_xs[2478]), .rectangle1_y(rectangle1_ys[2478]), .rectangle1_width(rectangle1_widths[2478]), .rectangle1_height(rectangle1_heights[2478]), .rectangle1_weight(rectangle1_weights[2478]), .rectangle2_x(rectangle2_xs[2478]), .rectangle2_y(rectangle2_ys[2478]), .rectangle2_width(rectangle2_widths[2478]), .rectangle2_height(rectangle2_heights[2478]), .rectangle2_weight(rectangle2_weights[2478]), .rectangle3_x(rectangle3_xs[2478]), .rectangle3_y(rectangle3_ys[2478]), .rectangle3_width(rectangle3_widths[2478]), .rectangle3_height(rectangle3_heights[2478]), .rectangle3_weight(rectangle3_weights[2478]), .feature_threshold(feature_thresholds[2478]), .feature_above(feature_aboves[2478]), .feature_below(feature_belows[2478]), .scan_win_std_dev(scan_win_std_dev[2478]), .feature_accum(feature_accums[2478]));
  accum_calculator ac2479(.scan_win(scan_win2479), .rectangle1_x(rectangle1_xs[2479]), .rectangle1_y(rectangle1_ys[2479]), .rectangle1_width(rectangle1_widths[2479]), .rectangle1_height(rectangle1_heights[2479]), .rectangle1_weight(rectangle1_weights[2479]), .rectangle2_x(rectangle2_xs[2479]), .rectangle2_y(rectangle2_ys[2479]), .rectangle2_width(rectangle2_widths[2479]), .rectangle2_height(rectangle2_heights[2479]), .rectangle2_weight(rectangle2_weights[2479]), .rectangle3_x(rectangle3_xs[2479]), .rectangle3_y(rectangle3_ys[2479]), .rectangle3_width(rectangle3_widths[2479]), .rectangle3_height(rectangle3_heights[2479]), .rectangle3_weight(rectangle3_weights[2479]), .feature_threshold(feature_thresholds[2479]), .feature_above(feature_aboves[2479]), .feature_below(feature_belows[2479]), .scan_win_std_dev(scan_win_std_dev[2479]), .feature_accum(feature_accums[2479]));
  accum_calculator ac2480(.scan_win(scan_win2480), .rectangle1_x(rectangle1_xs[2480]), .rectangle1_y(rectangle1_ys[2480]), .rectangle1_width(rectangle1_widths[2480]), .rectangle1_height(rectangle1_heights[2480]), .rectangle1_weight(rectangle1_weights[2480]), .rectangle2_x(rectangle2_xs[2480]), .rectangle2_y(rectangle2_ys[2480]), .rectangle2_width(rectangle2_widths[2480]), .rectangle2_height(rectangle2_heights[2480]), .rectangle2_weight(rectangle2_weights[2480]), .rectangle3_x(rectangle3_xs[2480]), .rectangle3_y(rectangle3_ys[2480]), .rectangle3_width(rectangle3_widths[2480]), .rectangle3_height(rectangle3_heights[2480]), .rectangle3_weight(rectangle3_weights[2480]), .feature_threshold(feature_thresholds[2480]), .feature_above(feature_aboves[2480]), .feature_below(feature_belows[2480]), .scan_win_std_dev(scan_win_std_dev[2480]), .feature_accum(feature_accums[2480]));
  accum_calculator ac2481(.scan_win(scan_win2481), .rectangle1_x(rectangle1_xs[2481]), .rectangle1_y(rectangle1_ys[2481]), .rectangle1_width(rectangle1_widths[2481]), .rectangle1_height(rectangle1_heights[2481]), .rectangle1_weight(rectangle1_weights[2481]), .rectangle2_x(rectangle2_xs[2481]), .rectangle2_y(rectangle2_ys[2481]), .rectangle2_width(rectangle2_widths[2481]), .rectangle2_height(rectangle2_heights[2481]), .rectangle2_weight(rectangle2_weights[2481]), .rectangle3_x(rectangle3_xs[2481]), .rectangle3_y(rectangle3_ys[2481]), .rectangle3_width(rectangle3_widths[2481]), .rectangle3_height(rectangle3_heights[2481]), .rectangle3_weight(rectangle3_weights[2481]), .feature_threshold(feature_thresholds[2481]), .feature_above(feature_aboves[2481]), .feature_below(feature_belows[2481]), .scan_win_std_dev(scan_win_std_dev[2481]), .feature_accum(feature_accums[2481]));
  accum_calculator ac2482(.scan_win(scan_win2482), .rectangle1_x(rectangle1_xs[2482]), .rectangle1_y(rectangle1_ys[2482]), .rectangle1_width(rectangle1_widths[2482]), .rectangle1_height(rectangle1_heights[2482]), .rectangle1_weight(rectangle1_weights[2482]), .rectangle2_x(rectangle2_xs[2482]), .rectangle2_y(rectangle2_ys[2482]), .rectangle2_width(rectangle2_widths[2482]), .rectangle2_height(rectangle2_heights[2482]), .rectangle2_weight(rectangle2_weights[2482]), .rectangle3_x(rectangle3_xs[2482]), .rectangle3_y(rectangle3_ys[2482]), .rectangle3_width(rectangle3_widths[2482]), .rectangle3_height(rectangle3_heights[2482]), .rectangle3_weight(rectangle3_weights[2482]), .feature_threshold(feature_thresholds[2482]), .feature_above(feature_aboves[2482]), .feature_below(feature_belows[2482]), .scan_win_std_dev(scan_win_std_dev[2482]), .feature_accum(feature_accums[2482]));
  accum_calculator ac2483(.scan_win(scan_win2483), .rectangle1_x(rectangle1_xs[2483]), .rectangle1_y(rectangle1_ys[2483]), .rectangle1_width(rectangle1_widths[2483]), .rectangle1_height(rectangle1_heights[2483]), .rectangle1_weight(rectangle1_weights[2483]), .rectangle2_x(rectangle2_xs[2483]), .rectangle2_y(rectangle2_ys[2483]), .rectangle2_width(rectangle2_widths[2483]), .rectangle2_height(rectangle2_heights[2483]), .rectangle2_weight(rectangle2_weights[2483]), .rectangle3_x(rectangle3_xs[2483]), .rectangle3_y(rectangle3_ys[2483]), .rectangle3_width(rectangle3_widths[2483]), .rectangle3_height(rectangle3_heights[2483]), .rectangle3_weight(rectangle3_weights[2483]), .feature_threshold(feature_thresholds[2483]), .feature_above(feature_aboves[2483]), .feature_below(feature_belows[2483]), .scan_win_std_dev(scan_win_std_dev[2483]), .feature_accum(feature_accums[2483]));
  accum_calculator ac2484(.scan_win(scan_win2484), .rectangle1_x(rectangle1_xs[2484]), .rectangle1_y(rectangle1_ys[2484]), .rectangle1_width(rectangle1_widths[2484]), .rectangle1_height(rectangle1_heights[2484]), .rectangle1_weight(rectangle1_weights[2484]), .rectangle2_x(rectangle2_xs[2484]), .rectangle2_y(rectangle2_ys[2484]), .rectangle2_width(rectangle2_widths[2484]), .rectangle2_height(rectangle2_heights[2484]), .rectangle2_weight(rectangle2_weights[2484]), .rectangle3_x(rectangle3_xs[2484]), .rectangle3_y(rectangle3_ys[2484]), .rectangle3_width(rectangle3_widths[2484]), .rectangle3_height(rectangle3_heights[2484]), .rectangle3_weight(rectangle3_weights[2484]), .feature_threshold(feature_thresholds[2484]), .feature_above(feature_aboves[2484]), .feature_below(feature_belows[2484]), .scan_win_std_dev(scan_win_std_dev[2484]), .feature_accum(feature_accums[2484]));
  accum_calculator ac2485(.scan_win(scan_win2485), .rectangle1_x(rectangle1_xs[2485]), .rectangle1_y(rectangle1_ys[2485]), .rectangle1_width(rectangle1_widths[2485]), .rectangle1_height(rectangle1_heights[2485]), .rectangle1_weight(rectangle1_weights[2485]), .rectangle2_x(rectangle2_xs[2485]), .rectangle2_y(rectangle2_ys[2485]), .rectangle2_width(rectangle2_widths[2485]), .rectangle2_height(rectangle2_heights[2485]), .rectangle2_weight(rectangle2_weights[2485]), .rectangle3_x(rectangle3_xs[2485]), .rectangle3_y(rectangle3_ys[2485]), .rectangle3_width(rectangle3_widths[2485]), .rectangle3_height(rectangle3_heights[2485]), .rectangle3_weight(rectangle3_weights[2485]), .feature_threshold(feature_thresholds[2485]), .feature_above(feature_aboves[2485]), .feature_below(feature_belows[2485]), .scan_win_std_dev(scan_win_std_dev[2485]), .feature_accum(feature_accums[2485]));
  accum_calculator ac2486(.scan_win(scan_win2486), .rectangle1_x(rectangle1_xs[2486]), .rectangle1_y(rectangle1_ys[2486]), .rectangle1_width(rectangle1_widths[2486]), .rectangle1_height(rectangle1_heights[2486]), .rectangle1_weight(rectangle1_weights[2486]), .rectangle2_x(rectangle2_xs[2486]), .rectangle2_y(rectangle2_ys[2486]), .rectangle2_width(rectangle2_widths[2486]), .rectangle2_height(rectangle2_heights[2486]), .rectangle2_weight(rectangle2_weights[2486]), .rectangle3_x(rectangle3_xs[2486]), .rectangle3_y(rectangle3_ys[2486]), .rectangle3_width(rectangle3_widths[2486]), .rectangle3_height(rectangle3_heights[2486]), .rectangle3_weight(rectangle3_weights[2486]), .feature_threshold(feature_thresholds[2486]), .feature_above(feature_aboves[2486]), .feature_below(feature_belows[2486]), .scan_win_std_dev(scan_win_std_dev[2486]), .feature_accum(feature_accums[2486]));
  accum_calculator ac2487(.scan_win(scan_win2487), .rectangle1_x(rectangle1_xs[2487]), .rectangle1_y(rectangle1_ys[2487]), .rectangle1_width(rectangle1_widths[2487]), .rectangle1_height(rectangle1_heights[2487]), .rectangle1_weight(rectangle1_weights[2487]), .rectangle2_x(rectangle2_xs[2487]), .rectangle2_y(rectangle2_ys[2487]), .rectangle2_width(rectangle2_widths[2487]), .rectangle2_height(rectangle2_heights[2487]), .rectangle2_weight(rectangle2_weights[2487]), .rectangle3_x(rectangle3_xs[2487]), .rectangle3_y(rectangle3_ys[2487]), .rectangle3_width(rectangle3_widths[2487]), .rectangle3_height(rectangle3_heights[2487]), .rectangle3_weight(rectangle3_weights[2487]), .feature_threshold(feature_thresholds[2487]), .feature_above(feature_aboves[2487]), .feature_below(feature_belows[2487]), .scan_win_std_dev(scan_win_std_dev[2487]), .feature_accum(feature_accums[2487]));
  accum_calculator ac2488(.scan_win(scan_win2488), .rectangle1_x(rectangle1_xs[2488]), .rectangle1_y(rectangle1_ys[2488]), .rectangle1_width(rectangle1_widths[2488]), .rectangle1_height(rectangle1_heights[2488]), .rectangle1_weight(rectangle1_weights[2488]), .rectangle2_x(rectangle2_xs[2488]), .rectangle2_y(rectangle2_ys[2488]), .rectangle2_width(rectangle2_widths[2488]), .rectangle2_height(rectangle2_heights[2488]), .rectangle2_weight(rectangle2_weights[2488]), .rectangle3_x(rectangle3_xs[2488]), .rectangle3_y(rectangle3_ys[2488]), .rectangle3_width(rectangle3_widths[2488]), .rectangle3_height(rectangle3_heights[2488]), .rectangle3_weight(rectangle3_weights[2488]), .feature_threshold(feature_thresholds[2488]), .feature_above(feature_aboves[2488]), .feature_below(feature_belows[2488]), .scan_win_std_dev(scan_win_std_dev[2488]), .feature_accum(feature_accums[2488]));
  accum_calculator ac2489(.scan_win(scan_win2489), .rectangle1_x(rectangle1_xs[2489]), .rectangle1_y(rectangle1_ys[2489]), .rectangle1_width(rectangle1_widths[2489]), .rectangle1_height(rectangle1_heights[2489]), .rectangle1_weight(rectangle1_weights[2489]), .rectangle2_x(rectangle2_xs[2489]), .rectangle2_y(rectangle2_ys[2489]), .rectangle2_width(rectangle2_widths[2489]), .rectangle2_height(rectangle2_heights[2489]), .rectangle2_weight(rectangle2_weights[2489]), .rectangle3_x(rectangle3_xs[2489]), .rectangle3_y(rectangle3_ys[2489]), .rectangle3_width(rectangle3_widths[2489]), .rectangle3_height(rectangle3_heights[2489]), .rectangle3_weight(rectangle3_weights[2489]), .feature_threshold(feature_thresholds[2489]), .feature_above(feature_aboves[2489]), .feature_below(feature_belows[2489]), .scan_win_std_dev(scan_win_std_dev[2489]), .feature_accum(feature_accums[2489]));
  accum_calculator ac2490(.scan_win(scan_win2490), .rectangle1_x(rectangle1_xs[2490]), .rectangle1_y(rectangle1_ys[2490]), .rectangle1_width(rectangle1_widths[2490]), .rectangle1_height(rectangle1_heights[2490]), .rectangle1_weight(rectangle1_weights[2490]), .rectangle2_x(rectangle2_xs[2490]), .rectangle2_y(rectangle2_ys[2490]), .rectangle2_width(rectangle2_widths[2490]), .rectangle2_height(rectangle2_heights[2490]), .rectangle2_weight(rectangle2_weights[2490]), .rectangle3_x(rectangle3_xs[2490]), .rectangle3_y(rectangle3_ys[2490]), .rectangle3_width(rectangle3_widths[2490]), .rectangle3_height(rectangle3_heights[2490]), .rectangle3_weight(rectangle3_weights[2490]), .feature_threshold(feature_thresholds[2490]), .feature_above(feature_aboves[2490]), .feature_below(feature_belows[2490]), .scan_win_std_dev(scan_win_std_dev[2490]), .feature_accum(feature_accums[2490]));
  accum_calculator ac2491(.scan_win(scan_win2491), .rectangle1_x(rectangle1_xs[2491]), .rectangle1_y(rectangle1_ys[2491]), .rectangle1_width(rectangle1_widths[2491]), .rectangle1_height(rectangle1_heights[2491]), .rectangle1_weight(rectangle1_weights[2491]), .rectangle2_x(rectangle2_xs[2491]), .rectangle2_y(rectangle2_ys[2491]), .rectangle2_width(rectangle2_widths[2491]), .rectangle2_height(rectangle2_heights[2491]), .rectangle2_weight(rectangle2_weights[2491]), .rectangle3_x(rectangle3_xs[2491]), .rectangle3_y(rectangle3_ys[2491]), .rectangle3_width(rectangle3_widths[2491]), .rectangle3_height(rectangle3_heights[2491]), .rectangle3_weight(rectangle3_weights[2491]), .feature_threshold(feature_thresholds[2491]), .feature_above(feature_aboves[2491]), .feature_below(feature_belows[2491]), .scan_win_std_dev(scan_win_std_dev[2491]), .feature_accum(feature_accums[2491]));
  accum_calculator ac2492(.scan_win(scan_win2492), .rectangle1_x(rectangle1_xs[2492]), .rectangle1_y(rectangle1_ys[2492]), .rectangle1_width(rectangle1_widths[2492]), .rectangle1_height(rectangle1_heights[2492]), .rectangle1_weight(rectangle1_weights[2492]), .rectangle2_x(rectangle2_xs[2492]), .rectangle2_y(rectangle2_ys[2492]), .rectangle2_width(rectangle2_widths[2492]), .rectangle2_height(rectangle2_heights[2492]), .rectangle2_weight(rectangle2_weights[2492]), .rectangle3_x(rectangle3_xs[2492]), .rectangle3_y(rectangle3_ys[2492]), .rectangle3_width(rectangle3_widths[2492]), .rectangle3_height(rectangle3_heights[2492]), .rectangle3_weight(rectangle3_weights[2492]), .feature_threshold(feature_thresholds[2492]), .feature_above(feature_aboves[2492]), .feature_below(feature_belows[2492]), .scan_win_std_dev(scan_win_std_dev[2492]), .feature_accum(feature_accums[2492]));
  accum_calculator ac2493(.scan_win(scan_win2493), .rectangle1_x(rectangle1_xs[2493]), .rectangle1_y(rectangle1_ys[2493]), .rectangle1_width(rectangle1_widths[2493]), .rectangle1_height(rectangle1_heights[2493]), .rectangle1_weight(rectangle1_weights[2493]), .rectangle2_x(rectangle2_xs[2493]), .rectangle2_y(rectangle2_ys[2493]), .rectangle2_width(rectangle2_widths[2493]), .rectangle2_height(rectangle2_heights[2493]), .rectangle2_weight(rectangle2_weights[2493]), .rectangle3_x(rectangle3_xs[2493]), .rectangle3_y(rectangle3_ys[2493]), .rectangle3_width(rectangle3_widths[2493]), .rectangle3_height(rectangle3_heights[2493]), .rectangle3_weight(rectangle3_weights[2493]), .feature_threshold(feature_thresholds[2493]), .feature_above(feature_aboves[2493]), .feature_below(feature_belows[2493]), .scan_win_std_dev(scan_win_std_dev[2493]), .feature_accum(feature_accums[2493]));
  accum_calculator ac2494(.scan_win(scan_win2494), .rectangle1_x(rectangle1_xs[2494]), .rectangle1_y(rectangle1_ys[2494]), .rectangle1_width(rectangle1_widths[2494]), .rectangle1_height(rectangle1_heights[2494]), .rectangle1_weight(rectangle1_weights[2494]), .rectangle2_x(rectangle2_xs[2494]), .rectangle2_y(rectangle2_ys[2494]), .rectangle2_width(rectangle2_widths[2494]), .rectangle2_height(rectangle2_heights[2494]), .rectangle2_weight(rectangle2_weights[2494]), .rectangle3_x(rectangle3_xs[2494]), .rectangle3_y(rectangle3_ys[2494]), .rectangle3_width(rectangle3_widths[2494]), .rectangle3_height(rectangle3_heights[2494]), .rectangle3_weight(rectangle3_weights[2494]), .feature_threshold(feature_thresholds[2494]), .feature_above(feature_aboves[2494]), .feature_below(feature_belows[2494]), .scan_win_std_dev(scan_win_std_dev[2494]), .feature_accum(feature_accums[2494]));
  accum_calculator ac2495(.scan_win(scan_win2495), .rectangle1_x(rectangle1_xs[2495]), .rectangle1_y(rectangle1_ys[2495]), .rectangle1_width(rectangle1_widths[2495]), .rectangle1_height(rectangle1_heights[2495]), .rectangle1_weight(rectangle1_weights[2495]), .rectangle2_x(rectangle2_xs[2495]), .rectangle2_y(rectangle2_ys[2495]), .rectangle2_width(rectangle2_widths[2495]), .rectangle2_height(rectangle2_heights[2495]), .rectangle2_weight(rectangle2_weights[2495]), .rectangle3_x(rectangle3_xs[2495]), .rectangle3_y(rectangle3_ys[2495]), .rectangle3_width(rectangle3_widths[2495]), .rectangle3_height(rectangle3_heights[2495]), .rectangle3_weight(rectangle3_weights[2495]), .feature_threshold(feature_thresholds[2495]), .feature_above(feature_aboves[2495]), .feature_below(feature_belows[2495]), .scan_win_std_dev(scan_win_std_dev[2495]), .feature_accum(feature_accums[2495]));
  accum_calculator ac2496(.scan_win(scan_win2496), .rectangle1_x(rectangle1_xs[2496]), .rectangle1_y(rectangle1_ys[2496]), .rectangle1_width(rectangle1_widths[2496]), .rectangle1_height(rectangle1_heights[2496]), .rectangle1_weight(rectangle1_weights[2496]), .rectangle2_x(rectangle2_xs[2496]), .rectangle2_y(rectangle2_ys[2496]), .rectangle2_width(rectangle2_widths[2496]), .rectangle2_height(rectangle2_heights[2496]), .rectangle2_weight(rectangle2_weights[2496]), .rectangle3_x(rectangle3_xs[2496]), .rectangle3_y(rectangle3_ys[2496]), .rectangle3_width(rectangle3_widths[2496]), .rectangle3_height(rectangle3_heights[2496]), .rectangle3_weight(rectangle3_weights[2496]), .feature_threshold(feature_thresholds[2496]), .feature_above(feature_aboves[2496]), .feature_below(feature_belows[2496]), .scan_win_std_dev(scan_win_std_dev[2496]), .feature_accum(feature_accums[2496]));
  accum_calculator ac2497(.scan_win(scan_win2497), .rectangle1_x(rectangle1_xs[2497]), .rectangle1_y(rectangle1_ys[2497]), .rectangle1_width(rectangle1_widths[2497]), .rectangle1_height(rectangle1_heights[2497]), .rectangle1_weight(rectangle1_weights[2497]), .rectangle2_x(rectangle2_xs[2497]), .rectangle2_y(rectangle2_ys[2497]), .rectangle2_width(rectangle2_widths[2497]), .rectangle2_height(rectangle2_heights[2497]), .rectangle2_weight(rectangle2_weights[2497]), .rectangle3_x(rectangle3_xs[2497]), .rectangle3_y(rectangle3_ys[2497]), .rectangle3_width(rectangle3_widths[2497]), .rectangle3_height(rectangle3_heights[2497]), .rectangle3_weight(rectangle3_weights[2497]), .feature_threshold(feature_thresholds[2497]), .feature_above(feature_aboves[2497]), .feature_below(feature_belows[2497]), .scan_win_std_dev(scan_win_std_dev[2497]), .feature_accum(feature_accums[2497]));
  accum_calculator ac2498(.scan_win(scan_win2498), .rectangle1_x(rectangle1_xs[2498]), .rectangle1_y(rectangle1_ys[2498]), .rectangle1_width(rectangle1_widths[2498]), .rectangle1_height(rectangle1_heights[2498]), .rectangle1_weight(rectangle1_weights[2498]), .rectangle2_x(rectangle2_xs[2498]), .rectangle2_y(rectangle2_ys[2498]), .rectangle2_width(rectangle2_widths[2498]), .rectangle2_height(rectangle2_heights[2498]), .rectangle2_weight(rectangle2_weights[2498]), .rectangle3_x(rectangle3_xs[2498]), .rectangle3_y(rectangle3_ys[2498]), .rectangle3_width(rectangle3_widths[2498]), .rectangle3_height(rectangle3_heights[2498]), .rectangle3_weight(rectangle3_weights[2498]), .feature_threshold(feature_thresholds[2498]), .feature_above(feature_aboves[2498]), .feature_below(feature_belows[2498]), .scan_win_std_dev(scan_win_std_dev[2498]), .feature_accum(feature_accums[2498]));
  accum_calculator ac2499(.scan_win(scan_win2499), .rectangle1_x(rectangle1_xs[2499]), .rectangle1_y(rectangle1_ys[2499]), .rectangle1_width(rectangle1_widths[2499]), .rectangle1_height(rectangle1_heights[2499]), .rectangle1_weight(rectangle1_weights[2499]), .rectangle2_x(rectangle2_xs[2499]), .rectangle2_y(rectangle2_ys[2499]), .rectangle2_width(rectangle2_widths[2499]), .rectangle2_height(rectangle2_heights[2499]), .rectangle2_weight(rectangle2_weights[2499]), .rectangle3_x(rectangle3_xs[2499]), .rectangle3_y(rectangle3_ys[2499]), .rectangle3_width(rectangle3_widths[2499]), .rectangle3_height(rectangle3_heights[2499]), .rectangle3_weight(rectangle3_weights[2499]), .feature_threshold(feature_thresholds[2499]), .feature_above(feature_aboves[2499]), .feature_below(feature_belows[2499]), .scan_win_std_dev(scan_win_std_dev[2499]), .feature_accum(feature_accums[2499]));
  accum_calculator ac2500(.scan_win(scan_win2500), .rectangle1_x(rectangle1_xs[2500]), .rectangle1_y(rectangle1_ys[2500]), .rectangle1_width(rectangle1_widths[2500]), .rectangle1_height(rectangle1_heights[2500]), .rectangle1_weight(rectangle1_weights[2500]), .rectangle2_x(rectangle2_xs[2500]), .rectangle2_y(rectangle2_ys[2500]), .rectangle2_width(rectangle2_widths[2500]), .rectangle2_height(rectangle2_heights[2500]), .rectangle2_weight(rectangle2_weights[2500]), .rectangle3_x(rectangle3_xs[2500]), .rectangle3_y(rectangle3_ys[2500]), .rectangle3_width(rectangle3_widths[2500]), .rectangle3_height(rectangle3_heights[2500]), .rectangle3_weight(rectangle3_weights[2500]), .feature_threshold(feature_thresholds[2500]), .feature_above(feature_aboves[2500]), .feature_below(feature_belows[2500]), .scan_win_std_dev(scan_win_std_dev[2500]), .feature_accum(feature_accums[2500]));
  accum_calculator ac2501(.scan_win(scan_win2501), .rectangle1_x(rectangle1_xs[2501]), .rectangle1_y(rectangle1_ys[2501]), .rectangle1_width(rectangle1_widths[2501]), .rectangle1_height(rectangle1_heights[2501]), .rectangle1_weight(rectangle1_weights[2501]), .rectangle2_x(rectangle2_xs[2501]), .rectangle2_y(rectangle2_ys[2501]), .rectangle2_width(rectangle2_widths[2501]), .rectangle2_height(rectangle2_heights[2501]), .rectangle2_weight(rectangle2_weights[2501]), .rectangle3_x(rectangle3_xs[2501]), .rectangle3_y(rectangle3_ys[2501]), .rectangle3_width(rectangle3_widths[2501]), .rectangle3_height(rectangle3_heights[2501]), .rectangle3_weight(rectangle3_weights[2501]), .feature_threshold(feature_thresholds[2501]), .feature_above(feature_aboves[2501]), .feature_below(feature_belows[2501]), .scan_win_std_dev(scan_win_std_dev[2501]), .feature_accum(feature_accums[2501]));
  accum_calculator ac2502(.scan_win(scan_win2502), .rectangle1_x(rectangle1_xs[2502]), .rectangle1_y(rectangle1_ys[2502]), .rectangle1_width(rectangle1_widths[2502]), .rectangle1_height(rectangle1_heights[2502]), .rectangle1_weight(rectangle1_weights[2502]), .rectangle2_x(rectangle2_xs[2502]), .rectangle2_y(rectangle2_ys[2502]), .rectangle2_width(rectangle2_widths[2502]), .rectangle2_height(rectangle2_heights[2502]), .rectangle2_weight(rectangle2_weights[2502]), .rectangle3_x(rectangle3_xs[2502]), .rectangle3_y(rectangle3_ys[2502]), .rectangle3_width(rectangle3_widths[2502]), .rectangle3_height(rectangle3_heights[2502]), .rectangle3_weight(rectangle3_weights[2502]), .feature_threshold(feature_thresholds[2502]), .feature_above(feature_aboves[2502]), .feature_below(feature_belows[2502]), .scan_win_std_dev(scan_win_std_dev[2502]), .feature_accum(feature_accums[2502]));
  accum_calculator ac2503(.scan_win(scan_win2503), .rectangle1_x(rectangle1_xs[2503]), .rectangle1_y(rectangle1_ys[2503]), .rectangle1_width(rectangle1_widths[2503]), .rectangle1_height(rectangle1_heights[2503]), .rectangle1_weight(rectangle1_weights[2503]), .rectangle2_x(rectangle2_xs[2503]), .rectangle2_y(rectangle2_ys[2503]), .rectangle2_width(rectangle2_widths[2503]), .rectangle2_height(rectangle2_heights[2503]), .rectangle2_weight(rectangle2_weights[2503]), .rectangle3_x(rectangle3_xs[2503]), .rectangle3_y(rectangle3_ys[2503]), .rectangle3_width(rectangle3_widths[2503]), .rectangle3_height(rectangle3_heights[2503]), .rectangle3_weight(rectangle3_weights[2503]), .feature_threshold(feature_thresholds[2503]), .feature_above(feature_aboves[2503]), .feature_below(feature_belows[2503]), .scan_win_std_dev(scan_win_std_dev[2503]), .feature_accum(feature_accums[2503]));
  accum_calculator ac2504(.scan_win(scan_win2504), .rectangle1_x(rectangle1_xs[2504]), .rectangle1_y(rectangle1_ys[2504]), .rectangle1_width(rectangle1_widths[2504]), .rectangle1_height(rectangle1_heights[2504]), .rectangle1_weight(rectangle1_weights[2504]), .rectangle2_x(rectangle2_xs[2504]), .rectangle2_y(rectangle2_ys[2504]), .rectangle2_width(rectangle2_widths[2504]), .rectangle2_height(rectangle2_heights[2504]), .rectangle2_weight(rectangle2_weights[2504]), .rectangle3_x(rectangle3_xs[2504]), .rectangle3_y(rectangle3_ys[2504]), .rectangle3_width(rectangle3_widths[2504]), .rectangle3_height(rectangle3_heights[2504]), .rectangle3_weight(rectangle3_weights[2504]), .feature_threshold(feature_thresholds[2504]), .feature_above(feature_aboves[2504]), .feature_below(feature_belows[2504]), .scan_win_std_dev(scan_win_std_dev[2504]), .feature_accum(feature_accums[2504]));
  accum_calculator ac2505(.scan_win(scan_win2505), .rectangle1_x(rectangle1_xs[2505]), .rectangle1_y(rectangle1_ys[2505]), .rectangle1_width(rectangle1_widths[2505]), .rectangle1_height(rectangle1_heights[2505]), .rectangle1_weight(rectangle1_weights[2505]), .rectangle2_x(rectangle2_xs[2505]), .rectangle2_y(rectangle2_ys[2505]), .rectangle2_width(rectangle2_widths[2505]), .rectangle2_height(rectangle2_heights[2505]), .rectangle2_weight(rectangle2_weights[2505]), .rectangle3_x(rectangle3_xs[2505]), .rectangle3_y(rectangle3_ys[2505]), .rectangle3_width(rectangle3_widths[2505]), .rectangle3_height(rectangle3_heights[2505]), .rectangle3_weight(rectangle3_weights[2505]), .feature_threshold(feature_thresholds[2505]), .feature_above(feature_aboves[2505]), .feature_below(feature_belows[2505]), .scan_win_std_dev(scan_win_std_dev[2505]), .feature_accum(feature_accums[2505]));
  accum_calculator ac2506(.scan_win(scan_win2506), .rectangle1_x(rectangle1_xs[2506]), .rectangle1_y(rectangle1_ys[2506]), .rectangle1_width(rectangle1_widths[2506]), .rectangle1_height(rectangle1_heights[2506]), .rectangle1_weight(rectangle1_weights[2506]), .rectangle2_x(rectangle2_xs[2506]), .rectangle2_y(rectangle2_ys[2506]), .rectangle2_width(rectangle2_widths[2506]), .rectangle2_height(rectangle2_heights[2506]), .rectangle2_weight(rectangle2_weights[2506]), .rectangle3_x(rectangle3_xs[2506]), .rectangle3_y(rectangle3_ys[2506]), .rectangle3_width(rectangle3_widths[2506]), .rectangle3_height(rectangle3_heights[2506]), .rectangle3_weight(rectangle3_weights[2506]), .feature_threshold(feature_thresholds[2506]), .feature_above(feature_aboves[2506]), .feature_below(feature_belows[2506]), .scan_win_std_dev(scan_win_std_dev[2506]), .feature_accum(feature_accums[2506]));
  accum_calculator ac2507(.scan_win(scan_win2507), .rectangle1_x(rectangle1_xs[2507]), .rectangle1_y(rectangle1_ys[2507]), .rectangle1_width(rectangle1_widths[2507]), .rectangle1_height(rectangle1_heights[2507]), .rectangle1_weight(rectangle1_weights[2507]), .rectangle2_x(rectangle2_xs[2507]), .rectangle2_y(rectangle2_ys[2507]), .rectangle2_width(rectangle2_widths[2507]), .rectangle2_height(rectangle2_heights[2507]), .rectangle2_weight(rectangle2_weights[2507]), .rectangle3_x(rectangle3_xs[2507]), .rectangle3_y(rectangle3_ys[2507]), .rectangle3_width(rectangle3_widths[2507]), .rectangle3_height(rectangle3_heights[2507]), .rectangle3_weight(rectangle3_weights[2507]), .feature_threshold(feature_thresholds[2507]), .feature_above(feature_aboves[2507]), .feature_below(feature_belows[2507]), .scan_win_std_dev(scan_win_std_dev[2507]), .feature_accum(feature_accums[2507]));
  accum_calculator ac2508(.scan_win(scan_win2508), .rectangle1_x(rectangle1_xs[2508]), .rectangle1_y(rectangle1_ys[2508]), .rectangle1_width(rectangle1_widths[2508]), .rectangle1_height(rectangle1_heights[2508]), .rectangle1_weight(rectangle1_weights[2508]), .rectangle2_x(rectangle2_xs[2508]), .rectangle2_y(rectangle2_ys[2508]), .rectangle2_width(rectangle2_widths[2508]), .rectangle2_height(rectangle2_heights[2508]), .rectangle2_weight(rectangle2_weights[2508]), .rectangle3_x(rectangle3_xs[2508]), .rectangle3_y(rectangle3_ys[2508]), .rectangle3_width(rectangle3_widths[2508]), .rectangle3_height(rectangle3_heights[2508]), .rectangle3_weight(rectangle3_weights[2508]), .feature_threshold(feature_thresholds[2508]), .feature_above(feature_aboves[2508]), .feature_below(feature_belows[2508]), .scan_win_std_dev(scan_win_std_dev[2508]), .feature_accum(feature_accums[2508]));
  accum_calculator ac2509(.scan_win(scan_win2509), .rectangle1_x(rectangle1_xs[2509]), .rectangle1_y(rectangle1_ys[2509]), .rectangle1_width(rectangle1_widths[2509]), .rectangle1_height(rectangle1_heights[2509]), .rectangle1_weight(rectangle1_weights[2509]), .rectangle2_x(rectangle2_xs[2509]), .rectangle2_y(rectangle2_ys[2509]), .rectangle2_width(rectangle2_widths[2509]), .rectangle2_height(rectangle2_heights[2509]), .rectangle2_weight(rectangle2_weights[2509]), .rectangle3_x(rectangle3_xs[2509]), .rectangle3_y(rectangle3_ys[2509]), .rectangle3_width(rectangle3_widths[2509]), .rectangle3_height(rectangle3_heights[2509]), .rectangle3_weight(rectangle3_weights[2509]), .feature_threshold(feature_thresholds[2509]), .feature_above(feature_aboves[2509]), .feature_below(feature_belows[2509]), .scan_win_std_dev(scan_win_std_dev[2509]), .feature_accum(feature_accums[2509]));
  accum_calculator ac2510(.scan_win(scan_win2510), .rectangle1_x(rectangle1_xs[2510]), .rectangle1_y(rectangle1_ys[2510]), .rectangle1_width(rectangle1_widths[2510]), .rectangle1_height(rectangle1_heights[2510]), .rectangle1_weight(rectangle1_weights[2510]), .rectangle2_x(rectangle2_xs[2510]), .rectangle2_y(rectangle2_ys[2510]), .rectangle2_width(rectangle2_widths[2510]), .rectangle2_height(rectangle2_heights[2510]), .rectangle2_weight(rectangle2_weights[2510]), .rectangle3_x(rectangle3_xs[2510]), .rectangle3_y(rectangle3_ys[2510]), .rectangle3_width(rectangle3_widths[2510]), .rectangle3_height(rectangle3_heights[2510]), .rectangle3_weight(rectangle3_weights[2510]), .feature_threshold(feature_thresholds[2510]), .feature_above(feature_aboves[2510]), .feature_below(feature_belows[2510]), .scan_win_std_dev(scan_win_std_dev[2510]), .feature_accum(feature_accums[2510]));
  accum_calculator ac2511(.scan_win(scan_win2511), .rectangle1_x(rectangle1_xs[2511]), .rectangle1_y(rectangle1_ys[2511]), .rectangle1_width(rectangle1_widths[2511]), .rectangle1_height(rectangle1_heights[2511]), .rectangle1_weight(rectangle1_weights[2511]), .rectangle2_x(rectangle2_xs[2511]), .rectangle2_y(rectangle2_ys[2511]), .rectangle2_width(rectangle2_widths[2511]), .rectangle2_height(rectangle2_heights[2511]), .rectangle2_weight(rectangle2_weights[2511]), .rectangle3_x(rectangle3_xs[2511]), .rectangle3_y(rectangle3_ys[2511]), .rectangle3_width(rectangle3_widths[2511]), .rectangle3_height(rectangle3_heights[2511]), .rectangle3_weight(rectangle3_weights[2511]), .feature_threshold(feature_thresholds[2511]), .feature_above(feature_aboves[2511]), .feature_below(feature_belows[2511]), .scan_win_std_dev(scan_win_std_dev[2511]), .feature_accum(feature_accums[2511]));
  accum_calculator ac2512(.scan_win(scan_win2512), .rectangle1_x(rectangle1_xs[2512]), .rectangle1_y(rectangle1_ys[2512]), .rectangle1_width(rectangle1_widths[2512]), .rectangle1_height(rectangle1_heights[2512]), .rectangle1_weight(rectangle1_weights[2512]), .rectangle2_x(rectangle2_xs[2512]), .rectangle2_y(rectangle2_ys[2512]), .rectangle2_width(rectangle2_widths[2512]), .rectangle2_height(rectangle2_heights[2512]), .rectangle2_weight(rectangle2_weights[2512]), .rectangle3_x(rectangle3_xs[2512]), .rectangle3_y(rectangle3_ys[2512]), .rectangle3_width(rectangle3_widths[2512]), .rectangle3_height(rectangle3_heights[2512]), .rectangle3_weight(rectangle3_weights[2512]), .feature_threshold(feature_thresholds[2512]), .feature_above(feature_aboves[2512]), .feature_below(feature_belows[2512]), .scan_win_std_dev(scan_win_std_dev[2512]), .feature_accum(feature_accums[2512]));
  accum_calculator ac2513(.scan_win(scan_win2513), .rectangle1_x(rectangle1_xs[2513]), .rectangle1_y(rectangle1_ys[2513]), .rectangle1_width(rectangle1_widths[2513]), .rectangle1_height(rectangle1_heights[2513]), .rectangle1_weight(rectangle1_weights[2513]), .rectangle2_x(rectangle2_xs[2513]), .rectangle2_y(rectangle2_ys[2513]), .rectangle2_width(rectangle2_widths[2513]), .rectangle2_height(rectangle2_heights[2513]), .rectangle2_weight(rectangle2_weights[2513]), .rectangle3_x(rectangle3_xs[2513]), .rectangle3_y(rectangle3_ys[2513]), .rectangle3_width(rectangle3_widths[2513]), .rectangle3_height(rectangle3_heights[2513]), .rectangle3_weight(rectangle3_weights[2513]), .feature_threshold(feature_thresholds[2513]), .feature_above(feature_aboves[2513]), .feature_below(feature_belows[2513]), .scan_win_std_dev(scan_win_std_dev[2513]), .feature_accum(feature_accums[2513]));
  accum_calculator ac2514(.scan_win(scan_win2514), .rectangle1_x(rectangle1_xs[2514]), .rectangle1_y(rectangle1_ys[2514]), .rectangle1_width(rectangle1_widths[2514]), .rectangle1_height(rectangle1_heights[2514]), .rectangle1_weight(rectangle1_weights[2514]), .rectangle2_x(rectangle2_xs[2514]), .rectangle2_y(rectangle2_ys[2514]), .rectangle2_width(rectangle2_widths[2514]), .rectangle2_height(rectangle2_heights[2514]), .rectangle2_weight(rectangle2_weights[2514]), .rectangle3_x(rectangle3_xs[2514]), .rectangle3_y(rectangle3_ys[2514]), .rectangle3_width(rectangle3_widths[2514]), .rectangle3_height(rectangle3_heights[2514]), .rectangle3_weight(rectangle3_weights[2514]), .feature_threshold(feature_thresholds[2514]), .feature_above(feature_aboves[2514]), .feature_below(feature_belows[2514]), .scan_win_std_dev(scan_win_std_dev[2514]), .feature_accum(feature_accums[2514]));
  accum_calculator ac2515(.scan_win(scan_win2515), .rectangle1_x(rectangle1_xs[2515]), .rectangle1_y(rectangle1_ys[2515]), .rectangle1_width(rectangle1_widths[2515]), .rectangle1_height(rectangle1_heights[2515]), .rectangle1_weight(rectangle1_weights[2515]), .rectangle2_x(rectangle2_xs[2515]), .rectangle2_y(rectangle2_ys[2515]), .rectangle2_width(rectangle2_widths[2515]), .rectangle2_height(rectangle2_heights[2515]), .rectangle2_weight(rectangle2_weights[2515]), .rectangle3_x(rectangle3_xs[2515]), .rectangle3_y(rectangle3_ys[2515]), .rectangle3_width(rectangle3_widths[2515]), .rectangle3_height(rectangle3_heights[2515]), .rectangle3_weight(rectangle3_weights[2515]), .feature_threshold(feature_thresholds[2515]), .feature_above(feature_aboves[2515]), .feature_below(feature_belows[2515]), .scan_win_std_dev(scan_win_std_dev[2515]), .feature_accum(feature_accums[2515]));
  accum_calculator ac2516(.scan_win(scan_win2516), .rectangle1_x(rectangle1_xs[2516]), .rectangle1_y(rectangle1_ys[2516]), .rectangle1_width(rectangle1_widths[2516]), .rectangle1_height(rectangle1_heights[2516]), .rectangle1_weight(rectangle1_weights[2516]), .rectangle2_x(rectangle2_xs[2516]), .rectangle2_y(rectangle2_ys[2516]), .rectangle2_width(rectangle2_widths[2516]), .rectangle2_height(rectangle2_heights[2516]), .rectangle2_weight(rectangle2_weights[2516]), .rectangle3_x(rectangle3_xs[2516]), .rectangle3_y(rectangle3_ys[2516]), .rectangle3_width(rectangle3_widths[2516]), .rectangle3_height(rectangle3_heights[2516]), .rectangle3_weight(rectangle3_weights[2516]), .feature_threshold(feature_thresholds[2516]), .feature_above(feature_aboves[2516]), .feature_below(feature_belows[2516]), .scan_win_std_dev(scan_win_std_dev[2516]), .feature_accum(feature_accums[2516]));
  accum_calculator ac2517(.scan_win(scan_win2517), .rectangle1_x(rectangle1_xs[2517]), .rectangle1_y(rectangle1_ys[2517]), .rectangle1_width(rectangle1_widths[2517]), .rectangle1_height(rectangle1_heights[2517]), .rectangle1_weight(rectangle1_weights[2517]), .rectangle2_x(rectangle2_xs[2517]), .rectangle2_y(rectangle2_ys[2517]), .rectangle2_width(rectangle2_widths[2517]), .rectangle2_height(rectangle2_heights[2517]), .rectangle2_weight(rectangle2_weights[2517]), .rectangle3_x(rectangle3_xs[2517]), .rectangle3_y(rectangle3_ys[2517]), .rectangle3_width(rectangle3_widths[2517]), .rectangle3_height(rectangle3_heights[2517]), .rectangle3_weight(rectangle3_weights[2517]), .feature_threshold(feature_thresholds[2517]), .feature_above(feature_aboves[2517]), .feature_below(feature_belows[2517]), .scan_win_std_dev(scan_win_std_dev[2517]), .feature_accum(feature_accums[2517]));
  accum_calculator ac2518(.scan_win(scan_win2518), .rectangle1_x(rectangle1_xs[2518]), .rectangle1_y(rectangle1_ys[2518]), .rectangle1_width(rectangle1_widths[2518]), .rectangle1_height(rectangle1_heights[2518]), .rectangle1_weight(rectangle1_weights[2518]), .rectangle2_x(rectangle2_xs[2518]), .rectangle2_y(rectangle2_ys[2518]), .rectangle2_width(rectangle2_widths[2518]), .rectangle2_height(rectangle2_heights[2518]), .rectangle2_weight(rectangle2_weights[2518]), .rectangle3_x(rectangle3_xs[2518]), .rectangle3_y(rectangle3_ys[2518]), .rectangle3_width(rectangle3_widths[2518]), .rectangle3_height(rectangle3_heights[2518]), .rectangle3_weight(rectangle3_weights[2518]), .feature_threshold(feature_thresholds[2518]), .feature_above(feature_aboves[2518]), .feature_below(feature_belows[2518]), .scan_win_std_dev(scan_win_std_dev[2518]), .feature_accum(feature_accums[2518]));
  accum_calculator ac2519(.scan_win(scan_win2519), .rectangle1_x(rectangle1_xs[2519]), .rectangle1_y(rectangle1_ys[2519]), .rectangle1_width(rectangle1_widths[2519]), .rectangle1_height(rectangle1_heights[2519]), .rectangle1_weight(rectangle1_weights[2519]), .rectangle2_x(rectangle2_xs[2519]), .rectangle2_y(rectangle2_ys[2519]), .rectangle2_width(rectangle2_widths[2519]), .rectangle2_height(rectangle2_heights[2519]), .rectangle2_weight(rectangle2_weights[2519]), .rectangle3_x(rectangle3_xs[2519]), .rectangle3_y(rectangle3_ys[2519]), .rectangle3_width(rectangle3_widths[2519]), .rectangle3_height(rectangle3_heights[2519]), .rectangle3_weight(rectangle3_weights[2519]), .feature_threshold(feature_thresholds[2519]), .feature_above(feature_aboves[2519]), .feature_below(feature_belows[2519]), .scan_win_std_dev(scan_win_std_dev[2519]), .feature_accum(feature_accums[2519]));
  accum_calculator ac2520(.scan_win(scan_win2520), .rectangle1_x(rectangle1_xs[2520]), .rectangle1_y(rectangle1_ys[2520]), .rectangle1_width(rectangle1_widths[2520]), .rectangle1_height(rectangle1_heights[2520]), .rectangle1_weight(rectangle1_weights[2520]), .rectangle2_x(rectangle2_xs[2520]), .rectangle2_y(rectangle2_ys[2520]), .rectangle2_width(rectangle2_widths[2520]), .rectangle2_height(rectangle2_heights[2520]), .rectangle2_weight(rectangle2_weights[2520]), .rectangle3_x(rectangle3_xs[2520]), .rectangle3_y(rectangle3_ys[2520]), .rectangle3_width(rectangle3_widths[2520]), .rectangle3_height(rectangle3_heights[2520]), .rectangle3_weight(rectangle3_weights[2520]), .feature_threshold(feature_thresholds[2520]), .feature_above(feature_aboves[2520]), .feature_below(feature_belows[2520]), .scan_win_std_dev(scan_win_std_dev[2520]), .feature_accum(feature_accums[2520]));
  accum_calculator ac2521(.scan_win(scan_win2521), .rectangle1_x(rectangle1_xs[2521]), .rectangle1_y(rectangle1_ys[2521]), .rectangle1_width(rectangle1_widths[2521]), .rectangle1_height(rectangle1_heights[2521]), .rectangle1_weight(rectangle1_weights[2521]), .rectangle2_x(rectangle2_xs[2521]), .rectangle2_y(rectangle2_ys[2521]), .rectangle2_width(rectangle2_widths[2521]), .rectangle2_height(rectangle2_heights[2521]), .rectangle2_weight(rectangle2_weights[2521]), .rectangle3_x(rectangle3_xs[2521]), .rectangle3_y(rectangle3_ys[2521]), .rectangle3_width(rectangle3_widths[2521]), .rectangle3_height(rectangle3_heights[2521]), .rectangle3_weight(rectangle3_weights[2521]), .feature_threshold(feature_thresholds[2521]), .feature_above(feature_aboves[2521]), .feature_below(feature_belows[2521]), .scan_win_std_dev(scan_win_std_dev[2521]), .feature_accum(feature_accums[2521]));
  accum_calculator ac2522(.scan_win(scan_win2522), .rectangle1_x(rectangle1_xs[2522]), .rectangle1_y(rectangle1_ys[2522]), .rectangle1_width(rectangle1_widths[2522]), .rectangle1_height(rectangle1_heights[2522]), .rectangle1_weight(rectangle1_weights[2522]), .rectangle2_x(rectangle2_xs[2522]), .rectangle2_y(rectangle2_ys[2522]), .rectangle2_width(rectangle2_widths[2522]), .rectangle2_height(rectangle2_heights[2522]), .rectangle2_weight(rectangle2_weights[2522]), .rectangle3_x(rectangle3_xs[2522]), .rectangle3_y(rectangle3_ys[2522]), .rectangle3_width(rectangle3_widths[2522]), .rectangle3_height(rectangle3_heights[2522]), .rectangle3_weight(rectangle3_weights[2522]), .feature_threshold(feature_thresholds[2522]), .feature_above(feature_aboves[2522]), .feature_below(feature_belows[2522]), .scan_win_std_dev(scan_win_std_dev[2522]), .feature_accum(feature_accums[2522]));
  accum_calculator ac2523(.scan_win(scan_win2523), .rectangle1_x(rectangle1_xs[2523]), .rectangle1_y(rectangle1_ys[2523]), .rectangle1_width(rectangle1_widths[2523]), .rectangle1_height(rectangle1_heights[2523]), .rectangle1_weight(rectangle1_weights[2523]), .rectangle2_x(rectangle2_xs[2523]), .rectangle2_y(rectangle2_ys[2523]), .rectangle2_width(rectangle2_widths[2523]), .rectangle2_height(rectangle2_heights[2523]), .rectangle2_weight(rectangle2_weights[2523]), .rectangle3_x(rectangle3_xs[2523]), .rectangle3_y(rectangle3_ys[2523]), .rectangle3_width(rectangle3_widths[2523]), .rectangle3_height(rectangle3_heights[2523]), .rectangle3_weight(rectangle3_weights[2523]), .feature_threshold(feature_thresholds[2523]), .feature_above(feature_aboves[2523]), .feature_below(feature_belows[2523]), .scan_win_std_dev(scan_win_std_dev[2523]), .feature_accum(feature_accums[2523]));
  accum_calculator ac2524(.scan_win(scan_win2524), .rectangle1_x(rectangle1_xs[2524]), .rectangle1_y(rectangle1_ys[2524]), .rectangle1_width(rectangle1_widths[2524]), .rectangle1_height(rectangle1_heights[2524]), .rectangle1_weight(rectangle1_weights[2524]), .rectangle2_x(rectangle2_xs[2524]), .rectangle2_y(rectangle2_ys[2524]), .rectangle2_width(rectangle2_widths[2524]), .rectangle2_height(rectangle2_heights[2524]), .rectangle2_weight(rectangle2_weights[2524]), .rectangle3_x(rectangle3_xs[2524]), .rectangle3_y(rectangle3_ys[2524]), .rectangle3_width(rectangle3_widths[2524]), .rectangle3_height(rectangle3_heights[2524]), .rectangle3_weight(rectangle3_weights[2524]), .feature_threshold(feature_thresholds[2524]), .feature_above(feature_aboves[2524]), .feature_below(feature_belows[2524]), .scan_win_std_dev(scan_win_std_dev[2524]), .feature_accum(feature_accums[2524]));
  accum_calculator ac2525(.scan_win(scan_win2525), .rectangle1_x(rectangle1_xs[2525]), .rectangle1_y(rectangle1_ys[2525]), .rectangle1_width(rectangle1_widths[2525]), .rectangle1_height(rectangle1_heights[2525]), .rectangle1_weight(rectangle1_weights[2525]), .rectangle2_x(rectangle2_xs[2525]), .rectangle2_y(rectangle2_ys[2525]), .rectangle2_width(rectangle2_widths[2525]), .rectangle2_height(rectangle2_heights[2525]), .rectangle2_weight(rectangle2_weights[2525]), .rectangle3_x(rectangle3_xs[2525]), .rectangle3_y(rectangle3_ys[2525]), .rectangle3_width(rectangle3_widths[2525]), .rectangle3_height(rectangle3_heights[2525]), .rectangle3_weight(rectangle3_weights[2525]), .feature_threshold(feature_thresholds[2525]), .feature_above(feature_aboves[2525]), .feature_below(feature_belows[2525]), .scan_win_std_dev(scan_win_std_dev[2525]), .feature_accum(feature_accums[2525]));
  accum_calculator ac2526(.scan_win(scan_win2526), .rectangle1_x(rectangle1_xs[2526]), .rectangle1_y(rectangle1_ys[2526]), .rectangle1_width(rectangle1_widths[2526]), .rectangle1_height(rectangle1_heights[2526]), .rectangle1_weight(rectangle1_weights[2526]), .rectangle2_x(rectangle2_xs[2526]), .rectangle2_y(rectangle2_ys[2526]), .rectangle2_width(rectangle2_widths[2526]), .rectangle2_height(rectangle2_heights[2526]), .rectangle2_weight(rectangle2_weights[2526]), .rectangle3_x(rectangle3_xs[2526]), .rectangle3_y(rectangle3_ys[2526]), .rectangle3_width(rectangle3_widths[2526]), .rectangle3_height(rectangle3_heights[2526]), .rectangle3_weight(rectangle3_weights[2526]), .feature_threshold(feature_thresholds[2526]), .feature_above(feature_aboves[2526]), .feature_below(feature_belows[2526]), .scan_win_std_dev(scan_win_std_dev[2526]), .feature_accum(feature_accums[2526]));
  accum_calculator ac2527(.scan_win(scan_win2527), .rectangle1_x(rectangle1_xs[2527]), .rectangle1_y(rectangle1_ys[2527]), .rectangle1_width(rectangle1_widths[2527]), .rectangle1_height(rectangle1_heights[2527]), .rectangle1_weight(rectangle1_weights[2527]), .rectangle2_x(rectangle2_xs[2527]), .rectangle2_y(rectangle2_ys[2527]), .rectangle2_width(rectangle2_widths[2527]), .rectangle2_height(rectangle2_heights[2527]), .rectangle2_weight(rectangle2_weights[2527]), .rectangle3_x(rectangle3_xs[2527]), .rectangle3_y(rectangle3_ys[2527]), .rectangle3_width(rectangle3_widths[2527]), .rectangle3_height(rectangle3_heights[2527]), .rectangle3_weight(rectangle3_weights[2527]), .feature_threshold(feature_thresholds[2527]), .feature_above(feature_aboves[2527]), .feature_below(feature_belows[2527]), .scan_win_std_dev(scan_win_std_dev[2527]), .feature_accum(feature_accums[2527]));
  accum_calculator ac2528(.scan_win(scan_win2528), .rectangle1_x(rectangle1_xs[2528]), .rectangle1_y(rectangle1_ys[2528]), .rectangle1_width(rectangle1_widths[2528]), .rectangle1_height(rectangle1_heights[2528]), .rectangle1_weight(rectangle1_weights[2528]), .rectangle2_x(rectangle2_xs[2528]), .rectangle2_y(rectangle2_ys[2528]), .rectangle2_width(rectangle2_widths[2528]), .rectangle2_height(rectangle2_heights[2528]), .rectangle2_weight(rectangle2_weights[2528]), .rectangle3_x(rectangle3_xs[2528]), .rectangle3_y(rectangle3_ys[2528]), .rectangle3_width(rectangle3_widths[2528]), .rectangle3_height(rectangle3_heights[2528]), .rectangle3_weight(rectangle3_weights[2528]), .feature_threshold(feature_thresholds[2528]), .feature_above(feature_aboves[2528]), .feature_below(feature_belows[2528]), .scan_win_std_dev(scan_win_std_dev[2528]), .feature_accum(feature_accums[2528]));
  accum_calculator ac2529(.scan_win(scan_win2529), .rectangle1_x(rectangle1_xs[2529]), .rectangle1_y(rectangle1_ys[2529]), .rectangle1_width(rectangle1_widths[2529]), .rectangle1_height(rectangle1_heights[2529]), .rectangle1_weight(rectangle1_weights[2529]), .rectangle2_x(rectangle2_xs[2529]), .rectangle2_y(rectangle2_ys[2529]), .rectangle2_width(rectangle2_widths[2529]), .rectangle2_height(rectangle2_heights[2529]), .rectangle2_weight(rectangle2_weights[2529]), .rectangle3_x(rectangle3_xs[2529]), .rectangle3_y(rectangle3_ys[2529]), .rectangle3_width(rectangle3_widths[2529]), .rectangle3_height(rectangle3_heights[2529]), .rectangle3_weight(rectangle3_weights[2529]), .feature_threshold(feature_thresholds[2529]), .feature_above(feature_aboves[2529]), .feature_below(feature_belows[2529]), .scan_win_std_dev(scan_win_std_dev[2529]), .feature_accum(feature_accums[2529]));
  accum_calculator ac2530(.scan_win(scan_win2530), .rectangle1_x(rectangle1_xs[2530]), .rectangle1_y(rectangle1_ys[2530]), .rectangle1_width(rectangle1_widths[2530]), .rectangle1_height(rectangle1_heights[2530]), .rectangle1_weight(rectangle1_weights[2530]), .rectangle2_x(rectangle2_xs[2530]), .rectangle2_y(rectangle2_ys[2530]), .rectangle2_width(rectangle2_widths[2530]), .rectangle2_height(rectangle2_heights[2530]), .rectangle2_weight(rectangle2_weights[2530]), .rectangle3_x(rectangle3_xs[2530]), .rectangle3_y(rectangle3_ys[2530]), .rectangle3_width(rectangle3_widths[2530]), .rectangle3_height(rectangle3_heights[2530]), .rectangle3_weight(rectangle3_weights[2530]), .feature_threshold(feature_thresholds[2530]), .feature_above(feature_aboves[2530]), .feature_below(feature_belows[2530]), .scan_win_std_dev(scan_win_std_dev[2530]), .feature_accum(feature_accums[2530]));
  accum_calculator ac2531(.scan_win(scan_win2531), .rectangle1_x(rectangle1_xs[2531]), .rectangle1_y(rectangle1_ys[2531]), .rectangle1_width(rectangle1_widths[2531]), .rectangle1_height(rectangle1_heights[2531]), .rectangle1_weight(rectangle1_weights[2531]), .rectangle2_x(rectangle2_xs[2531]), .rectangle2_y(rectangle2_ys[2531]), .rectangle2_width(rectangle2_widths[2531]), .rectangle2_height(rectangle2_heights[2531]), .rectangle2_weight(rectangle2_weights[2531]), .rectangle3_x(rectangle3_xs[2531]), .rectangle3_y(rectangle3_ys[2531]), .rectangle3_width(rectangle3_widths[2531]), .rectangle3_height(rectangle3_heights[2531]), .rectangle3_weight(rectangle3_weights[2531]), .feature_threshold(feature_thresholds[2531]), .feature_above(feature_aboves[2531]), .feature_below(feature_belows[2531]), .scan_win_std_dev(scan_win_std_dev[2531]), .feature_accum(feature_accums[2531]));
  accum_calculator ac2532(.scan_win(scan_win2532), .rectangle1_x(rectangle1_xs[2532]), .rectangle1_y(rectangle1_ys[2532]), .rectangle1_width(rectangle1_widths[2532]), .rectangle1_height(rectangle1_heights[2532]), .rectangle1_weight(rectangle1_weights[2532]), .rectangle2_x(rectangle2_xs[2532]), .rectangle2_y(rectangle2_ys[2532]), .rectangle2_width(rectangle2_widths[2532]), .rectangle2_height(rectangle2_heights[2532]), .rectangle2_weight(rectangle2_weights[2532]), .rectangle3_x(rectangle3_xs[2532]), .rectangle3_y(rectangle3_ys[2532]), .rectangle3_width(rectangle3_widths[2532]), .rectangle3_height(rectangle3_heights[2532]), .rectangle3_weight(rectangle3_weights[2532]), .feature_threshold(feature_thresholds[2532]), .feature_above(feature_aboves[2532]), .feature_below(feature_belows[2532]), .scan_win_std_dev(scan_win_std_dev[2532]), .feature_accum(feature_accums[2532]));
  accum_calculator ac2533(.scan_win(scan_win2533), .rectangle1_x(rectangle1_xs[2533]), .rectangle1_y(rectangle1_ys[2533]), .rectangle1_width(rectangle1_widths[2533]), .rectangle1_height(rectangle1_heights[2533]), .rectangle1_weight(rectangle1_weights[2533]), .rectangle2_x(rectangle2_xs[2533]), .rectangle2_y(rectangle2_ys[2533]), .rectangle2_width(rectangle2_widths[2533]), .rectangle2_height(rectangle2_heights[2533]), .rectangle2_weight(rectangle2_weights[2533]), .rectangle3_x(rectangle3_xs[2533]), .rectangle3_y(rectangle3_ys[2533]), .rectangle3_width(rectangle3_widths[2533]), .rectangle3_height(rectangle3_heights[2533]), .rectangle3_weight(rectangle3_weights[2533]), .feature_threshold(feature_thresholds[2533]), .feature_above(feature_aboves[2533]), .feature_below(feature_belows[2533]), .scan_win_std_dev(scan_win_std_dev[2533]), .feature_accum(feature_accums[2533]));
  accum_calculator ac2534(.scan_win(scan_win2534), .rectangle1_x(rectangle1_xs[2534]), .rectangle1_y(rectangle1_ys[2534]), .rectangle1_width(rectangle1_widths[2534]), .rectangle1_height(rectangle1_heights[2534]), .rectangle1_weight(rectangle1_weights[2534]), .rectangle2_x(rectangle2_xs[2534]), .rectangle2_y(rectangle2_ys[2534]), .rectangle2_width(rectangle2_widths[2534]), .rectangle2_height(rectangle2_heights[2534]), .rectangle2_weight(rectangle2_weights[2534]), .rectangle3_x(rectangle3_xs[2534]), .rectangle3_y(rectangle3_ys[2534]), .rectangle3_width(rectangle3_widths[2534]), .rectangle3_height(rectangle3_heights[2534]), .rectangle3_weight(rectangle3_weights[2534]), .feature_threshold(feature_thresholds[2534]), .feature_above(feature_aboves[2534]), .feature_below(feature_belows[2534]), .scan_win_std_dev(scan_win_std_dev[2534]), .feature_accum(feature_accums[2534]));
  accum_calculator ac2535(.scan_win(scan_win2535), .rectangle1_x(rectangle1_xs[2535]), .rectangle1_y(rectangle1_ys[2535]), .rectangle1_width(rectangle1_widths[2535]), .rectangle1_height(rectangle1_heights[2535]), .rectangle1_weight(rectangle1_weights[2535]), .rectangle2_x(rectangle2_xs[2535]), .rectangle2_y(rectangle2_ys[2535]), .rectangle2_width(rectangle2_widths[2535]), .rectangle2_height(rectangle2_heights[2535]), .rectangle2_weight(rectangle2_weights[2535]), .rectangle3_x(rectangle3_xs[2535]), .rectangle3_y(rectangle3_ys[2535]), .rectangle3_width(rectangle3_widths[2535]), .rectangle3_height(rectangle3_heights[2535]), .rectangle3_weight(rectangle3_weights[2535]), .feature_threshold(feature_thresholds[2535]), .feature_above(feature_aboves[2535]), .feature_below(feature_belows[2535]), .scan_win_std_dev(scan_win_std_dev[2535]), .feature_accum(feature_accums[2535]));
  accum_calculator ac2536(.scan_win(scan_win2536), .rectangle1_x(rectangle1_xs[2536]), .rectangle1_y(rectangle1_ys[2536]), .rectangle1_width(rectangle1_widths[2536]), .rectangle1_height(rectangle1_heights[2536]), .rectangle1_weight(rectangle1_weights[2536]), .rectangle2_x(rectangle2_xs[2536]), .rectangle2_y(rectangle2_ys[2536]), .rectangle2_width(rectangle2_widths[2536]), .rectangle2_height(rectangle2_heights[2536]), .rectangle2_weight(rectangle2_weights[2536]), .rectangle3_x(rectangle3_xs[2536]), .rectangle3_y(rectangle3_ys[2536]), .rectangle3_width(rectangle3_widths[2536]), .rectangle3_height(rectangle3_heights[2536]), .rectangle3_weight(rectangle3_weights[2536]), .feature_threshold(feature_thresholds[2536]), .feature_above(feature_aboves[2536]), .feature_below(feature_belows[2536]), .scan_win_std_dev(scan_win_std_dev[2536]), .feature_accum(feature_accums[2536]));
  accum_calculator ac2537(.scan_win(scan_win2537), .rectangle1_x(rectangle1_xs[2537]), .rectangle1_y(rectangle1_ys[2537]), .rectangle1_width(rectangle1_widths[2537]), .rectangle1_height(rectangle1_heights[2537]), .rectangle1_weight(rectangle1_weights[2537]), .rectangle2_x(rectangle2_xs[2537]), .rectangle2_y(rectangle2_ys[2537]), .rectangle2_width(rectangle2_widths[2537]), .rectangle2_height(rectangle2_heights[2537]), .rectangle2_weight(rectangle2_weights[2537]), .rectangle3_x(rectangle3_xs[2537]), .rectangle3_y(rectangle3_ys[2537]), .rectangle3_width(rectangle3_widths[2537]), .rectangle3_height(rectangle3_heights[2537]), .rectangle3_weight(rectangle3_weights[2537]), .feature_threshold(feature_thresholds[2537]), .feature_above(feature_aboves[2537]), .feature_below(feature_belows[2537]), .scan_win_std_dev(scan_win_std_dev[2537]), .feature_accum(feature_accums[2537]));
  accum_calculator ac2538(.scan_win(scan_win2538), .rectangle1_x(rectangle1_xs[2538]), .rectangle1_y(rectangle1_ys[2538]), .rectangle1_width(rectangle1_widths[2538]), .rectangle1_height(rectangle1_heights[2538]), .rectangle1_weight(rectangle1_weights[2538]), .rectangle2_x(rectangle2_xs[2538]), .rectangle2_y(rectangle2_ys[2538]), .rectangle2_width(rectangle2_widths[2538]), .rectangle2_height(rectangle2_heights[2538]), .rectangle2_weight(rectangle2_weights[2538]), .rectangle3_x(rectangle3_xs[2538]), .rectangle3_y(rectangle3_ys[2538]), .rectangle3_width(rectangle3_widths[2538]), .rectangle3_height(rectangle3_heights[2538]), .rectangle3_weight(rectangle3_weights[2538]), .feature_threshold(feature_thresholds[2538]), .feature_above(feature_aboves[2538]), .feature_below(feature_belows[2538]), .scan_win_std_dev(scan_win_std_dev[2538]), .feature_accum(feature_accums[2538]));
  accum_calculator ac2539(.scan_win(scan_win2539), .rectangle1_x(rectangle1_xs[2539]), .rectangle1_y(rectangle1_ys[2539]), .rectangle1_width(rectangle1_widths[2539]), .rectangle1_height(rectangle1_heights[2539]), .rectangle1_weight(rectangle1_weights[2539]), .rectangle2_x(rectangle2_xs[2539]), .rectangle2_y(rectangle2_ys[2539]), .rectangle2_width(rectangle2_widths[2539]), .rectangle2_height(rectangle2_heights[2539]), .rectangle2_weight(rectangle2_weights[2539]), .rectangle3_x(rectangle3_xs[2539]), .rectangle3_y(rectangle3_ys[2539]), .rectangle3_width(rectangle3_widths[2539]), .rectangle3_height(rectangle3_heights[2539]), .rectangle3_weight(rectangle3_weights[2539]), .feature_threshold(feature_thresholds[2539]), .feature_above(feature_aboves[2539]), .feature_below(feature_belows[2539]), .scan_win_std_dev(scan_win_std_dev[2539]), .feature_accum(feature_accums[2539]));
  accum_calculator ac2540(.scan_win(scan_win2540), .rectangle1_x(rectangle1_xs[2540]), .rectangle1_y(rectangle1_ys[2540]), .rectangle1_width(rectangle1_widths[2540]), .rectangle1_height(rectangle1_heights[2540]), .rectangle1_weight(rectangle1_weights[2540]), .rectangle2_x(rectangle2_xs[2540]), .rectangle2_y(rectangle2_ys[2540]), .rectangle2_width(rectangle2_widths[2540]), .rectangle2_height(rectangle2_heights[2540]), .rectangle2_weight(rectangle2_weights[2540]), .rectangle3_x(rectangle3_xs[2540]), .rectangle3_y(rectangle3_ys[2540]), .rectangle3_width(rectangle3_widths[2540]), .rectangle3_height(rectangle3_heights[2540]), .rectangle3_weight(rectangle3_weights[2540]), .feature_threshold(feature_thresholds[2540]), .feature_above(feature_aboves[2540]), .feature_below(feature_belows[2540]), .scan_win_std_dev(scan_win_std_dev[2540]), .feature_accum(feature_accums[2540]));
  accum_calculator ac2541(.scan_win(scan_win2541), .rectangle1_x(rectangle1_xs[2541]), .rectangle1_y(rectangle1_ys[2541]), .rectangle1_width(rectangle1_widths[2541]), .rectangle1_height(rectangle1_heights[2541]), .rectangle1_weight(rectangle1_weights[2541]), .rectangle2_x(rectangle2_xs[2541]), .rectangle2_y(rectangle2_ys[2541]), .rectangle2_width(rectangle2_widths[2541]), .rectangle2_height(rectangle2_heights[2541]), .rectangle2_weight(rectangle2_weights[2541]), .rectangle3_x(rectangle3_xs[2541]), .rectangle3_y(rectangle3_ys[2541]), .rectangle3_width(rectangle3_widths[2541]), .rectangle3_height(rectangle3_heights[2541]), .rectangle3_weight(rectangle3_weights[2541]), .feature_threshold(feature_thresholds[2541]), .feature_above(feature_aboves[2541]), .feature_below(feature_belows[2541]), .scan_win_std_dev(scan_win_std_dev[2541]), .feature_accum(feature_accums[2541]));
  accum_calculator ac2542(.scan_win(scan_win2542), .rectangle1_x(rectangle1_xs[2542]), .rectangle1_y(rectangle1_ys[2542]), .rectangle1_width(rectangle1_widths[2542]), .rectangle1_height(rectangle1_heights[2542]), .rectangle1_weight(rectangle1_weights[2542]), .rectangle2_x(rectangle2_xs[2542]), .rectangle2_y(rectangle2_ys[2542]), .rectangle2_width(rectangle2_widths[2542]), .rectangle2_height(rectangle2_heights[2542]), .rectangle2_weight(rectangle2_weights[2542]), .rectangle3_x(rectangle3_xs[2542]), .rectangle3_y(rectangle3_ys[2542]), .rectangle3_width(rectangle3_widths[2542]), .rectangle3_height(rectangle3_heights[2542]), .rectangle3_weight(rectangle3_weights[2542]), .feature_threshold(feature_thresholds[2542]), .feature_above(feature_aboves[2542]), .feature_below(feature_belows[2542]), .scan_win_std_dev(scan_win_std_dev[2542]), .feature_accum(feature_accums[2542]));
  accum_calculator ac2543(.scan_win(scan_win2543), .rectangle1_x(rectangle1_xs[2543]), .rectangle1_y(rectangle1_ys[2543]), .rectangle1_width(rectangle1_widths[2543]), .rectangle1_height(rectangle1_heights[2543]), .rectangle1_weight(rectangle1_weights[2543]), .rectangle2_x(rectangle2_xs[2543]), .rectangle2_y(rectangle2_ys[2543]), .rectangle2_width(rectangle2_widths[2543]), .rectangle2_height(rectangle2_heights[2543]), .rectangle2_weight(rectangle2_weights[2543]), .rectangle3_x(rectangle3_xs[2543]), .rectangle3_y(rectangle3_ys[2543]), .rectangle3_width(rectangle3_widths[2543]), .rectangle3_height(rectangle3_heights[2543]), .rectangle3_weight(rectangle3_weights[2543]), .feature_threshold(feature_thresholds[2543]), .feature_above(feature_aboves[2543]), .feature_below(feature_belows[2543]), .scan_win_std_dev(scan_win_std_dev[2543]), .feature_accum(feature_accums[2543]));
  accum_calculator ac2544(.scan_win(scan_win2544), .rectangle1_x(rectangle1_xs[2544]), .rectangle1_y(rectangle1_ys[2544]), .rectangle1_width(rectangle1_widths[2544]), .rectangle1_height(rectangle1_heights[2544]), .rectangle1_weight(rectangle1_weights[2544]), .rectangle2_x(rectangle2_xs[2544]), .rectangle2_y(rectangle2_ys[2544]), .rectangle2_width(rectangle2_widths[2544]), .rectangle2_height(rectangle2_heights[2544]), .rectangle2_weight(rectangle2_weights[2544]), .rectangle3_x(rectangle3_xs[2544]), .rectangle3_y(rectangle3_ys[2544]), .rectangle3_width(rectangle3_widths[2544]), .rectangle3_height(rectangle3_heights[2544]), .rectangle3_weight(rectangle3_weights[2544]), .feature_threshold(feature_thresholds[2544]), .feature_above(feature_aboves[2544]), .feature_below(feature_belows[2544]), .scan_win_std_dev(scan_win_std_dev[2544]), .feature_accum(feature_accums[2544]));
  accum_calculator ac2545(.scan_win(scan_win2545), .rectangle1_x(rectangle1_xs[2545]), .rectangle1_y(rectangle1_ys[2545]), .rectangle1_width(rectangle1_widths[2545]), .rectangle1_height(rectangle1_heights[2545]), .rectangle1_weight(rectangle1_weights[2545]), .rectangle2_x(rectangle2_xs[2545]), .rectangle2_y(rectangle2_ys[2545]), .rectangle2_width(rectangle2_widths[2545]), .rectangle2_height(rectangle2_heights[2545]), .rectangle2_weight(rectangle2_weights[2545]), .rectangle3_x(rectangle3_xs[2545]), .rectangle3_y(rectangle3_ys[2545]), .rectangle3_width(rectangle3_widths[2545]), .rectangle3_height(rectangle3_heights[2545]), .rectangle3_weight(rectangle3_weights[2545]), .feature_threshold(feature_thresholds[2545]), .feature_above(feature_aboves[2545]), .feature_below(feature_belows[2545]), .scan_win_std_dev(scan_win_std_dev[2545]), .feature_accum(feature_accums[2545]));
  accum_calculator ac2546(.scan_win(scan_win2546), .rectangle1_x(rectangle1_xs[2546]), .rectangle1_y(rectangle1_ys[2546]), .rectangle1_width(rectangle1_widths[2546]), .rectangle1_height(rectangle1_heights[2546]), .rectangle1_weight(rectangle1_weights[2546]), .rectangle2_x(rectangle2_xs[2546]), .rectangle2_y(rectangle2_ys[2546]), .rectangle2_width(rectangle2_widths[2546]), .rectangle2_height(rectangle2_heights[2546]), .rectangle2_weight(rectangle2_weights[2546]), .rectangle3_x(rectangle3_xs[2546]), .rectangle3_y(rectangle3_ys[2546]), .rectangle3_width(rectangle3_widths[2546]), .rectangle3_height(rectangle3_heights[2546]), .rectangle3_weight(rectangle3_weights[2546]), .feature_threshold(feature_thresholds[2546]), .feature_above(feature_aboves[2546]), .feature_below(feature_belows[2546]), .scan_win_std_dev(scan_win_std_dev[2546]), .feature_accum(feature_accums[2546]));
  accum_calculator ac2547(.scan_win(scan_win2547), .rectangle1_x(rectangle1_xs[2547]), .rectangle1_y(rectangle1_ys[2547]), .rectangle1_width(rectangle1_widths[2547]), .rectangle1_height(rectangle1_heights[2547]), .rectangle1_weight(rectangle1_weights[2547]), .rectangle2_x(rectangle2_xs[2547]), .rectangle2_y(rectangle2_ys[2547]), .rectangle2_width(rectangle2_widths[2547]), .rectangle2_height(rectangle2_heights[2547]), .rectangle2_weight(rectangle2_weights[2547]), .rectangle3_x(rectangle3_xs[2547]), .rectangle3_y(rectangle3_ys[2547]), .rectangle3_width(rectangle3_widths[2547]), .rectangle3_height(rectangle3_heights[2547]), .rectangle3_weight(rectangle3_weights[2547]), .feature_threshold(feature_thresholds[2547]), .feature_above(feature_aboves[2547]), .feature_below(feature_belows[2547]), .scan_win_std_dev(scan_win_std_dev[2547]), .feature_accum(feature_accums[2547]));
  accum_calculator ac2548(.scan_win(scan_win2548), .rectangle1_x(rectangle1_xs[2548]), .rectangle1_y(rectangle1_ys[2548]), .rectangle1_width(rectangle1_widths[2548]), .rectangle1_height(rectangle1_heights[2548]), .rectangle1_weight(rectangle1_weights[2548]), .rectangle2_x(rectangle2_xs[2548]), .rectangle2_y(rectangle2_ys[2548]), .rectangle2_width(rectangle2_widths[2548]), .rectangle2_height(rectangle2_heights[2548]), .rectangle2_weight(rectangle2_weights[2548]), .rectangle3_x(rectangle3_xs[2548]), .rectangle3_y(rectangle3_ys[2548]), .rectangle3_width(rectangle3_widths[2548]), .rectangle3_height(rectangle3_heights[2548]), .rectangle3_weight(rectangle3_weights[2548]), .feature_threshold(feature_thresholds[2548]), .feature_above(feature_aboves[2548]), .feature_below(feature_belows[2548]), .scan_win_std_dev(scan_win_std_dev[2548]), .feature_accum(feature_accums[2548]));
  accum_calculator ac2549(.scan_win(scan_win2549), .rectangle1_x(rectangle1_xs[2549]), .rectangle1_y(rectangle1_ys[2549]), .rectangle1_width(rectangle1_widths[2549]), .rectangle1_height(rectangle1_heights[2549]), .rectangle1_weight(rectangle1_weights[2549]), .rectangle2_x(rectangle2_xs[2549]), .rectangle2_y(rectangle2_ys[2549]), .rectangle2_width(rectangle2_widths[2549]), .rectangle2_height(rectangle2_heights[2549]), .rectangle2_weight(rectangle2_weights[2549]), .rectangle3_x(rectangle3_xs[2549]), .rectangle3_y(rectangle3_ys[2549]), .rectangle3_width(rectangle3_widths[2549]), .rectangle3_height(rectangle3_heights[2549]), .rectangle3_weight(rectangle3_weights[2549]), .feature_threshold(feature_thresholds[2549]), .feature_above(feature_aboves[2549]), .feature_below(feature_belows[2549]), .scan_win_std_dev(scan_win_std_dev[2549]), .feature_accum(feature_accums[2549]));
  accum_calculator ac2550(.scan_win(scan_win2550), .rectangle1_x(rectangle1_xs[2550]), .rectangle1_y(rectangle1_ys[2550]), .rectangle1_width(rectangle1_widths[2550]), .rectangle1_height(rectangle1_heights[2550]), .rectangle1_weight(rectangle1_weights[2550]), .rectangle2_x(rectangle2_xs[2550]), .rectangle2_y(rectangle2_ys[2550]), .rectangle2_width(rectangle2_widths[2550]), .rectangle2_height(rectangle2_heights[2550]), .rectangle2_weight(rectangle2_weights[2550]), .rectangle3_x(rectangle3_xs[2550]), .rectangle3_y(rectangle3_ys[2550]), .rectangle3_width(rectangle3_widths[2550]), .rectangle3_height(rectangle3_heights[2550]), .rectangle3_weight(rectangle3_weights[2550]), .feature_threshold(feature_thresholds[2550]), .feature_above(feature_aboves[2550]), .feature_below(feature_belows[2550]), .scan_win_std_dev(scan_win_std_dev[2550]), .feature_accum(feature_accums[2550]));
  accum_calculator ac2551(.scan_win(scan_win2551), .rectangle1_x(rectangle1_xs[2551]), .rectangle1_y(rectangle1_ys[2551]), .rectangle1_width(rectangle1_widths[2551]), .rectangle1_height(rectangle1_heights[2551]), .rectangle1_weight(rectangle1_weights[2551]), .rectangle2_x(rectangle2_xs[2551]), .rectangle2_y(rectangle2_ys[2551]), .rectangle2_width(rectangle2_widths[2551]), .rectangle2_height(rectangle2_heights[2551]), .rectangle2_weight(rectangle2_weights[2551]), .rectangle3_x(rectangle3_xs[2551]), .rectangle3_y(rectangle3_ys[2551]), .rectangle3_width(rectangle3_widths[2551]), .rectangle3_height(rectangle3_heights[2551]), .rectangle3_weight(rectangle3_weights[2551]), .feature_threshold(feature_thresholds[2551]), .feature_above(feature_aboves[2551]), .feature_below(feature_belows[2551]), .scan_win_std_dev(scan_win_std_dev[2551]), .feature_accum(feature_accums[2551]));
  accum_calculator ac2552(.scan_win(scan_win2552), .rectangle1_x(rectangle1_xs[2552]), .rectangle1_y(rectangle1_ys[2552]), .rectangle1_width(rectangle1_widths[2552]), .rectangle1_height(rectangle1_heights[2552]), .rectangle1_weight(rectangle1_weights[2552]), .rectangle2_x(rectangle2_xs[2552]), .rectangle2_y(rectangle2_ys[2552]), .rectangle2_width(rectangle2_widths[2552]), .rectangle2_height(rectangle2_heights[2552]), .rectangle2_weight(rectangle2_weights[2552]), .rectangle3_x(rectangle3_xs[2552]), .rectangle3_y(rectangle3_ys[2552]), .rectangle3_width(rectangle3_widths[2552]), .rectangle3_height(rectangle3_heights[2552]), .rectangle3_weight(rectangle3_weights[2552]), .feature_threshold(feature_thresholds[2552]), .feature_above(feature_aboves[2552]), .feature_below(feature_belows[2552]), .scan_win_std_dev(scan_win_std_dev[2552]), .feature_accum(feature_accums[2552]));
  accum_calculator ac2553(.scan_win(scan_win2553), .rectangle1_x(rectangle1_xs[2553]), .rectangle1_y(rectangle1_ys[2553]), .rectangle1_width(rectangle1_widths[2553]), .rectangle1_height(rectangle1_heights[2553]), .rectangle1_weight(rectangle1_weights[2553]), .rectangle2_x(rectangle2_xs[2553]), .rectangle2_y(rectangle2_ys[2553]), .rectangle2_width(rectangle2_widths[2553]), .rectangle2_height(rectangle2_heights[2553]), .rectangle2_weight(rectangle2_weights[2553]), .rectangle3_x(rectangle3_xs[2553]), .rectangle3_y(rectangle3_ys[2553]), .rectangle3_width(rectangle3_widths[2553]), .rectangle3_height(rectangle3_heights[2553]), .rectangle3_weight(rectangle3_weights[2553]), .feature_threshold(feature_thresholds[2553]), .feature_above(feature_aboves[2553]), .feature_below(feature_belows[2553]), .scan_win_std_dev(scan_win_std_dev[2553]), .feature_accum(feature_accums[2553]));
  accum_calculator ac2554(.scan_win(scan_win2554), .rectangle1_x(rectangle1_xs[2554]), .rectangle1_y(rectangle1_ys[2554]), .rectangle1_width(rectangle1_widths[2554]), .rectangle1_height(rectangle1_heights[2554]), .rectangle1_weight(rectangle1_weights[2554]), .rectangle2_x(rectangle2_xs[2554]), .rectangle2_y(rectangle2_ys[2554]), .rectangle2_width(rectangle2_widths[2554]), .rectangle2_height(rectangle2_heights[2554]), .rectangle2_weight(rectangle2_weights[2554]), .rectangle3_x(rectangle3_xs[2554]), .rectangle3_y(rectangle3_ys[2554]), .rectangle3_width(rectangle3_widths[2554]), .rectangle3_height(rectangle3_heights[2554]), .rectangle3_weight(rectangle3_weights[2554]), .feature_threshold(feature_thresholds[2554]), .feature_above(feature_aboves[2554]), .feature_below(feature_belows[2554]), .scan_win_std_dev(scan_win_std_dev[2554]), .feature_accum(feature_accums[2554]));
  accum_calculator ac2555(.scan_win(scan_win2555), .rectangle1_x(rectangle1_xs[2555]), .rectangle1_y(rectangle1_ys[2555]), .rectangle1_width(rectangle1_widths[2555]), .rectangle1_height(rectangle1_heights[2555]), .rectangle1_weight(rectangle1_weights[2555]), .rectangle2_x(rectangle2_xs[2555]), .rectangle2_y(rectangle2_ys[2555]), .rectangle2_width(rectangle2_widths[2555]), .rectangle2_height(rectangle2_heights[2555]), .rectangle2_weight(rectangle2_weights[2555]), .rectangle3_x(rectangle3_xs[2555]), .rectangle3_y(rectangle3_ys[2555]), .rectangle3_width(rectangle3_widths[2555]), .rectangle3_height(rectangle3_heights[2555]), .rectangle3_weight(rectangle3_weights[2555]), .feature_threshold(feature_thresholds[2555]), .feature_above(feature_aboves[2555]), .feature_below(feature_belows[2555]), .scan_win_std_dev(scan_win_std_dev[2555]), .feature_accum(feature_accums[2555]));
  accum_calculator ac2556(.scan_win(scan_win2556), .rectangle1_x(rectangle1_xs[2556]), .rectangle1_y(rectangle1_ys[2556]), .rectangle1_width(rectangle1_widths[2556]), .rectangle1_height(rectangle1_heights[2556]), .rectangle1_weight(rectangle1_weights[2556]), .rectangle2_x(rectangle2_xs[2556]), .rectangle2_y(rectangle2_ys[2556]), .rectangle2_width(rectangle2_widths[2556]), .rectangle2_height(rectangle2_heights[2556]), .rectangle2_weight(rectangle2_weights[2556]), .rectangle3_x(rectangle3_xs[2556]), .rectangle3_y(rectangle3_ys[2556]), .rectangle3_width(rectangle3_widths[2556]), .rectangle3_height(rectangle3_heights[2556]), .rectangle3_weight(rectangle3_weights[2556]), .feature_threshold(feature_thresholds[2556]), .feature_above(feature_aboves[2556]), .feature_below(feature_belows[2556]), .scan_win_std_dev(scan_win_std_dev[2556]), .feature_accum(feature_accums[2556]));
  accum_calculator ac2557(.scan_win(scan_win2557), .rectangle1_x(rectangle1_xs[2557]), .rectangle1_y(rectangle1_ys[2557]), .rectangle1_width(rectangle1_widths[2557]), .rectangle1_height(rectangle1_heights[2557]), .rectangle1_weight(rectangle1_weights[2557]), .rectangle2_x(rectangle2_xs[2557]), .rectangle2_y(rectangle2_ys[2557]), .rectangle2_width(rectangle2_widths[2557]), .rectangle2_height(rectangle2_heights[2557]), .rectangle2_weight(rectangle2_weights[2557]), .rectangle3_x(rectangle3_xs[2557]), .rectangle3_y(rectangle3_ys[2557]), .rectangle3_width(rectangle3_widths[2557]), .rectangle3_height(rectangle3_heights[2557]), .rectangle3_weight(rectangle3_weights[2557]), .feature_threshold(feature_thresholds[2557]), .feature_above(feature_aboves[2557]), .feature_below(feature_belows[2557]), .scan_win_std_dev(scan_win_std_dev[2557]), .feature_accum(feature_accums[2557]));
  accum_calculator ac2558(.scan_win(scan_win2558), .rectangle1_x(rectangle1_xs[2558]), .rectangle1_y(rectangle1_ys[2558]), .rectangle1_width(rectangle1_widths[2558]), .rectangle1_height(rectangle1_heights[2558]), .rectangle1_weight(rectangle1_weights[2558]), .rectangle2_x(rectangle2_xs[2558]), .rectangle2_y(rectangle2_ys[2558]), .rectangle2_width(rectangle2_widths[2558]), .rectangle2_height(rectangle2_heights[2558]), .rectangle2_weight(rectangle2_weights[2558]), .rectangle3_x(rectangle3_xs[2558]), .rectangle3_y(rectangle3_ys[2558]), .rectangle3_width(rectangle3_widths[2558]), .rectangle3_height(rectangle3_heights[2558]), .rectangle3_weight(rectangle3_weights[2558]), .feature_threshold(feature_thresholds[2558]), .feature_above(feature_aboves[2558]), .feature_below(feature_belows[2558]), .scan_win_std_dev(scan_win_std_dev[2558]), .feature_accum(feature_accums[2558]));
  accum_calculator ac2559(.scan_win(scan_win2559), .rectangle1_x(rectangle1_xs[2559]), .rectangle1_y(rectangle1_ys[2559]), .rectangle1_width(rectangle1_widths[2559]), .rectangle1_height(rectangle1_heights[2559]), .rectangle1_weight(rectangle1_weights[2559]), .rectangle2_x(rectangle2_xs[2559]), .rectangle2_y(rectangle2_ys[2559]), .rectangle2_width(rectangle2_widths[2559]), .rectangle2_height(rectangle2_heights[2559]), .rectangle2_weight(rectangle2_weights[2559]), .rectangle3_x(rectangle3_xs[2559]), .rectangle3_y(rectangle3_ys[2559]), .rectangle3_width(rectangle3_widths[2559]), .rectangle3_height(rectangle3_heights[2559]), .rectangle3_weight(rectangle3_weights[2559]), .feature_threshold(feature_thresholds[2559]), .feature_above(feature_aboves[2559]), .feature_below(feature_belows[2559]), .scan_win_std_dev(scan_win_std_dev[2559]), .feature_accum(feature_accums[2559]));
  accum_calculator ac2560(.scan_win(scan_win2560), .rectangle1_x(rectangle1_xs[2560]), .rectangle1_y(rectangle1_ys[2560]), .rectangle1_width(rectangle1_widths[2560]), .rectangle1_height(rectangle1_heights[2560]), .rectangle1_weight(rectangle1_weights[2560]), .rectangle2_x(rectangle2_xs[2560]), .rectangle2_y(rectangle2_ys[2560]), .rectangle2_width(rectangle2_widths[2560]), .rectangle2_height(rectangle2_heights[2560]), .rectangle2_weight(rectangle2_weights[2560]), .rectangle3_x(rectangle3_xs[2560]), .rectangle3_y(rectangle3_ys[2560]), .rectangle3_width(rectangle3_widths[2560]), .rectangle3_height(rectangle3_heights[2560]), .rectangle3_weight(rectangle3_weights[2560]), .feature_threshold(feature_thresholds[2560]), .feature_above(feature_aboves[2560]), .feature_below(feature_belows[2560]), .scan_win_std_dev(scan_win_std_dev[2560]), .feature_accum(feature_accums[2560]));
  accum_calculator ac2561(.scan_win(scan_win2561), .rectangle1_x(rectangle1_xs[2561]), .rectangle1_y(rectangle1_ys[2561]), .rectangle1_width(rectangle1_widths[2561]), .rectangle1_height(rectangle1_heights[2561]), .rectangle1_weight(rectangle1_weights[2561]), .rectangle2_x(rectangle2_xs[2561]), .rectangle2_y(rectangle2_ys[2561]), .rectangle2_width(rectangle2_widths[2561]), .rectangle2_height(rectangle2_heights[2561]), .rectangle2_weight(rectangle2_weights[2561]), .rectangle3_x(rectangle3_xs[2561]), .rectangle3_y(rectangle3_ys[2561]), .rectangle3_width(rectangle3_widths[2561]), .rectangle3_height(rectangle3_heights[2561]), .rectangle3_weight(rectangle3_weights[2561]), .feature_threshold(feature_thresholds[2561]), .feature_above(feature_aboves[2561]), .feature_below(feature_belows[2561]), .scan_win_std_dev(scan_win_std_dev[2561]), .feature_accum(feature_accums[2561]));
  accum_calculator ac2562(.scan_win(scan_win2562), .rectangle1_x(rectangle1_xs[2562]), .rectangle1_y(rectangle1_ys[2562]), .rectangle1_width(rectangle1_widths[2562]), .rectangle1_height(rectangle1_heights[2562]), .rectangle1_weight(rectangle1_weights[2562]), .rectangle2_x(rectangle2_xs[2562]), .rectangle2_y(rectangle2_ys[2562]), .rectangle2_width(rectangle2_widths[2562]), .rectangle2_height(rectangle2_heights[2562]), .rectangle2_weight(rectangle2_weights[2562]), .rectangle3_x(rectangle3_xs[2562]), .rectangle3_y(rectangle3_ys[2562]), .rectangle3_width(rectangle3_widths[2562]), .rectangle3_height(rectangle3_heights[2562]), .rectangle3_weight(rectangle3_weights[2562]), .feature_threshold(feature_thresholds[2562]), .feature_above(feature_aboves[2562]), .feature_below(feature_belows[2562]), .scan_win_std_dev(scan_win_std_dev[2562]), .feature_accum(feature_accums[2562]));
  accum_calculator ac2563(.scan_win(scan_win2563), .rectangle1_x(rectangle1_xs[2563]), .rectangle1_y(rectangle1_ys[2563]), .rectangle1_width(rectangle1_widths[2563]), .rectangle1_height(rectangle1_heights[2563]), .rectangle1_weight(rectangle1_weights[2563]), .rectangle2_x(rectangle2_xs[2563]), .rectangle2_y(rectangle2_ys[2563]), .rectangle2_width(rectangle2_widths[2563]), .rectangle2_height(rectangle2_heights[2563]), .rectangle2_weight(rectangle2_weights[2563]), .rectangle3_x(rectangle3_xs[2563]), .rectangle3_y(rectangle3_ys[2563]), .rectangle3_width(rectangle3_widths[2563]), .rectangle3_height(rectangle3_heights[2563]), .rectangle3_weight(rectangle3_weights[2563]), .feature_threshold(feature_thresholds[2563]), .feature_above(feature_aboves[2563]), .feature_below(feature_belows[2563]), .scan_win_std_dev(scan_win_std_dev[2563]), .feature_accum(feature_accums[2563]));
  accum_calculator ac2564(.scan_win(scan_win2564), .rectangle1_x(rectangle1_xs[2564]), .rectangle1_y(rectangle1_ys[2564]), .rectangle1_width(rectangle1_widths[2564]), .rectangle1_height(rectangle1_heights[2564]), .rectangle1_weight(rectangle1_weights[2564]), .rectangle2_x(rectangle2_xs[2564]), .rectangle2_y(rectangle2_ys[2564]), .rectangle2_width(rectangle2_widths[2564]), .rectangle2_height(rectangle2_heights[2564]), .rectangle2_weight(rectangle2_weights[2564]), .rectangle3_x(rectangle3_xs[2564]), .rectangle3_y(rectangle3_ys[2564]), .rectangle3_width(rectangle3_widths[2564]), .rectangle3_height(rectangle3_heights[2564]), .rectangle3_weight(rectangle3_weights[2564]), .feature_threshold(feature_thresholds[2564]), .feature_above(feature_aboves[2564]), .feature_below(feature_belows[2564]), .scan_win_std_dev(scan_win_std_dev[2564]), .feature_accum(feature_accums[2564]));
  accum_calculator ac2565(.scan_win(scan_win2565), .rectangle1_x(rectangle1_xs[2565]), .rectangle1_y(rectangle1_ys[2565]), .rectangle1_width(rectangle1_widths[2565]), .rectangle1_height(rectangle1_heights[2565]), .rectangle1_weight(rectangle1_weights[2565]), .rectangle2_x(rectangle2_xs[2565]), .rectangle2_y(rectangle2_ys[2565]), .rectangle2_width(rectangle2_widths[2565]), .rectangle2_height(rectangle2_heights[2565]), .rectangle2_weight(rectangle2_weights[2565]), .rectangle3_x(rectangle3_xs[2565]), .rectangle3_y(rectangle3_ys[2565]), .rectangle3_width(rectangle3_widths[2565]), .rectangle3_height(rectangle3_heights[2565]), .rectangle3_weight(rectangle3_weights[2565]), .feature_threshold(feature_thresholds[2565]), .feature_above(feature_aboves[2565]), .feature_below(feature_belows[2565]), .scan_win_std_dev(scan_win_std_dev[2565]), .feature_accum(feature_accums[2565]));
  accum_calculator ac2566(.scan_win(scan_win2566), .rectangle1_x(rectangle1_xs[2566]), .rectangle1_y(rectangle1_ys[2566]), .rectangle1_width(rectangle1_widths[2566]), .rectangle1_height(rectangle1_heights[2566]), .rectangle1_weight(rectangle1_weights[2566]), .rectangle2_x(rectangle2_xs[2566]), .rectangle2_y(rectangle2_ys[2566]), .rectangle2_width(rectangle2_widths[2566]), .rectangle2_height(rectangle2_heights[2566]), .rectangle2_weight(rectangle2_weights[2566]), .rectangle3_x(rectangle3_xs[2566]), .rectangle3_y(rectangle3_ys[2566]), .rectangle3_width(rectangle3_widths[2566]), .rectangle3_height(rectangle3_heights[2566]), .rectangle3_weight(rectangle3_weights[2566]), .feature_threshold(feature_thresholds[2566]), .feature_above(feature_aboves[2566]), .feature_below(feature_belows[2566]), .scan_win_std_dev(scan_win_std_dev[2566]), .feature_accum(feature_accums[2566]));
  accum_calculator ac2567(.scan_win(scan_win2567), .rectangle1_x(rectangle1_xs[2567]), .rectangle1_y(rectangle1_ys[2567]), .rectangle1_width(rectangle1_widths[2567]), .rectangle1_height(rectangle1_heights[2567]), .rectangle1_weight(rectangle1_weights[2567]), .rectangle2_x(rectangle2_xs[2567]), .rectangle2_y(rectangle2_ys[2567]), .rectangle2_width(rectangle2_widths[2567]), .rectangle2_height(rectangle2_heights[2567]), .rectangle2_weight(rectangle2_weights[2567]), .rectangle3_x(rectangle3_xs[2567]), .rectangle3_y(rectangle3_ys[2567]), .rectangle3_width(rectangle3_widths[2567]), .rectangle3_height(rectangle3_heights[2567]), .rectangle3_weight(rectangle3_weights[2567]), .feature_threshold(feature_thresholds[2567]), .feature_above(feature_aboves[2567]), .feature_below(feature_belows[2567]), .scan_win_std_dev(scan_win_std_dev[2567]), .feature_accum(feature_accums[2567]));
  accum_calculator ac2568(.scan_win(scan_win2568), .rectangle1_x(rectangle1_xs[2568]), .rectangle1_y(rectangle1_ys[2568]), .rectangle1_width(rectangle1_widths[2568]), .rectangle1_height(rectangle1_heights[2568]), .rectangle1_weight(rectangle1_weights[2568]), .rectangle2_x(rectangle2_xs[2568]), .rectangle2_y(rectangle2_ys[2568]), .rectangle2_width(rectangle2_widths[2568]), .rectangle2_height(rectangle2_heights[2568]), .rectangle2_weight(rectangle2_weights[2568]), .rectangle3_x(rectangle3_xs[2568]), .rectangle3_y(rectangle3_ys[2568]), .rectangle3_width(rectangle3_widths[2568]), .rectangle3_height(rectangle3_heights[2568]), .rectangle3_weight(rectangle3_weights[2568]), .feature_threshold(feature_thresholds[2568]), .feature_above(feature_aboves[2568]), .feature_below(feature_belows[2568]), .scan_win_std_dev(scan_win_std_dev[2568]), .feature_accum(feature_accums[2568]));
  accum_calculator ac2569(.scan_win(scan_win2569), .rectangle1_x(rectangle1_xs[2569]), .rectangle1_y(rectangle1_ys[2569]), .rectangle1_width(rectangle1_widths[2569]), .rectangle1_height(rectangle1_heights[2569]), .rectangle1_weight(rectangle1_weights[2569]), .rectangle2_x(rectangle2_xs[2569]), .rectangle2_y(rectangle2_ys[2569]), .rectangle2_width(rectangle2_widths[2569]), .rectangle2_height(rectangle2_heights[2569]), .rectangle2_weight(rectangle2_weights[2569]), .rectangle3_x(rectangle3_xs[2569]), .rectangle3_y(rectangle3_ys[2569]), .rectangle3_width(rectangle3_widths[2569]), .rectangle3_height(rectangle3_heights[2569]), .rectangle3_weight(rectangle3_weights[2569]), .feature_threshold(feature_thresholds[2569]), .feature_above(feature_aboves[2569]), .feature_below(feature_belows[2569]), .scan_win_std_dev(scan_win_std_dev[2569]), .feature_accum(feature_accums[2569]));
  accum_calculator ac2570(.scan_win(scan_win2570), .rectangle1_x(rectangle1_xs[2570]), .rectangle1_y(rectangle1_ys[2570]), .rectangle1_width(rectangle1_widths[2570]), .rectangle1_height(rectangle1_heights[2570]), .rectangle1_weight(rectangle1_weights[2570]), .rectangle2_x(rectangle2_xs[2570]), .rectangle2_y(rectangle2_ys[2570]), .rectangle2_width(rectangle2_widths[2570]), .rectangle2_height(rectangle2_heights[2570]), .rectangle2_weight(rectangle2_weights[2570]), .rectangle3_x(rectangle3_xs[2570]), .rectangle3_y(rectangle3_ys[2570]), .rectangle3_width(rectangle3_widths[2570]), .rectangle3_height(rectangle3_heights[2570]), .rectangle3_weight(rectangle3_weights[2570]), .feature_threshold(feature_thresholds[2570]), .feature_above(feature_aboves[2570]), .feature_below(feature_belows[2570]), .scan_win_std_dev(scan_win_std_dev[2570]), .feature_accum(feature_accums[2570]));
  accum_calculator ac2571(.scan_win(scan_win2571), .rectangle1_x(rectangle1_xs[2571]), .rectangle1_y(rectangle1_ys[2571]), .rectangle1_width(rectangle1_widths[2571]), .rectangle1_height(rectangle1_heights[2571]), .rectangle1_weight(rectangle1_weights[2571]), .rectangle2_x(rectangle2_xs[2571]), .rectangle2_y(rectangle2_ys[2571]), .rectangle2_width(rectangle2_widths[2571]), .rectangle2_height(rectangle2_heights[2571]), .rectangle2_weight(rectangle2_weights[2571]), .rectangle3_x(rectangle3_xs[2571]), .rectangle3_y(rectangle3_ys[2571]), .rectangle3_width(rectangle3_widths[2571]), .rectangle3_height(rectangle3_heights[2571]), .rectangle3_weight(rectangle3_weights[2571]), .feature_threshold(feature_thresholds[2571]), .feature_above(feature_aboves[2571]), .feature_below(feature_belows[2571]), .scan_win_std_dev(scan_win_std_dev[2571]), .feature_accum(feature_accums[2571]));
  accum_calculator ac2572(.scan_win(scan_win2572), .rectangle1_x(rectangle1_xs[2572]), .rectangle1_y(rectangle1_ys[2572]), .rectangle1_width(rectangle1_widths[2572]), .rectangle1_height(rectangle1_heights[2572]), .rectangle1_weight(rectangle1_weights[2572]), .rectangle2_x(rectangle2_xs[2572]), .rectangle2_y(rectangle2_ys[2572]), .rectangle2_width(rectangle2_widths[2572]), .rectangle2_height(rectangle2_heights[2572]), .rectangle2_weight(rectangle2_weights[2572]), .rectangle3_x(rectangle3_xs[2572]), .rectangle3_y(rectangle3_ys[2572]), .rectangle3_width(rectangle3_widths[2572]), .rectangle3_height(rectangle3_heights[2572]), .rectangle3_weight(rectangle3_weights[2572]), .feature_threshold(feature_thresholds[2572]), .feature_above(feature_aboves[2572]), .feature_below(feature_belows[2572]), .scan_win_std_dev(scan_win_std_dev[2572]), .feature_accum(feature_accums[2572]));
  accum_calculator ac2573(.scan_win(scan_win2573), .rectangle1_x(rectangle1_xs[2573]), .rectangle1_y(rectangle1_ys[2573]), .rectangle1_width(rectangle1_widths[2573]), .rectangle1_height(rectangle1_heights[2573]), .rectangle1_weight(rectangle1_weights[2573]), .rectangle2_x(rectangle2_xs[2573]), .rectangle2_y(rectangle2_ys[2573]), .rectangle2_width(rectangle2_widths[2573]), .rectangle2_height(rectangle2_heights[2573]), .rectangle2_weight(rectangle2_weights[2573]), .rectangle3_x(rectangle3_xs[2573]), .rectangle3_y(rectangle3_ys[2573]), .rectangle3_width(rectangle3_widths[2573]), .rectangle3_height(rectangle3_heights[2573]), .rectangle3_weight(rectangle3_weights[2573]), .feature_threshold(feature_thresholds[2573]), .feature_above(feature_aboves[2573]), .feature_below(feature_belows[2573]), .scan_win_std_dev(scan_win_std_dev[2573]), .feature_accum(feature_accums[2573]));
  accum_calculator ac2574(.scan_win(scan_win2574), .rectangle1_x(rectangle1_xs[2574]), .rectangle1_y(rectangle1_ys[2574]), .rectangle1_width(rectangle1_widths[2574]), .rectangle1_height(rectangle1_heights[2574]), .rectangle1_weight(rectangle1_weights[2574]), .rectangle2_x(rectangle2_xs[2574]), .rectangle2_y(rectangle2_ys[2574]), .rectangle2_width(rectangle2_widths[2574]), .rectangle2_height(rectangle2_heights[2574]), .rectangle2_weight(rectangle2_weights[2574]), .rectangle3_x(rectangle3_xs[2574]), .rectangle3_y(rectangle3_ys[2574]), .rectangle3_width(rectangle3_widths[2574]), .rectangle3_height(rectangle3_heights[2574]), .rectangle3_weight(rectangle3_weights[2574]), .feature_threshold(feature_thresholds[2574]), .feature_above(feature_aboves[2574]), .feature_below(feature_belows[2574]), .scan_win_std_dev(scan_win_std_dev[2574]), .feature_accum(feature_accums[2574]));
  accum_calculator ac2575(.scan_win(scan_win2575), .rectangle1_x(rectangle1_xs[2575]), .rectangle1_y(rectangle1_ys[2575]), .rectangle1_width(rectangle1_widths[2575]), .rectangle1_height(rectangle1_heights[2575]), .rectangle1_weight(rectangle1_weights[2575]), .rectangle2_x(rectangle2_xs[2575]), .rectangle2_y(rectangle2_ys[2575]), .rectangle2_width(rectangle2_widths[2575]), .rectangle2_height(rectangle2_heights[2575]), .rectangle2_weight(rectangle2_weights[2575]), .rectangle3_x(rectangle3_xs[2575]), .rectangle3_y(rectangle3_ys[2575]), .rectangle3_width(rectangle3_widths[2575]), .rectangle3_height(rectangle3_heights[2575]), .rectangle3_weight(rectangle3_weights[2575]), .feature_threshold(feature_thresholds[2575]), .feature_above(feature_aboves[2575]), .feature_below(feature_belows[2575]), .scan_win_std_dev(scan_win_std_dev[2575]), .feature_accum(feature_accums[2575]));
  accum_calculator ac2576(.scan_win(scan_win2576), .rectangle1_x(rectangle1_xs[2576]), .rectangle1_y(rectangle1_ys[2576]), .rectangle1_width(rectangle1_widths[2576]), .rectangle1_height(rectangle1_heights[2576]), .rectangle1_weight(rectangle1_weights[2576]), .rectangle2_x(rectangle2_xs[2576]), .rectangle2_y(rectangle2_ys[2576]), .rectangle2_width(rectangle2_widths[2576]), .rectangle2_height(rectangle2_heights[2576]), .rectangle2_weight(rectangle2_weights[2576]), .rectangle3_x(rectangle3_xs[2576]), .rectangle3_y(rectangle3_ys[2576]), .rectangle3_width(rectangle3_widths[2576]), .rectangle3_height(rectangle3_heights[2576]), .rectangle3_weight(rectangle3_weights[2576]), .feature_threshold(feature_thresholds[2576]), .feature_above(feature_aboves[2576]), .feature_below(feature_belows[2576]), .scan_win_std_dev(scan_win_std_dev[2576]), .feature_accum(feature_accums[2576]));
  accum_calculator ac2577(.scan_win(scan_win2577), .rectangle1_x(rectangle1_xs[2577]), .rectangle1_y(rectangle1_ys[2577]), .rectangle1_width(rectangle1_widths[2577]), .rectangle1_height(rectangle1_heights[2577]), .rectangle1_weight(rectangle1_weights[2577]), .rectangle2_x(rectangle2_xs[2577]), .rectangle2_y(rectangle2_ys[2577]), .rectangle2_width(rectangle2_widths[2577]), .rectangle2_height(rectangle2_heights[2577]), .rectangle2_weight(rectangle2_weights[2577]), .rectangle3_x(rectangle3_xs[2577]), .rectangle3_y(rectangle3_ys[2577]), .rectangle3_width(rectangle3_widths[2577]), .rectangle3_height(rectangle3_heights[2577]), .rectangle3_weight(rectangle3_weights[2577]), .feature_threshold(feature_thresholds[2577]), .feature_above(feature_aboves[2577]), .feature_below(feature_belows[2577]), .scan_win_std_dev(scan_win_std_dev[2577]), .feature_accum(feature_accums[2577]));
  accum_calculator ac2578(.scan_win(scan_win2578), .rectangle1_x(rectangle1_xs[2578]), .rectangle1_y(rectangle1_ys[2578]), .rectangle1_width(rectangle1_widths[2578]), .rectangle1_height(rectangle1_heights[2578]), .rectangle1_weight(rectangle1_weights[2578]), .rectangle2_x(rectangle2_xs[2578]), .rectangle2_y(rectangle2_ys[2578]), .rectangle2_width(rectangle2_widths[2578]), .rectangle2_height(rectangle2_heights[2578]), .rectangle2_weight(rectangle2_weights[2578]), .rectangle3_x(rectangle3_xs[2578]), .rectangle3_y(rectangle3_ys[2578]), .rectangle3_width(rectangle3_widths[2578]), .rectangle3_height(rectangle3_heights[2578]), .rectangle3_weight(rectangle3_weights[2578]), .feature_threshold(feature_thresholds[2578]), .feature_above(feature_aboves[2578]), .feature_below(feature_belows[2578]), .scan_win_std_dev(scan_win_std_dev[2578]), .feature_accum(feature_accums[2578]));
  accum_calculator ac2579(.scan_win(scan_win2579), .rectangle1_x(rectangle1_xs[2579]), .rectangle1_y(rectangle1_ys[2579]), .rectangle1_width(rectangle1_widths[2579]), .rectangle1_height(rectangle1_heights[2579]), .rectangle1_weight(rectangle1_weights[2579]), .rectangle2_x(rectangle2_xs[2579]), .rectangle2_y(rectangle2_ys[2579]), .rectangle2_width(rectangle2_widths[2579]), .rectangle2_height(rectangle2_heights[2579]), .rectangle2_weight(rectangle2_weights[2579]), .rectangle3_x(rectangle3_xs[2579]), .rectangle3_y(rectangle3_ys[2579]), .rectangle3_width(rectangle3_widths[2579]), .rectangle3_height(rectangle3_heights[2579]), .rectangle3_weight(rectangle3_weights[2579]), .feature_threshold(feature_thresholds[2579]), .feature_above(feature_aboves[2579]), .feature_below(feature_belows[2579]), .scan_win_std_dev(scan_win_std_dev[2579]), .feature_accum(feature_accums[2579]));
  accum_calculator ac2580(.scan_win(scan_win2580), .rectangle1_x(rectangle1_xs[2580]), .rectangle1_y(rectangle1_ys[2580]), .rectangle1_width(rectangle1_widths[2580]), .rectangle1_height(rectangle1_heights[2580]), .rectangle1_weight(rectangle1_weights[2580]), .rectangle2_x(rectangle2_xs[2580]), .rectangle2_y(rectangle2_ys[2580]), .rectangle2_width(rectangle2_widths[2580]), .rectangle2_height(rectangle2_heights[2580]), .rectangle2_weight(rectangle2_weights[2580]), .rectangle3_x(rectangle3_xs[2580]), .rectangle3_y(rectangle3_ys[2580]), .rectangle3_width(rectangle3_widths[2580]), .rectangle3_height(rectangle3_heights[2580]), .rectangle3_weight(rectangle3_weights[2580]), .feature_threshold(feature_thresholds[2580]), .feature_above(feature_aboves[2580]), .feature_below(feature_belows[2580]), .scan_win_std_dev(scan_win_std_dev[2580]), .feature_accum(feature_accums[2580]));
  accum_calculator ac2581(.scan_win(scan_win2581), .rectangle1_x(rectangle1_xs[2581]), .rectangle1_y(rectangle1_ys[2581]), .rectangle1_width(rectangle1_widths[2581]), .rectangle1_height(rectangle1_heights[2581]), .rectangle1_weight(rectangle1_weights[2581]), .rectangle2_x(rectangle2_xs[2581]), .rectangle2_y(rectangle2_ys[2581]), .rectangle2_width(rectangle2_widths[2581]), .rectangle2_height(rectangle2_heights[2581]), .rectangle2_weight(rectangle2_weights[2581]), .rectangle3_x(rectangle3_xs[2581]), .rectangle3_y(rectangle3_ys[2581]), .rectangle3_width(rectangle3_widths[2581]), .rectangle3_height(rectangle3_heights[2581]), .rectangle3_weight(rectangle3_weights[2581]), .feature_threshold(feature_thresholds[2581]), .feature_above(feature_aboves[2581]), .feature_below(feature_belows[2581]), .scan_win_std_dev(scan_win_std_dev[2581]), .feature_accum(feature_accums[2581]));
  accum_calculator ac2582(.scan_win(scan_win2582), .rectangle1_x(rectangle1_xs[2582]), .rectangle1_y(rectangle1_ys[2582]), .rectangle1_width(rectangle1_widths[2582]), .rectangle1_height(rectangle1_heights[2582]), .rectangle1_weight(rectangle1_weights[2582]), .rectangle2_x(rectangle2_xs[2582]), .rectangle2_y(rectangle2_ys[2582]), .rectangle2_width(rectangle2_widths[2582]), .rectangle2_height(rectangle2_heights[2582]), .rectangle2_weight(rectangle2_weights[2582]), .rectangle3_x(rectangle3_xs[2582]), .rectangle3_y(rectangle3_ys[2582]), .rectangle3_width(rectangle3_widths[2582]), .rectangle3_height(rectangle3_heights[2582]), .rectangle3_weight(rectangle3_weights[2582]), .feature_threshold(feature_thresholds[2582]), .feature_above(feature_aboves[2582]), .feature_below(feature_belows[2582]), .scan_win_std_dev(scan_win_std_dev[2582]), .feature_accum(feature_accums[2582]));
  accum_calculator ac2583(.scan_win(scan_win2583), .rectangle1_x(rectangle1_xs[2583]), .rectangle1_y(rectangle1_ys[2583]), .rectangle1_width(rectangle1_widths[2583]), .rectangle1_height(rectangle1_heights[2583]), .rectangle1_weight(rectangle1_weights[2583]), .rectangle2_x(rectangle2_xs[2583]), .rectangle2_y(rectangle2_ys[2583]), .rectangle2_width(rectangle2_widths[2583]), .rectangle2_height(rectangle2_heights[2583]), .rectangle2_weight(rectangle2_weights[2583]), .rectangle3_x(rectangle3_xs[2583]), .rectangle3_y(rectangle3_ys[2583]), .rectangle3_width(rectangle3_widths[2583]), .rectangle3_height(rectangle3_heights[2583]), .rectangle3_weight(rectangle3_weights[2583]), .feature_threshold(feature_thresholds[2583]), .feature_above(feature_aboves[2583]), .feature_below(feature_belows[2583]), .scan_win_std_dev(scan_win_std_dev[2583]), .feature_accum(feature_accums[2583]));
  accum_calculator ac2584(.scan_win(scan_win2584), .rectangle1_x(rectangle1_xs[2584]), .rectangle1_y(rectangle1_ys[2584]), .rectangle1_width(rectangle1_widths[2584]), .rectangle1_height(rectangle1_heights[2584]), .rectangle1_weight(rectangle1_weights[2584]), .rectangle2_x(rectangle2_xs[2584]), .rectangle2_y(rectangle2_ys[2584]), .rectangle2_width(rectangle2_widths[2584]), .rectangle2_height(rectangle2_heights[2584]), .rectangle2_weight(rectangle2_weights[2584]), .rectangle3_x(rectangle3_xs[2584]), .rectangle3_y(rectangle3_ys[2584]), .rectangle3_width(rectangle3_widths[2584]), .rectangle3_height(rectangle3_heights[2584]), .rectangle3_weight(rectangle3_weights[2584]), .feature_threshold(feature_thresholds[2584]), .feature_above(feature_aboves[2584]), .feature_below(feature_belows[2584]), .scan_win_std_dev(scan_win_std_dev[2584]), .feature_accum(feature_accums[2584]));
  accum_calculator ac2585(.scan_win(scan_win2585), .rectangle1_x(rectangle1_xs[2585]), .rectangle1_y(rectangle1_ys[2585]), .rectangle1_width(rectangle1_widths[2585]), .rectangle1_height(rectangle1_heights[2585]), .rectangle1_weight(rectangle1_weights[2585]), .rectangle2_x(rectangle2_xs[2585]), .rectangle2_y(rectangle2_ys[2585]), .rectangle2_width(rectangle2_widths[2585]), .rectangle2_height(rectangle2_heights[2585]), .rectangle2_weight(rectangle2_weights[2585]), .rectangle3_x(rectangle3_xs[2585]), .rectangle3_y(rectangle3_ys[2585]), .rectangle3_width(rectangle3_widths[2585]), .rectangle3_height(rectangle3_heights[2585]), .rectangle3_weight(rectangle3_weights[2585]), .feature_threshold(feature_thresholds[2585]), .feature_above(feature_aboves[2585]), .feature_below(feature_belows[2585]), .scan_win_std_dev(scan_win_std_dev[2585]), .feature_accum(feature_accums[2585]));
  accum_calculator ac2586(.scan_win(scan_win2586), .rectangle1_x(rectangle1_xs[2586]), .rectangle1_y(rectangle1_ys[2586]), .rectangle1_width(rectangle1_widths[2586]), .rectangle1_height(rectangle1_heights[2586]), .rectangle1_weight(rectangle1_weights[2586]), .rectangle2_x(rectangle2_xs[2586]), .rectangle2_y(rectangle2_ys[2586]), .rectangle2_width(rectangle2_widths[2586]), .rectangle2_height(rectangle2_heights[2586]), .rectangle2_weight(rectangle2_weights[2586]), .rectangle3_x(rectangle3_xs[2586]), .rectangle3_y(rectangle3_ys[2586]), .rectangle3_width(rectangle3_widths[2586]), .rectangle3_height(rectangle3_heights[2586]), .rectangle3_weight(rectangle3_weights[2586]), .feature_threshold(feature_thresholds[2586]), .feature_above(feature_aboves[2586]), .feature_below(feature_belows[2586]), .scan_win_std_dev(scan_win_std_dev[2586]), .feature_accum(feature_accums[2586]));
  accum_calculator ac2587(.scan_win(scan_win2587), .rectangle1_x(rectangle1_xs[2587]), .rectangle1_y(rectangle1_ys[2587]), .rectangle1_width(rectangle1_widths[2587]), .rectangle1_height(rectangle1_heights[2587]), .rectangle1_weight(rectangle1_weights[2587]), .rectangle2_x(rectangle2_xs[2587]), .rectangle2_y(rectangle2_ys[2587]), .rectangle2_width(rectangle2_widths[2587]), .rectangle2_height(rectangle2_heights[2587]), .rectangle2_weight(rectangle2_weights[2587]), .rectangle3_x(rectangle3_xs[2587]), .rectangle3_y(rectangle3_ys[2587]), .rectangle3_width(rectangle3_widths[2587]), .rectangle3_height(rectangle3_heights[2587]), .rectangle3_weight(rectangle3_weights[2587]), .feature_threshold(feature_thresholds[2587]), .feature_above(feature_aboves[2587]), .feature_below(feature_belows[2587]), .scan_win_std_dev(scan_win_std_dev[2587]), .feature_accum(feature_accums[2587]));
  accum_calculator ac2588(.scan_win(scan_win2588), .rectangle1_x(rectangle1_xs[2588]), .rectangle1_y(rectangle1_ys[2588]), .rectangle1_width(rectangle1_widths[2588]), .rectangle1_height(rectangle1_heights[2588]), .rectangle1_weight(rectangle1_weights[2588]), .rectangle2_x(rectangle2_xs[2588]), .rectangle2_y(rectangle2_ys[2588]), .rectangle2_width(rectangle2_widths[2588]), .rectangle2_height(rectangle2_heights[2588]), .rectangle2_weight(rectangle2_weights[2588]), .rectangle3_x(rectangle3_xs[2588]), .rectangle3_y(rectangle3_ys[2588]), .rectangle3_width(rectangle3_widths[2588]), .rectangle3_height(rectangle3_heights[2588]), .rectangle3_weight(rectangle3_weights[2588]), .feature_threshold(feature_thresholds[2588]), .feature_above(feature_aboves[2588]), .feature_below(feature_belows[2588]), .scan_win_std_dev(scan_win_std_dev[2588]), .feature_accum(feature_accums[2588]));
  accum_calculator ac2589(.scan_win(scan_win2589), .rectangle1_x(rectangle1_xs[2589]), .rectangle1_y(rectangle1_ys[2589]), .rectangle1_width(rectangle1_widths[2589]), .rectangle1_height(rectangle1_heights[2589]), .rectangle1_weight(rectangle1_weights[2589]), .rectangle2_x(rectangle2_xs[2589]), .rectangle2_y(rectangle2_ys[2589]), .rectangle2_width(rectangle2_widths[2589]), .rectangle2_height(rectangle2_heights[2589]), .rectangle2_weight(rectangle2_weights[2589]), .rectangle3_x(rectangle3_xs[2589]), .rectangle3_y(rectangle3_ys[2589]), .rectangle3_width(rectangle3_widths[2589]), .rectangle3_height(rectangle3_heights[2589]), .rectangle3_weight(rectangle3_weights[2589]), .feature_threshold(feature_thresholds[2589]), .feature_above(feature_aboves[2589]), .feature_below(feature_belows[2589]), .scan_win_std_dev(scan_win_std_dev[2589]), .feature_accum(feature_accums[2589]));
  accum_calculator ac2590(.scan_win(scan_win2590), .rectangle1_x(rectangle1_xs[2590]), .rectangle1_y(rectangle1_ys[2590]), .rectangle1_width(rectangle1_widths[2590]), .rectangle1_height(rectangle1_heights[2590]), .rectangle1_weight(rectangle1_weights[2590]), .rectangle2_x(rectangle2_xs[2590]), .rectangle2_y(rectangle2_ys[2590]), .rectangle2_width(rectangle2_widths[2590]), .rectangle2_height(rectangle2_heights[2590]), .rectangle2_weight(rectangle2_weights[2590]), .rectangle3_x(rectangle3_xs[2590]), .rectangle3_y(rectangle3_ys[2590]), .rectangle3_width(rectangle3_widths[2590]), .rectangle3_height(rectangle3_heights[2590]), .rectangle3_weight(rectangle3_weights[2590]), .feature_threshold(feature_thresholds[2590]), .feature_above(feature_aboves[2590]), .feature_below(feature_belows[2590]), .scan_win_std_dev(scan_win_std_dev[2590]), .feature_accum(feature_accums[2590]));
  accum_calculator ac2591(.scan_win(scan_win2591), .rectangle1_x(rectangle1_xs[2591]), .rectangle1_y(rectangle1_ys[2591]), .rectangle1_width(rectangle1_widths[2591]), .rectangle1_height(rectangle1_heights[2591]), .rectangle1_weight(rectangle1_weights[2591]), .rectangle2_x(rectangle2_xs[2591]), .rectangle2_y(rectangle2_ys[2591]), .rectangle2_width(rectangle2_widths[2591]), .rectangle2_height(rectangle2_heights[2591]), .rectangle2_weight(rectangle2_weights[2591]), .rectangle3_x(rectangle3_xs[2591]), .rectangle3_y(rectangle3_ys[2591]), .rectangle3_width(rectangle3_widths[2591]), .rectangle3_height(rectangle3_heights[2591]), .rectangle3_weight(rectangle3_weights[2591]), .feature_threshold(feature_thresholds[2591]), .feature_above(feature_aboves[2591]), .feature_below(feature_belows[2591]), .scan_win_std_dev(scan_win_std_dev[2591]), .feature_accum(feature_accums[2591]));
  accum_calculator ac2592(.scan_win(scan_win2592), .rectangle1_x(rectangle1_xs[2592]), .rectangle1_y(rectangle1_ys[2592]), .rectangle1_width(rectangle1_widths[2592]), .rectangle1_height(rectangle1_heights[2592]), .rectangle1_weight(rectangle1_weights[2592]), .rectangle2_x(rectangle2_xs[2592]), .rectangle2_y(rectangle2_ys[2592]), .rectangle2_width(rectangle2_widths[2592]), .rectangle2_height(rectangle2_heights[2592]), .rectangle2_weight(rectangle2_weights[2592]), .rectangle3_x(rectangle3_xs[2592]), .rectangle3_y(rectangle3_ys[2592]), .rectangle3_width(rectangle3_widths[2592]), .rectangle3_height(rectangle3_heights[2592]), .rectangle3_weight(rectangle3_weights[2592]), .feature_threshold(feature_thresholds[2592]), .feature_above(feature_aboves[2592]), .feature_below(feature_belows[2592]), .scan_win_std_dev(scan_win_std_dev[2592]), .feature_accum(feature_accums[2592]));
  accum_calculator ac2593(.scan_win(scan_win2593), .rectangle1_x(rectangle1_xs[2593]), .rectangle1_y(rectangle1_ys[2593]), .rectangle1_width(rectangle1_widths[2593]), .rectangle1_height(rectangle1_heights[2593]), .rectangle1_weight(rectangle1_weights[2593]), .rectangle2_x(rectangle2_xs[2593]), .rectangle2_y(rectangle2_ys[2593]), .rectangle2_width(rectangle2_widths[2593]), .rectangle2_height(rectangle2_heights[2593]), .rectangle2_weight(rectangle2_weights[2593]), .rectangle3_x(rectangle3_xs[2593]), .rectangle3_y(rectangle3_ys[2593]), .rectangle3_width(rectangle3_widths[2593]), .rectangle3_height(rectangle3_heights[2593]), .rectangle3_weight(rectangle3_weights[2593]), .feature_threshold(feature_thresholds[2593]), .feature_above(feature_aboves[2593]), .feature_below(feature_belows[2593]), .scan_win_std_dev(scan_win_std_dev[2593]), .feature_accum(feature_accums[2593]));
  accum_calculator ac2594(.scan_win(scan_win2594), .rectangle1_x(rectangle1_xs[2594]), .rectangle1_y(rectangle1_ys[2594]), .rectangle1_width(rectangle1_widths[2594]), .rectangle1_height(rectangle1_heights[2594]), .rectangle1_weight(rectangle1_weights[2594]), .rectangle2_x(rectangle2_xs[2594]), .rectangle2_y(rectangle2_ys[2594]), .rectangle2_width(rectangle2_widths[2594]), .rectangle2_height(rectangle2_heights[2594]), .rectangle2_weight(rectangle2_weights[2594]), .rectangle3_x(rectangle3_xs[2594]), .rectangle3_y(rectangle3_ys[2594]), .rectangle3_width(rectangle3_widths[2594]), .rectangle3_height(rectangle3_heights[2594]), .rectangle3_weight(rectangle3_weights[2594]), .feature_threshold(feature_thresholds[2594]), .feature_above(feature_aboves[2594]), .feature_below(feature_belows[2594]), .scan_win_std_dev(scan_win_std_dev[2594]), .feature_accum(feature_accums[2594]));
  accum_calculator ac2595(.scan_win(scan_win2595), .rectangle1_x(rectangle1_xs[2595]), .rectangle1_y(rectangle1_ys[2595]), .rectangle1_width(rectangle1_widths[2595]), .rectangle1_height(rectangle1_heights[2595]), .rectangle1_weight(rectangle1_weights[2595]), .rectangle2_x(rectangle2_xs[2595]), .rectangle2_y(rectangle2_ys[2595]), .rectangle2_width(rectangle2_widths[2595]), .rectangle2_height(rectangle2_heights[2595]), .rectangle2_weight(rectangle2_weights[2595]), .rectangle3_x(rectangle3_xs[2595]), .rectangle3_y(rectangle3_ys[2595]), .rectangle3_width(rectangle3_widths[2595]), .rectangle3_height(rectangle3_heights[2595]), .rectangle3_weight(rectangle3_weights[2595]), .feature_threshold(feature_thresholds[2595]), .feature_above(feature_aboves[2595]), .feature_below(feature_belows[2595]), .scan_win_std_dev(scan_win_std_dev[2595]), .feature_accum(feature_accums[2595]));
  accum_calculator ac2596(.scan_win(scan_win2596), .rectangle1_x(rectangle1_xs[2596]), .rectangle1_y(rectangle1_ys[2596]), .rectangle1_width(rectangle1_widths[2596]), .rectangle1_height(rectangle1_heights[2596]), .rectangle1_weight(rectangle1_weights[2596]), .rectangle2_x(rectangle2_xs[2596]), .rectangle2_y(rectangle2_ys[2596]), .rectangle2_width(rectangle2_widths[2596]), .rectangle2_height(rectangle2_heights[2596]), .rectangle2_weight(rectangle2_weights[2596]), .rectangle3_x(rectangle3_xs[2596]), .rectangle3_y(rectangle3_ys[2596]), .rectangle3_width(rectangle3_widths[2596]), .rectangle3_height(rectangle3_heights[2596]), .rectangle3_weight(rectangle3_weights[2596]), .feature_threshold(feature_thresholds[2596]), .feature_above(feature_aboves[2596]), .feature_below(feature_belows[2596]), .scan_win_std_dev(scan_win_std_dev[2596]), .feature_accum(feature_accums[2596]));
  accum_calculator ac2597(.scan_win(scan_win2597), .rectangle1_x(rectangle1_xs[2597]), .rectangle1_y(rectangle1_ys[2597]), .rectangle1_width(rectangle1_widths[2597]), .rectangle1_height(rectangle1_heights[2597]), .rectangle1_weight(rectangle1_weights[2597]), .rectangle2_x(rectangle2_xs[2597]), .rectangle2_y(rectangle2_ys[2597]), .rectangle2_width(rectangle2_widths[2597]), .rectangle2_height(rectangle2_heights[2597]), .rectangle2_weight(rectangle2_weights[2597]), .rectangle3_x(rectangle3_xs[2597]), .rectangle3_y(rectangle3_ys[2597]), .rectangle3_width(rectangle3_widths[2597]), .rectangle3_height(rectangle3_heights[2597]), .rectangle3_weight(rectangle3_weights[2597]), .feature_threshold(feature_thresholds[2597]), .feature_above(feature_aboves[2597]), .feature_below(feature_belows[2597]), .scan_win_std_dev(scan_win_std_dev[2597]), .feature_accum(feature_accums[2597]));
  accum_calculator ac2598(.scan_win(scan_win2598), .rectangle1_x(rectangle1_xs[2598]), .rectangle1_y(rectangle1_ys[2598]), .rectangle1_width(rectangle1_widths[2598]), .rectangle1_height(rectangle1_heights[2598]), .rectangle1_weight(rectangle1_weights[2598]), .rectangle2_x(rectangle2_xs[2598]), .rectangle2_y(rectangle2_ys[2598]), .rectangle2_width(rectangle2_widths[2598]), .rectangle2_height(rectangle2_heights[2598]), .rectangle2_weight(rectangle2_weights[2598]), .rectangle3_x(rectangle3_xs[2598]), .rectangle3_y(rectangle3_ys[2598]), .rectangle3_width(rectangle3_widths[2598]), .rectangle3_height(rectangle3_heights[2598]), .rectangle3_weight(rectangle3_weights[2598]), .feature_threshold(feature_thresholds[2598]), .feature_above(feature_aboves[2598]), .feature_below(feature_belows[2598]), .scan_win_std_dev(scan_win_std_dev[2598]), .feature_accum(feature_accums[2598]));
  accum_calculator ac2599(.scan_win(scan_win2599), .rectangle1_x(rectangle1_xs[2599]), .rectangle1_y(rectangle1_ys[2599]), .rectangle1_width(rectangle1_widths[2599]), .rectangle1_height(rectangle1_heights[2599]), .rectangle1_weight(rectangle1_weights[2599]), .rectangle2_x(rectangle2_xs[2599]), .rectangle2_y(rectangle2_ys[2599]), .rectangle2_width(rectangle2_widths[2599]), .rectangle2_height(rectangle2_heights[2599]), .rectangle2_weight(rectangle2_weights[2599]), .rectangle3_x(rectangle3_xs[2599]), .rectangle3_y(rectangle3_ys[2599]), .rectangle3_width(rectangle3_widths[2599]), .rectangle3_height(rectangle3_heights[2599]), .rectangle3_weight(rectangle3_weights[2599]), .feature_threshold(feature_thresholds[2599]), .feature_above(feature_aboves[2599]), .feature_below(feature_belows[2599]), .scan_win_std_dev(scan_win_std_dev[2599]), .feature_accum(feature_accums[2599]));
  accum_calculator ac2600(.scan_win(scan_win2600), .rectangle1_x(rectangle1_xs[2600]), .rectangle1_y(rectangle1_ys[2600]), .rectangle1_width(rectangle1_widths[2600]), .rectangle1_height(rectangle1_heights[2600]), .rectangle1_weight(rectangle1_weights[2600]), .rectangle2_x(rectangle2_xs[2600]), .rectangle2_y(rectangle2_ys[2600]), .rectangle2_width(rectangle2_widths[2600]), .rectangle2_height(rectangle2_heights[2600]), .rectangle2_weight(rectangle2_weights[2600]), .rectangle3_x(rectangle3_xs[2600]), .rectangle3_y(rectangle3_ys[2600]), .rectangle3_width(rectangle3_widths[2600]), .rectangle3_height(rectangle3_heights[2600]), .rectangle3_weight(rectangle3_weights[2600]), .feature_threshold(feature_thresholds[2600]), .feature_above(feature_aboves[2600]), .feature_below(feature_belows[2600]), .scan_win_std_dev(scan_win_std_dev[2600]), .feature_accum(feature_accums[2600]));
  accum_calculator ac2601(.scan_win(scan_win2601), .rectangle1_x(rectangle1_xs[2601]), .rectangle1_y(rectangle1_ys[2601]), .rectangle1_width(rectangle1_widths[2601]), .rectangle1_height(rectangle1_heights[2601]), .rectangle1_weight(rectangle1_weights[2601]), .rectangle2_x(rectangle2_xs[2601]), .rectangle2_y(rectangle2_ys[2601]), .rectangle2_width(rectangle2_widths[2601]), .rectangle2_height(rectangle2_heights[2601]), .rectangle2_weight(rectangle2_weights[2601]), .rectangle3_x(rectangle3_xs[2601]), .rectangle3_y(rectangle3_ys[2601]), .rectangle3_width(rectangle3_widths[2601]), .rectangle3_height(rectangle3_heights[2601]), .rectangle3_weight(rectangle3_weights[2601]), .feature_threshold(feature_thresholds[2601]), .feature_above(feature_aboves[2601]), .feature_below(feature_belows[2601]), .scan_win_std_dev(scan_win_std_dev[2601]), .feature_accum(feature_accums[2601]));
  accum_calculator ac2602(.scan_win(scan_win2602), .rectangle1_x(rectangle1_xs[2602]), .rectangle1_y(rectangle1_ys[2602]), .rectangle1_width(rectangle1_widths[2602]), .rectangle1_height(rectangle1_heights[2602]), .rectangle1_weight(rectangle1_weights[2602]), .rectangle2_x(rectangle2_xs[2602]), .rectangle2_y(rectangle2_ys[2602]), .rectangle2_width(rectangle2_widths[2602]), .rectangle2_height(rectangle2_heights[2602]), .rectangle2_weight(rectangle2_weights[2602]), .rectangle3_x(rectangle3_xs[2602]), .rectangle3_y(rectangle3_ys[2602]), .rectangle3_width(rectangle3_widths[2602]), .rectangle3_height(rectangle3_heights[2602]), .rectangle3_weight(rectangle3_weights[2602]), .feature_threshold(feature_thresholds[2602]), .feature_above(feature_aboves[2602]), .feature_below(feature_belows[2602]), .scan_win_std_dev(scan_win_std_dev[2602]), .feature_accum(feature_accums[2602]));
  accum_calculator ac2603(.scan_win(scan_win2603), .rectangle1_x(rectangle1_xs[2603]), .rectangle1_y(rectangle1_ys[2603]), .rectangle1_width(rectangle1_widths[2603]), .rectangle1_height(rectangle1_heights[2603]), .rectangle1_weight(rectangle1_weights[2603]), .rectangle2_x(rectangle2_xs[2603]), .rectangle2_y(rectangle2_ys[2603]), .rectangle2_width(rectangle2_widths[2603]), .rectangle2_height(rectangle2_heights[2603]), .rectangle2_weight(rectangle2_weights[2603]), .rectangle3_x(rectangle3_xs[2603]), .rectangle3_y(rectangle3_ys[2603]), .rectangle3_width(rectangle3_widths[2603]), .rectangle3_height(rectangle3_heights[2603]), .rectangle3_weight(rectangle3_weights[2603]), .feature_threshold(feature_thresholds[2603]), .feature_above(feature_aboves[2603]), .feature_below(feature_belows[2603]), .scan_win_std_dev(scan_win_std_dev[2603]), .feature_accum(feature_accums[2603]));
  accum_calculator ac2604(.scan_win(scan_win2604), .rectangle1_x(rectangle1_xs[2604]), .rectangle1_y(rectangle1_ys[2604]), .rectangle1_width(rectangle1_widths[2604]), .rectangle1_height(rectangle1_heights[2604]), .rectangle1_weight(rectangle1_weights[2604]), .rectangle2_x(rectangle2_xs[2604]), .rectangle2_y(rectangle2_ys[2604]), .rectangle2_width(rectangle2_widths[2604]), .rectangle2_height(rectangle2_heights[2604]), .rectangle2_weight(rectangle2_weights[2604]), .rectangle3_x(rectangle3_xs[2604]), .rectangle3_y(rectangle3_ys[2604]), .rectangle3_width(rectangle3_widths[2604]), .rectangle3_height(rectangle3_heights[2604]), .rectangle3_weight(rectangle3_weights[2604]), .feature_threshold(feature_thresholds[2604]), .feature_above(feature_aboves[2604]), .feature_below(feature_belows[2604]), .scan_win_std_dev(scan_win_std_dev[2604]), .feature_accum(feature_accums[2604]));
  accum_calculator ac2605(.scan_win(scan_win2605), .rectangle1_x(rectangle1_xs[2605]), .rectangle1_y(rectangle1_ys[2605]), .rectangle1_width(rectangle1_widths[2605]), .rectangle1_height(rectangle1_heights[2605]), .rectangle1_weight(rectangle1_weights[2605]), .rectangle2_x(rectangle2_xs[2605]), .rectangle2_y(rectangle2_ys[2605]), .rectangle2_width(rectangle2_widths[2605]), .rectangle2_height(rectangle2_heights[2605]), .rectangle2_weight(rectangle2_weights[2605]), .rectangle3_x(rectangle3_xs[2605]), .rectangle3_y(rectangle3_ys[2605]), .rectangle3_width(rectangle3_widths[2605]), .rectangle3_height(rectangle3_heights[2605]), .rectangle3_weight(rectangle3_weights[2605]), .feature_threshold(feature_thresholds[2605]), .feature_above(feature_aboves[2605]), .feature_below(feature_belows[2605]), .scan_win_std_dev(scan_win_std_dev[2605]), .feature_accum(feature_accums[2605]));
  accum_calculator ac2606(.scan_win(scan_win2606), .rectangle1_x(rectangle1_xs[2606]), .rectangle1_y(rectangle1_ys[2606]), .rectangle1_width(rectangle1_widths[2606]), .rectangle1_height(rectangle1_heights[2606]), .rectangle1_weight(rectangle1_weights[2606]), .rectangle2_x(rectangle2_xs[2606]), .rectangle2_y(rectangle2_ys[2606]), .rectangle2_width(rectangle2_widths[2606]), .rectangle2_height(rectangle2_heights[2606]), .rectangle2_weight(rectangle2_weights[2606]), .rectangle3_x(rectangle3_xs[2606]), .rectangle3_y(rectangle3_ys[2606]), .rectangle3_width(rectangle3_widths[2606]), .rectangle3_height(rectangle3_heights[2606]), .rectangle3_weight(rectangle3_weights[2606]), .feature_threshold(feature_thresholds[2606]), .feature_above(feature_aboves[2606]), .feature_below(feature_belows[2606]), .scan_win_std_dev(scan_win_std_dev[2606]), .feature_accum(feature_accums[2606]));
  accum_calculator ac2607(.scan_win(scan_win2607), .rectangle1_x(rectangle1_xs[2607]), .rectangle1_y(rectangle1_ys[2607]), .rectangle1_width(rectangle1_widths[2607]), .rectangle1_height(rectangle1_heights[2607]), .rectangle1_weight(rectangle1_weights[2607]), .rectangle2_x(rectangle2_xs[2607]), .rectangle2_y(rectangle2_ys[2607]), .rectangle2_width(rectangle2_widths[2607]), .rectangle2_height(rectangle2_heights[2607]), .rectangle2_weight(rectangle2_weights[2607]), .rectangle3_x(rectangle3_xs[2607]), .rectangle3_y(rectangle3_ys[2607]), .rectangle3_width(rectangle3_widths[2607]), .rectangle3_height(rectangle3_heights[2607]), .rectangle3_weight(rectangle3_weights[2607]), .feature_threshold(feature_thresholds[2607]), .feature_above(feature_aboves[2607]), .feature_below(feature_belows[2607]), .scan_win_std_dev(scan_win_std_dev[2607]), .feature_accum(feature_accums[2607]));
  accum_calculator ac2608(.scan_win(scan_win2608), .rectangle1_x(rectangle1_xs[2608]), .rectangle1_y(rectangle1_ys[2608]), .rectangle1_width(rectangle1_widths[2608]), .rectangle1_height(rectangle1_heights[2608]), .rectangle1_weight(rectangle1_weights[2608]), .rectangle2_x(rectangle2_xs[2608]), .rectangle2_y(rectangle2_ys[2608]), .rectangle2_width(rectangle2_widths[2608]), .rectangle2_height(rectangle2_heights[2608]), .rectangle2_weight(rectangle2_weights[2608]), .rectangle3_x(rectangle3_xs[2608]), .rectangle3_y(rectangle3_ys[2608]), .rectangle3_width(rectangle3_widths[2608]), .rectangle3_height(rectangle3_heights[2608]), .rectangle3_weight(rectangle3_weights[2608]), .feature_threshold(feature_thresholds[2608]), .feature_above(feature_aboves[2608]), .feature_below(feature_belows[2608]), .scan_win_std_dev(scan_win_std_dev[2608]), .feature_accum(feature_accums[2608]));
  accum_calculator ac2609(.scan_win(scan_win2609), .rectangle1_x(rectangle1_xs[2609]), .rectangle1_y(rectangle1_ys[2609]), .rectangle1_width(rectangle1_widths[2609]), .rectangle1_height(rectangle1_heights[2609]), .rectangle1_weight(rectangle1_weights[2609]), .rectangle2_x(rectangle2_xs[2609]), .rectangle2_y(rectangle2_ys[2609]), .rectangle2_width(rectangle2_widths[2609]), .rectangle2_height(rectangle2_heights[2609]), .rectangle2_weight(rectangle2_weights[2609]), .rectangle3_x(rectangle3_xs[2609]), .rectangle3_y(rectangle3_ys[2609]), .rectangle3_width(rectangle3_widths[2609]), .rectangle3_height(rectangle3_heights[2609]), .rectangle3_weight(rectangle3_weights[2609]), .feature_threshold(feature_thresholds[2609]), .feature_above(feature_aboves[2609]), .feature_below(feature_belows[2609]), .scan_win_std_dev(scan_win_std_dev[2609]), .feature_accum(feature_accums[2609]));
  accum_calculator ac2610(.scan_win(scan_win2610), .rectangle1_x(rectangle1_xs[2610]), .rectangle1_y(rectangle1_ys[2610]), .rectangle1_width(rectangle1_widths[2610]), .rectangle1_height(rectangle1_heights[2610]), .rectangle1_weight(rectangle1_weights[2610]), .rectangle2_x(rectangle2_xs[2610]), .rectangle2_y(rectangle2_ys[2610]), .rectangle2_width(rectangle2_widths[2610]), .rectangle2_height(rectangle2_heights[2610]), .rectangle2_weight(rectangle2_weights[2610]), .rectangle3_x(rectangle3_xs[2610]), .rectangle3_y(rectangle3_ys[2610]), .rectangle3_width(rectangle3_widths[2610]), .rectangle3_height(rectangle3_heights[2610]), .rectangle3_weight(rectangle3_weights[2610]), .feature_threshold(feature_thresholds[2610]), .feature_above(feature_aboves[2610]), .feature_below(feature_belows[2610]), .scan_win_std_dev(scan_win_std_dev[2610]), .feature_accum(feature_accums[2610]));
  accum_calculator ac2611(.scan_win(scan_win2611), .rectangle1_x(rectangle1_xs[2611]), .rectangle1_y(rectangle1_ys[2611]), .rectangle1_width(rectangle1_widths[2611]), .rectangle1_height(rectangle1_heights[2611]), .rectangle1_weight(rectangle1_weights[2611]), .rectangle2_x(rectangle2_xs[2611]), .rectangle2_y(rectangle2_ys[2611]), .rectangle2_width(rectangle2_widths[2611]), .rectangle2_height(rectangle2_heights[2611]), .rectangle2_weight(rectangle2_weights[2611]), .rectangle3_x(rectangle3_xs[2611]), .rectangle3_y(rectangle3_ys[2611]), .rectangle3_width(rectangle3_widths[2611]), .rectangle3_height(rectangle3_heights[2611]), .rectangle3_weight(rectangle3_weights[2611]), .feature_threshold(feature_thresholds[2611]), .feature_above(feature_aboves[2611]), .feature_below(feature_belows[2611]), .scan_win_std_dev(scan_win_std_dev[2611]), .feature_accum(feature_accums[2611]));
  accum_calculator ac2612(.scan_win(scan_win2612), .rectangle1_x(rectangle1_xs[2612]), .rectangle1_y(rectangle1_ys[2612]), .rectangle1_width(rectangle1_widths[2612]), .rectangle1_height(rectangle1_heights[2612]), .rectangle1_weight(rectangle1_weights[2612]), .rectangle2_x(rectangle2_xs[2612]), .rectangle2_y(rectangle2_ys[2612]), .rectangle2_width(rectangle2_widths[2612]), .rectangle2_height(rectangle2_heights[2612]), .rectangle2_weight(rectangle2_weights[2612]), .rectangle3_x(rectangle3_xs[2612]), .rectangle3_y(rectangle3_ys[2612]), .rectangle3_width(rectangle3_widths[2612]), .rectangle3_height(rectangle3_heights[2612]), .rectangle3_weight(rectangle3_weights[2612]), .feature_threshold(feature_thresholds[2612]), .feature_above(feature_aboves[2612]), .feature_below(feature_belows[2612]), .scan_win_std_dev(scan_win_std_dev[2612]), .feature_accum(feature_accums[2612]));
  accum_calculator ac2613(.scan_win(scan_win2613), .rectangle1_x(rectangle1_xs[2613]), .rectangle1_y(rectangle1_ys[2613]), .rectangle1_width(rectangle1_widths[2613]), .rectangle1_height(rectangle1_heights[2613]), .rectangle1_weight(rectangle1_weights[2613]), .rectangle2_x(rectangle2_xs[2613]), .rectangle2_y(rectangle2_ys[2613]), .rectangle2_width(rectangle2_widths[2613]), .rectangle2_height(rectangle2_heights[2613]), .rectangle2_weight(rectangle2_weights[2613]), .rectangle3_x(rectangle3_xs[2613]), .rectangle3_y(rectangle3_ys[2613]), .rectangle3_width(rectangle3_widths[2613]), .rectangle3_height(rectangle3_heights[2613]), .rectangle3_weight(rectangle3_weights[2613]), .feature_threshold(feature_thresholds[2613]), .feature_above(feature_aboves[2613]), .feature_below(feature_belows[2613]), .scan_win_std_dev(scan_win_std_dev[2613]), .feature_accum(feature_accums[2613]));
  accum_calculator ac2614(.scan_win(scan_win2614), .rectangle1_x(rectangle1_xs[2614]), .rectangle1_y(rectangle1_ys[2614]), .rectangle1_width(rectangle1_widths[2614]), .rectangle1_height(rectangle1_heights[2614]), .rectangle1_weight(rectangle1_weights[2614]), .rectangle2_x(rectangle2_xs[2614]), .rectangle2_y(rectangle2_ys[2614]), .rectangle2_width(rectangle2_widths[2614]), .rectangle2_height(rectangle2_heights[2614]), .rectangle2_weight(rectangle2_weights[2614]), .rectangle3_x(rectangle3_xs[2614]), .rectangle3_y(rectangle3_ys[2614]), .rectangle3_width(rectangle3_widths[2614]), .rectangle3_height(rectangle3_heights[2614]), .rectangle3_weight(rectangle3_weights[2614]), .feature_threshold(feature_thresholds[2614]), .feature_above(feature_aboves[2614]), .feature_below(feature_belows[2614]), .scan_win_std_dev(scan_win_std_dev[2614]), .feature_accum(feature_accums[2614]));
  accum_calculator ac2615(.scan_win(scan_win2615), .rectangle1_x(rectangle1_xs[2615]), .rectangle1_y(rectangle1_ys[2615]), .rectangle1_width(rectangle1_widths[2615]), .rectangle1_height(rectangle1_heights[2615]), .rectangle1_weight(rectangle1_weights[2615]), .rectangle2_x(rectangle2_xs[2615]), .rectangle2_y(rectangle2_ys[2615]), .rectangle2_width(rectangle2_widths[2615]), .rectangle2_height(rectangle2_heights[2615]), .rectangle2_weight(rectangle2_weights[2615]), .rectangle3_x(rectangle3_xs[2615]), .rectangle3_y(rectangle3_ys[2615]), .rectangle3_width(rectangle3_widths[2615]), .rectangle3_height(rectangle3_heights[2615]), .rectangle3_weight(rectangle3_weights[2615]), .feature_threshold(feature_thresholds[2615]), .feature_above(feature_aboves[2615]), .feature_below(feature_belows[2615]), .scan_win_std_dev(scan_win_std_dev[2615]), .feature_accum(feature_accums[2615]));
  accum_calculator ac2616(.scan_win(scan_win2616), .rectangle1_x(rectangle1_xs[2616]), .rectangle1_y(rectangle1_ys[2616]), .rectangle1_width(rectangle1_widths[2616]), .rectangle1_height(rectangle1_heights[2616]), .rectangle1_weight(rectangle1_weights[2616]), .rectangle2_x(rectangle2_xs[2616]), .rectangle2_y(rectangle2_ys[2616]), .rectangle2_width(rectangle2_widths[2616]), .rectangle2_height(rectangle2_heights[2616]), .rectangle2_weight(rectangle2_weights[2616]), .rectangle3_x(rectangle3_xs[2616]), .rectangle3_y(rectangle3_ys[2616]), .rectangle3_width(rectangle3_widths[2616]), .rectangle3_height(rectangle3_heights[2616]), .rectangle3_weight(rectangle3_weights[2616]), .feature_threshold(feature_thresholds[2616]), .feature_above(feature_aboves[2616]), .feature_below(feature_belows[2616]), .scan_win_std_dev(scan_win_std_dev[2616]), .feature_accum(feature_accums[2616]));
  accum_calculator ac2617(.scan_win(scan_win2617), .rectangle1_x(rectangle1_xs[2617]), .rectangle1_y(rectangle1_ys[2617]), .rectangle1_width(rectangle1_widths[2617]), .rectangle1_height(rectangle1_heights[2617]), .rectangle1_weight(rectangle1_weights[2617]), .rectangle2_x(rectangle2_xs[2617]), .rectangle2_y(rectangle2_ys[2617]), .rectangle2_width(rectangle2_widths[2617]), .rectangle2_height(rectangle2_heights[2617]), .rectangle2_weight(rectangle2_weights[2617]), .rectangle3_x(rectangle3_xs[2617]), .rectangle3_y(rectangle3_ys[2617]), .rectangle3_width(rectangle3_widths[2617]), .rectangle3_height(rectangle3_heights[2617]), .rectangle3_weight(rectangle3_weights[2617]), .feature_threshold(feature_thresholds[2617]), .feature_above(feature_aboves[2617]), .feature_below(feature_belows[2617]), .scan_win_std_dev(scan_win_std_dev[2617]), .feature_accum(feature_accums[2617]));
  accum_calculator ac2618(.scan_win(scan_win2618), .rectangle1_x(rectangle1_xs[2618]), .rectangle1_y(rectangle1_ys[2618]), .rectangle1_width(rectangle1_widths[2618]), .rectangle1_height(rectangle1_heights[2618]), .rectangle1_weight(rectangle1_weights[2618]), .rectangle2_x(rectangle2_xs[2618]), .rectangle2_y(rectangle2_ys[2618]), .rectangle2_width(rectangle2_widths[2618]), .rectangle2_height(rectangle2_heights[2618]), .rectangle2_weight(rectangle2_weights[2618]), .rectangle3_x(rectangle3_xs[2618]), .rectangle3_y(rectangle3_ys[2618]), .rectangle3_width(rectangle3_widths[2618]), .rectangle3_height(rectangle3_heights[2618]), .rectangle3_weight(rectangle3_weights[2618]), .feature_threshold(feature_thresholds[2618]), .feature_above(feature_aboves[2618]), .feature_below(feature_belows[2618]), .scan_win_std_dev(scan_win_std_dev[2618]), .feature_accum(feature_accums[2618]));
  accum_calculator ac2619(.scan_win(scan_win2619), .rectangle1_x(rectangle1_xs[2619]), .rectangle1_y(rectangle1_ys[2619]), .rectangle1_width(rectangle1_widths[2619]), .rectangle1_height(rectangle1_heights[2619]), .rectangle1_weight(rectangle1_weights[2619]), .rectangle2_x(rectangle2_xs[2619]), .rectangle2_y(rectangle2_ys[2619]), .rectangle2_width(rectangle2_widths[2619]), .rectangle2_height(rectangle2_heights[2619]), .rectangle2_weight(rectangle2_weights[2619]), .rectangle3_x(rectangle3_xs[2619]), .rectangle3_y(rectangle3_ys[2619]), .rectangle3_width(rectangle3_widths[2619]), .rectangle3_height(rectangle3_heights[2619]), .rectangle3_weight(rectangle3_weights[2619]), .feature_threshold(feature_thresholds[2619]), .feature_above(feature_aboves[2619]), .feature_below(feature_belows[2619]), .scan_win_std_dev(scan_win_std_dev[2619]), .feature_accum(feature_accums[2619]));
  accum_calculator ac2620(.scan_win(scan_win2620), .rectangle1_x(rectangle1_xs[2620]), .rectangle1_y(rectangle1_ys[2620]), .rectangle1_width(rectangle1_widths[2620]), .rectangle1_height(rectangle1_heights[2620]), .rectangle1_weight(rectangle1_weights[2620]), .rectangle2_x(rectangle2_xs[2620]), .rectangle2_y(rectangle2_ys[2620]), .rectangle2_width(rectangle2_widths[2620]), .rectangle2_height(rectangle2_heights[2620]), .rectangle2_weight(rectangle2_weights[2620]), .rectangle3_x(rectangle3_xs[2620]), .rectangle3_y(rectangle3_ys[2620]), .rectangle3_width(rectangle3_widths[2620]), .rectangle3_height(rectangle3_heights[2620]), .rectangle3_weight(rectangle3_weights[2620]), .feature_threshold(feature_thresholds[2620]), .feature_above(feature_aboves[2620]), .feature_below(feature_belows[2620]), .scan_win_std_dev(scan_win_std_dev[2620]), .feature_accum(feature_accums[2620]));
  accum_calculator ac2621(.scan_win(scan_win2621), .rectangle1_x(rectangle1_xs[2621]), .rectangle1_y(rectangle1_ys[2621]), .rectangle1_width(rectangle1_widths[2621]), .rectangle1_height(rectangle1_heights[2621]), .rectangle1_weight(rectangle1_weights[2621]), .rectangle2_x(rectangle2_xs[2621]), .rectangle2_y(rectangle2_ys[2621]), .rectangle2_width(rectangle2_widths[2621]), .rectangle2_height(rectangle2_heights[2621]), .rectangle2_weight(rectangle2_weights[2621]), .rectangle3_x(rectangle3_xs[2621]), .rectangle3_y(rectangle3_ys[2621]), .rectangle3_width(rectangle3_widths[2621]), .rectangle3_height(rectangle3_heights[2621]), .rectangle3_weight(rectangle3_weights[2621]), .feature_threshold(feature_thresholds[2621]), .feature_above(feature_aboves[2621]), .feature_below(feature_belows[2621]), .scan_win_std_dev(scan_win_std_dev[2621]), .feature_accum(feature_accums[2621]));
  accum_calculator ac2622(.scan_win(scan_win2622), .rectangle1_x(rectangle1_xs[2622]), .rectangle1_y(rectangle1_ys[2622]), .rectangle1_width(rectangle1_widths[2622]), .rectangle1_height(rectangle1_heights[2622]), .rectangle1_weight(rectangle1_weights[2622]), .rectangle2_x(rectangle2_xs[2622]), .rectangle2_y(rectangle2_ys[2622]), .rectangle2_width(rectangle2_widths[2622]), .rectangle2_height(rectangle2_heights[2622]), .rectangle2_weight(rectangle2_weights[2622]), .rectangle3_x(rectangle3_xs[2622]), .rectangle3_y(rectangle3_ys[2622]), .rectangle3_width(rectangle3_widths[2622]), .rectangle3_height(rectangle3_heights[2622]), .rectangle3_weight(rectangle3_weights[2622]), .feature_threshold(feature_thresholds[2622]), .feature_above(feature_aboves[2622]), .feature_below(feature_belows[2622]), .scan_win_std_dev(scan_win_std_dev[2622]), .feature_accum(feature_accums[2622]));
  accum_calculator ac2623(.scan_win(scan_win2623), .rectangle1_x(rectangle1_xs[2623]), .rectangle1_y(rectangle1_ys[2623]), .rectangle1_width(rectangle1_widths[2623]), .rectangle1_height(rectangle1_heights[2623]), .rectangle1_weight(rectangle1_weights[2623]), .rectangle2_x(rectangle2_xs[2623]), .rectangle2_y(rectangle2_ys[2623]), .rectangle2_width(rectangle2_widths[2623]), .rectangle2_height(rectangle2_heights[2623]), .rectangle2_weight(rectangle2_weights[2623]), .rectangle3_x(rectangle3_xs[2623]), .rectangle3_y(rectangle3_ys[2623]), .rectangle3_width(rectangle3_widths[2623]), .rectangle3_height(rectangle3_heights[2623]), .rectangle3_weight(rectangle3_weights[2623]), .feature_threshold(feature_thresholds[2623]), .feature_above(feature_aboves[2623]), .feature_below(feature_belows[2623]), .scan_win_std_dev(scan_win_std_dev[2623]), .feature_accum(feature_accums[2623]));
  accum_calculator ac2624(.scan_win(scan_win2624), .rectangle1_x(rectangle1_xs[2624]), .rectangle1_y(rectangle1_ys[2624]), .rectangle1_width(rectangle1_widths[2624]), .rectangle1_height(rectangle1_heights[2624]), .rectangle1_weight(rectangle1_weights[2624]), .rectangle2_x(rectangle2_xs[2624]), .rectangle2_y(rectangle2_ys[2624]), .rectangle2_width(rectangle2_widths[2624]), .rectangle2_height(rectangle2_heights[2624]), .rectangle2_weight(rectangle2_weights[2624]), .rectangle3_x(rectangle3_xs[2624]), .rectangle3_y(rectangle3_ys[2624]), .rectangle3_width(rectangle3_widths[2624]), .rectangle3_height(rectangle3_heights[2624]), .rectangle3_weight(rectangle3_weights[2624]), .feature_threshold(feature_thresholds[2624]), .feature_above(feature_aboves[2624]), .feature_below(feature_belows[2624]), .scan_win_std_dev(scan_win_std_dev[2624]), .feature_accum(feature_accums[2624]));
  accum_calculator ac2625(.scan_win(scan_win2625), .rectangle1_x(rectangle1_xs[2625]), .rectangle1_y(rectangle1_ys[2625]), .rectangle1_width(rectangle1_widths[2625]), .rectangle1_height(rectangle1_heights[2625]), .rectangle1_weight(rectangle1_weights[2625]), .rectangle2_x(rectangle2_xs[2625]), .rectangle2_y(rectangle2_ys[2625]), .rectangle2_width(rectangle2_widths[2625]), .rectangle2_height(rectangle2_heights[2625]), .rectangle2_weight(rectangle2_weights[2625]), .rectangle3_x(rectangle3_xs[2625]), .rectangle3_y(rectangle3_ys[2625]), .rectangle3_width(rectangle3_widths[2625]), .rectangle3_height(rectangle3_heights[2625]), .rectangle3_weight(rectangle3_weights[2625]), .feature_threshold(feature_thresholds[2625]), .feature_above(feature_aboves[2625]), .feature_below(feature_belows[2625]), .scan_win_std_dev(scan_win_std_dev[2625]), .feature_accum(feature_accums[2625]));
  accum_calculator ac2626(.scan_win(scan_win2626), .rectangle1_x(rectangle1_xs[2626]), .rectangle1_y(rectangle1_ys[2626]), .rectangle1_width(rectangle1_widths[2626]), .rectangle1_height(rectangle1_heights[2626]), .rectangle1_weight(rectangle1_weights[2626]), .rectangle2_x(rectangle2_xs[2626]), .rectangle2_y(rectangle2_ys[2626]), .rectangle2_width(rectangle2_widths[2626]), .rectangle2_height(rectangle2_heights[2626]), .rectangle2_weight(rectangle2_weights[2626]), .rectangle3_x(rectangle3_xs[2626]), .rectangle3_y(rectangle3_ys[2626]), .rectangle3_width(rectangle3_widths[2626]), .rectangle3_height(rectangle3_heights[2626]), .rectangle3_weight(rectangle3_weights[2626]), .feature_threshold(feature_thresholds[2626]), .feature_above(feature_aboves[2626]), .feature_below(feature_belows[2626]), .scan_win_std_dev(scan_win_std_dev[2626]), .feature_accum(feature_accums[2626]));
  accum_calculator ac2627(.scan_win(scan_win2627), .rectangle1_x(rectangle1_xs[2627]), .rectangle1_y(rectangle1_ys[2627]), .rectangle1_width(rectangle1_widths[2627]), .rectangle1_height(rectangle1_heights[2627]), .rectangle1_weight(rectangle1_weights[2627]), .rectangle2_x(rectangle2_xs[2627]), .rectangle2_y(rectangle2_ys[2627]), .rectangle2_width(rectangle2_widths[2627]), .rectangle2_height(rectangle2_heights[2627]), .rectangle2_weight(rectangle2_weights[2627]), .rectangle3_x(rectangle3_xs[2627]), .rectangle3_y(rectangle3_ys[2627]), .rectangle3_width(rectangle3_widths[2627]), .rectangle3_height(rectangle3_heights[2627]), .rectangle3_weight(rectangle3_weights[2627]), .feature_threshold(feature_thresholds[2627]), .feature_above(feature_aboves[2627]), .feature_below(feature_belows[2627]), .scan_win_std_dev(scan_win_std_dev[2627]), .feature_accum(feature_accums[2627]));
  accum_calculator ac2628(.scan_win(scan_win2628), .rectangle1_x(rectangle1_xs[2628]), .rectangle1_y(rectangle1_ys[2628]), .rectangle1_width(rectangle1_widths[2628]), .rectangle1_height(rectangle1_heights[2628]), .rectangle1_weight(rectangle1_weights[2628]), .rectangle2_x(rectangle2_xs[2628]), .rectangle2_y(rectangle2_ys[2628]), .rectangle2_width(rectangle2_widths[2628]), .rectangle2_height(rectangle2_heights[2628]), .rectangle2_weight(rectangle2_weights[2628]), .rectangle3_x(rectangle3_xs[2628]), .rectangle3_y(rectangle3_ys[2628]), .rectangle3_width(rectangle3_widths[2628]), .rectangle3_height(rectangle3_heights[2628]), .rectangle3_weight(rectangle3_weights[2628]), .feature_threshold(feature_thresholds[2628]), .feature_above(feature_aboves[2628]), .feature_below(feature_belows[2628]), .scan_win_std_dev(scan_win_std_dev[2628]), .feature_accum(feature_accums[2628]));
  accum_calculator ac2629(.scan_win(scan_win2629), .rectangle1_x(rectangle1_xs[2629]), .rectangle1_y(rectangle1_ys[2629]), .rectangle1_width(rectangle1_widths[2629]), .rectangle1_height(rectangle1_heights[2629]), .rectangle1_weight(rectangle1_weights[2629]), .rectangle2_x(rectangle2_xs[2629]), .rectangle2_y(rectangle2_ys[2629]), .rectangle2_width(rectangle2_widths[2629]), .rectangle2_height(rectangle2_heights[2629]), .rectangle2_weight(rectangle2_weights[2629]), .rectangle3_x(rectangle3_xs[2629]), .rectangle3_y(rectangle3_ys[2629]), .rectangle3_width(rectangle3_widths[2629]), .rectangle3_height(rectangle3_heights[2629]), .rectangle3_weight(rectangle3_weights[2629]), .feature_threshold(feature_thresholds[2629]), .feature_above(feature_aboves[2629]), .feature_below(feature_belows[2629]), .scan_win_std_dev(scan_win_std_dev[2629]), .feature_accum(feature_accums[2629]));
  accum_calculator ac2630(.scan_win(scan_win2630), .rectangle1_x(rectangle1_xs[2630]), .rectangle1_y(rectangle1_ys[2630]), .rectangle1_width(rectangle1_widths[2630]), .rectangle1_height(rectangle1_heights[2630]), .rectangle1_weight(rectangle1_weights[2630]), .rectangle2_x(rectangle2_xs[2630]), .rectangle2_y(rectangle2_ys[2630]), .rectangle2_width(rectangle2_widths[2630]), .rectangle2_height(rectangle2_heights[2630]), .rectangle2_weight(rectangle2_weights[2630]), .rectangle3_x(rectangle3_xs[2630]), .rectangle3_y(rectangle3_ys[2630]), .rectangle3_width(rectangle3_widths[2630]), .rectangle3_height(rectangle3_heights[2630]), .rectangle3_weight(rectangle3_weights[2630]), .feature_threshold(feature_thresholds[2630]), .feature_above(feature_aboves[2630]), .feature_below(feature_belows[2630]), .scan_win_std_dev(scan_win_std_dev[2630]), .feature_accum(feature_accums[2630]));
  accum_calculator ac2631(.scan_win(scan_win2631), .rectangle1_x(rectangle1_xs[2631]), .rectangle1_y(rectangle1_ys[2631]), .rectangle1_width(rectangle1_widths[2631]), .rectangle1_height(rectangle1_heights[2631]), .rectangle1_weight(rectangle1_weights[2631]), .rectangle2_x(rectangle2_xs[2631]), .rectangle2_y(rectangle2_ys[2631]), .rectangle2_width(rectangle2_widths[2631]), .rectangle2_height(rectangle2_heights[2631]), .rectangle2_weight(rectangle2_weights[2631]), .rectangle3_x(rectangle3_xs[2631]), .rectangle3_y(rectangle3_ys[2631]), .rectangle3_width(rectangle3_widths[2631]), .rectangle3_height(rectangle3_heights[2631]), .rectangle3_weight(rectangle3_weights[2631]), .feature_threshold(feature_thresholds[2631]), .feature_above(feature_aboves[2631]), .feature_below(feature_belows[2631]), .scan_win_std_dev(scan_win_std_dev[2631]), .feature_accum(feature_accums[2631]));
  accum_calculator ac2632(.scan_win(scan_win2632), .rectangle1_x(rectangle1_xs[2632]), .rectangle1_y(rectangle1_ys[2632]), .rectangle1_width(rectangle1_widths[2632]), .rectangle1_height(rectangle1_heights[2632]), .rectangle1_weight(rectangle1_weights[2632]), .rectangle2_x(rectangle2_xs[2632]), .rectangle2_y(rectangle2_ys[2632]), .rectangle2_width(rectangle2_widths[2632]), .rectangle2_height(rectangle2_heights[2632]), .rectangle2_weight(rectangle2_weights[2632]), .rectangle3_x(rectangle3_xs[2632]), .rectangle3_y(rectangle3_ys[2632]), .rectangle3_width(rectangle3_widths[2632]), .rectangle3_height(rectangle3_heights[2632]), .rectangle3_weight(rectangle3_weights[2632]), .feature_threshold(feature_thresholds[2632]), .feature_above(feature_aboves[2632]), .feature_below(feature_belows[2632]), .scan_win_std_dev(scan_win_std_dev[2632]), .feature_accum(feature_accums[2632]));
  accum_calculator ac2633(.scan_win(scan_win2633), .rectangle1_x(rectangle1_xs[2633]), .rectangle1_y(rectangle1_ys[2633]), .rectangle1_width(rectangle1_widths[2633]), .rectangle1_height(rectangle1_heights[2633]), .rectangle1_weight(rectangle1_weights[2633]), .rectangle2_x(rectangle2_xs[2633]), .rectangle2_y(rectangle2_ys[2633]), .rectangle2_width(rectangle2_widths[2633]), .rectangle2_height(rectangle2_heights[2633]), .rectangle2_weight(rectangle2_weights[2633]), .rectangle3_x(rectangle3_xs[2633]), .rectangle3_y(rectangle3_ys[2633]), .rectangle3_width(rectangle3_widths[2633]), .rectangle3_height(rectangle3_heights[2633]), .rectangle3_weight(rectangle3_weights[2633]), .feature_threshold(feature_thresholds[2633]), .feature_above(feature_aboves[2633]), .feature_below(feature_belows[2633]), .scan_win_std_dev(scan_win_std_dev[2633]), .feature_accum(feature_accums[2633]));
  accum_calculator ac2634(.scan_win(scan_win2634), .rectangle1_x(rectangle1_xs[2634]), .rectangle1_y(rectangle1_ys[2634]), .rectangle1_width(rectangle1_widths[2634]), .rectangle1_height(rectangle1_heights[2634]), .rectangle1_weight(rectangle1_weights[2634]), .rectangle2_x(rectangle2_xs[2634]), .rectangle2_y(rectangle2_ys[2634]), .rectangle2_width(rectangle2_widths[2634]), .rectangle2_height(rectangle2_heights[2634]), .rectangle2_weight(rectangle2_weights[2634]), .rectangle3_x(rectangle3_xs[2634]), .rectangle3_y(rectangle3_ys[2634]), .rectangle3_width(rectangle3_widths[2634]), .rectangle3_height(rectangle3_heights[2634]), .rectangle3_weight(rectangle3_weights[2634]), .feature_threshold(feature_thresholds[2634]), .feature_above(feature_aboves[2634]), .feature_below(feature_belows[2634]), .scan_win_std_dev(scan_win_std_dev[2634]), .feature_accum(feature_accums[2634]));
  accum_calculator ac2635(.scan_win(scan_win2635), .rectangle1_x(rectangle1_xs[2635]), .rectangle1_y(rectangle1_ys[2635]), .rectangle1_width(rectangle1_widths[2635]), .rectangle1_height(rectangle1_heights[2635]), .rectangle1_weight(rectangle1_weights[2635]), .rectangle2_x(rectangle2_xs[2635]), .rectangle2_y(rectangle2_ys[2635]), .rectangle2_width(rectangle2_widths[2635]), .rectangle2_height(rectangle2_heights[2635]), .rectangle2_weight(rectangle2_weights[2635]), .rectangle3_x(rectangle3_xs[2635]), .rectangle3_y(rectangle3_ys[2635]), .rectangle3_width(rectangle3_widths[2635]), .rectangle3_height(rectangle3_heights[2635]), .rectangle3_weight(rectangle3_weights[2635]), .feature_threshold(feature_thresholds[2635]), .feature_above(feature_aboves[2635]), .feature_below(feature_belows[2635]), .scan_win_std_dev(scan_win_std_dev[2635]), .feature_accum(feature_accums[2635]));
  accum_calculator ac2636(.scan_win(scan_win2636), .rectangle1_x(rectangle1_xs[2636]), .rectangle1_y(rectangle1_ys[2636]), .rectangle1_width(rectangle1_widths[2636]), .rectangle1_height(rectangle1_heights[2636]), .rectangle1_weight(rectangle1_weights[2636]), .rectangle2_x(rectangle2_xs[2636]), .rectangle2_y(rectangle2_ys[2636]), .rectangle2_width(rectangle2_widths[2636]), .rectangle2_height(rectangle2_heights[2636]), .rectangle2_weight(rectangle2_weights[2636]), .rectangle3_x(rectangle3_xs[2636]), .rectangle3_y(rectangle3_ys[2636]), .rectangle3_width(rectangle3_widths[2636]), .rectangle3_height(rectangle3_heights[2636]), .rectangle3_weight(rectangle3_weights[2636]), .feature_threshold(feature_thresholds[2636]), .feature_above(feature_aboves[2636]), .feature_below(feature_belows[2636]), .scan_win_std_dev(scan_win_std_dev[2636]), .feature_accum(feature_accums[2636]));
  accum_calculator ac2637(.scan_win(scan_win2637), .rectangle1_x(rectangle1_xs[2637]), .rectangle1_y(rectangle1_ys[2637]), .rectangle1_width(rectangle1_widths[2637]), .rectangle1_height(rectangle1_heights[2637]), .rectangle1_weight(rectangle1_weights[2637]), .rectangle2_x(rectangle2_xs[2637]), .rectangle2_y(rectangle2_ys[2637]), .rectangle2_width(rectangle2_widths[2637]), .rectangle2_height(rectangle2_heights[2637]), .rectangle2_weight(rectangle2_weights[2637]), .rectangle3_x(rectangle3_xs[2637]), .rectangle3_y(rectangle3_ys[2637]), .rectangle3_width(rectangle3_widths[2637]), .rectangle3_height(rectangle3_heights[2637]), .rectangle3_weight(rectangle3_weights[2637]), .feature_threshold(feature_thresholds[2637]), .feature_above(feature_aboves[2637]), .feature_below(feature_belows[2637]), .scan_win_std_dev(scan_win_std_dev[2637]), .feature_accum(feature_accums[2637]));
  accum_calculator ac2638(.scan_win(scan_win2638), .rectangle1_x(rectangle1_xs[2638]), .rectangle1_y(rectangle1_ys[2638]), .rectangle1_width(rectangle1_widths[2638]), .rectangle1_height(rectangle1_heights[2638]), .rectangle1_weight(rectangle1_weights[2638]), .rectangle2_x(rectangle2_xs[2638]), .rectangle2_y(rectangle2_ys[2638]), .rectangle2_width(rectangle2_widths[2638]), .rectangle2_height(rectangle2_heights[2638]), .rectangle2_weight(rectangle2_weights[2638]), .rectangle3_x(rectangle3_xs[2638]), .rectangle3_y(rectangle3_ys[2638]), .rectangle3_width(rectangle3_widths[2638]), .rectangle3_height(rectangle3_heights[2638]), .rectangle3_weight(rectangle3_weights[2638]), .feature_threshold(feature_thresholds[2638]), .feature_above(feature_aboves[2638]), .feature_below(feature_belows[2638]), .scan_win_std_dev(scan_win_std_dev[2638]), .feature_accum(feature_accums[2638]));
  accum_calculator ac2639(.scan_win(scan_win2639), .rectangle1_x(rectangle1_xs[2639]), .rectangle1_y(rectangle1_ys[2639]), .rectangle1_width(rectangle1_widths[2639]), .rectangle1_height(rectangle1_heights[2639]), .rectangle1_weight(rectangle1_weights[2639]), .rectangle2_x(rectangle2_xs[2639]), .rectangle2_y(rectangle2_ys[2639]), .rectangle2_width(rectangle2_widths[2639]), .rectangle2_height(rectangle2_heights[2639]), .rectangle2_weight(rectangle2_weights[2639]), .rectangle3_x(rectangle3_xs[2639]), .rectangle3_y(rectangle3_ys[2639]), .rectangle3_width(rectangle3_widths[2639]), .rectangle3_height(rectangle3_heights[2639]), .rectangle3_weight(rectangle3_weights[2639]), .feature_threshold(feature_thresholds[2639]), .feature_above(feature_aboves[2639]), .feature_below(feature_belows[2639]), .scan_win_std_dev(scan_win_std_dev[2639]), .feature_accum(feature_accums[2639]));
  accum_calculator ac2640(.scan_win(scan_win2640), .rectangle1_x(rectangle1_xs[2640]), .rectangle1_y(rectangle1_ys[2640]), .rectangle1_width(rectangle1_widths[2640]), .rectangle1_height(rectangle1_heights[2640]), .rectangle1_weight(rectangle1_weights[2640]), .rectangle2_x(rectangle2_xs[2640]), .rectangle2_y(rectangle2_ys[2640]), .rectangle2_width(rectangle2_widths[2640]), .rectangle2_height(rectangle2_heights[2640]), .rectangle2_weight(rectangle2_weights[2640]), .rectangle3_x(rectangle3_xs[2640]), .rectangle3_y(rectangle3_ys[2640]), .rectangle3_width(rectangle3_widths[2640]), .rectangle3_height(rectangle3_heights[2640]), .rectangle3_weight(rectangle3_weights[2640]), .feature_threshold(feature_thresholds[2640]), .feature_above(feature_aboves[2640]), .feature_below(feature_belows[2640]), .scan_win_std_dev(scan_win_std_dev[2640]), .feature_accum(feature_accums[2640]));
  accum_calculator ac2641(.scan_win(scan_win2641), .rectangle1_x(rectangle1_xs[2641]), .rectangle1_y(rectangle1_ys[2641]), .rectangle1_width(rectangle1_widths[2641]), .rectangle1_height(rectangle1_heights[2641]), .rectangle1_weight(rectangle1_weights[2641]), .rectangle2_x(rectangle2_xs[2641]), .rectangle2_y(rectangle2_ys[2641]), .rectangle2_width(rectangle2_widths[2641]), .rectangle2_height(rectangle2_heights[2641]), .rectangle2_weight(rectangle2_weights[2641]), .rectangle3_x(rectangle3_xs[2641]), .rectangle3_y(rectangle3_ys[2641]), .rectangle3_width(rectangle3_widths[2641]), .rectangle3_height(rectangle3_heights[2641]), .rectangle3_weight(rectangle3_weights[2641]), .feature_threshold(feature_thresholds[2641]), .feature_above(feature_aboves[2641]), .feature_below(feature_belows[2641]), .scan_win_std_dev(scan_win_std_dev[2641]), .feature_accum(feature_accums[2641]));
  accum_calculator ac2642(.scan_win(scan_win2642), .rectangle1_x(rectangle1_xs[2642]), .rectangle1_y(rectangle1_ys[2642]), .rectangle1_width(rectangle1_widths[2642]), .rectangle1_height(rectangle1_heights[2642]), .rectangle1_weight(rectangle1_weights[2642]), .rectangle2_x(rectangle2_xs[2642]), .rectangle2_y(rectangle2_ys[2642]), .rectangle2_width(rectangle2_widths[2642]), .rectangle2_height(rectangle2_heights[2642]), .rectangle2_weight(rectangle2_weights[2642]), .rectangle3_x(rectangle3_xs[2642]), .rectangle3_y(rectangle3_ys[2642]), .rectangle3_width(rectangle3_widths[2642]), .rectangle3_height(rectangle3_heights[2642]), .rectangle3_weight(rectangle3_weights[2642]), .feature_threshold(feature_thresholds[2642]), .feature_above(feature_aboves[2642]), .feature_below(feature_belows[2642]), .scan_win_std_dev(scan_win_std_dev[2642]), .feature_accum(feature_accums[2642]));
  accum_calculator ac2643(.scan_win(scan_win2643), .rectangle1_x(rectangle1_xs[2643]), .rectangle1_y(rectangle1_ys[2643]), .rectangle1_width(rectangle1_widths[2643]), .rectangle1_height(rectangle1_heights[2643]), .rectangle1_weight(rectangle1_weights[2643]), .rectangle2_x(rectangle2_xs[2643]), .rectangle2_y(rectangle2_ys[2643]), .rectangle2_width(rectangle2_widths[2643]), .rectangle2_height(rectangle2_heights[2643]), .rectangle2_weight(rectangle2_weights[2643]), .rectangle3_x(rectangle3_xs[2643]), .rectangle3_y(rectangle3_ys[2643]), .rectangle3_width(rectangle3_widths[2643]), .rectangle3_height(rectangle3_heights[2643]), .rectangle3_weight(rectangle3_weights[2643]), .feature_threshold(feature_thresholds[2643]), .feature_above(feature_aboves[2643]), .feature_below(feature_belows[2643]), .scan_win_std_dev(scan_win_std_dev[2643]), .feature_accum(feature_accums[2643]));
  accum_calculator ac2644(.scan_win(scan_win2644), .rectangle1_x(rectangle1_xs[2644]), .rectangle1_y(rectangle1_ys[2644]), .rectangle1_width(rectangle1_widths[2644]), .rectangle1_height(rectangle1_heights[2644]), .rectangle1_weight(rectangle1_weights[2644]), .rectangle2_x(rectangle2_xs[2644]), .rectangle2_y(rectangle2_ys[2644]), .rectangle2_width(rectangle2_widths[2644]), .rectangle2_height(rectangle2_heights[2644]), .rectangle2_weight(rectangle2_weights[2644]), .rectangle3_x(rectangle3_xs[2644]), .rectangle3_y(rectangle3_ys[2644]), .rectangle3_width(rectangle3_widths[2644]), .rectangle3_height(rectangle3_heights[2644]), .rectangle3_weight(rectangle3_weights[2644]), .feature_threshold(feature_thresholds[2644]), .feature_above(feature_aboves[2644]), .feature_below(feature_belows[2644]), .scan_win_std_dev(scan_win_std_dev[2644]), .feature_accum(feature_accums[2644]));
  accum_calculator ac2645(.scan_win(scan_win2645), .rectangle1_x(rectangle1_xs[2645]), .rectangle1_y(rectangle1_ys[2645]), .rectangle1_width(rectangle1_widths[2645]), .rectangle1_height(rectangle1_heights[2645]), .rectangle1_weight(rectangle1_weights[2645]), .rectangle2_x(rectangle2_xs[2645]), .rectangle2_y(rectangle2_ys[2645]), .rectangle2_width(rectangle2_widths[2645]), .rectangle2_height(rectangle2_heights[2645]), .rectangle2_weight(rectangle2_weights[2645]), .rectangle3_x(rectangle3_xs[2645]), .rectangle3_y(rectangle3_ys[2645]), .rectangle3_width(rectangle3_widths[2645]), .rectangle3_height(rectangle3_heights[2645]), .rectangle3_weight(rectangle3_weights[2645]), .feature_threshold(feature_thresholds[2645]), .feature_above(feature_aboves[2645]), .feature_below(feature_belows[2645]), .scan_win_std_dev(scan_win_std_dev[2645]), .feature_accum(feature_accums[2645]));
  accum_calculator ac2646(.scan_win(scan_win2646), .rectangle1_x(rectangle1_xs[2646]), .rectangle1_y(rectangle1_ys[2646]), .rectangle1_width(rectangle1_widths[2646]), .rectangle1_height(rectangle1_heights[2646]), .rectangle1_weight(rectangle1_weights[2646]), .rectangle2_x(rectangle2_xs[2646]), .rectangle2_y(rectangle2_ys[2646]), .rectangle2_width(rectangle2_widths[2646]), .rectangle2_height(rectangle2_heights[2646]), .rectangle2_weight(rectangle2_weights[2646]), .rectangle3_x(rectangle3_xs[2646]), .rectangle3_y(rectangle3_ys[2646]), .rectangle3_width(rectangle3_widths[2646]), .rectangle3_height(rectangle3_heights[2646]), .rectangle3_weight(rectangle3_weights[2646]), .feature_threshold(feature_thresholds[2646]), .feature_above(feature_aboves[2646]), .feature_below(feature_belows[2646]), .scan_win_std_dev(scan_win_std_dev[2646]), .feature_accum(feature_accums[2646]));
  accum_calculator ac2647(.scan_win(scan_win2647), .rectangle1_x(rectangle1_xs[2647]), .rectangle1_y(rectangle1_ys[2647]), .rectangle1_width(rectangle1_widths[2647]), .rectangle1_height(rectangle1_heights[2647]), .rectangle1_weight(rectangle1_weights[2647]), .rectangle2_x(rectangle2_xs[2647]), .rectangle2_y(rectangle2_ys[2647]), .rectangle2_width(rectangle2_widths[2647]), .rectangle2_height(rectangle2_heights[2647]), .rectangle2_weight(rectangle2_weights[2647]), .rectangle3_x(rectangle3_xs[2647]), .rectangle3_y(rectangle3_ys[2647]), .rectangle3_width(rectangle3_widths[2647]), .rectangle3_height(rectangle3_heights[2647]), .rectangle3_weight(rectangle3_weights[2647]), .feature_threshold(feature_thresholds[2647]), .feature_above(feature_aboves[2647]), .feature_below(feature_belows[2647]), .scan_win_std_dev(scan_win_std_dev[2647]), .feature_accum(feature_accums[2647]));
  accum_calculator ac2648(.scan_win(scan_win2648), .rectangle1_x(rectangle1_xs[2648]), .rectangle1_y(rectangle1_ys[2648]), .rectangle1_width(rectangle1_widths[2648]), .rectangle1_height(rectangle1_heights[2648]), .rectangle1_weight(rectangle1_weights[2648]), .rectangle2_x(rectangle2_xs[2648]), .rectangle2_y(rectangle2_ys[2648]), .rectangle2_width(rectangle2_widths[2648]), .rectangle2_height(rectangle2_heights[2648]), .rectangle2_weight(rectangle2_weights[2648]), .rectangle3_x(rectangle3_xs[2648]), .rectangle3_y(rectangle3_ys[2648]), .rectangle3_width(rectangle3_widths[2648]), .rectangle3_height(rectangle3_heights[2648]), .rectangle3_weight(rectangle3_weights[2648]), .feature_threshold(feature_thresholds[2648]), .feature_above(feature_aboves[2648]), .feature_below(feature_belows[2648]), .scan_win_std_dev(scan_win_std_dev[2648]), .feature_accum(feature_accums[2648]));
  accum_calculator ac2649(.scan_win(scan_win2649), .rectangle1_x(rectangle1_xs[2649]), .rectangle1_y(rectangle1_ys[2649]), .rectangle1_width(rectangle1_widths[2649]), .rectangle1_height(rectangle1_heights[2649]), .rectangle1_weight(rectangle1_weights[2649]), .rectangle2_x(rectangle2_xs[2649]), .rectangle2_y(rectangle2_ys[2649]), .rectangle2_width(rectangle2_widths[2649]), .rectangle2_height(rectangle2_heights[2649]), .rectangle2_weight(rectangle2_weights[2649]), .rectangle3_x(rectangle3_xs[2649]), .rectangle3_y(rectangle3_ys[2649]), .rectangle3_width(rectangle3_widths[2649]), .rectangle3_height(rectangle3_heights[2649]), .rectangle3_weight(rectangle3_weights[2649]), .feature_threshold(feature_thresholds[2649]), .feature_above(feature_aboves[2649]), .feature_below(feature_belows[2649]), .scan_win_std_dev(scan_win_std_dev[2649]), .feature_accum(feature_accums[2649]));
  accum_calculator ac2650(.scan_win(scan_win2650), .rectangle1_x(rectangle1_xs[2650]), .rectangle1_y(rectangle1_ys[2650]), .rectangle1_width(rectangle1_widths[2650]), .rectangle1_height(rectangle1_heights[2650]), .rectangle1_weight(rectangle1_weights[2650]), .rectangle2_x(rectangle2_xs[2650]), .rectangle2_y(rectangle2_ys[2650]), .rectangle2_width(rectangle2_widths[2650]), .rectangle2_height(rectangle2_heights[2650]), .rectangle2_weight(rectangle2_weights[2650]), .rectangle3_x(rectangle3_xs[2650]), .rectangle3_y(rectangle3_ys[2650]), .rectangle3_width(rectangle3_widths[2650]), .rectangle3_height(rectangle3_heights[2650]), .rectangle3_weight(rectangle3_weights[2650]), .feature_threshold(feature_thresholds[2650]), .feature_above(feature_aboves[2650]), .feature_below(feature_belows[2650]), .scan_win_std_dev(scan_win_std_dev[2650]), .feature_accum(feature_accums[2650]));
  accum_calculator ac2651(.scan_win(scan_win2651), .rectangle1_x(rectangle1_xs[2651]), .rectangle1_y(rectangle1_ys[2651]), .rectangle1_width(rectangle1_widths[2651]), .rectangle1_height(rectangle1_heights[2651]), .rectangle1_weight(rectangle1_weights[2651]), .rectangle2_x(rectangle2_xs[2651]), .rectangle2_y(rectangle2_ys[2651]), .rectangle2_width(rectangle2_widths[2651]), .rectangle2_height(rectangle2_heights[2651]), .rectangle2_weight(rectangle2_weights[2651]), .rectangle3_x(rectangle3_xs[2651]), .rectangle3_y(rectangle3_ys[2651]), .rectangle3_width(rectangle3_widths[2651]), .rectangle3_height(rectangle3_heights[2651]), .rectangle3_weight(rectangle3_weights[2651]), .feature_threshold(feature_thresholds[2651]), .feature_above(feature_aboves[2651]), .feature_below(feature_belows[2651]), .scan_win_std_dev(scan_win_std_dev[2651]), .feature_accum(feature_accums[2651]));
  accum_calculator ac2652(.scan_win(scan_win2652), .rectangle1_x(rectangle1_xs[2652]), .rectangle1_y(rectangle1_ys[2652]), .rectangle1_width(rectangle1_widths[2652]), .rectangle1_height(rectangle1_heights[2652]), .rectangle1_weight(rectangle1_weights[2652]), .rectangle2_x(rectangle2_xs[2652]), .rectangle2_y(rectangle2_ys[2652]), .rectangle2_width(rectangle2_widths[2652]), .rectangle2_height(rectangle2_heights[2652]), .rectangle2_weight(rectangle2_weights[2652]), .rectangle3_x(rectangle3_xs[2652]), .rectangle3_y(rectangle3_ys[2652]), .rectangle3_width(rectangle3_widths[2652]), .rectangle3_height(rectangle3_heights[2652]), .rectangle3_weight(rectangle3_weights[2652]), .feature_threshold(feature_thresholds[2652]), .feature_above(feature_aboves[2652]), .feature_below(feature_belows[2652]), .scan_win_std_dev(scan_win_std_dev[2652]), .feature_accum(feature_accums[2652]));
  accum_calculator ac2653(.scan_win(scan_win2653), .rectangle1_x(rectangle1_xs[2653]), .rectangle1_y(rectangle1_ys[2653]), .rectangle1_width(rectangle1_widths[2653]), .rectangle1_height(rectangle1_heights[2653]), .rectangle1_weight(rectangle1_weights[2653]), .rectangle2_x(rectangle2_xs[2653]), .rectangle2_y(rectangle2_ys[2653]), .rectangle2_width(rectangle2_widths[2653]), .rectangle2_height(rectangle2_heights[2653]), .rectangle2_weight(rectangle2_weights[2653]), .rectangle3_x(rectangle3_xs[2653]), .rectangle3_y(rectangle3_ys[2653]), .rectangle3_width(rectangle3_widths[2653]), .rectangle3_height(rectangle3_heights[2653]), .rectangle3_weight(rectangle3_weights[2653]), .feature_threshold(feature_thresholds[2653]), .feature_above(feature_aboves[2653]), .feature_below(feature_belows[2653]), .scan_win_std_dev(scan_win_std_dev[2653]), .feature_accum(feature_accums[2653]));
  accum_calculator ac2654(.scan_win(scan_win2654), .rectangle1_x(rectangle1_xs[2654]), .rectangle1_y(rectangle1_ys[2654]), .rectangle1_width(rectangle1_widths[2654]), .rectangle1_height(rectangle1_heights[2654]), .rectangle1_weight(rectangle1_weights[2654]), .rectangle2_x(rectangle2_xs[2654]), .rectangle2_y(rectangle2_ys[2654]), .rectangle2_width(rectangle2_widths[2654]), .rectangle2_height(rectangle2_heights[2654]), .rectangle2_weight(rectangle2_weights[2654]), .rectangle3_x(rectangle3_xs[2654]), .rectangle3_y(rectangle3_ys[2654]), .rectangle3_width(rectangle3_widths[2654]), .rectangle3_height(rectangle3_heights[2654]), .rectangle3_weight(rectangle3_weights[2654]), .feature_threshold(feature_thresholds[2654]), .feature_above(feature_aboves[2654]), .feature_below(feature_belows[2654]), .scan_win_std_dev(scan_win_std_dev[2654]), .feature_accum(feature_accums[2654]));
  accum_calculator ac2655(.scan_win(scan_win2655), .rectangle1_x(rectangle1_xs[2655]), .rectangle1_y(rectangle1_ys[2655]), .rectangle1_width(rectangle1_widths[2655]), .rectangle1_height(rectangle1_heights[2655]), .rectangle1_weight(rectangle1_weights[2655]), .rectangle2_x(rectangle2_xs[2655]), .rectangle2_y(rectangle2_ys[2655]), .rectangle2_width(rectangle2_widths[2655]), .rectangle2_height(rectangle2_heights[2655]), .rectangle2_weight(rectangle2_weights[2655]), .rectangle3_x(rectangle3_xs[2655]), .rectangle3_y(rectangle3_ys[2655]), .rectangle3_width(rectangle3_widths[2655]), .rectangle3_height(rectangle3_heights[2655]), .rectangle3_weight(rectangle3_weights[2655]), .feature_threshold(feature_thresholds[2655]), .feature_above(feature_aboves[2655]), .feature_below(feature_belows[2655]), .scan_win_std_dev(scan_win_std_dev[2655]), .feature_accum(feature_accums[2655]));
  accum_calculator ac2656(.scan_win(scan_win2656), .rectangle1_x(rectangle1_xs[2656]), .rectangle1_y(rectangle1_ys[2656]), .rectangle1_width(rectangle1_widths[2656]), .rectangle1_height(rectangle1_heights[2656]), .rectangle1_weight(rectangle1_weights[2656]), .rectangle2_x(rectangle2_xs[2656]), .rectangle2_y(rectangle2_ys[2656]), .rectangle2_width(rectangle2_widths[2656]), .rectangle2_height(rectangle2_heights[2656]), .rectangle2_weight(rectangle2_weights[2656]), .rectangle3_x(rectangle3_xs[2656]), .rectangle3_y(rectangle3_ys[2656]), .rectangle3_width(rectangle3_widths[2656]), .rectangle3_height(rectangle3_heights[2656]), .rectangle3_weight(rectangle3_weights[2656]), .feature_threshold(feature_thresholds[2656]), .feature_above(feature_aboves[2656]), .feature_below(feature_belows[2656]), .scan_win_std_dev(scan_win_std_dev[2656]), .feature_accum(feature_accums[2656]));
  accum_calculator ac2657(.scan_win(scan_win2657), .rectangle1_x(rectangle1_xs[2657]), .rectangle1_y(rectangle1_ys[2657]), .rectangle1_width(rectangle1_widths[2657]), .rectangle1_height(rectangle1_heights[2657]), .rectangle1_weight(rectangle1_weights[2657]), .rectangle2_x(rectangle2_xs[2657]), .rectangle2_y(rectangle2_ys[2657]), .rectangle2_width(rectangle2_widths[2657]), .rectangle2_height(rectangle2_heights[2657]), .rectangle2_weight(rectangle2_weights[2657]), .rectangle3_x(rectangle3_xs[2657]), .rectangle3_y(rectangle3_ys[2657]), .rectangle3_width(rectangle3_widths[2657]), .rectangle3_height(rectangle3_heights[2657]), .rectangle3_weight(rectangle3_weights[2657]), .feature_threshold(feature_thresholds[2657]), .feature_above(feature_aboves[2657]), .feature_below(feature_belows[2657]), .scan_win_std_dev(scan_win_std_dev[2657]), .feature_accum(feature_accums[2657]));
  accum_calculator ac2658(.scan_win(scan_win2658), .rectangle1_x(rectangle1_xs[2658]), .rectangle1_y(rectangle1_ys[2658]), .rectangle1_width(rectangle1_widths[2658]), .rectangle1_height(rectangle1_heights[2658]), .rectangle1_weight(rectangle1_weights[2658]), .rectangle2_x(rectangle2_xs[2658]), .rectangle2_y(rectangle2_ys[2658]), .rectangle2_width(rectangle2_widths[2658]), .rectangle2_height(rectangle2_heights[2658]), .rectangle2_weight(rectangle2_weights[2658]), .rectangle3_x(rectangle3_xs[2658]), .rectangle3_y(rectangle3_ys[2658]), .rectangle3_width(rectangle3_widths[2658]), .rectangle3_height(rectangle3_heights[2658]), .rectangle3_weight(rectangle3_weights[2658]), .feature_threshold(feature_thresholds[2658]), .feature_above(feature_aboves[2658]), .feature_below(feature_belows[2658]), .scan_win_std_dev(scan_win_std_dev[2658]), .feature_accum(feature_accums[2658]));
  accum_calculator ac2659(.scan_win(scan_win2659), .rectangle1_x(rectangle1_xs[2659]), .rectangle1_y(rectangle1_ys[2659]), .rectangle1_width(rectangle1_widths[2659]), .rectangle1_height(rectangle1_heights[2659]), .rectangle1_weight(rectangle1_weights[2659]), .rectangle2_x(rectangle2_xs[2659]), .rectangle2_y(rectangle2_ys[2659]), .rectangle2_width(rectangle2_widths[2659]), .rectangle2_height(rectangle2_heights[2659]), .rectangle2_weight(rectangle2_weights[2659]), .rectangle3_x(rectangle3_xs[2659]), .rectangle3_y(rectangle3_ys[2659]), .rectangle3_width(rectangle3_widths[2659]), .rectangle3_height(rectangle3_heights[2659]), .rectangle3_weight(rectangle3_weights[2659]), .feature_threshold(feature_thresholds[2659]), .feature_above(feature_aboves[2659]), .feature_below(feature_belows[2659]), .scan_win_std_dev(scan_win_std_dev[2659]), .feature_accum(feature_accums[2659]));
  accum_calculator ac2660(.scan_win(scan_win2660), .rectangle1_x(rectangle1_xs[2660]), .rectangle1_y(rectangle1_ys[2660]), .rectangle1_width(rectangle1_widths[2660]), .rectangle1_height(rectangle1_heights[2660]), .rectangle1_weight(rectangle1_weights[2660]), .rectangle2_x(rectangle2_xs[2660]), .rectangle2_y(rectangle2_ys[2660]), .rectangle2_width(rectangle2_widths[2660]), .rectangle2_height(rectangle2_heights[2660]), .rectangle2_weight(rectangle2_weights[2660]), .rectangle3_x(rectangle3_xs[2660]), .rectangle3_y(rectangle3_ys[2660]), .rectangle3_width(rectangle3_widths[2660]), .rectangle3_height(rectangle3_heights[2660]), .rectangle3_weight(rectangle3_weights[2660]), .feature_threshold(feature_thresholds[2660]), .feature_above(feature_aboves[2660]), .feature_below(feature_belows[2660]), .scan_win_std_dev(scan_win_std_dev[2660]), .feature_accum(feature_accums[2660]));
  accum_calculator ac2661(.scan_win(scan_win2661), .rectangle1_x(rectangle1_xs[2661]), .rectangle1_y(rectangle1_ys[2661]), .rectangle1_width(rectangle1_widths[2661]), .rectangle1_height(rectangle1_heights[2661]), .rectangle1_weight(rectangle1_weights[2661]), .rectangle2_x(rectangle2_xs[2661]), .rectangle2_y(rectangle2_ys[2661]), .rectangle2_width(rectangle2_widths[2661]), .rectangle2_height(rectangle2_heights[2661]), .rectangle2_weight(rectangle2_weights[2661]), .rectangle3_x(rectangle3_xs[2661]), .rectangle3_y(rectangle3_ys[2661]), .rectangle3_width(rectangle3_widths[2661]), .rectangle3_height(rectangle3_heights[2661]), .rectangle3_weight(rectangle3_weights[2661]), .feature_threshold(feature_thresholds[2661]), .feature_above(feature_aboves[2661]), .feature_below(feature_belows[2661]), .scan_win_std_dev(scan_win_std_dev[2661]), .feature_accum(feature_accums[2661]));
  accum_calculator ac2662(.scan_win(scan_win2662), .rectangle1_x(rectangle1_xs[2662]), .rectangle1_y(rectangle1_ys[2662]), .rectangle1_width(rectangle1_widths[2662]), .rectangle1_height(rectangle1_heights[2662]), .rectangle1_weight(rectangle1_weights[2662]), .rectangle2_x(rectangle2_xs[2662]), .rectangle2_y(rectangle2_ys[2662]), .rectangle2_width(rectangle2_widths[2662]), .rectangle2_height(rectangle2_heights[2662]), .rectangle2_weight(rectangle2_weights[2662]), .rectangle3_x(rectangle3_xs[2662]), .rectangle3_y(rectangle3_ys[2662]), .rectangle3_width(rectangle3_widths[2662]), .rectangle3_height(rectangle3_heights[2662]), .rectangle3_weight(rectangle3_weights[2662]), .feature_threshold(feature_thresholds[2662]), .feature_above(feature_aboves[2662]), .feature_below(feature_belows[2662]), .scan_win_std_dev(scan_win_std_dev[2662]), .feature_accum(feature_accums[2662]));
  accum_calculator ac2663(.scan_win(scan_win2663), .rectangle1_x(rectangle1_xs[2663]), .rectangle1_y(rectangle1_ys[2663]), .rectangle1_width(rectangle1_widths[2663]), .rectangle1_height(rectangle1_heights[2663]), .rectangle1_weight(rectangle1_weights[2663]), .rectangle2_x(rectangle2_xs[2663]), .rectangle2_y(rectangle2_ys[2663]), .rectangle2_width(rectangle2_widths[2663]), .rectangle2_height(rectangle2_heights[2663]), .rectangle2_weight(rectangle2_weights[2663]), .rectangle3_x(rectangle3_xs[2663]), .rectangle3_y(rectangle3_ys[2663]), .rectangle3_width(rectangle3_widths[2663]), .rectangle3_height(rectangle3_heights[2663]), .rectangle3_weight(rectangle3_weights[2663]), .feature_threshold(feature_thresholds[2663]), .feature_above(feature_aboves[2663]), .feature_below(feature_belows[2663]), .scan_win_std_dev(scan_win_std_dev[2663]), .feature_accum(feature_accums[2663]));
  accum_calculator ac2664(.scan_win(scan_win2664), .rectangle1_x(rectangle1_xs[2664]), .rectangle1_y(rectangle1_ys[2664]), .rectangle1_width(rectangle1_widths[2664]), .rectangle1_height(rectangle1_heights[2664]), .rectangle1_weight(rectangle1_weights[2664]), .rectangle2_x(rectangle2_xs[2664]), .rectangle2_y(rectangle2_ys[2664]), .rectangle2_width(rectangle2_widths[2664]), .rectangle2_height(rectangle2_heights[2664]), .rectangle2_weight(rectangle2_weights[2664]), .rectangle3_x(rectangle3_xs[2664]), .rectangle3_y(rectangle3_ys[2664]), .rectangle3_width(rectangle3_widths[2664]), .rectangle3_height(rectangle3_heights[2664]), .rectangle3_weight(rectangle3_weights[2664]), .feature_threshold(feature_thresholds[2664]), .feature_above(feature_aboves[2664]), .feature_below(feature_belows[2664]), .scan_win_std_dev(scan_win_std_dev[2664]), .feature_accum(feature_accums[2664]));
  accum_calculator ac2665(.scan_win(scan_win2665), .rectangle1_x(rectangle1_xs[2665]), .rectangle1_y(rectangle1_ys[2665]), .rectangle1_width(rectangle1_widths[2665]), .rectangle1_height(rectangle1_heights[2665]), .rectangle1_weight(rectangle1_weights[2665]), .rectangle2_x(rectangle2_xs[2665]), .rectangle2_y(rectangle2_ys[2665]), .rectangle2_width(rectangle2_widths[2665]), .rectangle2_height(rectangle2_heights[2665]), .rectangle2_weight(rectangle2_weights[2665]), .rectangle3_x(rectangle3_xs[2665]), .rectangle3_y(rectangle3_ys[2665]), .rectangle3_width(rectangle3_widths[2665]), .rectangle3_height(rectangle3_heights[2665]), .rectangle3_weight(rectangle3_weights[2665]), .feature_threshold(feature_thresholds[2665]), .feature_above(feature_aboves[2665]), .feature_below(feature_belows[2665]), .scan_win_std_dev(scan_win_std_dev[2665]), .feature_accum(feature_accums[2665]));
  accum_calculator ac2666(.scan_win(scan_win2666), .rectangle1_x(rectangle1_xs[2666]), .rectangle1_y(rectangle1_ys[2666]), .rectangle1_width(rectangle1_widths[2666]), .rectangle1_height(rectangle1_heights[2666]), .rectangle1_weight(rectangle1_weights[2666]), .rectangle2_x(rectangle2_xs[2666]), .rectangle2_y(rectangle2_ys[2666]), .rectangle2_width(rectangle2_widths[2666]), .rectangle2_height(rectangle2_heights[2666]), .rectangle2_weight(rectangle2_weights[2666]), .rectangle3_x(rectangle3_xs[2666]), .rectangle3_y(rectangle3_ys[2666]), .rectangle3_width(rectangle3_widths[2666]), .rectangle3_height(rectangle3_heights[2666]), .rectangle3_weight(rectangle3_weights[2666]), .feature_threshold(feature_thresholds[2666]), .feature_above(feature_aboves[2666]), .feature_below(feature_belows[2666]), .scan_win_std_dev(scan_win_std_dev[2666]), .feature_accum(feature_accums[2666]));
  accum_calculator ac2667(.scan_win(scan_win2667), .rectangle1_x(rectangle1_xs[2667]), .rectangle1_y(rectangle1_ys[2667]), .rectangle1_width(rectangle1_widths[2667]), .rectangle1_height(rectangle1_heights[2667]), .rectangle1_weight(rectangle1_weights[2667]), .rectangle2_x(rectangle2_xs[2667]), .rectangle2_y(rectangle2_ys[2667]), .rectangle2_width(rectangle2_widths[2667]), .rectangle2_height(rectangle2_heights[2667]), .rectangle2_weight(rectangle2_weights[2667]), .rectangle3_x(rectangle3_xs[2667]), .rectangle3_y(rectangle3_ys[2667]), .rectangle3_width(rectangle3_widths[2667]), .rectangle3_height(rectangle3_heights[2667]), .rectangle3_weight(rectangle3_weights[2667]), .feature_threshold(feature_thresholds[2667]), .feature_above(feature_aboves[2667]), .feature_below(feature_belows[2667]), .scan_win_std_dev(scan_win_std_dev[2667]), .feature_accum(feature_accums[2667]));
  accum_calculator ac2668(.scan_win(scan_win2668), .rectangle1_x(rectangle1_xs[2668]), .rectangle1_y(rectangle1_ys[2668]), .rectangle1_width(rectangle1_widths[2668]), .rectangle1_height(rectangle1_heights[2668]), .rectangle1_weight(rectangle1_weights[2668]), .rectangle2_x(rectangle2_xs[2668]), .rectangle2_y(rectangle2_ys[2668]), .rectangle2_width(rectangle2_widths[2668]), .rectangle2_height(rectangle2_heights[2668]), .rectangle2_weight(rectangle2_weights[2668]), .rectangle3_x(rectangle3_xs[2668]), .rectangle3_y(rectangle3_ys[2668]), .rectangle3_width(rectangle3_widths[2668]), .rectangle3_height(rectangle3_heights[2668]), .rectangle3_weight(rectangle3_weights[2668]), .feature_threshold(feature_thresholds[2668]), .feature_above(feature_aboves[2668]), .feature_below(feature_belows[2668]), .scan_win_std_dev(scan_win_std_dev[2668]), .feature_accum(feature_accums[2668]));
  accum_calculator ac2669(.scan_win(scan_win2669), .rectangle1_x(rectangle1_xs[2669]), .rectangle1_y(rectangle1_ys[2669]), .rectangle1_width(rectangle1_widths[2669]), .rectangle1_height(rectangle1_heights[2669]), .rectangle1_weight(rectangle1_weights[2669]), .rectangle2_x(rectangle2_xs[2669]), .rectangle2_y(rectangle2_ys[2669]), .rectangle2_width(rectangle2_widths[2669]), .rectangle2_height(rectangle2_heights[2669]), .rectangle2_weight(rectangle2_weights[2669]), .rectangle3_x(rectangle3_xs[2669]), .rectangle3_y(rectangle3_ys[2669]), .rectangle3_width(rectangle3_widths[2669]), .rectangle3_height(rectangle3_heights[2669]), .rectangle3_weight(rectangle3_weights[2669]), .feature_threshold(feature_thresholds[2669]), .feature_above(feature_aboves[2669]), .feature_below(feature_belows[2669]), .scan_win_std_dev(scan_win_std_dev[2669]), .feature_accum(feature_accums[2669]));
  accum_calculator ac2670(.scan_win(scan_win2670), .rectangle1_x(rectangle1_xs[2670]), .rectangle1_y(rectangle1_ys[2670]), .rectangle1_width(rectangle1_widths[2670]), .rectangle1_height(rectangle1_heights[2670]), .rectangle1_weight(rectangle1_weights[2670]), .rectangle2_x(rectangle2_xs[2670]), .rectangle2_y(rectangle2_ys[2670]), .rectangle2_width(rectangle2_widths[2670]), .rectangle2_height(rectangle2_heights[2670]), .rectangle2_weight(rectangle2_weights[2670]), .rectangle3_x(rectangle3_xs[2670]), .rectangle3_y(rectangle3_ys[2670]), .rectangle3_width(rectangle3_widths[2670]), .rectangle3_height(rectangle3_heights[2670]), .rectangle3_weight(rectangle3_weights[2670]), .feature_threshold(feature_thresholds[2670]), .feature_above(feature_aboves[2670]), .feature_below(feature_belows[2670]), .scan_win_std_dev(scan_win_std_dev[2670]), .feature_accum(feature_accums[2670]));
  accum_calculator ac2671(.scan_win(scan_win2671), .rectangle1_x(rectangle1_xs[2671]), .rectangle1_y(rectangle1_ys[2671]), .rectangle1_width(rectangle1_widths[2671]), .rectangle1_height(rectangle1_heights[2671]), .rectangle1_weight(rectangle1_weights[2671]), .rectangle2_x(rectangle2_xs[2671]), .rectangle2_y(rectangle2_ys[2671]), .rectangle2_width(rectangle2_widths[2671]), .rectangle2_height(rectangle2_heights[2671]), .rectangle2_weight(rectangle2_weights[2671]), .rectangle3_x(rectangle3_xs[2671]), .rectangle3_y(rectangle3_ys[2671]), .rectangle3_width(rectangle3_widths[2671]), .rectangle3_height(rectangle3_heights[2671]), .rectangle3_weight(rectangle3_weights[2671]), .feature_threshold(feature_thresholds[2671]), .feature_above(feature_aboves[2671]), .feature_below(feature_belows[2671]), .scan_win_std_dev(scan_win_std_dev[2671]), .feature_accum(feature_accums[2671]));
  accum_calculator ac2672(.scan_win(scan_win2672), .rectangle1_x(rectangle1_xs[2672]), .rectangle1_y(rectangle1_ys[2672]), .rectangle1_width(rectangle1_widths[2672]), .rectangle1_height(rectangle1_heights[2672]), .rectangle1_weight(rectangle1_weights[2672]), .rectangle2_x(rectangle2_xs[2672]), .rectangle2_y(rectangle2_ys[2672]), .rectangle2_width(rectangle2_widths[2672]), .rectangle2_height(rectangle2_heights[2672]), .rectangle2_weight(rectangle2_weights[2672]), .rectangle3_x(rectangle3_xs[2672]), .rectangle3_y(rectangle3_ys[2672]), .rectangle3_width(rectangle3_widths[2672]), .rectangle3_height(rectangle3_heights[2672]), .rectangle3_weight(rectangle3_weights[2672]), .feature_threshold(feature_thresholds[2672]), .feature_above(feature_aboves[2672]), .feature_below(feature_belows[2672]), .scan_win_std_dev(scan_win_std_dev[2672]), .feature_accum(feature_accums[2672]));
  accum_calculator ac2673(.scan_win(scan_win2673), .rectangle1_x(rectangle1_xs[2673]), .rectangle1_y(rectangle1_ys[2673]), .rectangle1_width(rectangle1_widths[2673]), .rectangle1_height(rectangle1_heights[2673]), .rectangle1_weight(rectangle1_weights[2673]), .rectangle2_x(rectangle2_xs[2673]), .rectangle2_y(rectangle2_ys[2673]), .rectangle2_width(rectangle2_widths[2673]), .rectangle2_height(rectangle2_heights[2673]), .rectangle2_weight(rectangle2_weights[2673]), .rectangle3_x(rectangle3_xs[2673]), .rectangle3_y(rectangle3_ys[2673]), .rectangle3_width(rectangle3_widths[2673]), .rectangle3_height(rectangle3_heights[2673]), .rectangle3_weight(rectangle3_weights[2673]), .feature_threshold(feature_thresholds[2673]), .feature_above(feature_aboves[2673]), .feature_below(feature_belows[2673]), .scan_win_std_dev(scan_win_std_dev[2673]), .feature_accum(feature_accums[2673]));
  accum_calculator ac2674(.scan_win(scan_win2674), .rectangle1_x(rectangle1_xs[2674]), .rectangle1_y(rectangle1_ys[2674]), .rectangle1_width(rectangle1_widths[2674]), .rectangle1_height(rectangle1_heights[2674]), .rectangle1_weight(rectangle1_weights[2674]), .rectangle2_x(rectangle2_xs[2674]), .rectangle2_y(rectangle2_ys[2674]), .rectangle2_width(rectangle2_widths[2674]), .rectangle2_height(rectangle2_heights[2674]), .rectangle2_weight(rectangle2_weights[2674]), .rectangle3_x(rectangle3_xs[2674]), .rectangle3_y(rectangle3_ys[2674]), .rectangle3_width(rectangle3_widths[2674]), .rectangle3_height(rectangle3_heights[2674]), .rectangle3_weight(rectangle3_weights[2674]), .feature_threshold(feature_thresholds[2674]), .feature_above(feature_aboves[2674]), .feature_below(feature_belows[2674]), .scan_win_std_dev(scan_win_std_dev[2674]), .feature_accum(feature_accums[2674]));
  accum_calculator ac2675(.scan_win(scan_win2675), .rectangle1_x(rectangle1_xs[2675]), .rectangle1_y(rectangle1_ys[2675]), .rectangle1_width(rectangle1_widths[2675]), .rectangle1_height(rectangle1_heights[2675]), .rectangle1_weight(rectangle1_weights[2675]), .rectangle2_x(rectangle2_xs[2675]), .rectangle2_y(rectangle2_ys[2675]), .rectangle2_width(rectangle2_widths[2675]), .rectangle2_height(rectangle2_heights[2675]), .rectangle2_weight(rectangle2_weights[2675]), .rectangle3_x(rectangle3_xs[2675]), .rectangle3_y(rectangle3_ys[2675]), .rectangle3_width(rectangle3_widths[2675]), .rectangle3_height(rectangle3_heights[2675]), .rectangle3_weight(rectangle3_weights[2675]), .feature_threshold(feature_thresholds[2675]), .feature_above(feature_aboves[2675]), .feature_below(feature_belows[2675]), .scan_win_std_dev(scan_win_std_dev[2675]), .feature_accum(feature_accums[2675]));
  accum_calculator ac2676(.scan_win(scan_win2676), .rectangle1_x(rectangle1_xs[2676]), .rectangle1_y(rectangle1_ys[2676]), .rectangle1_width(rectangle1_widths[2676]), .rectangle1_height(rectangle1_heights[2676]), .rectangle1_weight(rectangle1_weights[2676]), .rectangle2_x(rectangle2_xs[2676]), .rectangle2_y(rectangle2_ys[2676]), .rectangle2_width(rectangle2_widths[2676]), .rectangle2_height(rectangle2_heights[2676]), .rectangle2_weight(rectangle2_weights[2676]), .rectangle3_x(rectangle3_xs[2676]), .rectangle3_y(rectangle3_ys[2676]), .rectangle3_width(rectangle3_widths[2676]), .rectangle3_height(rectangle3_heights[2676]), .rectangle3_weight(rectangle3_weights[2676]), .feature_threshold(feature_thresholds[2676]), .feature_above(feature_aboves[2676]), .feature_below(feature_belows[2676]), .scan_win_std_dev(scan_win_std_dev[2676]), .feature_accum(feature_accums[2676]));
  accum_calculator ac2677(.scan_win(scan_win2677), .rectangle1_x(rectangle1_xs[2677]), .rectangle1_y(rectangle1_ys[2677]), .rectangle1_width(rectangle1_widths[2677]), .rectangle1_height(rectangle1_heights[2677]), .rectangle1_weight(rectangle1_weights[2677]), .rectangle2_x(rectangle2_xs[2677]), .rectangle2_y(rectangle2_ys[2677]), .rectangle2_width(rectangle2_widths[2677]), .rectangle2_height(rectangle2_heights[2677]), .rectangle2_weight(rectangle2_weights[2677]), .rectangle3_x(rectangle3_xs[2677]), .rectangle3_y(rectangle3_ys[2677]), .rectangle3_width(rectangle3_widths[2677]), .rectangle3_height(rectangle3_heights[2677]), .rectangle3_weight(rectangle3_weights[2677]), .feature_threshold(feature_thresholds[2677]), .feature_above(feature_aboves[2677]), .feature_below(feature_belows[2677]), .scan_win_std_dev(scan_win_std_dev[2677]), .feature_accum(feature_accums[2677]));
  accum_calculator ac2678(.scan_win(scan_win2678), .rectangle1_x(rectangle1_xs[2678]), .rectangle1_y(rectangle1_ys[2678]), .rectangle1_width(rectangle1_widths[2678]), .rectangle1_height(rectangle1_heights[2678]), .rectangle1_weight(rectangle1_weights[2678]), .rectangle2_x(rectangle2_xs[2678]), .rectangle2_y(rectangle2_ys[2678]), .rectangle2_width(rectangle2_widths[2678]), .rectangle2_height(rectangle2_heights[2678]), .rectangle2_weight(rectangle2_weights[2678]), .rectangle3_x(rectangle3_xs[2678]), .rectangle3_y(rectangle3_ys[2678]), .rectangle3_width(rectangle3_widths[2678]), .rectangle3_height(rectangle3_heights[2678]), .rectangle3_weight(rectangle3_weights[2678]), .feature_threshold(feature_thresholds[2678]), .feature_above(feature_aboves[2678]), .feature_below(feature_belows[2678]), .scan_win_std_dev(scan_win_std_dev[2678]), .feature_accum(feature_accums[2678]));
  accum_calculator ac2679(.scan_win(scan_win2679), .rectangle1_x(rectangle1_xs[2679]), .rectangle1_y(rectangle1_ys[2679]), .rectangle1_width(rectangle1_widths[2679]), .rectangle1_height(rectangle1_heights[2679]), .rectangle1_weight(rectangle1_weights[2679]), .rectangle2_x(rectangle2_xs[2679]), .rectangle2_y(rectangle2_ys[2679]), .rectangle2_width(rectangle2_widths[2679]), .rectangle2_height(rectangle2_heights[2679]), .rectangle2_weight(rectangle2_weights[2679]), .rectangle3_x(rectangle3_xs[2679]), .rectangle3_y(rectangle3_ys[2679]), .rectangle3_width(rectangle3_widths[2679]), .rectangle3_height(rectangle3_heights[2679]), .rectangle3_weight(rectangle3_weights[2679]), .feature_threshold(feature_thresholds[2679]), .feature_above(feature_aboves[2679]), .feature_below(feature_belows[2679]), .scan_win_std_dev(scan_win_std_dev[2679]), .feature_accum(feature_accums[2679]));
  accum_calculator ac2680(.scan_win(scan_win2680), .rectangle1_x(rectangle1_xs[2680]), .rectangle1_y(rectangle1_ys[2680]), .rectangle1_width(rectangle1_widths[2680]), .rectangle1_height(rectangle1_heights[2680]), .rectangle1_weight(rectangle1_weights[2680]), .rectangle2_x(rectangle2_xs[2680]), .rectangle2_y(rectangle2_ys[2680]), .rectangle2_width(rectangle2_widths[2680]), .rectangle2_height(rectangle2_heights[2680]), .rectangle2_weight(rectangle2_weights[2680]), .rectangle3_x(rectangle3_xs[2680]), .rectangle3_y(rectangle3_ys[2680]), .rectangle3_width(rectangle3_widths[2680]), .rectangle3_height(rectangle3_heights[2680]), .rectangle3_weight(rectangle3_weights[2680]), .feature_threshold(feature_thresholds[2680]), .feature_above(feature_aboves[2680]), .feature_below(feature_belows[2680]), .scan_win_std_dev(scan_win_std_dev[2680]), .feature_accum(feature_accums[2680]));
  accum_calculator ac2681(.scan_win(scan_win2681), .rectangle1_x(rectangle1_xs[2681]), .rectangle1_y(rectangle1_ys[2681]), .rectangle1_width(rectangle1_widths[2681]), .rectangle1_height(rectangle1_heights[2681]), .rectangle1_weight(rectangle1_weights[2681]), .rectangle2_x(rectangle2_xs[2681]), .rectangle2_y(rectangle2_ys[2681]), .rectangle2_width(rectangle2_widths[2681]), .rectangle2_height(rectangle2_heights[2681]), .rectangle2_weight(rectangle2_weights[2681]), .rectangle3_x(rectangle3_xs[2681]), .rectangle3_y(rectangle3_ys[2681]), .rectangle3_width(rectangle3_widths[2681]), .rectangle3_height(rectangle3_heights[2681]), .rectangle3_weight(rectangle3_weights[2681]), .feature_threshold(feature_thresholds[2681]), .feature_above(feature_aboves[2681]), .feature_below(feature_belows[2681]), .scan_win_std_dev(scan_win_std_dev[2681]), .feature_accum(feature_accums[2681]));
  accum_calculator ac2682(.scan_win(scan_win2682), .rectangle1_x(rectangle1_xs[2682]), .rectangle1_y(rectangle1_ys[2682]), .rectangle1_width(rectangle1_widths[2682]), .rectangle1_height(rectangle1_heights[2682]), .rectangle1_weight(rectangle1_weights[2682]), .rectangle2_x(rectangle2_xs[2682]), .rectangle2_y(rectangle2_ys[2682]), .rectangle2_width(rectangle2_widths[2682]), .rectangle2_height(rectangle2_heights[2682]), .rectangle2_weight(rectangle2_weights[2682]), .rectangle3_x(rectangle3_xs[2682]), .rectangle3_y(rectangle3_ys[2682]), .rectangle3_width(rectangle3_widths[2682]), .rectangle3_height(rectangle3_heights[2682]), .rectangle3_weight(rectangle3_weights[2682]), .feature_threshold(feature_thresholds[2682]), .feature_above(feature_aboves[2682]), .feature_below(feature_belows[2682]), .scan_win_std_dev(scan_win_std_dev[2682]), .feature_accum(feature_accums[2682]));
  accum_calculator ac2683(.scan_win(scan_win2683), .rectangle1_x(rectangle1_xs[2683]), .rectangle1_y(rectangle1_ys[2683]), .rectangle1_width(rectangle1_widths[2683]), .rectangle1_height(rectangle1_heights[2683]), .rectangle1_weight(rectangle1_weights[2683]), .rectangle2_x(rectangle2_xs[2683]), .rectangle2_y(rectangle2_ys[2683]), .rectangle2_width(rectangle2_widths[2683]), .rectangle2_height(rectangle2_heights[2683]), .rectangle2_weight(rectangle2_weights[2683]), .rectangle3_x(rectangle3_xs[2683]), .rectangle3_y(rectangle3_ys[2683]), .rectangle3_width(rectangle3_widths[2683]), .rectangle3_height(rectangle3_heights[2683]), .rectangle3_weight(rectangle3_weights[2683]), .feature_threshold(feature_thresholds[2683]), .feature_above(feature_aboves[2683]), .feature_below(feature_belows[2683]), .scan_win_std_dev(scan_win_std_dev[2683]), .feature_accum(feature_accums[2683]));
  accum_calculator ac2684(.scan_win(scan_win2684), .rectangle1_x(rectangle1_xs[2684]), .rectangle1_y(rectangle1_ys[2684]), .rectangle1_width(rectangle1_widths[2684]), .rectangle1_height(rectangle1_heights[2684]), .rectangle1_weight(rectangle1_weights[2684]), .rectangle2_x(rectangle2_xs[2684]), .rectangle2_y(rectangle2_ys[2684]), .rectangle2_width(rectangle2_widths[2684]), .rectangle2_height(rectangle2_heights[2684]), .rectangle2_weight(rectangle2_weights[2684]), .rectangle3_x(rectangle3_xs[2684]), .rectangle3_y(rectangle3_ys[2684]), .rectangle3_width(rectangle3_widths[2684]), .rectangle3_height(rectangle3_heights[2684]), .rectangle3_weight(rectangle3_weights[2684]), .feature_threshold(feature_thresholds[2684]), .feature_above(feature_aboves[2684]), .feature_below(feature_belows[2684]), .scan_win_std_dev(scan_win_std_dev[2684]), .feature_accum(feature_accums[2684]));
  accum_calculator ac2685(.scan_win(scan_win2685), .rectangle1_x(rectangle1_xs[2685]), .rectangle1_y(rectangle1_ys[2685]), .rectangle1_width(rectangle1_widths[2685]), .rectangle1_height(rectangle1_heights[2685]), .rectangle1_weight(rectangle1_weights[2685]), .rectangle2_x(rectangle2_xs[2685]), .rectangle2_y(rectangle2_ys[2685]), .rectangle2_width(rectangle2_widths[2685]), .rectangle2_height(rectangle2_heights[2685]), .rectangle2_weight(rectangle2_weights[2685]), .rectangle3_x(rectangle3_xs[2685]), .rectangle3_y(rectangle3_ys[2685]), .rectangle3_width(rectangle3_widths[2685]), .rectangle3_height(rectangle3_heights[2685]), .rectangle3_weight(rectangle3_weights[2685]), .feature_threshold(feature_thresholds[2685]), .feature_above(feature_aboves[2685]), .feature_below(feature_belows[2685]), .scan_win_std_dev(scan_win_std_dev[2685]), .feature_accum(feature_accums[2685]));
  accum_calculator ac2686(.scan_win(scan_win2686), .rectangle1_x(rectangle1_xs[2686]), .rectangle1_y(rectangle1_ys[2686]), .rectangle1_width(rectangle1_widths[2686]), .rectangle1_height(rectangle1_heights[2686]), .rectangle1_weight(rectangle1_weights[2686]), .rectangle2_x(rectangle2_xs[2686]), .rectangle2_y(rectangle2_ys[2686]), .rectangle2_width(rectangle2_widths[2686]), .rectangle2_height(rectangle2_heights[2686]), .rectangle2_weight(rectangle2_weights[2686]), .rectangle3_x(rectangle3_xs[2686]), .rectangle3_y(rectangle3_ys[2686]), .rectangle3_width(rectangle3_widths[2686]), .rectangle3_height(rectangle3_heights[2686]), .rectangle3_weight(rectangle3_weights[2686]), .feature_threshold(feature_thresholds[2686]), .feature_above(feature_aboves[2686]), .feature_below(feature_belows[2686]), .scan_win_std_dev(scan_win_std_dev[2686]), .feature_accum(feature_accums[2686]));
  accum_calculator ac2687(.scan_win(scan_win2687), .rectangle1_x(rectangle1_xs[2687]), .rectangle1_y(rectangle1_ys[2687]), .rectangle1_width(rectangle1_widths[2687]), .rectangle1_height(rectangle1_heights[2687]), .rectangle1_weight(rectangle1_weights[2687]), .rectangle2_x(rectangle2_xs[2687]), .rectangle2_y(rectangle2_ys[2687]), .rectangle2_width(rectangle2_widths[2687]), .rectangle2_height(rectangle2_heights[2687]), .rectangle2_weight(rectangle2_weights[2687]), .rectangle3_x(rectangle3_xs[2687]), .rectangle3_y(rectangle3_ys[2687]), .rectangle3_width(rectangle3_widths[2687]), .rectangle3_height(rectangle3_heights[2687]), .rectangle3_weight(rectangle3_weights[2687]), .feature_threshold(feature_thresholds[2687]), .feature_above(feature_aboves[2687]), .feature_below(feature_belows[2687]), .scan_win_std_dev(scan_win_std_dev[2687]), .feature_accum(feature_accums[2687]));
  accum_calculator ac2688(.scan_win(scan_win2688), .rectangle1_x(rectangle1_xs[2688]), .rectangle1_y(rectangle1_ys[2688]), .rectangle1_width(rectangle1_widths[2688]), .rectangle1_height(rectangle1_heights[2688]), .rectangle1_weight(rectangle1_weights[2688]), .rectangle2_x(rectangle2_xs[2688]), .rectangle2_y(rectangle2_ys[2688]), .rectangle2_width(rectangle2_widths[2688]), .rectangle2_height(rectangle2_heights[2688]), .rectangle2_weight(rectangle2_weights[2688]), .rectangle3_x(rectangle3_xs[2688]), .rectangle3_y(rectangle3_ys[2688]), .rectangle3_width(rectangle3_widths[2688]), .rectangle3_height(rectangle3_heights[2688]), .rectangle3_weight(rectangle3_weights[2688]), .feature_threshold(feature_thresholds[2688]), .feature_above(feature_aboves[2688]), .feature_below(feature_belows[2688]), .scan_win_std_dev(scan_win_std_dev[2688]), .feature_accum(feature_accums[2688]));
  accum_calculator ac2689(.scan_win(scan_win2689), .rectangle1_x(rectangle1_xs[2689]), .rectangle1_y(rectangle1_ys[2689]), .rectangle1_width(rectangle1_widths[2689]), .rectangle1_height(rectangle1_heights[2689]), .rectangle1_weight(rectangle1_weights[2689]), .rectangle2_x(rectangle2_xs[2689]), .rectangle2_y(rectangle2_ys[2689]), .rectangle2_width(rectangle2_widths[2689]), .rectangle2_height(rectangle2_heights[2689]), .rectangle2_weight(rectangle2_weights[2689]), .rectangle3_x(rectangle3_xs[2689]), .rectangle3_y(rectangle3_ys[2689]), .rectangle3_width(rectangle3_widths[2689]), .rectangle3_height(rectangle3_heights[2689]), .rectangle3_weight(rectangle3_weights[2689]), .feature_threshold(feature_thresholds[2689]), .feature_above(feature_aboves[2689]), .feature_below(feature_belows[2689]), .scan_win_std_dev(scan_win_std_dev[2689]), .feature_accum(feature_accums[2689]));
  accum_calculator ac2690(.scan_win(scan_win2690), .rectangle1_x(rectangle1_xs[2690]), .rectangle1_y(rectangle1_ys[2690]), .rectangle1_width(rectangle1_widths[2690]), .rectangle1_height(rectangle1_heights[2690]), .rectangle1_weight(rectangle1_weights[2690]), .rectangle2_x(rectangle2_xs[2690]), .rectangle2_y(rectangle2_ys[2690]), .rectangle2_width(rectangle2_widths[2690]), .rectangle2_height(rectangle2_heights[2690]), .rectangle2_weight(rectangle2_weights[2690]), .rectangle3_x(rectangle3_xs[2690]), .rectangle3_y(rectangle3_ys[2690]), .rectangle3_width(rectangle3_widths[2690]), .rectangle3_height(rectangle3_heights[2690]), .rectangle3_weight(rectangle3_weights[2690]), .feature_threshold(feature_thresholds[2690]), .feature_above(feature_aboves[2690]), .feature_below(feature_belows[2690]), .scan_win_std_dev(scan_win_std_dev[2690]), .feature_accum(feature_accums[2690]));
  accum_calculator ac2691(.scan_win(scan_win2691), .rectangle1_x(rectangle1_xs[2691]), .rectangle1_y(rectangle1_ys[2691]), .rectangle1_width(rectangle1_widths[2691]), .rectangle1_height(rectangle1_heights[2691]), .rectangle1_weight(rectangle1_weights[2691]), .rectangle2_x(rectangle2_xs[2691]), .rectangle2_y(rectangle2_ys[2691]), .rectangle2_width(rectangle2_widths[2691]), .rectangle2_height(rectangle2_heights[2691]), .rectangle2_weight(rectangle2_weights[2691]), .rectangle3_x(rectangle3_xs[2691]), .rectangle3_y(rectangle3_ys[2691]), .rectangle3_width(rectangle3_widths[2691]), .rectangle3_height(rectangle3_heights[2691]), .rectangle3_weight(rectangle3_weights[2691]), .feature_threshold(feature_thresholds[2691]), .feature_above(feature_aboves[2691]), .feature_below(feature_belows[2691]), .scan_win_std_dev(scan_win_std_dev[2691]), .feature_accum(feature_accums[2691]));
  accum_calculator ac2692(.scan_win(scan_win2692), .rectangle1_x(rectangle1_xs[2692]), .rectangle1_y(rectangle1_ys[2692]), .rectangle1_width(rectangle1_widths[2692]), .rectangle1_height(rectangle1_heights[2692]), .rectangle1_weight(rectangle1_weights[2692]), .rectangle2_x(rectangle2_xs[2692]), .rectangle2_y(rectangle2_ys[2692]), .rectangle2_width(rectangle2_widths[2692]), .rectangle2_height(rectangle2_heights[2692]), .rectangle2_weight(rectangle2_weights[2692]), .rectangle3_x(rectangle3_xs[2692]), .rectangle3_y(rectangle3_ys[2692]), .rectangle3_width(rectangle3_widths[2692]), .rectangle3_height(rectangle3_heights[2692]), .rectangle3_weight(rectangle3_weights[2692]), .feature_threshold(feature_thresholds[2692]), .feature_above(feature_aboves[2692]), .feature_below(feature_belows[2692]), .scan_win_std_dev(scan_win_std_dev[2692]), .feature_accum(feature_accums[2692]));
  accum_calculator ac2693(.scan_win(scan_win2693), .rectangle1_x(rectangle1_xs[2693]), .rectangle1_y(rectangle1_ys[2693]), .rectangle1_width(rectangle1_widths[2693]), .rectangle1_height(rectangle1_heights[2693]), .rectangle1_weight(rectangle1_weights[2693]), .rectangle2_x(rectangle2_xs[2693]), .rectangle2_y(rectangle2_ys[2693]), .rectangle2_width(rectangle2_widths[2693]), .rectangle2_height(rectangle2_heights[2693]), .rectangle2_weight(rectangle2_weights[2693]), .rectangle3_x(rectangle3_xs[2693]), .rectangle3_y(rectangle3_ys[2693]), .rectangle3_width(rectangle3_widths[2693]), .rectangle3_height(rectangle3_heights[2693]), .rectangle3_weight(rectangle3_weights[2693]), .feature_threshold(feature_thresholds[2693]), .feature_above(feature_aboves[2693]), .feature_below(feature_belows[2693]), .scan_win_std_dev(scan_win_std_dev[2693]), .feature_accum(feature_accums[2693]));
  accum_calculator ac2694(.scan_win(scan_win2694), .rectangle1_x(rectangle1_xs[2694]), .rectangle1_y(rectangle1_ys[2694]), .rectangle1_width(rectangle1_widths[2694]), .rectangle1_height(rectangle1_heights[2694]), .rectangle1_weight(rectangle1_weights[2694]), .rectangle2_x(rectangle2_xs[2694]), .rectangle2_y(rectangle2_ys[2694]), .rectangle2_width(rectangle2_widths[2694]), .rectangle2_height(rectangle2_heights[2694]), .rectangle2_weight(rectangle2_weights[2694]), .rectangle3_x(rectangle3_xs[2694]), .rectangle3_y(rectangle3_ys[2694]), .rectangle3_width(rectangle3_widths[2694]), .rectangle3_height(rectangle3_heights[2694]), .rectangle3_weight(rectangle3_weights[2694]), .feature_threshold(feature_thresholds[2694]), .feature_above(feature_aboves[2694]), .feature_below(feature_belows[2694]), .scan_win_std_dev(scan_win_std_dev[2694]), .feature_accum(feature_accums[2694]));
  accum_calculator ac2695(.scan_win(scan_win2695), .rectangle1_x(rectangle1_xs[2695]), .rectangle1_y(rectangle1_ys[2695]), .rectangle1_width(rectangle1_widths[2695]), .rectangle1_height(rectangle1_heights[2695]), .rectangle1_weight(rectangle1_weights[2695]), .rectangle2_x(rectangle2_xs[2695]), .rectangle2_y(rectangle2_ys[2695]), .rectangle2_width(rectangle2_widths[2695]), .rectangle2_height(rectangle2_heights[2695]), .rectangle2_weight(rectangle2_weights[2695]), .rectangle3_x(rectangle3_xs[2695]), .rectangle3_y(rectangle3_ys[2695]), .rectangle3_width(rectangle3_widths[2695]), .rectangle3_height(rectangle3_heights[2695]), .rectangle3_weight(rectangle3_weights[2695]), .feature_threshold(feature_thresholds[2695]), .feature_above(feature_aboves[2695]), .feature_below(feature_belows[2695]), .scan_win_std_dev(scan_win_std_dev[2695]), .feature_accum(feature_accums[2695]));
  accum_calculator ac2696(.scan_win(scan_win2696), .rectangle1_x(rectangle1_xs[2696]), .rectangle1_y(rectangle1_ys[2696]), .rectangle1_width(rectangle1_widths[2696]), .rectangle1_height(rectangle1_heights[2696]), .rectangle1_weight(rectangle1_weights[2696]), .rectangle2_x(rectangle2_xs[2696]), .rectangle2_y(rectangle2_ys[2696]), .rectangle2_width(rectangle2_widths[2696]), .rectangle2_height(rectangle2_heights[2696]), .rectangle2_weight(rectangle2_weights[2696]), .rectangle3_x(rectangle3_xs[2696]), .rectangle3_y(rectangle3_ys[2696]), .rectangle3_width(rectangle3_widths[2696]), .rectangle3_height(rectangle3_heights[2696]), .rectangle3_weight(rectangle3_weights[2696]), .feature_threshold(feature_thresholds[2696]), .feature_above(feature_aboves[2696]), .feature_below(feature_belows[2696]), .scan_win_std_dev(scan_win_std_dev[2696]), .feature_accum(feature_accums[2696]));
  accum_calculator ac2697(.scan_win(scan_win2697), .rectangle1_x(rectangle1_xs[2697]), .rectangle1_y(rectangle1_ys[2697]), .rectangle1_width(rectangle1_widths[2697]), .rectangle1_height(rectangle1_heights[2697]), .rectangle1_weight(rectangle1_weights[2697]), .rectangle2_x(rectangle2_xs[2697]), .rectangle2_y(rectangle2_ys[2697]), .rectangle2_width(rectangle2_widths[2697]), .rectangle2_height(rectangle2_heights[2697]), .rectangle2_weight(rectangle2_weights[2697]), .rectangle3_x(rectangle3_xs[2697]), .rectangle3_y(rectangle3_ys[2697]), .rectangle3_width(rectangle3_widths[2697]), .rectangle3_height(rectangle3_heights[2697]), .rectangle3_weight(rectangle3_weights[2697]), .feature_threshold(feature_thresholds[2697]), .feature_above(feature_aboves[2697]), .feature_below(feature_belows[2697]), .scan_win_std_dev(scan_win_std_dev[2697]), .feature_accum(feature_accums[2697]));
  accum_calculator ac2698(.scan_win(scan_win2698), .rectangle1_x(rectangle1_xs[2698]), .rectangle1_y(rectangle1_ys[2698]), .rectangle1_width(rectangle1_widths[2698]), .rectangle1_height(rectangle1_heights[2698]), .rectangle1_weight(rectangle1_weights[2698]), .rectangle2_x(rectangle2_xs[2698]), .rectangle2_y(rectangle2_ys[2698]), .rectangle2_width(rectangle2_widths[2698]), .rectangle2_height(rectangle2_heights[2698]), .rectangle2_weight(rectangle2_weights[2698]), .rectangle3_x(rectangle3_xs[2698]), .rectangle3_y(rectangle3_ys[2698]), .rectangle3_width(rectangle3_widths[2698]), .rectangle3_height(rectangle3_heights[2698]), .rectangle3_weight(rectangle3_weights[2698]), .feature_threshold(feature_thresholds[2698]), .feature_above(feature_aboves[2698]), .feature_below(feature_belows[2698]), .scan_win_std_dev(scan_win_std_dev[2698]), .feature_accum(feature_accums[2698]));
  accum_calculator ac2699(.scan_win(scan_win2699), .rectangle1_x(rectangle1_xs[2699]), .rectangle1_y(rectangle1_ys[2699]), .rectangle1_width(rectangle1_widths[2699]), .rectangle1_height(rectangle1_heights[2699]), .rectangle1_weight(rectangle1_weights[2699]), .rectangle2_x(rectangle2_xs[2699]), .rectangle2_y(rectangle2_ys[2699]), .rectangle2_width(rectangle2_widths[2699]), .rectangle2_height(rectangle2_heights[2699]), .rectangle2_weight(rectangle2_weights[2699]), .rectangle3_x(rectangle3_xs[2699]), .rectangle3_y(rectangle3_ys[2699]), .rectangle3_width(rectangle3_widths[2699]), .rectangle3_height(rectangle3_heights[2699]), .rectangle3_weight(rectangle3_weights[2699]), .feature_threshold(feature_thresholds[2699]), .feature_above(feature_aboves[2699]), .feature_below(feature_belows[2699]), .scan_win_std_dev(scan_win_std_dev[2699]), .feature_accum(feature_accums[2699]));
  accum_calculator ac2700(.scan_win(scan_win2700), .rectangle1_x(rectangle1_xs[2700]), .rectangle1_y(rectangle1_ys[2700]), .rectangle1_width(rectangle1_widths[2700]), .rectangle1_height(rectangle1_heights[2700]), .rectangle1_weight(rectangle1_weights[2700]), .rectangle2_x(rectangle2_xs[2700]), .rectangle2_y(rectangle2_ys[2700]), .rectangle2_width(rectangle2_widths[2700]), .rectangle2_height(rectangle2_heights[2700]), .rectangle2_weight(rectangle2_weights[2700]), .rectangle3_x(rectangle3_xs[2700]), .rectangle3_y(rectangle3_ys[2700]), .rectangle3_width(rectangle3_widths[2700]), .rectangle3_height(rectangle3_heights[2700]), .rectangle3_weight(rectangle3_weights[2700]), .feature_threshold(feature_thresholds[2700]), .feature_above(feature_aboves[2700]), .feature_below(feature_belows[2700]), .scan_win_std_dev(scan_win_std_dev[2700]), .feature_accum(feature_accums[2700]));
  accum_calculator ac2701(.scan_win(scan_win2701), .rectangle1_x(rectangle1_xs[2701]), .rectangle1_y(rectangle1_ys[2701]), .rectangle1_width(rectangle1_widths[2701]), .rectangle1_height(rectangle1_heights[2701]), .rectangle1_weight(rectangle1_weights[2701]), .rectangle2_x(rectangle2_xs[2701]), .rectangle2_y(rectangle2_ys[2701]), .rectangle2_width(rectangle2_widths[2701]), .rectangle2_height(rectangle2_heights[2701]), .rectangle2_weight(rectangle2_weights[2701]), .rectangle3_x(rectangle3_xs[2701]), .rectangle3_y(rectangle3_ys[2701]), .rectangle3_width(rectangle3_widths[2701]), .rectangle3_height(rectangle3_heights[2701]), .rectangle3_weight(rectangle3_weights[2701]), .feature_threshold(feature_thresholds[2701]), .feature_above(feature_aboves[2701]), .feature_below(feature_belows[2701]), .scan_win_std_dev(scan_win_std_dev[2701]), .feature_accum(feature_accums[2701]));
  accum_calculator ac2702(.scan_win(scan_win2702), .rectangle1_x(rectangle1_xs[2702]), .rectangle1_y(rectangle1_ys[2702]), .rectangle1_width(rectangle1_widths[2702]), .rectangle1_height(rectangle1_heights[2702]), .rectangle1_weight(rectangle1_weights[2702]), .rectangle2_x(rectangle2_xs[2702]), .rectangle2_y(rectangle2_ys[2702]), .rectangle2_width(rectangle2_widths[2702]), .rectangle2_height(rectangle2_heights[2702]), .rectangle2_weight(rectangle2_weights[2702]), .rectangle3_x(rectangle3_xs[2702]), .rectangle3_y(rectangle3_ys[2702]), .rectangle3_width(rectangle3_widths[2702]), .rectangle3_height(rectangle3_heights[2702]), .rectangle3_weight(rectangle3_weights[2702]), .feature_threshold(feature_thresholds[2702]), .feature_above(feature_aboves[2702]), .feature_below(feature_belows[2702]), .scan_win_std_dev(scan_win_std_dev[2702]), .feature_accum(feature_accums[2702]));
  accum_calculator ac2703(.scan_win(scan_win2703), .rectangle1_x(rectangle1_xs[2703]), .rectangle1_y(rectangle1_ys[2703]), .rectangle1_width(rectangle1_widths[2703]), .rectangle1_height(rectangle1_heights[2703]), .rectangle1_weight(rectangle1_weights[2703]), .rectangle2_x(rectangle2_xs[2703]), .rectangle2_y(rectangle2_ys[2703]), .rectangle2_width(rectangle2_widths[2703]), .rectangle2_height(rectangle2_heights[2703]), .rectangle2_weight(rectangle2_weights[2703]), .rectangle3_x(rectangle3_xs[2703]), .rectangle3_y(rectangle3_ys[2703]), .rectangle3_width(rectangle3_widths[2703]), .rectangle3_height(rectangle3_heights[2703]), .rectangle3_weight(rectangle3_weights[2703]), .feature_threshold(feature_thresholds[2703]), .feature_above(feature_aboves[2703]), .feature_below(feature_belows[2703]), .scan_win_std_dev(scan_win_std_dev[2703]), .feature_accum(feature_accums[2703]));
  accum_calculator ac2704(.scan_win(scan_win2704), .rectangle1_x(rectangle1_xs[2704]), .rectangle1_y(rectangle1_ys[2704]), .rectangle1_width(rectangle1_widths[2704]), .rectangle1_height(rectangle1_heights[2704]), .rectangle1_weight(rectangle1_weights[2704]), .rectangle2_x(rectangle2_xs[2704]), .rectangle2_y(rectangle2_ys[2704]), .rectangle2_width(rectangle2_widths[2704]), .rectangle2_height(rectangle2_heights[2704]), .rectangle2_weight(rectangle2_weights[2704]), .rectangle3_x(rectangle3_xs[2704]), .rectangle3_y(rectangle3_ys[2704]), .rectangle3_width(rectangle3_widths[2704]), .rectangle3_height(rectangle3_heights[2704]), .rectangle3_weight(rectangle3_weights[2704]), .feature_threshold(feature_thresholds[2704]), .feature_above(feature_aboves[2704]), .feature_below(feature_belows[2704]), .scan_win_std_dev(scan_win_std_dev[2704]), .feature_accum(feature_accums[2704]));
  accum_calculator ac2705(.scan_win(scan_win2705), .rectangle1_x(rectangle1_xs[2705]), .rectangle1_y(rectangle1_ys[2705]), .rectangle1_width(rectangle1_widths[2705]), .rectangle1_height(rectangle1_heights[2705]), .rectangle1_weight(rectangle1_weights[2705]), .rectangle2_x(rectangle2_xs[2705]), .rectangle2_y(rectangle2_ys[2705]), .rectangle2_width(rectangle2_widths[2705]), .rectangle2_height(rectangle2_heights[2705]), .rectangle2_weight(rectangle2_weights[2705]), .rectangle3_x(rectangle3_xs[2705]), .rectangle3_y(rectangle3_ys[2705]), .rectangle3_width(rectangle3_widths[2705]), .rectangle3_height(rectangle3_heights[2705]), .rectangle3_weight(rectangle3_weights[2705]), .feature_threshold(feature_thresholds[2705]), .feature_above(feature_aboves[2705]), .feature_below(feature_belows[2705]), .scan_win_std_dev(scan_win_std_dev[2705]), .feature_accum(feature_accums[2705]));
  accum_calculator ac2706(.scan_win(scan_win2706), .rectangle1_x(rectangle1_xs[2706]), .rectangle1_y(rectangle1_ys[2706]), .rectangle1_width(rectangle1_widths[2706]), .rectangle1_height(rectangle1_heights[2706]), .rectangle1_weight(rectangle1_weights[2706]), .rectangle2_x(rectangle2_xs[2706]), .rectangle2_y(rectangle2_ys[2706]), .rectangle2_width(rectangle2_widths[2706]), .rectangle2_height(rectangle2_heights[2706]), .rectangle2_weight(rectangle2_weights[2706]), .rectangle3_x(rectangle3_xs[2706]), .rectangle3_y(rectangle3_ys[2706]), .rectangle3_width(rectangle3_widths[2706]), .rectangle3_height(rectangle3_heights[2706]), .rectangle3_weight(rectangle3_weights[2706]), .feature_threshold(feature_thresholds[2706]), .feature_above(feature_aboves[2706]), .feature_below(feature_belows[2706]), .scan_win_std_dev(scan_win_std_dev[2706]), .feature_accum(feature_accums[2706]));
  accum_calculator ac2707(.scan_win(scan_win2707), .rectangle1_x(rectangle1_xs[2707]), .rectangle1_y(rectangle1_ys[2707]), .rectangle1_width(rectangle1_widths[2707]), .rectangle1_height(rectangle1_heights[2707]), .rectangle1_weight(rectangle1_weights[2707]), .rectangle2_x(rectangle2_xs[2707]), .rectangle2_y(rectangle2_ys[2707]), .rectangle2_width(rectangle2_widths[2707]), .rectangle2_height(rectangle2_heights[2707]), .rectangle2_weight(rectangle2_weights[2707]), .rectangle3_x(rectangle3_xs[2707]), .rectangle3_y(rectangle3_ys[2707]), .rectangle3_width(rectangle3_widths[2707]), .rectangle3_height(rectangle3_heights[2707]), .rectangle3_weight(rectangle3_weights[2707]), .feature_threshold(feature_thresholds[2707]), .feature_above(feature_aboves[2707]), .feature_below(feature_belows[2707]), .scan_win_std_dev(scan_win_std_dev[2707]), .feature_accum(feature_accums[2707]));
  accum_calculator ac2708(.scan_win(scan_win2708), .rectangle1_x(rectangle1_xs[2708]), .rectangle1_y(rectangle1_ys[2708]), .rectangle1_width(rectangle1_widths[2708]), .rectangle1_height(rectangle1_heights[2708]), .rectangle1_weight(rectangle1_weights[2708]), .rectangle2_x(rectangle2_xs[2708]), .rectangle2_y(rectangle2_ys[2708]), .rectangle2_width(rectangle2_widths[2708]), .rectangle2_height(rectangle2_heights[2708]), .rectangle2_weight(rectangle2_weights[2708]), .rectangle3_x(rectangle3_xs[2708]), .rectangle3_y(rectangle3_ys[2708]), .rectangle3_width(rectangle3_widths[2708]), .rectangle3_height(rectangle3_heights[2708]), .rectangle3_weight(rectangle3_weights[2708]), .feature_threshold(feature_thresholds[2708]), .feature_above(feature_aboves[2708]), .feature_below(feature_belows[2708]), .scan_win_std_dev(scan_win_std_dev[2708]), .feature_accum(feature_accums[2708]));
  accum_calculator ac2709(.scan_win(scan_win2709), .rectangle1_x(rectangle1_xs[2709]), .rectangle1_y(rectangle1_ys[2709]), .rectangle1_width(rectangle1_widths[2709]), .rectangle1_height(rectangle1_heights[2709]), .rectangle1_weight(rectangle1_weights[2709]), .rectangle2_x(rectangle2_xs[2709]), .rectangle2_y(rectangle2_ys[2709]), .rectangle2_width(rectangle2_widths[2709]), .rectangle2_height(rectangle2_heights[2709]), .rectangle2_weight(rectangle2_weights[2709]), .rectangle3_x(rectangle3_xs[2709]), .rectangle3_y(rectangle3_ys[2709]), .rectangle3_width(rectangle3_widths[2709]), .rectangle3_height(rectangle3_heights[2709]), .rectangle3_weight(rectangle3_weights[2709]), .feature_threshold(feature_thresholds[2709]), .feature_above(feature_aboves[2709]), .feature_below(feature_belows[2709]), .scan_win_std_dev(scan_win_std_dev[2709]), .feature_accum(feature_accums[2709]));
  accum_calculator ac2710(.scan_win(scan_win2710), .rectangle1_x(rectangle1_xs[2710]), .rectangle1_y(rectangle1_ys[2710]), .rectangle1_width(rectangle1_widths[2710]), .rectangle1_height(rectangle1_heights[2710]), .rectangle1_weight(rectangle1_weights[2710]), .rectangle2_x(rectangle2_xs[2710]), .rectangle2_y(rectangle2_ys[2710]), .rectangle2_width(rectangle2_widths[2710]), .rectangle2_height(rectangle2_heights[2710]), .rectangle2_weight(rectangle2_weights[2710]), .rectangle3_x(rectangle3_xs[2710]), .rectangle3_y(rectangle3_ys[2710]), .rectangle3_width(rectangle3_widths[2710]), .rectangle3_height(rectangle3_heights[2710]), .rectangle3_weight(rectangle3_weights[2710]), .feature_threshold(feature_thresholds[2710]), .feature_above(feature_aboves[2710]), .feature_below(feature_belows[2710]), .scan_win_std_dev(scan_win_std_dev[2710]), .feature_accum(feature_accums[2710]));
  accum_calculator ac2711(.scan_win(scan_win2711), .rectangle1_x(rectangle1_xs[2711]), .rectangle1_y(rectangle1_ys[2711]), .rectangle1_width(rectangle1_widths[2711]), .rectangle1_height(rectangle1_heights[2711]), .rectangle1_weight(rectangle1_weights[2711]), .rectangle2_x(rectangle2_xs[2711]), .rectangle2_y(rectangle2_ys[2711]), .rectangle2_width(rectangle2_widths[2711]), .rectangle2_height(rectangle2_heights[2711]), .rectangle2_weight(rectangle2_weights[2711]), .rectangle3_x(rectangle3_xs[2711]), .rectangle3_y(rectangle3_ys[2711]), .rectangle3_width(rectangle3_widths[2711]), .rectangle3_height(rectangle3_heights[2711]), .rectangle3_weight(rectangle3_weights[2711]), .feature_threshold(feature_thresholds[2711]), .feature_above(feature_aboves[2711]), .feature_below(feature_belows[2711]), .scan_win_std_dev(scan_win_std_dev[2711]), .feature_accum(feature_accums[2711]));
  accum_calculator ac2712(.scan_win(scan_win2712), .rectangle1_x(rectangle1_xs[2712]), .rectangle1_y(rectangle1_ys[2712]), .rectangle1_width(rectangle1_widths[2712]), .rectangle1_height(rectangle1_heights[2712]), .rectangle1_weight(rectangle1_weights[2712]), .rectangle2_x(rectangle2_xs[2712]), .rectangle2_y(rectangle2_ys[2712]), .rectangle2_width(rectangle2_widths[2712]), .rectangle2_height(rectangle2_heights[2712]), .rectangle2_weight(rectangle2_weights[2712]), .rectangle3_x(rectangle3_xs[2712]), .rectangle3_y(rectangle3_ys[2712]), .rectangle3_width(rectangle3_widths[2712]), .rectangle3_height(rectangle3_heights[2712]), .rectangle3_weight(rectangle3_weights[2712]), .feature_threshold(feature_thresholds[2712]), .feature_above(feature_aboves[2712]), .feature_below(feature_belows[2712]), .scan_win_std_dev(scan_win_std_dev[2712]), .feature_accum(feature_accums[2712]));
  accum_calculator ac2713(.scan_win(scan_win2713), .rectangle1_x(rectangle1_xs[2713]), .rectangle1_y(rectangle1_ys[2713]), .rectangle1_width(rectangle1_widths[2713]), .rectangle1_height(rectangle1_heights[2713]), .rectangle1_weight(rectangle1_weights[2713]), .rectangle2_x(rectangle2_xs[2713]), .rectangle2_y(rectangle2_ys[2713]), .rectangle2_width(rectangle2_widths[2713]), .rectangle2_height(rectangle2_heights[2713]), .rectangle2_weight(rectangle2_weights[2713]), .rectangle3_x(rectangle3_xs[2713]), .rectangle3_y(rectangle3_ys[2713]), .rectangle3_width(rectangle3_widths[2713]), .rectangle3_height(rectangle3_heights[2713]), .rectangle3_weight(rectangle3_weights[2713]), .feature_threshold(feature_thresholds[2713]), .feature_above(feature_aboves[2713]), .feature_below(feature_belows[2713]), .scan_win_std_dev(scan_win_std_dev[2713]), .feature_accum(feature_accums[2713]));
  accum_calculator ac2714(.scan_win(scan_win2714), .rectangle1_x(rectangle1_xs[2714]), .rectangle1_y(rectangle1_ys[2714]), .rectangle1_width(rectangle1_widths[2714]), .rectangle1_height(rectangle1_heights[2714]), .rectangle1_weight(rectangle1_weights[2714]), .rectangle2_x(rectangle2_xs[2714]), .rectangle2_y(rectangle2_ys[2714]), .rectangle2_width(rectangle2_widths[2714]), .rectangle2_height(rectangle2_heights[2714]), .rectangle2_weight(rectangle2_weights[2714]), .rectangle3_x(rectangle3_xs[2714]), .rectangle3_y(rectangle3_ys[2714]), .rectangle3_width(rectangle3_widths[2714]), .rectangle3_height(rectangle3_heights[2714]), .rectangle3_weight(rectangle3_weights[2714]), .feature_threshold(feature_thresholds[2714]), .feature_above(feature_aboves[2714]), .feature_below(feature_belows[2714]), .scan_win_std_dev(scan_win_std_dev[2714]), .feature_accum(feature_accums[2714]));
  accum_calculator ac2715(.scan_win(scan_win2715), .rectangle1_x(rectangle1_xs[2715]), .rectangle1_y(rectangle1_ys[2715]), .rectangle1_width(rectangle1_widths[2715]), .rectangle1_height(rectangle1_heights[2715]), .rectangle1_weight(rectangle1_weights[2715]), .rectangle2_x(rectangle2_xs[2715]), .rectangle2_y(rectangle2_ys[2715]), .rectangle2_width(rectangle2_widths[2715]), .rectangle2_height(rectangle2_heights[2715]), .rectangle2_weight(rectangle2_weights[2715]), .rectangle3_x(rectangle3_xs[2715]), .rectangle3_y(rectangle3_ys[2715]), .rectangle3_width(rectangle3_widths[2715]), .rectangle3_height(rectangle3_heights[2715]), .rectangle3_weight(rectangle3_weights[2715]), .feature_threshold(feature_thresholds[2715]), .feature_above(feature_aboves[2715]), .feature_below(feature_belows[2715]), .scan_win_std_dev(scan_win_std_dev[2715]), .feature_accum(feature_accums[2715]));
  accum_calculator ac2716(.scan_win(scan_win2716), .rectangle1_x(rectangle1_xs[2716]), .rectangle1_y(rectangle1_ys[2716]), .rectangle1_width(rectangle1_widths[2716]), .rectangle1_height(rectangle1_heights[2716]), .rectangle1_weight(rectangle1_weights[2716]), .rectangle2_x(rectangle2_xs[2716]), .rectangle2_y(rectangle2_ys[2716]), .rectangle2_width(rectangle2_widths[2716]), .rectangle2_height(rectangle2_heights[2716]), .rectangle2_weight(rectangle2_weights[2716]), .rectangle3_x(rectangle3_xs[2716]), .rectangle3_y(rectangle3_ys[2716]), .rectangle3_width(rectangle3_widths[2716]), .rectangle3_height(rectangle3_heights[2716]), .rectangle3_weight(rectangle3_weights[2716]), .feature_threshold(feature_thresholds[2716]), .feature_above(feature_aboves[2716]), .feature_below(feature_belows[2716]), .scan_win_std_dev(scan_win_std_dev[2716]), .feature_accum(feature_accums[2716]));
  accum_calculator ac2717(.scan_win(scan_win2717), .rectangle1_x(rectangle1_xs[2717]), .rectangle1_y(rectangle1_ys[2717]), .rectangle1_width(rectangle1_widths[2717]), .rectangle1_height(rectangle1_heights[2717]), .rectangle1_weight(rectangle1_weights[2717]), .rectangle2_x(rectangle2_xs[2717]), .rectangle2_y(rectangle2_ys[2717]), .rectangle2_width(rectangle2_widths[2717]), .rectangle2_height(rectangle2_heights[2717]), .rectangle2_weight(rectangle2_weights[2717]), .rectangle3_x(rectangle3_xs[2717]), .rectangle3_y(rectangle3_ys[2717]), .rectangle3_width(rectangle3_widths[2717]), .rectangle3_height(rectangle3_heights[2717]), .rectangle3_weight(rectangle3_weights[2717]), .feature_threshold(feature_thresholds[2717]), .feature_above(feature_aboves[2717]), .feature_below(feature_belows[2717]), .scan_win_std_dev(scan_win_std_dev[2717]), .feature_accum(feature_accums[2717]));
  accum_calculator ac2718(.scan_win(scan_win2718), .rectangle1_x(rectangle1_xs[2718]), .rectangle1_y(rectangle1_ys[2718]), .rectangle1_width(rectangle1_widths[2718]), .rectangle1_height(rectangle1_heights[2718]), .rectangle1_weight(rectangle1_weights[2718]), .rectangle2_x(rectangle2_xs[2718]), .rectangle2_y(rectangle2_ys[2718]), .rectangle2_width(rectangle2_widths[2718]), .rectangle2_height(rectangle2_heights[2718]), .rectangle2_weight(rectangle2_weights[2718]), .rectangle3_x(rectangle3_xs[2718]), .rectangle3_y(rectangle3_ys[2718]), .rectangle3_width(rectangle3_widths[2718]), .rectangle3_height(rectangle3_heights[2718]), .rectangle3_weight(rectangle3_weights[2718]), .feature_threshold(feature_thresholds[2718]), .feature_above(feature_aboves[2718]), .feature_below(feature_belows[2718]), .scan_win_std_dev(scan_win_std_dev[2718]), .feature_accum(feature_accums[2718]));
  accum_calculator ac2719(.scan_win(scan_win2719), .rectangle1_x(rectangle1_xs[2719]), .rectangle1_y(rectangle1_ys[2719]), .rectangle1_width(rectangle1_widths[2719]), .rectangle1_height(rectangle1_heights[2719]), .rectangle1_weight(rectangle1_weights[2719]), .rectangle2_x(rectangle2_xs[2719]), .rectangle2_y(rectangle2_ys[2719]), .rectangle2_width(rectangle2_widths[2719]), .rectangle2_height(rectangle2_heights[2719]), .rectangle2_weight(rectangle2_weights[2719]), .rectangle3_x(rectangle3_xs[2719]), .rectangle3_y(rectangle3_ys[2719]), .rectangle3_width(rectangle3_widths[2719]), .rectangle3_height(rectangle3_heights[2719]), .rectangle3_weight(rectangle3_weights[2719]), .feature_threshold(feature_thresholds[2719]), .feature_above(feature_aboves[2719]), .feature_below(feature_belows[2719]), .scan_win_std_dev(scan_win_std_dev[2719]), .feature_accum(feature_accums[2719]));
  accum_calculator ac2720(.scan_win(scan_win2720), .rectangle1_x(rectangle1_xs[2720]), .rectangle1_y(rectangle1_ys[2720]), .rectangle1_width(rectangle1_widths[2720]), .rectangle1_height(rectangle1_heights[2720]), .rectangle1_weight(rectangle1_weights[2720]), .rectangle2_x(rectangle2_xs[2720]), .rectangle2_y(rectangle2_ys[2720]), .rectangle2_width(rectangle2_widths[2720]), .rectangle2_height(rectangle2_heights[2720]), .rectangle2_weight(rectangle2_weights[2720]), .rectangle3_x(rectangle3_xs[2720]), .rectangle3_y(rectangle3_ys[2720]), .rectangle3_width(rectangle3_widths[2720]), .rectangle3_height(rectangle3_heights[2720]), .rectangle3_weight(rectangle3_weights[2720]), .feature_threshold(feature_thresholds[2720]), .feature_above(feature_aboves[2720]), .feature_below(feature_belows[2720]), .scan_win_std_dev(scan_win_std_dev[2720]), .feature_accum(feature_accums[2720]));
  accum_calculator ac2721(.scan_win(scan_win2721), .rectangle1_x(rectangle1_xs[2721]), .rectangle1_y(rectangle1_ys[2721]), .rectangle1_width(rectangle1_widths[2721]), .rectangle1_height(rectangle1_heights[2721]), .rectangle1_weight(rectangle1_weights[2721]), .rectangle2_x(rectangle2_xs[2721]), .rectangle2_y(rectangle2_ys[2721]), .rectangle2_width(rectangle2_widths[2721]), .rectangle2_height(rectangle2_heights[2721]), .rectangle2_weight(rectangle2_weights[2721]), .rectangle3_x(rectangle3_xs[2721]), .rectangle3_y(rectangle3_ys[2721]), .rectangle3_width(rectangle3_widths[2721]), .rectangle3_height(rectangle3_heights[2721]), .rectangle3_weight(rectangle3_weights[2721]), .feature_threshold(feature_thresholds[2721]), .feature_above(feature_aboves[2721]), .feature_below(feature_belows[2721]), .scan_win_std_dev(scan_win_std_dev[2721]), .feature_accum(feature_accums[2721]));
  accum_calculator ac2722(.scan_win(scan_win2722), .rectangle1_x(rectangle1_xs[2722]), .rectangle1_y(rectangle1_ys[2722]), .rectangle1_width(rectangle1_widths[2722]), .rectangle1_height(rectangle1_heights[2722]), .rectangle1_weight(rectangle1_weights[2722]), .rectangle2_x(rectangle2_xs[2722]), .rectangle2_y(rectangle2_ys[2722]), .rectangle2_width(rectangle2_widths[2722]), .rectangle2_height(rectangle2_heights[2722]), .rectangle2_weight(rectangle2_weights[2722]), .rectangle3_x(rectangle3_xs[2722]), .rectangle3_y(rectangle3_ys[2722]), .rectangle3_width(rectangle3_widths[2722]), .rectangle3_height(rectangle3_heights[2722]), .rectangle3_weight(rectangle3_weights[2722]), .feature_threshold(feature_thresholds[2722]), .feature_above(feature_aboves[2722]), .feature_below(feature_belows[2722]), .scan_win_std_dev(scan_win_std_dev[2722]), .feature_accum(feature_accums[2722]));
  accum_calculator ac2723(.scan_win(scan_win2723), .rectangle1_x(rectangle1_xs[2723]), .rectangle1_y(rectangle1_ys[2723]), .rectangle1_width(rectangle1_widths[2723]), .rectangle1_height(rectangle1_heights[2723]), .rectangle1_weight(rectangle1_weights[2723]), .rectangle2_x(rectangle2_xs[2723]), .rectangle2_y(rectangle2_ys[2723]), .rectangle2_width(rectangle2_widths[2723]), .rectangle2_height(rectangle2_heights[2723]), .rectangle2_weight(rectangle2_weights[2723]), .rectangle3_x(rectangle3_xs[2723]), .rectangle3_y(rectangle3_ys[2723]), .rectangle3_width(rectangle3_widths[2723]), .rectangle3_height(rectangle3_heights[2723]), .rectangle3_weight(rectangle3_weights[2723]), .feature_threshold(feature_thresholds[2723]), .feature_above(feature_aboves[2723]), .feature_below(feature_belows[2723]), .scan_win_std_dev(scan_win_std_dev[2723]), .feature_accum(feature_accums[2723]));
  accum_calculator ac2724(.scan_win(scan_win2724), .rectangle1_x(rectangle1_xs[2724]), .rectangle1_y(rectangle1_ys[2724]), .rectangle1_width(rectangle1_widths[2724]), .rectangle1_height(rectangle1_heights[2724]), .rectangle1_weight(rectangle1_weights[2724]), .rectangle2_x(rectangle2_xs[2724]), .rectangle2_y(rectangle2_ys[2724]), .rectangle2_width(rectangle2_widths[2724]), .rectangle2_height(rectangle2_heights[2724]), .rectangle2_weight(rectangle2_weights[2724]), .rectangle3_x(rectangle3_xs[2724]), .rectangle3_y(rectangle3_ys[2724]), .rectangle3_width(rectangle3_widths[2724]), .rectangle3_height(rectangle3_heights[2724]), .rectangle3_weight(rectangle3_weights[2724]), .feature_threshold(feature_thresholds[2724]), .feature_above(feature_aboves[2724]), .feature_below(feature_belows[2724]), .scan_win_std_dev(scan_win_std_dev[2724]), .feature_accum(feature_accums[2724]));
  accum_calculator ac2725(.scan_win(scan_win2725), .rectangle1_x(rectangle1_xs[2725]), .rectangle1_y(rectangle1_ys[2725]), .rectangle1_width(rectangle1_widths[2725]), .rectangle1_height(rectangle1_heights[2725]), .rectangle1_weight(rectangle1_weights[2725]), .rectangle2_x(rectangle2_xs[2725]), .rectangle2_y(rectangle2_ys[2725]), .rectangle2_width(rectangle2_widths[2725]), .rectangle2_height(rectangle2_heights[2725]), .rectangle2_weight(rectangle2_weights[2725]), .rectangle3_x(rectangle3_xs[2725]), .rectangle3_y(rectangle3_ys[2725]), .rectangle3_width(rectangle3_widths[2725]), .rectangle3_height(rectangle3_heights[2725]), .rectangle3_weight(rectangle3_weights[2725]), .feature_threshold(feature_thresholds[2725]), .feature_above(feature_aboves[2725]), .feature_below(feature_belows[2725]), .scan_win_std_dev(scan_win_std_dev[2725]), .feature_accum(feature_accums[2725]));
  accum_calculator ac2726(.scan_win(scan_win2726), .rectangle1_x(rectangle1_xs[2726]), .rectangle1_y(rectangle1_ys[2726]), .rectangle1_width(rectangle1_widths[2726]), .rectangle1_height(rectangle1_heights[2726]), .rectangle1_weight(rectangle1_weights[2726]), .rectangle2_x(rectangle2_xs[2726]), .rectangle2_y(rectangle2_ys[2726]), .rectangle2_width(rectangle2_widths[2726]), .rectangle2_height(rectangle2_heights[2726]), .rectangle2_weight(rectangle2_weights[2726]), .rectangle3_x(rectangle3_xs[2726]), .rectangle3_y(rectangle3_ys[2726]), .rectangle3_width(rectangle3_widths[2726]), .rectangle3_height(rectangle3_heights[2726]), .rectangle3_weight(rectangle3_weights[2726]), .feature_threshold(feature_thresholds[2726]), .feature_above(feature_aboves[2726]), .feature_below(feature_belows[2726]), .scan_win_std_dev(scan_win_std_dev[2726]), .feature_accum(feature_accums[2726]));
  accum_calculator ac2727(.scan_win(scan_win2727), .rectangle1_x(rectangle1_xs[2727]), .rectangle1_y(rectangle1_ys[2727]), .rectangle1_width(rectangle1_widths[2727]), .rectangle1_height(rectangle1_heights[2727]), .rectangle1_weight(rectangle1_weights[2727]), .rectangle2_x(rectangle2_xs[2727]), .rectangle2_y(rectangle2_ys[2727]), .rectangle2_width(rectangle2_widths[2727]), .rectangle2_height(rectangle2_heights[2727]), .rectangle2_weight(rectangle2_weights[2727]), .rectangle3_x(rectangle3_xs[2727]), .rectangle3_y(rectangle3_ys[2727]), .rectangle3_width(rectangle3_widths[2727]), .rectangle3_height(rectangle3_heights[2727]), .rectangle3_weight(rectangle3_weights[2727]), .feature_threshold(feature_thresholds[2727]), .feature_above(feature_aboves[2727]), .feature_below(feature_belows[2727]), .scan_win_std_dev(scan_win_std_dev[2727]), .feature_accum(feature_accums[2727]));
  accum_calculator ac2728(.scan_win(scan_win2728), .rectangle1_x(rectangle1_xs[2728]), .rectangle1_y(rectangle1_ys[2728]), .rectangle1_width(rectangle1_widths[2728]), .rectangle1_height(rectangle1_heights[2728]), .rectangle1_weight(rectangle1_weights[2728]), .rectangle2_x(rectangle2_xs[2728]), .rectangle2_y(rectangle2_ys[2728]), .rectangle2_width(rectangle2_widths[2728]), .rectangle2_height(rectangle2_heights[2728]), .rectangle2_weight(rectangle2_weights[2728]), .rectangle3_x(rectangle3_xs[2728]), .rectangle3_y(rectangle3_ys[2728]), .rectangle3_width(rectangle3_widths[2728]), .rectangle3_height(rectangle3_heights[2728]), .rectangle3_weight(rectangle3_weights[2728]), .feature_threshold(feature_thresholds[2728]), .feature_above(feature_aboves[2728]), .feature_below(feature_belows[2728]), .scan_win_std_dev(scan_win_std_dev[2728]), .feature_accum(feature_accums[2728]));
  accum_calculator ac2729(.scan_win(scan_win2729), .rectangle1_x(rectangle1_xs[2729]), .rectangle1_y(rectangle1_ys[2729]), .rectangle1_width(rectangle1_widths[2729]), .rectangle1_height(rectangle1_heights[2729]), .rectangle1_weight(rectangle1_weights[2729]), .rectangle2_x(rectangle2_xs[2729]), .rectangle2_y(rectangle2_ys[2729]), .rectangle2_width(rectangle2_widths[2729]), .rectangle2_height(rectangle2_heights[2729]), .rectangle2_weight(rectangle2_weights[2729]), .rectangle3_x(rectangle3_xs[2729]), .rectangle3_y(rectangle3_ys[2729]), .rectangle3_width(rectangle3_widths[2729]), .rectangle3_height(rectangle3_heights[2729]), .rectangle3_weight(rectangle3_weights[2729]), .feature_threshold(feature_thresholds[2729]), .feature_above(feature_aboves[2729]), .feature_below(feature_belows[2729]), .scan_win_std_dev(scan_win_std_dev[2729]), .feature_accum(feature_accums[2729]));
  accum_calculator ac2730(.scan_win(scan_win2730), .rectangle1_x(rectangle1_xs[2730]), .rectangle1_y(rectangle1_ys[2730]), .rectangle1_width(rectangle1_widths[2730]), .rectangle1_height(rectangle1_heights[2730]), .rectangle1_weight(rectangle1_weights[2730]), .rectangle2_x(rectangle2_xs[2730]), .rectangle2_y(rectangle2_ys[2730]), .rectangle2_width(rectangle2_widths[2730]), .rectangle2_height(rectangle2_heights[2730]), .rectangle2_weight(rectangle2_weights[2730]), .rectangle3_x(rectangle3_xs[2730]), .rectangle3_y(rectangle3_ys[2730]), .rectangle3_width(rectangle3_widths[2730]), .rectangle3_height(rectangle3_heights[2730]), .rectangle3_weight(rectangle3_weights[2730]), .feature_threshold(feature_thresholds[2730]), .feature_above(feature_aboves[2730]), .feature_below(feature_belows[2730]), .scan_win_std_dev(scan_win_std_dev[2730]), .feature_accum(feature_accums[2730]));
  accum_calculator ac2731(.scan_win(scan_win2731), .rectangle1_x(rectangle1_xs[2731]), .rectangle1_y(rectangle1_ys[2731]), .rectangle1_width(rectangle1_widths[2731]), .rectangle1_height(rectangle1_heights[2731]), .rectangle1_weight(rectangle1_weights[2731]), .rectangle2_x(rectangle2_xs[2731]), .rectangle2_y(rectangle2_ys[2731]), .rectangle2_width(rectangle2_widths[2731]), .rectangle2_height(rectangle2_heights[2731]), .rectangle2_weight(rectangle2_weights[2731]), .rectangle3_x(rectangle3_xs[2731]), .rectangle3_y(rectangle3_ys[2731]), .rectangle3_width(rectangle3_widths[2731]), .rectangle3_height(rectangle3_heights[2731]), .rectangle3_weight(rectangle3_weights[2731]), .feature_threshold(feature_thresholds[2731]), .feature_above(feature_aboves[2731]), .feature_below(feature_belows[2731]), .scan_win_std_dev(scan_win_std_dev[2731]), .feature_accum(feature_accums[2731]));
  accum_calculator ac2732(.scan_win(scan_win2732), .rectangle1_x(rectangle1_xs[2732]), .rectangle1_y(rectangle1_ys[2732]), .rectangle1_width(rectangle1_widths[2732]), .rectangle1_height(rectangle1_heights[2732]), .rectangle1_weight(rectangle1_weights[2732]), .rectangle2_x(rectangle2_xs[2732]), .rectangle2_y(rectangle2_ys[2732]), .rectangle2_width(rectangle2_widths[2732]), .rectangle2_height(rectangle2_heights[2732]), .rectangle2_weight(rectangle2_weights[2732]), .rectangle3_x(rectangle3_xs[2732]), .rectangle3_y(rectangle3_ys[2732]), .rectangle3_width(rectangle3_widths[2732]), .rectangle3_height(rectangle3_heights[2732]), .rectangle3_weight(rectangle3_weights[2732]), .feature_threshold(feature_thresholds[2732]), .feature_above(feature_aboves[2732]), .feature_below(feature_belows[2732]), .scan_win_std_dev(scan_win_std_dev[2732]), .feature_accum(feature_accums[2732]));
  accum_calculator ac2733(.scan_win(scan_win2733), .rectangle1_x(rectangle1_xs[2733]), .rectangle1_y(rectangle1_ys[2733]), .rectangle1_width(rectangle1_widths[2733]), .rectangle1_height(rectangle1_heights[2733]), .rectangle1_weight(rectangle1_weights[2733]), .rectangle2_x(rectangle2_xs[2733]), .rectangle2_y(rectangle2_ys[2733]), .rectangle2_width(rectangle2_widths[2733]), .rectangle2_height(rectangle2_heights[2733]), .rectangle2_weight(rectangle2_weights[2733]), .rectangle3_x(rectangle3_xs[2733]), .rectangle3_y(rectangle3_ys[2733]), .rectangle3_width(rectangle3_widths[2733]), .rectangle3_height(rectangle3_heights[2733]), .rectangle3_weight(rectangle3_weights[2733]), .feature_threshold(feature_thresholds[2733]), .feature_above(feature_aboves[2733]), .feature_below(feature_belows[2733]), .scan_win_std_dev(scan_win_std_dev[2733]), .feature_accum(feature_accums[2733]));
  accum_calculator ac2734(.scan_win(scan_win2734), .rectangle1_x(rectangle1_xs[2734]), .rectangle1_y(rectangle1_ys[2734]), .rectangle1_width(rectangle1_widths[2734]), .rectangle1_height(rectangle1_heights[2734]), .rectangle1_weight(rectangle1_weights[2734]), .rectangle2_x(rectangle2_xs[2734]), .rectangle2_y(rectangle2_ys[2734]), .rectangle2_width(rectangle2_widths[2734]), .rectangle2_height(rectangle2_heights[2734]), .rectangle2_weight(rectangle2_weights[2734]), .rectangle3_x(rectangle3_xs[2734]), .rectangle3_y(rectangle3_ys[2734]), .rectangle3_width(rectangle3_widths[2734]), .rectangle3_height(rectangle3_heights[2734]), .rectangle3_weight(rectangle3_weights[2734]), .feature_threshold(feature_thresholds[2734]), .feature_above(feature_aboves[2734]), .feature_below(feature_belows[2734]), .scan_win_std_dev(scan_win_std_dev[2734]), .feature_accum(feature_accums[2734]));
  accum_calculator ac2735(.scan_win(scan_win2735), .rectangle1_x(rectangle1_xs[2735]), .rectangle1_y(rectangle1_ys[2735]), .rectangle1_width(rectangle1_widths[2735]), .rectangle1_height(rectangle1_heights[2735]), .rectangle1_weight(rectangle1_weights[2735]), .rectangle2_x(rectangle2_xs[2735]), .rectangle2_y(rectangle2_ys[2735]), .rectangle2_width(rectangle2_widths[2735]), .rectangle2_height(rectangle2_heights[2735]), .rectangle2_weight(rectangle2_weights[2735]), .rectangle3_x(rectangle3_xs[2735]), .rectangle3_y(rectangle3_ys[2735]), .rectangle3_width(rectangle3_widths[2735]), .rectangle3_height(rectangle3_heights[2735]), .rectangle3_weight(rectangle3_weights[2735]), .feature_threshold(feature_thresholds[2735]), .feature_above(feature_aboves[2735]), .feature_below(feature_belows[2735]), .scan_win_std_dev(scan_win_std_dev[2735]), .feature_accum(feature_accums[2735]));
  accum_calculator ac2736(.scan_win(scan_win2736), .rectangle1_x(rectangle1_xs[2736]), .rectangle1_y(rectangle1_ys[2736]), .rectangle1_width(rectangle1_widths[2736]), .rectangle1_height(rectangle1_heights[2736]), .rectangle1_weight(rectangle1_weights[2736]), .rectangle2_x(rectangle2_xs[2736]), .rectangle2_y(rectangle2_ys[2736]), .rectangle2_width(rectangle2_widths[2736]), .rectangle2_height(rectangle2_heights[2736]), .rectangle2_weight(rectangle2_weights[2736]), .rectangle3_x(rectangle3_xs[2736]), .rectangle3_y(rectangle3_ys[2736]), .rectangle3_width(rectangle3_widths[2736]), .rectangle3_height(rectangle3_heights[2736]), .rectangle3_weight(rectangle3_weights[2736]), .feature_threshold(feature_thresholds[2736]), .feature_above(feature_aboves[2736]), .feature_below(feature_belows[2736]), .scan_win_std_dev(scan_win_std_dev[2736]), .feature_accum(feature_accums[2736]));
  accum_calculator ac2737(.scan_win(scan_win2737), .rectangle1_x(rectangle1_xs[2737]), .rectangle1_y(rectangle1_ys[2737]), .rectangle1_width(rectangle1_widths[2737]), .rectangle1_height(rectangle1_heights[2737]), .rectangle1_weight(rectangle1_weights[2737]), .rectangle2_x(rectangle2_xs[2737]), .rectangle2_y(rectangle2_ys[2737]), .rectangle2_width(rectangle2_widths[2737]), .rectangle2_height(rectangle2_heights[2737]), .rectangle2_weight(rectangle2_weights[2737]), .rectangle3_x(rectangle3_xs[2737]), .rectangle3_y(rectangle3_ys[2737]), .rectangle3_width(rectangle3_widths[2737]), .rectangle3_height(rectangle3_heights[2737]), .rectangle3_weight(rectangle3_weights[2737]), .feature_threshold(feature_thresholds[2737]), .feature_above(feature_aboves[2737]), .feature_below(feature_belows[2737]), .scan_win_std_dev(scan_win_std_dev[2737]), .feature_accum(feature_accums[2737]));
  accum_calculator ac2738(.scan_win(scan_win2738), .rectangle1_x(rectangle1_xs[2738]), .rectangle1_y(rectangle1_ys[2738]), .rectangle1_width(rectangle1_widths[2738]), .rectangle1_height(rectangle1_heights[2738]), .rectangle1_weight(rectangle1_weights[2738]), .rectangle2_x(rectangle2_xs[2738]), .rectangle2_y(rectangle2_ys[2738]), .rectangle2_width(rectangle2_widths[2738]), .rectangle2_height(rectangle2_heights[2738]), .rectangle2_weight(rectangle2_weights[2738]), .rectangle3_x(rectangle3_xs[2738]), .rectangle3_y(rectangle3_ys[2738]), .rectangle3_width(rectangle3_widths[2738]), .rectangle3_height(rectangle3_heights[2738]), .rectangle3_weight(rectangle3_weights[2738]), .feature_threshold(feature_thresholds[2738]), .feature_above(feature_aboves[2738]), .feature_below(feature_belows[2738]), .scan_win_std_dev(scan_win_std_dev[2738]), .feature_accum(feature_accums[2738]));
  accum_calculator ac2739(.scan_win(scan_win2739), .rectangle1_x(rectangle1_xs[2739]), .rectangle1_y(rectangle1_ys[2739]), .rectangle1_width(rectangle1_widths[2739]), .rectangle1_height(rectangle1_heights[2739]), .rectangle1_weight(rectangle1_weights[2739]), .rectangle2_x(rectangle2_xs[2739]), .rectangle2_y(rectangle2_ys[2739]), .rectangle2_width(rectangle2_widths[2739]), .rectangle2_height(rectangle2_heights[2739]), .rectangle2_weight(rectangle2_weights[2739]), .rectangle3_x(rectangle3_xs[2739]), .rectangle3_y(rectangle3_ys[2739]), .rectangle3_width(rectangle3_widths[2739]), .rectangle3_height(rectangle3_heights[2739]), .rectangle3_weight(rectangle3_weights[2739]), .feature_threshold(feature_thresholds[2739]), .feature_above(feature_aboves[2739]), .feature_below(feature_belows[2739]), .scan_win_std_dev(scan_win_std_dev[2739]), .feature_accum(feature_accums[2739]));
  accum_calculator ac2740(.scan_win(scan_win2740), .rectangle1_x(rectangle1_xs[2740]), .rectangle1_y(rectangle1_ys[2740]), .rectangle1_width(rectangle1_widths[2740]), .rectangle1_height(rectangle1_heights[2740]), .rectangle1_weight(rectangle1_weights[2740]), .rectangle2_x(rectangle2_xs[2740]), .rectangle2_y(rectangle2_ys[2740]), .rectangle2_width(rectangle2_widths[2740]), .rectangle2_height(rectangle2_heights[2740]), .rectangle2_weight(rectangle2_weights[2740]), .rectangle3_x(rectangle3_xs[2740]), .rectangle3_y(rectangle3_ys[2740]), .rectangle3_width(rectangle3_widths[2740]), .rectangle3_height(rectangle3_heights[2740]), .rectangle3_weight(rectangle3_weights[2740]), .feature_threshold(feature_thresholds[2740]), .feature_above(feature_aboves[2740]), .feature_below(feature_belows[2740]), .scan_win_std_dev(scan_win_std_dev[2740]), .feature_accum(feature_accums[2740]));
  accum_calculator ac2741(.scan_win(scan_win2741), .rectangle1_x(rectangle1_xs[2741]), .rectangle1_y(rectangle1_ys[2741]), .rectangle1_width(rectangle1_widths[2741]), .rectangle1_height(rectangle1_heights[2741]), .rectangle1_weight(rectangle1_weights[2741]), .rectangle2_x(rectangle2_xs[2741]), .rectangle2_y(rectangle2_ys[2741]), .rectangle2_width(rectangle2_widths[2741]), .rectangle2_height(rectangle2_heights[2741]), .rectangle2_weight(rectangle2_weights[2741]), .rectangle3_x(rectangle3_xs[2741]), .rectangle3_y(rectangle3_ys[2741]), .rectangle3_width(rectangle3_widths[2741]), .rectangle3_height(rectangle3_heights[2741]), .rectangle3_weight(rectangle3_weights[2741]), .feature_threshold(feature_thresholds[2741]), .feature_above(feature_aboves[2741]), .feature_below(feature_belows[2741]), .scan_win_std_dev(scan_win_std_dev[2741]), .feature_accum(feature_accums[2741]));
  accum_calculator ac2742(.scan_win(scan_win2742), .rectangle1_x(rectangle1_xs[2742]), .rectangle1_y(rectangle1_ys[2742]), .rectangle1_width(rectangle1_widths[2742]), .rectangle1_height(rectangle1_heights[2742]), .rectangle1_weight(rectangle1_weights[2742]), .rectangle2_x(rectangle2_xs[2742]), .rectangle2_y(rectangle2_ys[2742]), .rectangle2_width(rectangle2_widths[2742]), .rectangle2_height(rectangle2_heights[2742]), .rectangle2_weight(rectangle2_weights[2742]), .rectangle3_x(rectangle3_xs[2742]), .rectangle3_y(rectangle3_ys[2742]), .rectangle3_width(rectangle3_widths[2742]), .rectangle3_height(rectangle3_heights[2742]), .rectangle3_weight(rectangle3_weights[2742]), .feature_threshold(feature_thresholds[2742]), .feature_above(feature_aboves[2742]), .feature_below(feature_belows[2742]), .scan_win_std_dev(scan_win_std_dev[2742]), .feature_accum(feature_accums[2742]));
  accum_calculator ac2743(.scan_win(scan_win2743), .rectangle1_x(rectangle1_xs[2743]), .rectangle1_y(rectangle1_ys[2743]), .rectangle1_width(rectangle1_widths[2743]), .rectangle1_height(rectangle1_heights[2743]), .rectangle1_weight(rectangle1_weights[2743]), .rectangle2_x(rectangle2_xs[2743]), .rectangle2_y(rectangle2_ys[2743]), .rectangle2_width(rectangle2_widths[2743]), .rectangle2_height(rectangle2_heights[2743]), .rectangle2_weight(rectangle2_weights[2743]), .rectangle3_x(rectangle3_xs[2743]), .rectangle3_y(rectangle3_ys[2743]), .rectangle3_width(rectangle3_widths[2743]), .rectangle3_height(rectangle3_heights[2743]), .rectangle3_weight(rectangle3_weights[2743]), .feature_threshold(feature_thresholds[2743]), .feature_above(feature_aboves[2743]), .feature_below(feature_belows[2743]), .scan_win_std_dev(scan_win_std_dev[2743]), .feature_accum(feature_accums[2743]));
  accum_calculator ac2744(.scan_win(scan_win2744), .rectangle1_x(rectangle1_xs[2744]), .rectangle1_y(rectangle1_ys[2744]), .rectangle1_width(rectangle1_widths[2744]), .rectangle1_height(rectangle1_heights[2744]), .rectangle1_weight(rectangle1_weights[2744]), .rectangle2_x(rectangle2_xs[2744]), .rectangle2_y(rectangle2_ys[2744]), .rectangle2_width(rectangle2_widths[2744]), .rectangle2_height(rectangle2_heights[2744]), .rectangle2_weight(rectangle2_weights[2744]), .rectangle3_x(rectangle3_xs[2744]), .rectangle3_y(rectangle3_ys[2744]), .rectangle3_width(rectangle3_widths[2744]), .rectangle3_height(rectangle3_heights[2744]), .rectangle3_weight(rectangle3_weights[2744]), .feature_threshold(feature_thresholds[2744]), .feature_above(feature_aboves[2744]), .feature_below(feature_belows[2744]), .scan_win_std_dev(scan_win_std_dev[2744]), .feature_accum(feature_accums[2744]));
  accum_calculator ac2745(.scan_win(scan_win2745), .rectangle1_x(rectangle1_xs[2745]), .rectangle1_y(rectangle1_ys[2745]), .rectangle1_width(rectangle1_widths[2745]), .rectangle1_height(rectangle1_heights[2745]), .rectangle1_weight(rectangle1_weights[2745]), .rectangle2_x(rectangle2_xs[2745]), .rectangle2_y(rectangle2_ys[2745]), .rectangle2_width(rectangle2_widths[2745]), .rectangle2_height(rectangle2_heights[2745]), .rectangle2_weight(rectangle2_weights[2745]), .rectangle3_x(rectangle3_xs[2745]), .rectangle3_y(rectangle3_ys[2745]), .rectangle3_width(rectangle3_widths[2745]), .rectangle3_height(rectangle3_heights[2745]), .rectangle3_weight(rectangle3_weights[2745]), .feature_threshold(feature_thresholds[2745]), .feature_above(feature_aboves[2745]), .feature_below(feature_belows[2745]), .scan_win_std_dev(scan_win_std_dev[2745]), .feature_accum(feature_accums[2745]));
  accum_calculator ac2746(.scan_win(scan_win2746), .rectangle1_x(rectangle1_xs[2746]), .rectangle1_y(rectangle1_ys[2746]), .rectangle1_width(rectangle1_widths[2746]), .rectangle1_height(rectangle1_heights[2746]), .rectangle1_weight(rectangle1_weights[2746]), .rectangle2_x(rectangle2_xs[2746]), .rectangle2_y(rectangle2_ys[2746]), .rectangle2_width(rectangle2_widths[2746]), .rectangle2_height(rectangle2_heights[2746]), .rectangle2_weight(rectangle2_weights[2746]), .rectangle3_x(rectangle3_xs[2746]), .rectangle3_y(rectangle3_ys[2746]), .rectangle3_width(rectangle3_widths[2746]), .rectangle3_height(rectangle3_heights[2746]), .rectangle3_weight(rectangle3_weights[2746]), .feature_threshold(feature_thresholds[2746]), .feature_above(feature_aboves[2746]), .feature_below(feature_belows[2746]), .scan_win_std_dev(scan_win_std_dev[2746]), .feature_accum(feature_accums[2746]));
  accum_calculator ac2747(.scan_win(scan_win2747), .rectangle1_x(rectangle1_xs[2747]), .rectangle1_y(rectangle1_ys[2747]), .rectangle1_width(rectangle1_widths[2747]), .rectangle1_height(rectangle1_heights[2747]), .rectangle1_weight(rectangle1_weights[2747]), .rectangle2_x(rectangle2_xs[2747]), .rectangle2_y(rectangle2_ys[2747]), .rectangle2_width(rectangle2_widths[2747]), .rectangle2_height(rectangle2_heights[2747]), .rectangle2_weight(rectangle2_weights[2747]), .rectangle3_x(rectangle3_xs[2747]), .rectangle3_y(rectangle3_ys[2747]), .rectangle3_width(rectangle3_widths[2747]), .rectangle3_height(rectangle3_heights[2747]), .rectangle3_weight(rectangle3_weights[2747]), .feature_threshold(feature_thresholds[2747]), .feature_above(feature_aboves[2747]), .feature_below(feature_belows[2747]), .scan_win_std_dev(scan_win_std_dev[2747]), .feature_accum(feature_accums[2747]));
  accum_calculator ac2748(.scan_win(scan_win2748), .rectangle1_x(rectangle1_xs[2748]), .rectangle1_y(rectangle1_ys[2748]), .rectangle1_width(rectangle1_widths[2748]), .rectangle1_height(rectangle1_heights[2748]), .rectangle1_weight(rectangle1_weights[2748]), .rectangle2_x(rectangle2_xs[2748]), .rectangle2_y(rectangle2_ys[2748]), .rectangle2_width(rectangle2_widths[2748]), .rectangle2_height(rectangle2_heights[2748]), .rectangle2_weight(rectangle2_weights[2748]), .rectangle3_x(rectangle3_xs[2748]), .rectangle3_y(rectangle3_ys[2748]), .rectangle3_width(rectangle3_widths[2748]), .rectangle3_height(rectangle3_heights[2748]), .rectangle3_weight(rectangle3_weights[2748]), .feature_threshold(feature_thresholds[2748]), .feature_above(feature_aboves[2748]), .feature_below(feature_belows[2748]), .scan_win_std_dev(scan_win_std_dev[2748]), .feature_accum(feature_accums[2748]));
  accum_calculator ac2749(.scan_win(scan_win2749), .rectangle1_x(rectangle1_xs[2749]), .rectangle1_y(rectangle1_ys[2749]), .rectangle1_width(rectangle1_widths[2749]), .rectangle1_height(rectangle1_heights[2749]), .rectangle1_weight(rectangle1_weights[2749]), .rectangle2_x(rectangle2_xs[2749]), .rectangle2_y(rectangle2_ys[2749]), .rectangle2_width(rectangle2_widths[2749]), .rectangle2_height(rectangle2_heights[2749]), .rectangle2_weight(rectangle2_weights[2749]), .rectangle3_x(rectangle3_xs[2749]), .rectangle3_y(rectangle3_ys[2749]), .rectangle3_width(rectangle3_widths[2749]), .rectangle3_height(rectangle3_heights[2749]), .rectangle3_weight(rectangle3_weights[2749]), .feature_threshold(feature_thresholds[2749]), .feature_above(feature_aboves[2749]), .feature_below(feature_belows[2749]), .scan_win_std_dev(scan_win_std_dev[2749]), .feature_accum(feature_accums[2749]));
  accum_calculator ac2750(.scan_win(scan_win2750), .rectangle1_x(rectangle1_xs[2750]), .rectangle1_y(rectangle1_ys[2750]), .rectangle1_width(rectangle1_widths[2750]), .rectangle1_height(rectangle1_heights[2750]), .rectangle1_weight(rectangle1_weights[2750]), .rectangle2_x(rectangle2_xs[2750]), .rectangle2_y(rectangle2_ys[2750]), .rectangle2_width(rectangle2_widths[2750]), .rectangle2_height(rectangle2_heights[2750]), .rectangle2_weight(rectangle2_weights[2750]), .rectangle3_x(rectangle3_xs[2750]), .rectangle3_y(rectangle3_ys[2750]), .rectangle3_width(rectangle3_widths[2750]), .rectangle3_height(rectangle3_heights[2750]), .rectangle3_weight(rectangle3_weights[2750]), .feature_threshold(feature_thresholds[2750]), .feature_above(feature_aboves[2750]), .feature_below(feature_belows[2750]), .scan_win_std_dev(scan_win_std_dev[2750]), .feature_accum(feature_accums[2750]));
  accum_calculator ac2751(.scan_win(scan_win2751), .rectangle1_x(rectangle1_xs[2751]), .rectangle1_y(rectangle1_ys[2751]), .rectangle1_width(rectangle1_widths[2751]), .rectangle1_height(rectangle1_heights[2751]), .rectangle1_weight(rectangle1_weights[2751]), .rectangle2_x(rectangle2_xs[2751]), .rectangle2_y(rectangle2_ys[2751]), .rectangle2_width(rectangle2_widths[2751]), .rectangle2_height(rectangle2_heights[2751]), .rectangle2_weight(rectangle2_weights[2751]), .rectangle3_x(rectangle3_xs[2751]), .rectangle3_y(rectangle3_ys[2751]), .rectangle3_width(rectangle3_widths[2751]), .rectangle3_height(rectangle3_heights[2751]), .rectangle3_weight(rectangle3_weights[2751]), .feature_threshold(feature_thresholds[2751]), .feature_above(feature_aboves[2751]), .feature_below(feature_belows[2751]), .scan_win_std_dev(scan_win_std_dev[2751]), .feature_accum(feature_accums[2751]));
  accum_calculator ac2752(.scan_win(scan_win2752), .rectangle1_x(rectangle1_xs[2752]), .rectangle1_y(rectangle1_ys[2752]), .rectangle1_width(rectangle1_widths[2752]), .rectangle1_height(rectangle1_heights[2752]), .rectangle1_weight(rectangle1_weights[2752]), .rectangle2_x(rectangle2_xs[2752]), .rectangle2_y(rectangle2_ys[2752]), .rectangle2_width(rectangle2_widths[2752]), .rectangle2_height(rectangle2_heights[2752]), .rectangle2_weight(rectangle2_weights[2752]), .rectangle3_x(rectangle3_xs[2752]), .rectangle3_y(rectangle3_ys[2752]), .rectangle3_width(rectangle3_widths[2752]), .rectangle3_height(rectangle3_heights[2752]), .rectangle3_weight(rectangle3_weights[2752]), .feature_threshold(feature_thresholds[2752]), .feature_above(feature_aboves[2752]), .feature_below(feature_belows[2752]), .scan_win_std_dev(scan_win_std_dev[2752]), .feature_accum(feature_accums[2752]));
  accum_calculator ac2753(.scan_win(scan_win2753), .rectangle1_x(rectangle1_xs[2753]), .rectangle1_y(rectangle1_ys[2753]), .rectangle1_width(rectangle1_widths[2753]), .rectangle1_height(rectangle1_heights[2753]), .rectangle1_weight(rectangle1_weights[2753]), .rectangle2_x(rectangle2_xs[2753]), .rectangle2_y(rectangle2_ys[2753]), .rectangle2_width(rectangle2_widths[2753]), .rectangle2_height(rectangle2_heights[2753]), .rectangle2_weight(rectangle2_weights[2753]), .rectangle3_x(rectangle3_xs[2753]), .rectangle3_y(rectangle3_ys[2753]), .rectangle3_width(rectangle3_widths[2753]), .rectangle3_height(rectangle3_heights[2753]), .rectangle3_weight(rectangle3_weights[2753]), .feature_threshold(feature_thresholds[2753]), .feature_above(feature_aboves[2753]), .feature_below(feature_belows[2753]), .scan_win_std_dev(scan_win_std_dev[2753]), .feature_accum(feature_accums[2753]));
  accum_calculator ac2754(.scan_win(scan_win2754), .rectangle1_x(rectangle1_xs[2754]), .rectangle1_y(rectangle1_ys[2754]), .rectangle1_width(rectangle1_widths[2754]), .rectangle1_height(rectangle1_heights[2754]), .rectangle1_weight(rectangle1_weights[2754]), .rectangle2_x(rectangle2_xs[2754]), .rectangle2_y(rectangle2_ys[2754]), .rectangle2_width(rectangle2_widths[2754]), .rectangle2_height(rectangle2_heights[2754]), .rectangle2_weight(rectangle2_weights[2754]), .rectangle3_x(rectangle3_xs[2754]), .rectangle3_y(rectangle3_ys[2754]), .rectangle3_width(rectangle3_widths[2754]), .rectangle3_height(rectangle3_heights[2754]), .rectangle3_weight(rectangle3_weights[2754]), .feature_threshold(feature_thresholds[2754]), .feature_above(feature_aboves[2754]), .feature_below(feature_belows[2754]), .scan_win_std_dev(scan_win_std_dev[2754]), .feature_accum(feature_accums[2754]));
  accum_calculator ac2755(.scan_win(scan_win2755), .rectangle1_x(rectangle1_xs[2755]), .rectangle1_y(rectangle1_ys[2755]), .rectangle1_width(rectangle1_widths[2755]), .rectangle1_height(rectangle1_heights[2755]), .rectangle1_weight(rectangle1_weights[2755]), .rectangle2_x(rectangle2_xs[2755]), .rectangle2_y(rectangle2_ys[2755]), .rectangle2_width(rectangle2_widths[2755]), .rectangle2_height(rectangle2_heights[2755]), .rectangle2_weight(rectangle2_weights[2755]), .rectangle3_x(rectangle3_xs[2755]), .rectangle3_y(rectangle3_ys[2755]), .rectangle3_width(rectangle3_widths[2755]), .rectangle3_height(rectangle3_heights[2755]), .rectangle3_weight(rectangle3_weights[2755]), .feature_threshold(feature_thresholds[2755]), .feature_above(feature_aboves[2755]), .feature_below(feature_belows[2755]), .scan_win_std_dev(scan_win_std_dev[2755]), .feature_accum(feature_accums[2755]));
  accum_calculator ac2756(.scan_win(scan_win2756), .rectangle1_x(rectangle1_xs[2756]), .rectangle1_y(rectangle1_ys[2756]), .rectangle1_width(rectangle1_widths[2756]), .rectangle1_height(rectangle1_heights[2756]), .rectangle1_weight(rectangle1_weights[2756]), .rectangle2_x(rectangle2_xs[2756]), .rectangle2_y(rectangle2_ys[2756]), .rectangle2_width(rectangle2_widths[2756]), .rectangle2_height(rectangle2_heights[2756]), .rectangle2_weight(rectangle2_weights[2756]), .rectangle3_x(rectangle3_xs[2756]), .rectangle3_y(rectangle3_ys[2756]), .rectangle3_width(rectangle3_widths[2756]), .rectangle3_height(rectangle3_heights[2756]), .rectangle3_weight(rectangle3_weights[2756]), .feature_threshold(feature_thresholds[2756]), .feature_above(feature_aboves[2756]), .feature_below(feature_belows[2756]), .scan_win_std_dev(scan_win_std_dev[2756]), .feature_accum(feature_accums[2756]));
  accum_calculator ac2757(.scan_win(scan_win2757), .rectangle1_x(rectangle1_xs[2757]), .rectangle1_y(rectangle1_ys[2757]), .rectangle1_width(rectangle1_widths[2757]), .rectangle1_height(rectangle1_heights[2757]), .rectangle1_weight(rectangle1_weights[2757]), .rectangle2_x(rectangle2_xs[2757]), .rectangle2_y(rectangle2_ys[2757]), .rectangle2_width(rectangle2_widths[2757]), .rectangle2_height(rectangle2_heights[2757]), .rectangle2_weight(rectangle2_weights[2757]), .rectangle3_x(rectangle3_xs[2757]), .rectangle3_y(rectangle3_ys[2757]), .rectangle3_width(rectangle3_widths[2757]), .rectangle3_height(rectangle3_heights[2757]), .rectangle3_weight(rectangle3_weights[2757]), .feature_threshold(feature_thresholds[2757]), .feature_above(feature_aboves[2757]), .feature_below(feature_belows[2757]), .scan_win_std_dev(scan_win_std_dev[2757]), .feature_accum(feature_accums[2757]));
  accum_calculator ac2758(.scan_win(scan_win2758), .rectangle1_x(rectangle1_xs[2758]), .rectangle1_y(rectangle1_ys[2758]), .rectangle1_width(rectangle1_widths[2758]), .rectangle1_height(rectangle1_heights[2758]), .rectangle1_weight(rectangle1_weights[2758]), .rectangle2_x(rectangle2_xs[2758]), .rectangle2_y(rectangle2_ys[2758]), .rectangle2_width(rectangle2_widths[2758]), .rectangle2_height(rectangle2_heights[2758]), .rectangle2_weight(rectangle2_weights[2758]), .rectangle3_x(rectangle3_xs[2758]), .rectangle3_y(rectangle3_ys[2758]), .rectangle3_width(rectangle3_widths[2758]), .rectangle3_height(rectangle3_heights[2758]), .rectangle3_weight(rectangle3_weights[2758]), .feature_threshold(feature_thresholds[2758]), .feature_above(feature_aboves[2758]), .feature_below(feature_belows[2758]), .scan_win_std_dev(scan_win_std_dev[2758]), .feature_accum(feature_accums[2758]));
  accum_calculator ac2759(.scan_win(scan_win2759), .rectangle1_x(rectangle1_xs[2759]), .rectangle1_y(rectangle1_ys[2759]), .rectangle1_width(rectangle1_widths[2759]), .rectangle1_height(rectangle1_heights[2759]), .rectangle1_weight(rectangle1_weights[2759]), .rectangle2_x(rectangle2_xs[2759]), .rectangle2_y(rectangle2_ys[2759]), .rectangle2_width(rectangle2_widths[2759]), .rectangle2_height(rectangle2_heights[2759]), .rectangle2_weight(rectangle2_weights[2759]), .rectangle3_x(rectangle3_xs[2759]), .rectangle3_y(rectangle3_ys[2759]), .rectangle3_width(rectangle3_widths[2759]), .rectangle3_height(rectangle3_heights[2759]), .rectangle3_weight(rectangle3_weights[2759]), .feature_threshold(feature_thresholds[2759]), .feature_above(feature_aboves[2759]), .feature_below(feature_belows[2759]), .scan_win_std_dev(scan_win_std_dev[2759]), .feature_accum(feature_accums[2759]));
  accum_calculator ac2760(.scan_win(scan_win2760), .rectangle1_x(rectangle1_xs[2760]), .rectangle1_y(rectangle1_ys[2760]), .rectangle1_width(rectangle1_widths[2760]), .rectangle1_height(rectangle1_heights[2760]), .rectangle1_weight(rectangle1_weights[2760]), .rectangle2_x(rectangle2_xs[2760]), .rectangle2_y(rectangle2_ys[2760]), .rectangle2_width(rectangle2_widths[2760]), .rectangle2_height(rectangle2_heights[2760]), .rectangle2_weight(rectangle2_weights[2760]), .rectangle3_x(rectangle3_xs[2760]), .rectangle3_y(rectangle3_ys[2760]), .rectangle3_width(rectangle3_widths[2760]), .rectangle3_height(rectangle3_heights[2760]), .rectangle3_weight(rectangle3_weights[2760]), .feature_threshold(feature_thresholds[2760]), .feature_above(feature_aboves[2760]), .feature_below(feature_belows[2760]), .scan_win_std_dev(scan_win_std_dev[2760]), .feature_accum(feature_accums[2760]));
  accum_calculator ac2761(.scan_win(scan_win2761), .rectangle1_x(rectangle1_xs[2761]), .rectangle1_y(rectangle1_ys[2761]), .rectangle1_width(rectangle1_widths[2761]), .rectangle1_height(rectangle1_heights[2761]), .rectangle1_weight(rectangle1_weights[2761]), .rectangle2_x(rectangle2_xs[2761]), .rectangle2_y(rectangle2_ys[2761]), .rectangle2_width(rectangle2_widths[2761]), .rectangle2_height(rectangle2_heights[2761]), .rectangle2_weight(rectangle2_weights[2761]), .rectangle3_x(rectangle3_xs[2761]), .rectangle3_y(rectangle3_ys[2761]), .rectangle3_width(rectangle3_widths[2761]), .rectangle3_height(rectangle3_heights[2761]), .rectangle3_weight(rectangle3_weights[2761]), .feature_threshold(feature_thresholds[2761]), .feature_above(feature_aboves[2761]), .feature_below(feature_belows[2761]), .scan_win_std_dev(scan_win_std_dev[2761]), .feature_accum(feature_accums[2761]));
  accum_calculator ac2762(.scan_win(scan_win2762), .rectangle1_x(rectangle1_xs[2762]), .rectangle1_y(rectangle1_ys[2762]), .rectangle1_width(rectangle1_widths[2762]), .rectangle1_height(rectangle1_heights[2762]), .rectangle1_weight(rectangle1_weights[2762]), .rectangle2_x(rectangle2_xs[2762]), .rectangle2_y(rectangle2_ys[2762]), .rectangle2_width(rectangle2_widths[2762]), .rectangle2_height(rectangle2_heights[2762]), .rectangle2_weight(rectangle2_weights[2762]), .rectangle3_x(rectangle3_xs[2762]), .rectangle3_y(rectangle3_ys[2762]), .rectangle3_width(rectangle3_widths[2762]), .rectangle3_height(rectangle3_heights[2762]), .rectangle3_weight(rectangle3_weights[2762]), .feature_threshold(feature_thresholds[2762]), .feature_above(feature_aboves[2762]), .feature_below(feature_belows[2762]), .scan_win_std_dev(scan_win_std_dev[2762]), .feature_accum(feature_accums[2762]));
  accum_calculator ac2763(.scan_win(scan_win2763), .rectangle1_x(rectangle1_xs[2763]), .rectangle1_y(rectangle1_ys[2763]), .rectangle1_width(rectangle1_widths[2763]), .rectangle1_height(rectangle1_heights[2763]), .rectangle1_weight(rectangle1_weights[2763]), .rectangle2_x(rectangle2_xs[2763]), .rectangle2_y(rectangle2_ys[2763]), .rectangle2_width(rectangle2_widths[2763]), .rectangle2_height(rectangle2_heights[2763]), .rectangle2_weight(rectangle2_weights[2763]), .rectangle3_x(rectangle3_xs[2763]), .rectangle3_y(rectangle3_ys[2763]), .rectangle3_width(rectangle3_widths[2763]), .rectangle3_height(rectangle3_heights[2763]), .rectangle3_weight(rectangle3_weights[2763]), .feature_threshold(feature_thresholds[2763]), .feature_above(feature_aboves[2763]), .feature_below(feature_belows[2763]), .scan_win_std_dev(scan_win_std_dev[2763]), .feature_accum(feature_accums[2763]));
  accum_calculator ac2764(.scan_win(scan_win2764), .rectangle1_x(rectangle1_xs[2764]), .rectangle1_y(rectangle1_ys[2764]), .rectangle1_width(rectangle1_widths[2764]), .rectangle1_height(rectangle1_heights[2764]), .rectangle1_weight(rectangle1_weights[2764]), .rectangle2_x(rectangle2_xs[2764]), .rectangle2_y(rectangle2_ys[2764]), .rectangle2_width(rectangle2_widths[2764]), .rectangle2_height(rectangle2_heights[2764]), .rectangle2_weight(rectangle2_weights[2764]), .rectangle3_x(rectangle3_xs[2764]), .rectangle3_y(rectangle3_ys[2764]), .rectangle3_width(rectangle3_widths[2764]), .rectangle3_height(rectangle3_heights[2764]), .rectangle3_weight(rectangle3_weights[2764]), .feature_threshold(feature_thresholds[2764]), .feature_above(feature_aboves[2764]), .feature_below(feature_belows[2764]), .scan_win_std_dev(scan_win_std_dev[2764]), .feature_accum(feature_accums[2764]));
  accum_calculator ac2765(.scan_win(scan_win2765), .rectangle1_x(rectangle1_xs[2765]), .rectangle1_y(rectangle1_ys[2765]), .rectangle1_width(rectangle1_widths[2765]), .rectangle1_height(rectangle1_heights[2765]), .rectangle1_weight(rectangle1_weights[2765]), .rectangle2_x(rectangle2_xs[2765]), .rectangle2_y(rectangle2_ys[2765]), .rectangle2_width(rectangle2_widths[2765]), .rectangle2_height(rectangle2_heights[2765]), .rectangle2_weight(rectangle2_weights[2765]), .rectangle3_x(rectangle3_xs[2765]), .rectangle3_y(rectangle3_ys[2765]), .rectangle3_width(rectangle3_widths[2765]), .rectangle3_height(rectangle3_heights[2765]), .rectangle3_weight(rectangle3_weights[2765]), .feature_threshold(feature_thresholds[2765]), .feature_above(feature_aboves[2765]), .feature_below(feature_belows[2765]), .scan_win_std_dev(scan_win_std_dev[2765]), .feature_accum(feature_accums[2765]));
  accum_calculator ac2766(.scan_win(scan_win2766), .rectangle1_x(rectangle1_xs[2766]), .rectangle1_y(rectangle1_ys[2766]), .rectangle1_width(rectangle1_widths[2766]), .rectangle1_height(rectangle1_heights[2766]), .rectangle1_weight(rectangle1_weights[2766]), .rectangle2_x(rectangle2_xs[2766]), .rectangle2_y(rectangle2_ys[2766]), .rectangle2_width(rectangle2_widths[2766]), .rectangle2_height(rectangle2_heights[2766]), .rectangle2_weight(rectangle2_weights[2766]), .rectangle3_x(rectangle3_xs[2766]), .rectangle3_y(rectangle3_ys[2766]), .rectangle3_width(rectangle3_widths[2766]), .rectangle3_height(rectangle3_heights[2766]), .rectangle3_weight(rectangle3_weights[2766]), .feature_threshold(feature_thresholds[2766]), .feature_above(feature_aboves[2766]), .feature_below(feature_belows[2766]), .scan_win_std_dev(scan_win_std_dev[2766]), .feature_accum(feature_accums[2766]));
  accum_calculator ac2767(.scan_win(scan_win2767), .rectangle1_x(rectangle1_xs[2767]), .rectangle1_y(rectangle1_ys[2767]), .rectangle1_width(rectangle1_widths[2767]), .rectangle1_height(rectangle1_heights[2767]), .rectangle1_weight(rectangle1_weights[2767]), .rectangle2_x(rectangle2_xs[2767]), .rectangle2_y(rectangle2_ys[2767]), .rectangle2_width(rectangle2_widths[2767]), .rectangle2_height(rectangle2_heights[2767]), .rectangle2_weight(rectangle2_weights[2767]), .rectangle3_x(rectangle3_xs[2767]), .rectangle3_y(rectangle3_ys[2767]), .rectangle3_width(rectangle3_widths[2767]), .rectangle3_height(rectangle3_heights[2767]), .rectangle3_weight(rectangle3_weights[2767]), .feature_threshold(feature_thresholds[2767]), .feature_above(feature_aboves[2767]), .feature_below(feature_belows[2767]), .scan_win_std_dev(scan_win_std_dev[2767]), .feature_accum(feature_accums[2767]));
  accum_calculator ac2768(.scan_win(scan_win2768), .rectangle1_x(rectangle1_xs[2768]), .rectangle1_y(rectangle1_ys[2768]), .rectangle1_width(rectangle1_widths[2768]), .rectangle1_height(rectangle1_heights[2768]), .rectangle1_weight(rectangle1_weights[2768]), .rectangle2_x(rectangle2_xs[2768]), .rectangle2_y(rectangle2_ys[2768]), .rectangle2_width(rectangle2_widths[2768]), .rectangle2_height(rectangle2_heights[2768]), .rectangle2_weight(rectangle2_weights[2768]), .rectangle3_x(rectangle3_xs[2768]), .rectangle3_y(rectangle3_ys[2768]), .rectangle3_width(rectangle3_widths[2768]), .rectangle3_height(rectangle3_heights[2768]), .rectangle3_weight(rectangle3_weights[2768]), .feature_threshold(feature_thresholds[2768]), .feature_above(feature_aboves[2768]), .feature_below(feature_belows[2768]), .scan_win_std_dev(scan_win_std_dev[2768]), .feature_accum(feature_accums[2768]));
  accum_calculator ac2769(.scan_win(scan_win2769), .rectangle1_x(rectangle1_xs[2769]), .rectangle1_y(rectangle1_ys[2769]), .rectangle1_width(rectangle1_widths[2769]), .rectangle1_height(rectangle1_heights[2769]), .rectangle1_weight(rectangle1_weights[2769]), .rectangle2_x(rectangle2_xs[2769]), .rectangle2_y(rectangle2_ys[2769]), .rectangle2_width(rectangle2_widths[2769]), .rectangle2_height(rectangle2_heights[2769]), .rectangle2_weight(rectangle2_weights[2769]), .rectangle3_x(rectangle3_xs[2769]), .rectangle3_y(rectangle3_ys[2769]), .rectangle3_width(rectangle3_widths[2769]), .rectangle3_height(rectangle3_heights[2769]), .rectangle3_weight(rectangle3_weights[2769]), .feature_threshold(feature_thresholds[2769]), .feature_above(feature_aboves[2769]), .feature_below(feature_belows[2769]), .scan_win_std_dev(scan_win_std_dev[2769]), .feature_accum(feature_accums[2769]));
  accum_calculator ac2770(.scan_win(scan_win2770), .rectangle1_x(rectangle1_xs[2770]), .rectangle1_y(rectangle1_ys[2770]), .rectangle1_width(rectangle1_widths[2770]), .rectangle1_height(rectangle1_heights[2770]), .rectangle1_weight(rectangle1_weights[2770]), .rectangle2_x(rectangle2_xs[2770]), .rectangle2_y(rectangle2_ys[2770]), .rectangle2_width(rectangle2_widths[2770]), .rectangle2_height(rectangle2_heights[2770]), .rectangle2_weight(rectangle2_weights[2770]), .rectangle3_x(rectangle3_xs[2770]), .rectangle3_y(rectangle3_ys[2770]), .rectangle3_width(rectangle3_widths[2770]), .rectangle3_height(rectangle3_heights[2770]), .rectangle3_weight(rectangle3_weights[2770]), .feature_threshold(feature_thresholds[2770]), .feature_above(feature_aboves[2770]), .feature_below(feature_belows[2770]), .scan_win_std_dev(scan_win_std_dev[2770]), .feature_accum(feature_accums[2770]));
  accum_calculator ac2771(.scan_win(scan_win2771), .rectangle1_x(rectangle1_xs[2771]), .rectangle1_y(rectangle1_ys[2771]), .rectangle1_width(rectangle1_widths[2771]), .rectangle1_height(rectangle1_heights[2771]), .rectangle1_weight(rectangle1_weights[2771]), .rectangle2_x(rectangle2_xs[2771]), .rectangle2_y(rectangle2_ys[2771]), .rectangle2_width(rectangle2_widths[2771]), .rectangle2_height(rectangle2_heights[2771]), .rectangle2_weight(rectangle2_weights[2771]), .rectangle3_x(rectangle3_xs[2771]), .rectangle3_y(rectangle3_ys[2771]), .rectangle3_width(rectangle3_widths[2771]), .rectangle3_height(rectangle3_heights[2771]), .rectangle3_weight(rectangle3_weights[2771]), .feature_threshold(feature_thresholds[2771]), .feature_above(feature_aboves[2771]), .feature_below(feature_belows[2771]), .scan_win_std_dev(scan_win_std_dev[2771]), .feature_accum(feature_accums[2771]));
  accum_calculator ac2772(.scan_win(scan_win2772), .rectangle1_x(rectangle1_xs[2772]), .rectangle1_y(rectangle1_ys[2772]), .rectangle1_width(rectangle1_widths[2772]), .rectangle1_height(rectangle1_heights[2772]), .rectangle1_weight(rectangle1_weights[2772]), .rectangle2_x(rectangle2_xs[2772]), .rectangle2_y(rectangle2_ys[2772]), .rectangle2_width(rectangle2_widths[2772]), .rectangle2_height(rectangle2_heights[2772]), .rectangle2_weight(rectangle2_weights[2772]), .rectangle3_x(rectangle3_xs[2772]), .rectangle3_y(rectangle3_ys[2772]), .rectangle3_width(rectangle3_widths[2772]), .rectangle3_height(rectangle3_heights[2772]), .rectangle3_weight(rectangle3_weights[2772]), .feature_threshold(feature_thresholds[2772]), .feature_above(feature_aboves[2772]), .feature_below(feature_belows[2772]), .scan_win_std_dev(scan_win_std_dev[2772]), .feature_accum(feature_accums[2772]));
  accum_calculator ac2773(.scan_win(scan_win2773), .rectangle1_x(rectangle1_xs[2773]), .rectangle1_y(rectangle1_ys[2773]), .rectangle1_width(rectangle1_widths[2773]), .rectangle1_height(rectangle1_heights[2773]), .rectangle1_weight(rectangle1_weights[2773]), .rectangle2_x(rectangle2_xs[2773]), .rectangle2_y(rectangle2_ys[2773]), .rectangle2_width(rectangle2_widths[2773]), .rectangle2_height(rectangle2_heights[2773]), .rectangle2_weight(rectangle2_weights[2773]), .rectangle3_x(rectangle3_xs[2773]), .rectangle3_y(rectangle3_ys[2773]), .rectangle3_width(rectangle3_widths[2773]), .rectangle3_height(rectangle3_heights[2773]), .rectangle3_weight(rectangle3_weights[2773]), .feature_threshold(feature_thresholds[2773]), .feature_above(feature_aboves[2773]), .feature_below(feature_belows[2773]), .scan_win_std_dev(scan_win_std_dev[2773]), .feature_accum(feature_accums[2773]));
  accum_calculator ac2774(.scan_win(scan_win2774), .rectangle1_x(rectangle1_xs[2774]), .rectangle1_y(rectangle1_ys[2774]), .rectangle1_width(rectangle1_widths[2774]), .rectangle1_height(rectangle1_heights[2774]), .rectangle1_weight(rectangle1_weights[2774]), .rectangle2_x(rectangle2_xs[2774]), .rectangle2_y(rectangle2_ys[2774]), .rectangle2_width(rectangle2_widths[2774]), .rectangle2_height(rectangle2_heights[2774]), .rectangle2_weight(rectangle2_weights[2774]), .rectangle3_x(rectangle3_xs[2774]), .rectangle3_y(rectangle3_ys[2774]), .rectangle3_width(rectangle3_widths[2774]), .rectangle3_height(rectangle3_heights[2774]), .rectangle3_weight(rectangle3_weights[2774]), .feature_threshold(feature_thresholds[2774]), .feature_above(feature_aboves[2774]), .feature_below(feature_belows[2774]), .scan_win_std_dev(scan_win_std_dev[2774]), .feature_accum(feature_accums[2774]));
  accum_calculator ac2775(.scan_win(scan_win2775), .rectangle1_x(rectangle1_xs[2775]), .rectangle1_y(rectangle1_ys[2775]), .rectangle1_width(rectangle1_widths[2775]), .rectangle1_height(rectangle1_heights[2775]), .rectangle1_weight(rectangle1_weights[2775]), .rectangle2_x(rectangle2_xs[2775]), .rectangle2_y(rectangle2_ys[2775]), .rectangle2_width(rectangle2_widths[2775]), .rectangle2_height(rectangle2_heights[2775]), .rectangle2_weight(rectangle2_weights[2775]), .rectangle3_x(rectangle3_xs[2775]), .rectangle3_y(rectangle3_ys[2775]), .rectangle3_width(rectangle3_widths[2775]), .rectangle3_height(rectangle3_heights[2775]), .rectangle3_weight(rectangle3_weights[2775]), .feature_threshold(feature_thresholds[2775]), .feature_above(feature_aboves[2775]), .feature_below(feature_belows[2775]), .scan_win_std_dev(scan_win_std_dev[2775]), .feature_accum(feature_accums[2775]));
  accum_calculator ac2776(.scan_win(scan_win2776), .rectangle1_x(rectangle1_xs[2776]), .rectangle1_y(rectangle1_ys[2776]), .rectangle1_width(rectangle1_widths[2776]), .rectangle1_height(rectangle1_heights[2776]), .rectangle1_weight(rectangle1_weights[2776]), .rectangle2_x(rectangle2_xs[2776]), .rectangle2_y(rectangle2_ys[2776]), .rectangle2_width(rectangle2_widths[2776]), .rectangle2_height(rectangle2_heights[2776]), .rectangle2_weight(rectangle2_weights[2776]), .rectangle3_x(rectangle3_xs[2776]), .rectangle3_y(rectangle3_ys[2776]), .rectangle3_width(rectangle3_widths[2776]), .rectangle3_height(rectangle3_heights[2776]), .rectangle3_weight(rectangle3_weights[2776]), .feature_threshold(feature_thresholds[2776]), .feature_above(feature_aboves[2776]), .feature_below(feature_belows[2776]), .scan_win_std_dev(scan_win_std_dev[2776]), .feature_accum(feature_accums[2776]));
  accum_calculator ac2777(.scan_win(scan_win2777), .rectangle1_x(rectangle1_xs[2777]), .rectangle1_y(rectangle1_ys[2777]), .rectangle1_width(rectangle1_widths[2777]), .rectangle1_height(rectangle1_heights[2777]), .rectangle1_weight(rectangle1_weights[2777]), .rectangle2_x(rectangle2_xs[2777]), .rectangle2_y(rectangle2_ys[2777]), .rectangle2_width(rectangle2_widths[2777]), .rectangle2_height(rectangle2_heights[2777]), .rectangle2_weight(rectangle2_weights[2777]), .rectangle3_x(rectangle3_xs[2777]), .rectangle3_y(rectangle3_ys[2777]), .rectangle3_width(rectangle3_widths[2777]), .rectangle3_height(rectangle3_heights[2777]), .rectangle3_weight(rectangle3_weights[2777]), .feature_threshold(feature_thresholds[2777]), .feature_above(feature_aboves[2777]), .feature_below(feature_belows[2777]), .scan_win_std_dev(scan_win_std_dev[2777]), .feature_accum(feature_accums[2777]));
  accum_calculator ac2778(.scan_win(scan_win2778), .rectangle1_x(rectangle1_xs[2778]), .rectangle1_y(rectangle1_ys[2778]), .rectangle1_width(rectangle1_widths[2778]), .rectangle1_height(rectangle1_heights[2778]), .rectangle1_weight(rectangle1_weights[2778]), .rectangle2_x(rectangle2_xs[2778]), .rectangle2_y(rectangle2_ys[2778]), .rectangle2_width(rectangle2_widths[2778]), .rectangle2_height(rectangle2_heights[2778]), .rectangle2_weight(rectangle2_weights[2778]), .rectangle3_x(rectangle3_xs[2778]), .rectangle3_y(rectangle3_ys[2778]), .rectangle3_width(rectangle3_widths[2778]), .rectangle3_height(rectangle3_heights[2778]), .rectangle3_weight(rectangle3_weights[2778]), .feature_threshold(feature_thresholds[2778]), .feature_above(feature_aboves[2778]), .feature_below(feature_belows[2778]), .scan_win_std_dev(scan_win_std_dev[2778]), .feature_accum(feature_accums[2778]));
  accum_calculator ac2779(.scan_win(scan_win2779), .rectangle1_x(rectangle1_xs[2779]), .rectangle1_y(rectangle1_ys[2779]), .rectangle1_width(rectangle1_widths[2779]), .rectangle1_height(rectangle1_heights[2779]), .rectangle1_weight(rectangle1_weights[2779]), .rectangle2_x(rectangle2_xs[2779]), .rectangle2_y(rectangle2_ys[2779]), .rectangle2_width(rectangle2_widths[2779]), .rectangle2_height(rectangle2_heights[2779]), .rectangle2_weight(rectangle2_weights[2779]), .rectangle3_x(rectangle3_xs[2779]), .rectangle3_y(rectangle3_ys[2779]), .rectangle3_width(rectangle3_widths[2779]), .rectangle3_height(rectangle3_heights[2779]), .rectangle3_weight(rectangle3_weights[2779]), .feature_threshold(feature_thresholds[2779]), .feature_above(feature_aboves[2779]), .feature_below(feature_belows[2779]), .scan_win_std_dev(scan_win_std_dev[2779]), .feature_accum(feature_accums[2779]));
  accum_calculator ac2780(.scan_win(scan_win2780), .rectangle1_x(rectangle1_xs[2780]), .rectangle1_y(rectangle1_ys[2780]), .rectangle1_width(rectangle1_widths[2780]), .rectangle1_height(rectangle1_heights[2780]), .rectangle1_weight(rectangle1_weights[2780]), .rectangle2_x(rectangle2_xs[2780]), .rectangle2_y(rectangle2_ys[2780]), .rectangle2_width(rectangle2_widths[2780]), .rectangle2_height(rectangle2_heights[2780]), .rectangle2_weight(rectangle2_weights[2780]), .rectangle3_x(rectangle3_xs[2780]), .rectangle3_y(rectangle3_ys[2780]), .rectangle3_width(rectangle3_widths[2780]), .rectangle3_height(rectangle3_heights[2780]), .rectangle3_weight(rectangle3_weights[2780]), .feature_threshold(feature_thresholds[2780]), .feature_above(feature_aboves[2780]), .feature_below(feature_belows[2780]), .scan_win_std_dev(scan_win_std_dev[2780]), .feature_accum(feature_accums[2780]));
  accum_calculator ac2781(.scan_win(scan_win2781), .rectangle1_x(rectangle1_xs[2781]), .rectangle1_y(rectangle1_ys[2781]), .rectangle1_width(rectangle1_widths[2781]), .rectangle1_height(rectangle1_heights[2781]), .rectangle1_weight(rectangle1_weights[2781]), .rectangle2_x(rectangle2_xs[2781]), .rectangle2_y(rectangle2_ys[2781]), .rectangle2_width(rectangle2_widths[2781]), .rectangle2_height(rectangle2_heights[2781]), .rectangle2_weight(rectangle2_weights[2781]), .rectangle3_x(rectangle3_xs[2781]), .rectangle3_y(rectangle3_ys[2781]), .rectangle3_width(rectangle3_widths[2781]), .rectangle3_height(rectangle3_heights[2781]), .rectangle3_weight(rectangle3_weights[2781]), .feature_threshold(feature_thresholds[2781]), .feature_above(feature_aboves[2781]), .feature_below(feature_belows[2781]), .scan_win_std_dev(scan_win_std_dev[2781]), .feature_accum(feature_accums[2781]));
  accum_calculator ac2782(.scan_win(scan_win2782), .rectangle1_x(rectangle1_xs[2782]), .rectangle1_y(rectangle1_ys[2782]), .rectangle1_width(rectangle1_widths[2782]), .rectangle1_height(rectangle1_heights[2782]), .rectangle1_weight(rectangle1_weights[2782]), .rectangle2_x(rectangle2_xs[2782]), .rectangle2_y(rectangle2_ys[2782]), .rectangle2_width(rectangle2_widths[2782]), .rectangle2_height(rectangle2_heights[2782]), .rectangle2_weight(rectangle2_weights[2782]), .rectangle3_x(rectangle3_xs[2782]), .rectangle3_y(rectangle3_ys[2782]), .rectangle3_width(rectangle3_widths[2782]), .rectangle3_height(rectangle3_heights[2782]), .rectangle3_weight(rectangle3_weights[2782]), .feature_threshold(feature_thresholds[2782]), .feature_above(feature_aboves[2782]), .feature_below(feature_belows[2782]), .scan_win_std_dev(scan_win_std_dev[2782]), .feature_accum(feature_accums[2782]));
  accum_calculator ac2783(.scan_win(scan_win2783), .rectangle1_x(rectangle1_xs[2783]), .rectangle1_y(rectangle1_ys[2783]), .rectangle1_width(rectangle1_widths[2783]), .rectangle1_height(rectangle1_heights[2783]), .rectangle1_weight(rectangle1_weights[2783]), .rectangle2_x(rectangle2_xs[2783]), .rectangle2_y(rectangle2_ys[2783]), .rectangle2_width(rectangle2_widths[2783]), .rectangle2_height(rectangle2_heights[2783]), .rectangle2_weight(rectangle2_weights[2783]), .rectangle3_x(rectangle3_xs[2783]), .rectangle3_y(rectangle3_ys[2783]), .rectangle3_width(rectangle3_widths[2783]), .rectangle3_height(rectangle3_heights[2783]), .rectangle3_weight(rectangle3_weights[2783]), .feature_threshold(feature_thresholds[2783]), .feature_above(feature_aboves[2783]), .feature_below(feature_belows[2783]), .scan_win_std_dev(scan_win_std_dev[2783]), .feature_accum(feature_accums[2783]));
  accum_calculator ac2784(.scan_win(scan_win2784), .rectangle1_x(rectangle1_xs[2784]), .rectangle1_y(rectangle1_ys[2784]), .rectangle1_width(rectangle1_widths[2784]), .rectangle1_height(rectangle1_heights[2784]), .rectangle1_weight(rectangle1_weights[2784]), .rectangle2_x(rectangle2_xs[2784]), .rectangle2_y(rectangle2_ys[2784]), .rectangle2_width(rectangle2_widths[2784]), .rectangle2_height(rectangle2_heights[2784]), .rectangle2_weight(rectangle2_weights[2784]), .rectangle3_x(rectangle3_xs[2784]), .rectangle3_y(rectangle3_ys[2784]), .rectangle3_width(rectangle3_widths[2784]), .rectangle3_height(rectangle3_heights[2784]), .rectangle3_weight(rectangle3_weights[2784]), .feature_threshold(feature_thresholds[2784]), .feature_above(feature_aboves[2784]), .feature_below(feature_belows[2784]), .scan_win_std_dev(scan_win_std_dev[2784]), .feature_accum(feature_accums[2784]));
  accum_calculator ac2785(.scan_win(scan_win2785), .rectangle1_x(rectangle1_xs[2785]), .rectangle1_y(rectangle1_ys[2785]), .rectangle1_width(rectangle1_widths[2785]), .rectangle1_height(rectangle1_heights[2785]), .rectangle1_weight(rectangle1_weights[2785]), .rectangle2_x(rectangle2_xs[2785]), .rectangle2_y(rectangle2_ys[2785]), .rectangle2_width(rectangle2_widths[2785]), .rectangle2_height(rectangle2_heights[2785]), .rectangle2_weight(rectangle2_weights[2785]), .rectangle3_x(rectangle3_xs[2785]), .rectangle3_y(rectangle3_ys[2785]), .rectangle3_width(rectangle3_widths[2785]), .rectangle3_height(rectangle3_heights[2785]), .rectangle3_weight(rectangle3_weights[2785]), .feature_threshold(feature_thresholds[2785]), .feature_above(feature_aboves[2785]), .feature_below(feature_belows[2785]), .scan_win_std_dev(scan_win_std_dev[2785]), .feature_accum(feature_accums[2785]));
  accum_calculator ac2786(.scan_win(scan_win2786), .rectangle1_x(rectangle1_xs[2786]), .rectangle1_y(rectangle1_ys[2786]), .rectangle1_width(rectangle1_widths[2786]), .rectangle1_height(rectangle1_heights[2786]), .rectangle1_weight(rectangle1_weights[2786]), .rectangle2_x(rectangle2_xs[2786]), .rectangle2_y(rectangle2_ys[2786]), .rectangle2_width(rectangle2_widths[2786]), .rectangle2_height(rectangle2_heights[2786]), .rectangle2_weight(rectangle2_weights[2786]), .rectangle3_x(rectangle3_xs[2786]), .rectangle3_y(rectangle3_ys[2786]), .rectangle3_width(rectangle3_widths[2786]), .rectangle3_height(rectangle3_heights[2786]), .rectangle3_weight(rectangle3_weights[2786]), .feature_threshold(feature_thresholds[2786]), .feature_above(feature_aboves[2786]), .feature_below(feature_belows[2786]), .scan_win_std_dev(scan_win_std_dev[2786]), .feature_accum(feature_accums[2786]));
  accum_calculator ac2787(.scan_win(scan_win2787), .rectangle1_x(rectangle1_xs[2787]), .rectangle1_y(rectangle1_ys[2787]), .rectangle1_width(rectangle1_widths[2787]), .rectangle1_height(rectangle1_heights[2787]), .rectangle1_weight(rectangle1_weights[2787]), .rectangle2_x(rectangle2_xs[2787]), .rectangle2_y(rectangle2_ys[2787]), .rectangle2_width(rectangle2_widths[2787]), .rectangle2_height(rectangle2_heights[2787]), .rectangle2_weight(rectangle2_weights[2787]), .rectangle3_x(rectangle3_xs[2787]), .rectangle3_y(rectangle3_ys[2787]), .rectangle3_width(rectangle3_widths[2787]), .rectangle3_height(rectangle3_heights[2787]), .rectangle3_weight(rectangle3_weights[2787]), .feature_threshold(feature_thresholds[2787]), .feature_above(feature_aboves[2787]), .feature_below(feature_belows[2787]), .scan_win_std_dev(scan_win_std_dev[2787]), .feature_accum(feature_accums[2787]));
  accum_calculator ac2788(.scan_win(scan_win2788), .rectangle1_x(rectangle1_xs[2788]), .rectangle1_y(rectangle1_ys[2788]), .rectangle1_width(rectangle1_widths[2788]), .rectangle1_height(rectangle1_heights[2788]), .rectangle1_weight(rectangle1_weights[2788]), .rectangle2_x(rectangle2_xs[2788]), .rectangle2_y(rectangle2_ys[2788]), .rectangle2_width(rectangle2_widths[2788]), .rectangle2_height(rectangle2_heights[2788]), .rectangle2_weight(rectangle2_weights[2788]), .rectangle3_x(rectangle3_xs[2788]), .rectangle3_y(rectangle3_ys[2788]), .rectangle3_width(rectangle3_widths[2788]), .rectangle3_height(rectangle3_heights[2788]), .rectangle3_weight(rectangle3_weights[2788]), .feature_threshold(feature_thresholds[2788]), .feature_above(feature_aboves[2788]), .feature_below(feature_belows[2788]), .scan_win_std_dev(scan_win_std_dev[2788]), .feature_accum(feature_accums[2788]));
  accum_calculator ac2789(.scan_win(scan_win2789), .rectangle1_x(rectangle1_xs[2789]), .rectangle1_y(rectangle1_ys[2789]), .rectangle1_width(rectangle1_widths[2789]), .rectangle1_height(rectangle1_heights[2789]), .rectangle1_weight(rectangle1_weights[2789]), .rectangle2_x(rectangle2_xs[2789]), .rectangle2_y(rectangle2_ys[2789]), .rectangle2_width(rectangle2_widths[2789]), .rectangle2_height(rectangle2_heights[2789]), .rectangle2_weight(rectangle2_weights[2789]), .rectangle3_x(rectangle3_xs[2789]), .rectangle3_y(rectangle3_ys[2789]), .rectangle3_width(rectangle3_widths[2789]), .rectangle3_height(rectangle3_heights[2789]), .rectangle3_weight(rectangle3_weights[2789]), .feature_threshold(feature_thresholds[2789]), .feature_above(feature_aboves[2789]), .feature_below(feature_belows[2789]), .scan_win_std_dev(scan_win_std_dev[2789]), .feature_accum(feature_accums[2789]));
  accum_calculator ac2790(.scan_win(scan_win2790), .rectangle1_x(rectangle1_xs[2790]), .rectangle1_y(rectangle1_ys[2790]), .rectangle1_width(rectangle1_widths[2790]), .rectangle1_height(rectangle1_heights[2790]), .rectangle1_weight(rectangle1_weights[2790]), .rectangle2_x(rectangle2_xs[2790]), .rectangle2_y(rectangle2_ys[2790]), .rectangle2_width(rectangle2_widths[2790]), .rectangle2_height(rectangle2_heights[2790]), .rectangle2_weight(rectangle2_weights[2790]), .rectangle3_x(rectangle3_xs[2790]), .rectangle3_y(rectangle3_ys[2790]), .rectangle3_width(rectangle3_widths[2790]), .rectangle3_height(rectangle3_heights[2790]), .rectangle3_weight(rectangle3_weights[2790]), .feature_threshold(feature_thresholds[2790]), .feature_above(feature_aboves[2790]), .feature_below(feature_belows[2790]), .scan_win_std_dev(scan_win_std_dev[2790]), .feature_accum(feature_accums[2790]));
  accum_calculator ac2791(.scan_win(scan_win2791), .rectangle1_x(rectangle1_xs[2791]), .rectangle1_y(rectangle1_ys[2791]), .rectangle1_width(rectangle1_widths[2791]), .rectangle1_height(rectangle1_heights[2791]), .rectangle1_weight(rectangle1_weights[2791]), .rectangle2_x(rectangle2_xs[2791]), .rectangle2_y(rectangle2_ys[2791]), .rectangle2_width(rectangle2_widths[2791]), .rectangle2_height(rectangle2_heights[2791]), .rectangle2_weight(rectangle2_weights[2791]), .rectangle3_x(rectangle3_xs[2791]), .rectangle3_y(rectangle3_ys[2791]), .rectangle3_width(rectangle3_widths[2791]), .rectangle3_height(rectangle3_heights[2791]), .rectangle3_weight(rectangle3_weights[2791]), .feature_threshold(feature_thresholds[2791]), .feature_above(feature_aboves[2791]), .feature_below(feature_belows[2791]), .scan_win_std_dev(scan_win_std_dev[2791]), .feature_accum(feature_accums[2791]));
  accum_calculator ac2792(.scan_win(scan_win2792), .rectangle1_x(rectangle1_xs[2792]), .rectangle1_y(rectangle1_ys[2792]), .rectangle1_width(rectangle1_widths[2792]), .rectangle1_height(rectangle1_heights[2792]), .rectangle1_weight(rectangle1_weights[2792]), .rectangle2_x(rectangle2_xs[2792]), .rectangle2_y(rectangle2_ys[2792]), .rectangle2_width(rectangle2_widths[2792]), .rectangle2_height(rectangle2_heights[2792]), .rectangle2_weight(rectangle2_weights[2792]), .rectangle3_x(rectangle3_xs[2792]), .rectangle3_y(rectangle3_ys[2792]), .rectangle3_width(rectangle3_widths[2792]), .rectangle3_height(rectangle3_heights[2792]), .rectangle3_weight(rectangle3_weights[2792]), .feature_threshold(feature_thresholds[2792]), .feature_above(feature_aboves[2792]), .feature_below(feature_belows[2792]), .scan_win_std_dev(scan_win_std_dev[2792]), .feature_accum(feature_accums[2792]));
  accum_calculator ac2793(.scan_win(scan_win2793), .rectangle1_x(rectangle1_xs[2793]), .rectangle1_y(rectangle1_ys[2793]), .rectangle1_width(rectangle1_widths[2793]), .rectangle1_height(rectangle1_heights[2793]), .rectangle1_weight(rectangle1_weights[2793]), .rectangle2_x(rectangle2_xs[2793]), .rectangle2_y(rectangle2_ys[2793]), .rectangle2_width(rectangle2_widths[2793]), .rectangle2_height(rectangle2_heights[2793]), .rectangle2_weight(rectangle2_weights[2793]), .rectangle3_x(rectangle3_xs[2793]), .rectangle3_y(rectangle3_ys[2793]), .rectangle3_width(rectangle3_widths[2793]), .rectangle3_height(rectangle3_heights[2793]), .rectangle3_weight(rectangle3_weights[2793]), .feature_threshold(feature_thresholds[2793]), .feature_above(feature_aboves[2793]), .feature_below(feature_belows[2793]), .scan_win_std_dev(scan_win_std_dev[2793]), .feature_accum(feature_accums[2793]));
  accum_calculator ac2794(.scan_win(scan_win2794), .rectangle1_x(rectangle1_xs[2794]), .rectangle1_y(rectangle1_ys[2794]), .rectangle1_width(rectangle1_widths[2794]), .rectangle1_height(rectangle1_heights[2794]), .rectangle1_weight(rectangle1_weights[2794]), .rectangle2_x(rectangle2_xs[2794]), .rectangle2_y(rectangle2_ys[2794]), .rectangle2_width(rectangle2_widths[2794]), .rectangle2_height(rectangle2_heights[2794]), .rectangle2_weight(rectangle2_weights[2794]), .rectangle3_x(rectangle3_xs[2794]), .rectangle3_y(rectangle3_ys[2794]), .rectangle3_width(rectangle3_widths[2794]), .rectangle3_height(rectangle3_heights[2794]), .rectangle3_weight(rectangle3_weights[2794]), .feature_threshold(feature_thresholds[2794]), .feature_above(feature_aboves[2794]), .feature_below(feature_belows[2794]), .scan_win_std_dev(scan_win_std_dev[2794]), .feature_accum(feature_accums[2794]));
  accum_calculator ac2795(.scan_win(scan_win2795), .rectangle1_x(rectangle1_xs[2795]), .rectangle1_y(rectangle1_ys[2795]), .rectangle1_width(rectangle1_widths[2795]), .rectangle1_height(rectangle1_heights[2795]), .rectangle1_weight(rectangle1_weights[2795]), .rectangle2_x(rectangle2_xs[2795]), .rectangle2_y(rectangle2_ys[2795]), .rectangle2_width(rectangle2_widths[2795]), .rectangle2_height(rectangle2_heights[2795]), .rectangle2_weight(rectangle2_weights[2795]), .rectangle3_x(rectangle3_xs[2795]), .rectangle3_y(rectangle3_ys[2795]), .rectangle3_width(rectangle3_widths[2795]), .rectangle3_height(rectangle3_heights[2795]), .rectangle3_weight(rectangle3_weights[2795]), .feature_threshold(feature_thresholds[2795]), .feature_above(feature_aboves[2795]), .feature_below(feature_belows[2795]), .scan_win_std_dev(scan_win_std_dev[2795]), .feature_accum(feature_accums[2795]));
  accum_calculator ac2796(.scan_win(scan_win2796), .rectangle1_x(rectangle1_xs[2796]), .rectangle1_y(rectangle1_ys[2796]), .rectangle1_width(rectangle1_widths[2796]), .rectangle1_height(rectangle1_heights[2796]), .rectangle1_weight(rectangle1_weights[2796]), .rectangle2_x(rectangle2_xs[2796]), .rectangle2_y(rectangle2_ys[2796]), .rectangle2_width(rectangle2_widths[2796]), .rectangle2_height(rectangle2_heights[2796]), .rectangle2_weight(rectangle2_weights[2796]), .rectangle3_x(rectangle3_xs[2796]), .rectangle3_y(rectangle3_ys[2796]), .rectangle3_width(rectangle3_widths[2796]), .rectangle3_height(rectangle3_heights[2796]), .rectangle3_weight(rectangle3_weights[2796]), .feature_threshold(feature_thresholds[2796]), .feature_above(feature_aboves[2796]), .feature_below(feature_belows[2796]), .scan_win_std_dev(scan_win_std_dev[2796]), .feature_accum(feature_accums[2796]));
  accum_calculator ac2797(.scan_win(scan_win2797), .rectangle1_x(rectangle1_xs[2797]), .rectangle1_y(rectangle1_ys[2797]), .rectangle1_width(rectangle1_widths[2797]), .rectangle1_height(rectangle1_heights[2797]), .rectangle1_weight(rectangle1_weights[2797]), .rectangle2_x(rectangle2_xs[2797]), .rectangle2_y(rectangle2_ys[2797]), .rectangle2_width(rectangle2_widths[2797]), .rectangle2_height(rectangle2_heights[2797]), .rectangle2_weight(rectangle2_weights[2797]), .rectangle3_x(rectangle3_xs[2797]), .rectangle3_y(rectangle3_ys[2797]), .rectangle3_width(rectangle3_widths[2797]), .rectangle3_height(rectangle3_heights[2797]), .rectangle3_weight(rectangle3_weights[2797]), .feature_threshold(feature_thresholds[2797]), .feature_above(feature_aboves[2797]), .feature_below(feature_belows[2797]), .scan_win_std_dev(scan_win_std_dev[2797]), .feature_accum(feature_accums[2797]));
  accum_calculator ac2798(.scan_win(scan_win2798), .rectangle1_x(rectangle1_xs[2798]), .rectangle1_y(rectangle1_ys[2798]), .rectangle1_width(rectangle1_widths[2798]), .rectangle1_height(rectangle1_heights[2798]), .rectangle1_weight(rectangle1_weights[2798]), .rectangle2_x(rectangle2_xs[2798]), .rectangle2_y(rectangle2_ys[2798]), .rectangle2_width(rectangle2_widths[2798]), .rectangle2_height(rectangle2_heights[2798]), .rectangle2_weight(rectangle2_weights[2798]), .rectangle3_x(rectangle3_xs[2798]), .rectangle3_y(rectangle3_ys[2798]), .rectangle3_width(rectangle3_widths[2798]), .rectangle3_height(rectangle3_heights[2798]), .rectangle3_weight(rectangle3_weights[2798]), .feature_threshold(feature_thresholds[2798]), .feature_above(feature_aboves[2798]), .feature_below(feature_belows[2798]), .scan_win_std_dev(scan_win_std_dev[2798]), .feature_accum(feature_accums[2798]));
  accum_calculator ac2799(.scan_win(scan_win2799), .rectangle1_x(rectangle1_xs[2799]), .rectangle1_y(rectangle1_ys[2799]), .rectangle1_width(rectangle1_widths[2799]), .rectangle1_height(rectangle1_heights[2799]), .rectangle1_weight(rectangle1_weights[2799]), .rectangle2_x(rectangle2_xs[2799]), .rectangle2_y(rectangle2_ys[2799]), .rectangle2_width(rectangle2_widths[2799]), .rectangle2_height(rectangle2_heights[2799]), .rectangle2_weight(rectangle2_weights[2799]), .rectangle3_x(rectangle3_xs[2799]), .rectangle3_y(rectangle3_ys[2799]), .rectangle3_width(rectangle3_widths[2799]), .rectangle3_height(rectangle3_heights[2799]), .rectangle3_weight(rectangle3_weights[2799]), .feature_threshold(feature_thresholds[2799]), .feature_above(feature_aboves[2799]), .feature_below(feature_belows[2799]), .scan_win_std_dev(scan_win_std_dev[2799]), .feature_accum(feature_accums[2799]));
  accum_calculator ac2800(.scan_win(scan_win2800), .rectangle1_x(rectangle1_xs[2800]), .rectangle1_y(rectangle1_ys[2800]), .rectangle1_width(rectangle1_widths[2800]), .rectangle1_height(rectangle1_heights[2800]), .rectangle1_weight(rectangle1_weights[2800]), .rectangle2_x(rectangle2_xs[2800]), .rectangle2_y(rectangle2_ys[2800]), .rectangle2_width(rectangle2_widths[2800]), .rectangle2_height(rectangle2_heights[2800]), .rectangle2_weight(rectangle2_weights[2800]), .rectangle3_x(rectangle3_xs[2800]), .rectangle3_y(rectangle3_ys[2800]), .rectangle3_width(rectangle3_widths[2800]), .rectangle3_height(rectangle3_heights[2800]), .rectangle3_weight(rectangle3_weights[2800]), .feature_threshold(feature_thresholds[2800]), .feature_above(feature_aboves[2800]), .feature_below(feature_belows[2800]), .scan_win_std_dev(scan_win_std_dev[2800]), .feature_accum(feature_accums[2800]));
  accum_calculator ac2801(.scan_win(scan_win2801), .rectangle1_x(rectangle1_xs[2801]), .rectangle1_y(rectangle1_ys[2801]), .rectangle1_width(rectangle1_widths[2801]), .rectangle1_height(rectangle1_heights[2801]), .rectangle1_weight(rectangle1_weights[2801]), .rectangle2_x(rectangle2_xs[2801]), .rectangle2_y(rectangle2_ys[2801]), .rectangle2_width(rectangle2_widths[2801]), .rectangle2_height(rectangle2_heights[2801]), .rectangle2_weight(rectangle2_weights[2801]), .rectangle3_x(rectangle3_xs[2801]), .rectangle3_y(rectangle3_ys[2801]), .rectangle3_width(rectangle3_widths[2801]), .rectangle3_height(rectangle3_heights[2801]), .rectangle3_weight(rectangle3_weights[2801]), .feature_threshold(feature_thresholds[2801]), .feature_above(feature_aboves[2801]), .feature_below(feature_belows[2801]), .scan_win_std_dev(scan_win_std_dev[2801]), .feature_accum(feature_accums[2801]));
  accum_calculator ac2802(.scan_win(scan_win2802), .rectangle1_x(rectangle1_xs[2802]), .rectangle1_y(rectangle1_ys[2802]), .rectangle1_width(rectangle1_widths[2802]), .rectangle1_height(rectangle1_heights[2802]), .rectangle1_weight(rectangle1_weights[2802]), .rectangle2_x(rectangle2_xs[2802]), .rectangle2_y(rectangle2_ys[2802]), .rectangle2_width(rectangle2_widths[2802]), .rectangle2_height(rectangle2_heights[2802]), .rectangle2_weight(rectangle2_weights[2802]), .rectangle3_x(rectangle3_xs[2802]), .rectangle3_y(rectangle3_ys[2802]), .rectangle3_width(rectangle3_widths[2802]), .rectangle3_height(rectangle3_heights[2802]), .rectangle3_weight(rectangle3_weights[2802]), .feature_threshold(feature_thresholds[2802]), .feature_above(feature_aboves[2802]), .feature_below(feature_belows[2802]), .scan_win_std_dev(scan_win_std_dev[2802]), .feature_accum(feature_accums[2802]));
  accum_calculator ac2803(.scan_win(scan_win2803), .rectangle1_x(rectangle1_xs[2803]), .rectangle1_y(rectangle1_ys[2803]), .rectangle1_width(rectangle1_widths[2803]), .rectangle1_height(rectangle1_heights[2803]), .rectangle1_weight(rectangle1_weights[2803]), .rectangle2_x(rectangle2_xs[2803]), .rectangle2_y(rectangle2_ys[2803]), .rectangle2_width(rectangle2_widths[2803]), .rectangle2_height(rectangle2_heights[2803]), .rectangle2_weight(rectangle2_weights[2803]), .rectangle3_x(rectangle3_xs[2803]), .rectangle3_y(rectangle3_ys[2803]), .rectangle3_width(rectangle3_widths[2803]), .rectangle3_height(rectangle3_heights[2803]), .rectangle3_weight(rectangle3_weights[2803]), .feature_threshold(feature_thresholds[2803]), .feature_above(feature_aboves[2803]), .feature_below(feature_belows[2803]), .scan_win_std_dev(scan_win_std_dev[2803]), .feature_accum(feature_accums[2803]));
  accum_calculator ac2804(.scan_win(scan_win2804), .rectangle1_x(rectangle1_xs[2804]), .rectangle1_y(rectangle1_ys[2804]), .rectangle1_width(rectangle1_widths[2804]), .rectangle1_height(rectangle1_heights[2804]), .rectangle1_weight(rectangle1_weights[2804]), .rectangle2_x(rectangle2_xs[2804]), .rectangle2_y(rectangle2_ys[2804]), .rectangle2_width(rectangle2_widths[2804]), .rectangle2_height(rectangle2_heights[2804]), .rectangle2_weight(rectangle2_weights[2804]), .rectangle3_x(rectangle3_xs[2804]), .rectangle3_y(rectangle3_ys[2804]), .rectangle3_width(rectangle3_widths[2804]), .rectangle3_height(rectangle3_heights[2804]), .rectangle3_weight(rectangle3_weights[2804]), .feature_threshold(feature_thresholds[2804]), .feature_above(feature_aboves[2804]), .feature_below(feature_belows[2804]), .scan_win_std_dev(scan_win_std_dev[2804]), .feature_accum(feature_accums[2804]));
  accum_calculator ac2805(.scan_win(scan_win2805), .rectangle1_x(rectangle1_xs[2805]), .rectangle1_y(rectangle1_ys[2805]), .rectangle1_width(rectangle1_widths[2805]), .rectangle1_height(rectangle1_heights[2805]), .rectangle1_weight(rectangle1_weights[2805]), .rectangle2_x(rectangle2_xs[2805]), .rectangle2_y(rectangle2_ys[2805]), .rectangle2_width(rectangle2_widths[2805]), .rectangle2_height(rectangle2_heights[2805]), .rectangle2_weight(rectangle2_weights[2805]), .rectangle3_x(rectangle3_xs[2805]), .rectangle3_y(rectangle3_ys[2805]), .rectangle3_width(rectangle3_widths[2805]), .rectangle3_height(rectangle3_heights[2805]), .rectangle3_weight(rectangle3_weights[2805]), .feature_threshold(feature_thresholds[2805]), .feature_above(feature_aboves[2805]), .feature_below(feature_belows[2805]), .scan_win_std_dev(scan_win_std_dev[2805]), .feature_accum(feature_accums[2805]));
  accum_calculator ac2806(.scan_win(scan_win2806), .rectangle1_x(rectangle1_xs[2806]), .rectangle1_y(rectangle1_ys[2806]), .rectangle1_width(rectangle1_widths[2806]), .rectangle1_height(rectangle1_heights[2806]), .rectangle1_weight(rectangle1_weights[2806]), .rectangle2_x(rectangle2_xs[2806]), .rectangle2_y(rectangle2_ys[2806]), .rectangle2_width(rectangle2_widths[2806]), .rectangle2_height(rectangle2_heights[2806]), .rectangle2_weight(rectangle2_weights[2806]), .rectangle3_x(rectangle3_xs[2806]), .rectangle3_y(rectangle3_ys[2806]), .rectangle3_width(rectangle3_widths[2806]), .rectangle3_height(rectangle3_heights[2806]), .rectangle3_weight(rectangle3_weights[2806]), .feature_threshold(feature_thresholds[2806]), .feature_above(feature_aboves[2806]), .feature_below(feature_belows[2806]), .scan_win_std_dev(scan_win_std_dev[2806]), .feature_accum(feature_accums[2806]));
  accum_calculator ac2807(.scan_win(scan_win2807), .rectangle1_x(rectangle1_xs[2807]), .rectangle1_y(rectangle1_ys[2807]), .rectangle1_width(rectangle1_widths[2807]), .rectangle1_height(rectangle1_heights[2807]), .rectangle1_weight(rectangle1_weights[2807]), .rectangle2_x(rectangle2_xs[2807]), .rectangle2_y(rectangle2_ys[2807]), .rectangle2_width(rectangle2_widths[2807]), .rectangle2_height(rectangle2_heights[2807]), .rectangle2_weight(rectangle2_weights[2807]), .rectangle3_x(rectangle3_xs[2807]), .rectangle3_y(rectangle3_ys[2807]), .rectangle3_width(rectangle3_widths[2807]), .rectangle3_height(rectangle3_heights[2807]), .rectangle3_weight(rectangle3_weights[2807]), .feature_threshold(feature_thresholds[2807]), .feature_above(feature_aboves[2807]), .feature_below(feature_belows[2807]), .scan_win_std_dev(scan_win_std_dev[2807]), .feature_accum(feature_accums[2807]));
  accum_calculator ac2808(.scan_win(scan_win2808), .rectangle1_x(rectangle1_xs[2808]), .rectangle1_y(rectangle1_ys[2808]), .rectangle1_width(rectangle1_widths[2808]), .rectangle1_height(rectangle1_heights[2808]), .rectangle1_weight(rectangle1_weights[2808]), .rectangle2_x(rectangle2_xs[2808]), .rectangle2_y(rectangle2_ys[2808]), .rectangle2_width(rectangle2_widths[2808]), .rectangle2_height(rectangle2_heights[2808]), .rectangle2_weight(rectangle2_weights[2808]), .rectangle3_x(rectangle3_xs[2808]), .rectangle3_y(rectangle3_ys[2808]), .rectangle3_width(rectangle3_widths[2808]), .rectangle3_height(rectangle3_heights[2808]), .rectangle3_weight(rectangle3_weights[2808]), .feature_threshold(feature_thresholds[2808]), .feature_above(feature_aboves[2808]), .feature_below(feature_belows[2808]), .scan_win_std_dev(scan_win_std_dev[2808]), .feature_accum(feature_accums[2808]));
  accum_calculator ac2809(.scan_win(scan_win2809), .rectangle1_x(rectangle1_xs[2809]), .rectangle1_y(rectangle1_ys[2809]), .rectangle1_width(rectangle1_widths[2809]), .rectangle1_height(rectangle1_heights[2809]), .rectangle1_weight(rectangle1_weights[2809]), .rectangle2_x(rectangle2_xs[2809]), .rectangle2_y(rectangle2_ys[2809]), .rectangle2_width(rectangle2_widths[2809]), .rectangle2_height(rectangle2_heights[2809]), .rectangle2_weight(rectangle2_weights[2809]), .rectangle3_x(rectangle3_xs[2809]), .rectangle3_y(rectangle3_ys[2809]), .rectangle3_width(rectangle3_widths[2809]), .rectangle3_height(rectangle3_heights[2809]), .rectangle3_weight(rectangle3_weights[2809]), .feature_threshold(feature_thresholds[2809]), .feature_above(feature_aboves[2809]), .feature_below(feature_belows[2809]), .scan_win_std_dev(scan_win_std_dev[2809]), .feature_accum(feature_accums[2809]));
  accum_calculator ac2810(.scan_win(scan_win2810), .rectangle1_x(rectangle1_xs[2810]), .rectangle1_y(rectangle1_ys[2810]), .rectangle1_width(rectangle1_widths[2810]), .rectangle1_height(rectangle1_heights[2810]), .rectangle1_weight(rectangle1_weights[2810]), .rectangle2_x(rectangle2_xs[2810]), .rectangle2_y(rectangle2_ys[2810]), .rectangle2_width(rectangle2_widths[2810]), .rectangle2_height(rectangle2_heights[2810]), .rectangle2_weight(rectangle2_weights[2810]), .rectangle3_x(rectangle3_xs[2810]), .rectangle3_y(rectangle3_ys[2810]), .rectangle3_width(rectangle3_widths[2810]), .rectangle3_height(rectangle3_heights[2810]), .rectangle3_weight(rectangle3_weights[2810]), .feature_threshold(feature_thresholds[2810]), .feature_above(feature_aboves[2810]), .feature_below(feature_belows[2810]), .scan_win_std_dev(scan_win_std_dev[2810]), .feature_accum(feature_accums[2810]));
  accum_calculator ac2811(.scan_win(scan_win2811), .rectangle1_x(rectangle1_xs[2811]), .rectangle1_y(rectangle1_ys[2811]), .rectangle1_width(rectangle1_widths[2811]), .rectangle1_height(rectangle1_heights[2811]), .rectangle1_weight(rectangle1_weights[2811]), .rectangle2_x(rectangle2_xs[2811]), .rectangle2_y(rectangle2_ys[2811]), .rectangle2_width(rectangle2_widths[2811]), .rectangle2_height(rectangle2_heights[2811]), .rectangle2_weight(rectangle2_weights[2811]), .rectangle3_x(rectangle3_xs[2811]), .rectangle3_y(rectangle3_ys[2811]), .rectangle3_width(rectangle3_widths[2811]), .rectangle3_height(rectangle3_heights[2811]), .rectangle3_weight(rectangle3_weights[2811]), .feature_threshold(feature_thresholds[2811]), .feature_above(feature_aboves[2811]), .feature_below(feature_belows[2811]), .scan_win_std_dev(scan_win_std_dev[2811]), .feature_accum(feature_accums[2811]));
  accum_calculator ac2812(.scan_win(scan_win2812), .rectangle1_x(rectangle1_xs[2812]), .rectangle1_y(rectangle1_ys[2812]), .rectangle1_width(rectangle1_widths[2812]), .rectangle1_height(rectangle1_heights[2812]), .rectangle1_weight(rectangle1_weights[2812]), .rectangle2_x(rectangle2_xs[2812]), .rectangle2_y(rectangle2_ys[2812]), .rectangle2_width(rectangle2_widths[2812]), .rectangle2_height(rectangle2_heights[2812]), .rectangle2_weight(rectangle2_weights[2812]), .rectangle3_x(rectangle3_xs[2812]), .rectangle3_y(rectangle3_ys[2812]), .rectangle3_width(rectangle3_widths[2812]), .rectangle3_height(rectangle3_heights[2812]), .rectangle3_weight(rectangle3_weights[2812]), .feature_threshold(feature_thresholds[2812]), .feature_above(feature_aboves[2812]), .feature_below(feature_belows[2812]), .scan_win_std_dev(scan_win_std_dev[2812]), .feature_accum(feature_accums[2812]));
  accum_calculator ac2813(.scan_win(scan_win2813), .rectangle1_x(rectangle1_xs[2813]), .rectangle1_y(rectangle1_ys[2813]), .rectangle1_width(rectangle1_widths[2813]), .rectangle1_height(rectangle1_heights[2813]), .rectangle1_weight(rectangle1_weights[2813]), .rectangle2_x(rectangle2_xs[2813]), .rectangle2_y(rectangle2_ys[2813]), .rectangle2_width(rectangle2_widths[2813]), .rectangle2_height(rectangle2_heights[2813]), .rectangle2_weight(rectangle2_weights[2813]), .rectangle3_x(rectangle3_xs[2813]), .rectangle3_y(rectangle3_ys[2813]), .rectangle3_width(rectangle3_widths[2813]), .rectangle3_height(rectangle3_heights[2813]), .rectangle3_weight(rectangle3_weights[2813]), .feature_threshold(feature_thresholds[2813]), .feature_above(feature_aboves[2813]), .feature_below(feature_belows[2813]), .scan_win_std_dev(scan_win_std_dev[2813]), .feature_accum(feature_accums[2813]));
  accum_calculator ac2814(.scan_win(scan_win2814), .rectangle1_x(rectangle1_xs[2814]), .rectangle1_y(rectangle1_ys[2814]), .rectangle1_width(rectangle1_widths[2814]), .rectangle1_height(rectangle1_heights[2814]), .rectangle1_weight(rectangle1_weights[2814]), .rectangle2_x(rectangle2_xs[2814]), .rectangle2_y(rectangle2_ys[2814]), .rectangle2_width(rectangle2_widths[2814]), .rectangle2_height(rectangle2_heights[2814]), .rectangle2_weight(rectangle2_weights[2814]), .rectangle3_x(rectangle3_xs[2814]), .rectangle3_y(rectangle3_ys[2814]), .rectangle3_width(rectangle3_widths[2814]), .rectangle3_height(rectangle3_heights[2814]), .rectangle3_weight(rectangle3_weights[2814]), .feature_threshold(feature_thresholds[2814]), .feature_above(feature_aboves[2814]), .feature_below(feature_belows[2814]), .scan_win_std_dev(scan_win_std_dev[2814]), .feature_accum(feature_accums[2814]));
  accum_calculator ac2815(.scan_win(scan_win2815), .rectangle1_x(rectangle1_xs[2815]), .rectangle1_y(rectangle1_ys[2815]), .rectangle1_width(rectangle1_widths[2815]), .rectangle1_height(rectangle1_heights[2815]), .rectangle1_weight(rectangle1_weights[2815]), .rectangle2_x(rectangle2_xs[2815]), .rectangle2_y(rectangle2_ys[2815]), .rectangle2_width(rectangle2_widths[2815]), .rectangle2_height(rectangle2_heights[2815]), .rectangle2_weight(rectangle2_weights[2815]), .rectangle3_x(rectangle3_xs[2815]), .rectangle3_y(rectangle3_ys[2815]), .rectangle3_width(rectangle3_widths[2815]), .rectangle3_height(rectangle3_heights[2815]), .rectangle3_weight(rectangle3_weights[2815]), .feature_threshold(feature_thresholds[2815]), .feature_above(feature_aboves[2815]), .feature_below(feature_belows[2815]), .scan_win_std_dev(scan_win_std_dev[2815]), .feature_accum(feature_accums[2815]));
  accum_calculator ac2816(.scan_win(scan_win2816), .rectangle1_x(rectangle1_xs[2816]), .rectangle1_y(rectangle1_ys[2816]), .rectangle1_width(rectangle1_widths[2816]), .rectangle1_height(rectangle1_heights[2816]), .rectangle1_weight(rectangle1_weights[2816]), .rectangle2_x(rectangle2_xs[2816]), .rectangle2_y(rectangle2_ys[2816]), .rectangle2_width(rectangle2_widths[2816]), .rectangle2_height(rectangle2_heights[2816]), .rectangle2_weight(rectangle2_weights[2816]), .rectangle3_x(rectangle3_xs[2816]), .rectangle3_y(rectangle3_ys[2816]), .rectangle3_width(rectangle3_widths[2816]), .rectangle3_height(rectangle3_heights[2816]), .rectangle3_weight(rectangle3_weights[2816]), .feature_threshold(feature_thresholds[2816]), .feature_above(feature_aboves[2816]), .feature_below(feature_belows[2816]), .scan_win_std_dev(scan_win_std_dev[2816]), .feature_accum(feature_accums[2816]));
  accum_calculator ac2817(.scan_win(scan_win2817), .rectangle1_x(rectangle1_xs[2817]), .rectangle1_y(rectangle1_ys[2817]), .rectangle1_width(rectangle1_widths[2817]), .rectangle1_height(rectangle1_heights[2817]), .rectangle1_weight(rectangle1_weights[2817]), .rectangle2_x(rectangle2_xs[2817]), .rectangle2_y(rectangle2_ys[2817]), .rectangle2_width(rectangle2_widths[2817]), .rectangle2_height(rectangle2_heights[2817]), .rectangle2_weight(rectangle2_weights[2817]), .rectangle3_x(rectangle3_xs[2817]), .rectangle3_y(rectangle3_ys[2817]), .rectangle3_width(rectangle3_widths[2817]), .rectangle3_height(rectangle3_heights[2817]), .rectangle3_weight(rectangle3_weights[2817]), .feature_threshold(feature_thresholds[2817]), .feature_above(feature_aboves[2817]), .feature_below(feature_belows[2817]), .scan_win_std_dev(scan_win_std_dev[2817]), .feature_accum(feature_accums[2817]));
  accum_calculator ac2818(.scan_win(scan_win2818), .rectangle1_x(rectangle1_xs[2818]), .rectangle1_y(rectangle1_ys[2818]), .rectangle1_width(rectangle1_widths[2818]), .rectangle1_height(rectangle1_heights[2818]), .rectangle1_weight(rectangle1_weights[2818]), .rectangle2_x(rectangle2_xs[2818]), .rectangle2_y(rectangle2_ys[2818]), .rectangle2_width(rectangle2_widths[2818]), .rectangle2_height(rectangle2_heights[2818]), .rectangle2_weight(rectangle2_weights[2818]), .rectangle3_x(rectangle3_xs[2818]), .rectangle3_y(rectangle3_ys[2818]), .rectangle3_width(rectangle3_widths[2818]), .rectangle3_height(rectangle3_heights[2818]), .rectangle3_weight(rectangle3_weights[2818]), .feature_threshold(feature_thresholds[2818]), .feature_above(feature_aboves[2818]), .feature_below(feature_belows[2818]), .scan_win_std_dev(scan_win_std_dev[2818]), .feature_accum(feature_accums[2818]));
  accum_calculator ac2819(.scan_win(scan_win2819), .rectangle1_x(rectangle1_xs[2819]), .rectangle1_y(rectangle1_ys[2819]), .rectangle1_width(rectangle1_widths[2819]), .rectangle1_height(rectangle1_heights[2819]), .rectangle1_weight(rectangle1_weights[2819]), .rectangle2_x(rectangle2_xs[2819]), .rectangle2_y(rectangle2_ys[2819]), .rectangle2_width(rectangle2_widths[2819]), .rectangle2_height(rectangle2_heights[2819]), .rectangle2_weight(rectangle2_weights[2819]), .rectangle3_x(rectangle3_xs[2819]), .rectangle3_y(rectangle3_ys[2819]), .rectangle3_width(rectangle3_widths[2819]), .rectangle3_height(rectangle3_heights[2819]), .rectangle3_weight(rectangle3_weights[2819]), .feature_threshold(feature_thresholds[2819]), .feature_above(feature_aboves[2819]), .feature_below(feature_belows[2819]), .scan_win_std_dev(scan_win_std_dev[2819]), .feature_accum(feature_accums[2819]));
  accum_calculator ac2820(.scan_win(scan_win2820), .rectangle1_x(rectangle1_xs[2820]), .rectangle1_y(rectangle1_ys[2820]), .rectangle1_width(rectangle1_widths[2820]), .rectangle1_height(rectangle1_heights[2820]), .rectangle1_weight(rectangle1_weights[2820]), .rectangle2_x(rectangle2_xs[2820]), .rectangle2_y(rectangle2_ys[2820]), .rectangle2_width(rectangle2_widths[2820]), .rectangle2_height(rectangle2_heights[2820]), .rectangle2_weight(rectangle2_weights[2820]), .rectangle3_x(rectangle3_xs[2820]), .rectangle3_y(rectangle3_ys[2820]), .rectangle3_width(rectangle3_widths[2820]), .rectangle3_height(rectangle3_heights[2820]), .rectangle3_weight(rectangle3_weights[2820]), .feature_threshold(feature_thresholds[2820]), .feature_above(feature_aboves[2820]), .feature_below(feature_belows[2820]), .scan_win_std_dev(scan_win_std_dev[2820]), .feature_accum(feature_accums[2820]));
  accum_calculator ac2821(.scan_win(scan_win2821), .rectangle1_x(rectangle1_xs[2821]), .rectangle1_y(rectangle1_ys[2821]), .rectangle1_width(rectangle1_widths[2821]), .rectangle1_height(rectangle1_heights[2821]), .rectangle1_weight(rectangle1_weights[2821]), .rectangle2_x(rectangle2_xs[2821]), .rectangle2_y(rectangle2_ys[2821]), .rectangle2_width(rectangle2_widths[2821]), .rectangle2_height(rectangle2_heights[2821]), .rectangle2_weight(rectangle2_weights[2821]), .rectangle3_x(rectangle3_xs[2821]), .rectangle3_y(rectangle3_ys[2821]), .rectangle3_width(rectangle3_widths[2821]), .rectangle3_height(rectangle3_heights[2821]), .rectangle3_weight(rectangle3_weights[2821]), .feature_threshold(feature_thresholds[2821]), .feature_above(feature_aboves[2821]), .feature_below(feature_belows[2821]), .scan_win_std_dev(scan_win_std_dev[2821]), .feature_accum(feature_accums[2821]));
  accum_calculator ac2822(.scan_win(scan_win2822), .rectangle1_x(rectangle1_xs[2822]), .rectangle1_y(rectangle1_ys[2822]), .rectangle1_width(rectangle1_widths[2822]), .rectangle1_height(rectangle1_heights[2822]), .rectangle1_weight(rectangle1_weights[2822]), .rectangle2_x(rectangle2_xs[2822]), .rectangle2_y(rectangle2_ys[2822]), .rectangle2_width(rectangle2_widths[2822]), .rectangle2_height(rectangle2_heights[2822]), .rectangle2_weight(rectangle2_weights[2822]), .rectangle3_x(rectangle3_xs[2822]), .rectangle3_y(rectangle3_ys[2822]), .rectangle3_width(rectangle3_widths[2822]), .rectangle3_height(rectangle3_heights[2822]), .rectangle3_weight(rectangle3_weights[2822]), .feature_threshold(feature_thresholds[2822]), .feature_above(feature_aboves[2822]), .feature_below(feature_belows[2822]), .scan_win_std_dev(scan_win_std_dev[2822]), .feature_accum(feature_accums[2822]));
  accum_calculator ac2823(.scan_win(scan_win2823), .rectangle1_x(rectangle1_xs[2823]), .rectangle1_y(rectangle1_ys[2823]), .rectangle1_width(rectangle1_widths[2823]), .rectangle1_height(rectangle1_heights[2823]), .rectangle1_weight(rectangle1_weights[2823]), .rectangle2_x(rectangle2_xs[2823]), .rectangle2_y(rectangle2_ys[2823]), .rectangle2_width(rectangle2_widths[2823]), .rectangle2_height(rectangle2_heights[2823]), .rectangle2_weight(rectangle2_weights[2823]), .rectangle3_x(rectangle3_xs[2823]), .rectangle3_y(rectangle3_ys[2823]), .rectangle3_width(rectangle3_widths[2823]), .rectangle3_height(rectangle3_heights[2823]), .rectangle3_weight(rectangle3_weights[2823]), .feature_threshold(feature_thresholds[2823]), .feature_above(feature_aboves[2823]), .feature_below(feature_belows[2823]), .scan_win_std_dev(scan_win_std_dev[2823]), .feature_accum(feature_accums[2823]));
  accum_calculator ac2824(.scan_win(scan_win2824), .rectangle1_x(rectangle1_xs[2824]), .rectangle1_y(rectangle1_ys[2824]), .rectangle1_width(rectangle1_widths[2824]), .rectangle1_height(rectangle1_heights[2824]), .rectangle1_weight(rectangle1_weights[2824]), .rectangle2_x(rectangle2_xs[2824]), .rectangle2_y(rectangle2_ys[2824]), .rectangle2_width(rectangle2_widths[2824]), .rectangle2_height(rectangle2_heights[2824]), .rectangle2_weight(rectangle2_weights[2824]), .rectangle3_x(rectangle3_xs[2824]), .rectangle3_y(rectangle3_ys[2824]), .rectangle3_width(rectangle3_widths[2824]), .rectangle3_height(rectangle3_heights[2824]), .rectangle3_weight(rectangle3_weights[2824]), .feature_threshold(feature_thresholds[2824]), .feature_above(feature_aboves[2824]), .feature_below(feature_belows[2824]), .scan_win_std_dev(scan_win_std_dev[2824]), .feature_accum(feature_accums[2824]));
  accum_calculator ac2825(.scan_win(scan_win2825), .rectangle1_x(rectangle1_xs[2825]), .rectangle1_y(rectangle1_ys[2825]), .rectangle1_width(rectangle1_widths[2825]), .rectangle1_height(rectangle1_heights[2825]), .rectangle1_weight(rectangle1_weights[2825]), .rectangle2_x(rectangle2_xs[2825]), .rectangle2_y(rectangle2_ys[2825]), .rectangle2_width(rectangle2_widths[2825]), .rectangle2_height(rectangle2_heights[2825]), .rectangle2_weight(rectangle2_weights[2825]), .rectangle3_x(rectangle3_xs[2825]), .rectangle3_y(rectangle3_ys[2825]), .rectangle3_width(rectangle3_widths[2825]), .rectangle3_height(rectangle3_heights[2825]), .rectangle3_weight(rectangle3_weights[2825]), .feature_threshold(feature_thresholds[2825]), .feature_above(feature_aboves[2825]), .feature_below(feature_belows[2825]), .scan_win_std_dev(scan_win_std_dev[2825]), .feature_accum(feature_accums[2825]));
  accum_calculator ac2826(.scan_win(scan_win2826), .rectangle1_x(rectangle1_xs[2826]), .rectangle1_y(rectangle1_ys[2826]), .rectangle1_width(rectangle1_widths[2826]), .rectangle1_height(rectangle1_heights[2826]), .rectangle1_weight(rectangle1_weights[2826]), .rectangle2_x(rectangle2_xs[2826]), .rectangle2_y(rectangle2_ys[2826]), .rectangle2_width(rectangle2_widths[2826]), .rectangle2_height(rectangle2_heights[2826]), .rectangle2_weight(rectangle2_weights[2826]), .rectangle3_x(rectangle3_xs[2826]), .rectangle3_y(rectangle3_ys[2826]), .rectangle3_width(rectangle3_widths[2826]), .rectangle3_height(rectangle3_heights[2826]), .rectangle3_weight(rectangle3_weights[2826]), .feature_threshold(feature_thresholds[2826]), .feature_above(feature_aboves[2826]), .feature_below(feature_belows[2826]), .scan_win_std_dev(scan_win_std_dev[2826]), .feature_accum(feature_accums[2826]));
  accum_calculator ac2827(.scan_win(scan_win2827), .rectangle1_x(rectangle1_xs[2827]), .rectangle1_y(rectangle1_ys[2827]), .rectangle1_width(rectangle1_widths[2827]), .rectangle1_height(rectangle1_heights[2827]), .rectangle1_weight(rectangle1_weights[2827]), .rectangle2_x(rectangle2_xs[2827]), .rectangle2_y(rectangle2_ys[2827]), .rectangle2_width(rectangle2_widths[2827]), .rectangle2_height(rectangle2_heights[2827]), .rectangle2_weight(rectangle2_weights[2827]), .rectangle3_x(rectangle3_xs[2827]), .rectangle3_y(rectangle3_ys[2827]), .rectangle3_width(rectangle3_widths[2827]), .rectangle3_height(rectangle3_heights[2827]), .rectangle3_weight(rectangle3_weights[2827]), .feature_threshold(feature_thresholds[2827]), .feature_above(feature_aboves[2827]), .feature_below(feature_belows[2827]), .scan_win_std_dev(scan_win_std_dev[2827]), .feature_accum(feature_accums[2827]));
  accum_calculator ac2828(.scan_win(scan_win2828), .rectangle1_x(rectangle1_xs[2828]), .rectangle1_y(rectangle1_ys[2828]), .rectangle1_width(rectangle1_widths[2828]), .rectangle1_height(rectangle1_heights[2828]), .rectangle1_weight(rectangle1_weights[2828]), .rectangle2_x(rectangle2_xs[2828]), .rectangle2_y(rectangle2_ys[2828]), .rectangle2_width(rectangle2_widths[2828]), .rectangle2_height(rectangle2_heights[2828]), .rectangle2_weight(rectangle2_weights[2828]), .rectangle3_x(rectangle3_xs[2828]), .rectangle3_y(rectangle3_ys[2828]), .rectangle3_width(rectangle3_widths[2828]), .rectangle3_height(rectangle3_heights[2828]), .rectangle3_weight(rectangle3_weights[2828]), .feature_threshold(feature_thresholds[2828]), .feature_above(feature_aboves[2828]), .feature_below(feature_belows[2828]), .scan_win_std_dev(scan_win_std_dev[2828]), .feature_accum(feature_accums[2828]));
  accum_calculator ac2829(.scan_win(scan_win2829), .rectangle1_x(rectangle1_xs[2829]), .rectangle1_y(rectangle1_ys[2829]), .rectangle1_width(rectangle1_widths[2829]), .rectangle1_height(rectangle1_heights[2829]), .rectangle1_weight(rectangle1_weights[2829]), .rectangle2_x(rectangle2_xs[2829]), .rectangle2_y(rectangle2_ys[2829]), .rectangle2_width(rectangle2_widths[2829]), .rectangle2_height(rectangle2_heights[2829]), .rectangle2_weight(rectangle2_weights[2829]), .rectangle3_x(rectangle3_xs[2829]), .rectangle3_y(rectangle3_ys[2829]), .rectangle3_width(rectangle3_widths[2829]), .rectangle3_height(rectangle3_heights[2829]), .rectangle3_weight(rectangle3_weights[2829]), .feature_threshold(feature_thresholds[2829]), .feature_above(feature_aboves[2829]), .feature_below(feature_belows[2829]), .scan_win_std_dev(scan_win_std_dev[2829]), .feature_accum(feature_accums[2829]));
  accum_calculator ac2830(.scan_win(scan_win2830), .rectangle1_x(rectangle1_xs[2830]), .rectangle1_y(rectangle1_ys[2830]), .rectangle1_width(rectangle1_widths[2830]), .rectangle1_height(rectangle1_heights[2830]), .rectangle1_weight(rectangle1_weights[2830]), .rectangle2_x(rectangle2_xs[2830]), .rectangle2_y(rectangle2_ys[2830]), .rectangle2_width(rectangle2_widths[2830]), .rectangle2_height(rectangle2_heights[2830]), .rectangle2_weight(rectangle2_weights[2830]), .rectangle3_x(rectangle3_xs[2830]), .rectangle3_y(rectangle3_ys[2830]), .rectangle3_width(rectangle3_widths[2830]), .rectangle3_height(rectangle3_heights[2830]), .rectangle3_weight(rectangle3_weights[2830]), .feature_threshold(feature_thresholds[2830]), .feature_above(feature_aboves[2830]), .feature_below(feature_belows[2830]), .scan_win_std_dev(scan_win_std_dev[2830]), .feature_accum(feature_accums[2830]));
  accum_calculator ac2831(.scan_win(scan_win2831), .rectangle1_x(rectangle1_xs[2831]), .rectangle1_y(rectangle1_ys[2831]), .rectangle1_width(rectangle1_widths[2831]), .rectangle1_height(rectangle1_heights[2831]), .rectangle1_weight(rectangle1_weights[2831]), .rectangle2_x(rectangle2_xs[2831]), .rectangle2_y(rectangle2_ys[2831]), .rectangle2_width(rectangle2_widths[2831]), .rectangle2_height(rectangle2_heights[2831]), .rectangle2_weight(rectangle2_weights[2831]), .rectangle3_x(rectangle3_xs[2831]), .rectangle3_y(rectangle3_ys[2831]), .rectangle3_width(rectangle3_widths[2831]), .rectangle3_height(rectangle3_heights[2831]), .rectangle3_weight(rectangle3_weights[2831]), .feature_threshold(feature_thresholds[2831]), .feature_above(feature_aboves[2831]), .feature_below(feature_belows[2831]), .scan_win_std_dev(scan_win_std_dev[2831]), .feature_accum(feature_accums[2831]));
  accum_calculator ac2832(.scan_win(scan_win2832), .rectangle1_x(rectangle1_xs[2832]), .rectangle1_y(rectangle1_ys[2832]), .rectangle1_width(rectangle1_widths[2832]), .rectangle1_height(rectangle1_heights[2832]), .rectangle1_weight(rectangle1_weights[2832]), .rectangle2_x(rectangle2_xs[2832]), .rectangle2_y(rectangle2_ys[2832]), .rectangle2_width(rectangle2_widths[2832]), .rectangle2_height(rectangle2_heights[2832]), .rectangle2_weight(rectangle2_weights[2832]), .rectangle3_x(rectangle3_xs[2832]), .rectangle3_y(rectangle3_ys[2832]), .rectangle3_width(rectangle3_widths[2832]), .rectangle3_height(rectangle3_heights[2832]), .rectangle3_weight(rectangle3_weights[2832]), .feature_threshold(feature_thresholds[2832]), .feature_above(feature_aboves[2832]), .feature_below(feature_belows[2832]), .scan_win_std_dev(scan_win_std_dev[2832]), .feature_accum(feature_accums[2832]));
  accum_calculator ac2833(.scan_win(scan_win2833), .rectangle1_x(rectangle1_xs[2833]), .rectangle1_y(rectangle1_ys[2833]), .rectangle1_width(rectangle1_widths[2833]), .rectangle1_height(rectangle1_heights[2833]), .rectangle1_weight(rectangle1_weights[2833]), .rectangle2_x(rectangle2_xs[2833]), .rectangle2_y(rectangle2_ys[2833]), .rectangle2_width(rectangle2_widths[2833]), .rectangle2_height(rectangle2_heights[2833]), .rectangle2_weight(rectangle2_weights[2833]), .rectangle3_x(rectangle3_xs[2833]), .rectangle3_y(rectangle3_ys[2833]), .rectangle3_width(rectangle3_widths[2833]), .rectangle3_height(rectangle3_heights[2833]), .rectangle3_weight(rectangle3_weights[2833]), .feature_threshold(feature_thresholds[2833]), .feature_above(feature_aboves[2833]), .feature_below(feature_belows[2833]), .scan_win_std_dev(scan_win_std_dev[2833]), .feature_accum(feature_accums[2833]));
  accum_calculator ac2834(.scan_win(scan_win2834), .rectangle1_x(rectangle1_xs[2834]), .rectangle1_y(rectangle1_ys[2834]), .rectangle1_width(rectangle1_widths[2834]), .rectangle1_height(rectangle1_heights[2834]), .rectangle1_weight(rectangle1_weights[2834]), .rectangle2_x(rectangle2_xs[2834]), .rectangle2_y(rectangle2_ys[2834]), .rectangle2_width(rectangle2_widths[2834]), .rectangle2_height(rectangle2_heights[2834]), .rectangle2_weight(rectangle2_weights[2834]), .rectangle3_x(rectangle3_xs[2834]), .rectangle3_y(rectangle3_ys[2834]), .rectangle3_width(rectangle3_widths[2834]), .rectangle3_height(rectangle3_heights[2834]), .rectangle3_weight(rectangle3_weights[2834]), .feature_threshold(feature_thresholds[2834]), .feature_above(feature_aboves[2834]), .feature_below(feature_belows[2834]), .scan_win_std_dev(scan_win_std_dev[2834]), .feature_accum(feature_accums[2834]));
  accum_calculator ac2835(.scan_win(scan_win2835), .rectangle1_x(rectangle1_xs[2835]), .rectangle1_y(rectangle1_ys[2835]), .rectangle1_width(rectangle1_widths[2835]), .rectangle1_height(rectangle1_heights[2835]), .rectangle1_weight(rectangle1_weights[2835]), .rectangle2_x(rectangle2_xs[2835]), .rectangle2_y(rectangle2_ys[2835]), .rectangle2_width(rectangle2_widths[2835]), .rectangle2_height(rectangle2_heights[2835]), .rectangle2_weight(rectangle2_weights[2835]), .rectangle3_x(rectangle3_xs[2835]), .rectangle3_y(rectangle3_ys[2835]), .rectangle3_width(rectangle3_widths[2835]), .rectangle3_height(rectangle3_heights[2835]), .rectangle3_weight(rectangle3_weights[2835]), .feature_threshold(feature_thresholds[2835]), .feature_above(feature_aboves[2835]), .feature_below(feature_belows[2835]), .scan_win_std_dev(scan_win_std_dev[2835]), .feature_accum(feature_accums[2835]));
  accum_calculator ac2836(.scan_win(scan_win2836), .rectangle1_x(rectangle1_xs[2836]), .rectangle1_y(rectangle1_ys[2836]), .rectangle1_width(rectangle1_widths[2836]), .rectangle1_height(rectangle1_heights[2836]), .rectangle1_weight(rectangle1_weights[2836]), .rectangle2_x(rectangle2_xs[2836]), .rectangle2_y(rectangle2_ys[2836]), .rectangle2_width(rectangle2_widths[2836]), .rectangle2_height(rectangle2_heights[2836]), .rectangle2_weight(rectangle2_weights[2836]), .rectangle3_x(rectangle3_xs[2836]), .rectangle3_y(rectangle3_ys[2836]), .rectangle3_width(rectangle3_widths[2836]), .rectangle3_height(rectangle3_heights[2836]), .rectangle3_weight(rectangle3_weights[2836]), .feature_threshold(feature_thresholds[2836]), .feature_above(feature_aboves[2836]), .feature_below(feature_belows[2836]), .scan_win_std_dev(scan_win_std_dev[2836]), .feature_accum(feature_accums[2836]));
  accum_calculator ac2837(.scan_win(scan_win2837), .rectangle1_x(rectangle1_xs[2837]), .rectangle1_y(rectangle1_ys[2837]), .rectangle1_width(rectangle1_widths[2837]), .rectangle1_height(rectangle1_heights[2837]), .rectangle1_weight(rectangle1_weights[2837]), .rectangle2_x(rectangle2_xs[2837]), .rectangle2_y(rectangle2_ys[2837]), .rectangle2_width(rectangle2_widths[2837]), .rectangle2_height(rectangle2_heights[2837]), .rectangle2_weight(rectangle2_weights[2837]), .rectangle3_x(rectangle3_xs[2837]), .rectangle3_y(rectangle3_ys[2837]), .rectangle3_width(rectangle3_widths[2837]), .rectangle3_height(rectangle3_heights[2837]), .rectangle3_weight(rectangle3_weights[2837]), .feature_threshold(feature_thresholds[2837]), .feature_above(feature_aboves[2837]), .feature_below(feature_belows[2837]), .scan_win_std_dev(scan_win_std_dev[2837]), .feature_accum(feature_accums[2837]));
  accum_calculator ac2838(.scan_win(scan_win2838), .rectangle1_x(rectangle1_xs[2838]), .rectangle1_y(rectangle1_ys[2838]), .rectangle1_width(rectangle1_widths[2838]), .rectangle1_height(rectangle1_heights[2838]), .rectangle1_weight(rectangle1_weights[2838]), .rectangle2_x(rectangle2_xs[2838]), .rectangle2_y(rectangle2_ys[2838]), .rectangle2_width(rectangle2_widths[2838]), .rectangle2_height(rectangle2_heights[2838]), .rectangle2_weight(rectangle2_weights[2838]), .rectangle3_x(rectangle3_xs[2838]), .rectangle3_y(rectangle3_ys[2838]), .rectangle3_width(rectangle3_widths[2838]), .rectangle3_height(rectangle3_heights[2838]), .rectangle3_weight(rectangle3_weights[2838]), .feature_threshold(feature_thresholds[2838]), .feature_above(feature_aboves[2838]), .feature_below(feature_belows[2838]), .scan_win_std_dev(scan_win_std_dev[2838]), .feature_accum(feature_accums[2838]));
  accum_calculator ac2839(.scan_win(scan_win2839), .rectangle1_x(rectangle1_xs[2839]), .rectangle1_y(rectangle1_ys[2839]), .rectangle1_width(rectangle1_widths[2839]), .rectangle1_height(rectangle1_heights[2839]), .rectangle1_weight(rectangle1_weights[2839]), .rectangle2_x(rectangle2_xs[2839]), .rectangle2_y(rectangle2_ys[2839]), .rectangle2_width(rectangle2_widths[2839]), .rectangle2_height(rectangle2_heights[2839]), .rectangle2_weight(rectangle2_weights[2839]), .rectangle3_x(rectangle3_xs[2839]), .rectangle3_y(rectangle3_ys[2839]), .rectangle3_width(rectangle3_widths[2839]), .rectangle3_height(rectangle3_heights[2839]), .rectangle3_weight(rectangle3_weights[2839]), .feature_threshold(feature_thresholds[2839]), .feature_above(feature_aboves[2839]), .feature_below(feature_belows[2839]), .scan_win_std_dev(scan_win_std_dev[2839]), .feature_accum(feature_accums[2839]));
  accum_calculator ac2840(.scan_win(scan_win2840), .rectangle1_x(rectangle1_xs[2840]), .rectangle1_y(rectangle1_ys[2840]), .rectangle1_width(rectangle1_widths[2840]), .rectangle1_height(rectangle1_heights[2840]), .rectangle1_weight(rectangle1_weights[2840]), .rectangle2_x(rectangle2_xs[2840]), .rectangle2_y(rectangle2_ys[2840]), .rectangle2_width(rectangle2_widths[2840]), .rectangle2_height(rectangle2_heights[2840]), .rectangle2_weight(rectangle2_weights[2840]), .rectangle3_x(rectangle3_xs[2840]), .rectangle3_y(rectangle3_ys[2840]), .rectangle3_width(rectangle3_widths[2840]), .rectangle3_height(rectangle3_heights[2840]), .rectangle3_weight(rectangle3_weights[2840]), .feature_threshold(feature_thresholds[2840]), .feature_above(feature_aboves[2840]), .feature_below(feature_belows[2840]), .scan_win_std_dev(scan_win_std_dev[2840]), .feature_accum(feature_accums[2840]));
  accum_calculator ac2841(.scan_win(scan_win2841), .rectangle1_x(rectangle1_xs[2841]), .rectangle1_y(rectangle1_ys[2841]), .rectangle1_width(rectangle1_widths[2841]), .rectangle1_height(rectangle1_heights[2841]), .rectangle1_weight(rectangle1_weights[2841]), .rectangle2_x(rectangle2_xs[2841]), .rectangle2_y(rectangle2_ys[2841]), .rectangle2_width(rectangle2_widths[2841]), .rectangle2_height(rectangle2_heights[2841]), .rectangle2_weight(rectangle2_weights[2841]), .rectangle3_x(rectangle3_xs[2841]), .rectangle3_y(rectangle3_ys[2841]), .rectangle3_width(rectangle3_widths[2841]), .rectangle3_height(rectangle3_heights[2841]), .rectangle3_weight(rectangle3_weights[2841]), .feature_threshold(feature_thresholds[2841]), .feature_above(feature_aboves[2841]), .feature_below(feature_belows[2841]), .scan_win_std_dev(scan_win_std_dev[2841]), .feature_accum(feature_accums[2841]));
  accum_calculator ac2842(.scan_win(scan_win2842), .rectangle1_x(rectangle1_xs[2842]), .rectangle1_y(rectangle1_ys[2842]), .rectangle1_width(rectangle1_widths[2842]), .rectangle1_height(rectangle1_heights[2842]), .rectangle1_weight(rectangle1_weights[2842]), .rectangle2_x(rectangle2_xs[2842]), .rectangle2_y(rectangle2_ys[2842]), .rectangle2_width(rectangle2_widths[2842]), .rectangle2_height(rectangle2_heights[2842]), .rectangle2_weight(rectangle2_weights[2842]), .rectangle3_x(rectangle3_xs[2842]), .rectangle3_y(rectangle3_ys[2842]), .rectangle3_width(rectangle3_widths[2842]), .rectangle3_height(rectangle3_heights[2842]), .rectangle3_weight(rectangle3_weights[2842]), .feature_threshold(feature_thresholds[2842]), .feature_above(feature_aboves[2842]), .feature_below(feature_belows[2842]), .scan_win_std_dev(scan_win_std_dev[2842]), .feature_accum(feature_accums[2842]));
  accum_calculator ac2843(.scan_win(scan_win2843), .rectangle1_x(rectangle1_xs[2843]), .rectangle1_y(rectangle1_ys[2843]), .rectangle1_width(rectangle1_widths[2843]), .rectangle1_height(rectangle1_heights[2843]), .rectangle1_weight(rectangle1_weights[2843]), .rectangle2_x(rectangle2_xs[2843]), .rectangle2_y(rectangle2_ys[2843]), .rectangle2_width(rectangle2_widths[2843]), .rectangle2_height(rectangle2_heights[2843]), .rectangle2_weight(rectangle2_weights[2843]), .rectangle3_x(rectangle3_xs[2843]), .rectangle3_y(rectangle3_ys[2843]), .rectangle3_width(rectangle3_widths[2843]), .rectangle3_height(rectangle3_heights[2843]), .rectangle3_weight(rectangle3_weights[2843]), .feature_threshold(feature_thresholds[2843]), .feature_above(feature_aboves[2843]), .feature_below(feature_belows[2843]), .scan_win_std_dev(scan_win_std_dev[2843]), .feature_accum(feature_accums[2843]));
  accum_calculator ac2844(.scan_win(scan_win2844), .rectangle1_x(rectangle1_xs[2844]), .rectangle1_y(rectangle1_ys[2844]), .rectangle1_width(rectangle1_widths[2844]), .rectangle1_height(rectangle1_heights[2844]), .rectangle1_weight(rectangle1_weights[2844]), .rectangle2_x(rectangle2_xs[2844]), .rectangle2_y(rectangle2_ys[2844]), .rectangle2_width(rectangle2_widths[2844]), .rectangle2_height(rectangle2_heights[2844]), .rectangle2_weight(rectangle2_weights[2844]), .rectangle3_x(rectangle3_xs[2844]), .rectangle3_y(rectangle3_ys[2844]), .rectangle3_width(rectangle3_widths[2844]), .rectangle3_height(rectangle3_heights[2844]), .rectangle3_weight(rectangle3_weights[2844]), .feature_threshold(feature_thresholds[2844]), .feature_above(feature_aboves[2844]), .feature_below(feature_belows[2844]), .scan_win_std_dev(scan_win_std_dev[2844]), .feature_accum(feature_accums[2844]));
  accum_calculator ac2845(.scan_win(scan_win2845), .rectangle1_x(rectangle1_xs[2845]), .rectangle1_y(rectangle1_ys[2845]), .rectangle1_width(rectangle1_widths[2845]), .rectangle1_height(rectangle1_heights[2845]), .rectangle1_weight(rectangle1_weights[2845]), .rectangle2_x(rectangle2_xs[2845]), .rectangle2_y(rectangle2_ys[2845]), .rectangle2_width(rectangle2_widths[2845]), .rectangle2_height(rectangle2_heights[2845]), .rectangle2_weight(rectangle2_weights[2845]), .rectangle3_x(rectangle3_xs[2845]), .rectangle3_y(rectangle3_ys[2845]), .rectangle3_width(rectangle3_widths[2845]), .rectangle3_height(rectangle3_heights[2845]), .rectangle3_weight(rectangle3_weights[2845]), .feature_threshold(feature_thresholds[2845]), .feature_above(feature_aboves[2845]), .feature_below(feature_belows[2845]), .scan_win_std_dev(scan_win_std_dev[2845]), .feature_accum(feature_accums[2845]));
  accum_calculator ac2846(.scan_win(scan_win2846), .rectangle1_x(rectangle1_xs[2846]), .rectangle1_y(rectangle1_ys[2846]), .rectangle1_width(rectangle1_widths[2846]), .rectangle1_height(rectangle1_heights[2846]), .rectangle1_weight(rectangle1_weights[2846]), .rectangle2_x(rectangle2_xs[2846]), .rectangle2_y(rectangle2_ys[2846]), .rectangle2_width(rectangle2_widths[2846]), .rectangle2_height(rectangle2_heights[2846]), .rectangle2_weight(rectangle2_weights[2846]), .rectangle3_x(rectangle3_xs[2846]), .rectangle3_y(rectangle3_ys[2846]), .rectangle3_width(rectangle3_widths[2846]), .rectangle3_height(rectangle3_heights[2846]), .rectangle3_weight(rectangle3_weights[2846]), .feature_threshold(feature_thresholds[2846]), .feature_above(feature_aboves[2846]), .feature_below(feature_belows[2846]), .scan_win_std_dev(scan_win_std_dev[2846]), .feature_accum(feature_accums[2846]));
  accum_calculator ac2847(.scan_win(scan_win2847), .rectangle1_x(rectangle1_xs[2847]), .rectangle1_y(rectangle1_ys[2847]), .rectangle1_width(rectangle1_widths[2847]), .rectangle1_height(rectangle1_heights[2847]), .rectangle1_weight(rectangle1_weights[2847]), .rectangle2_x(rectangle2_xs[2847]), .rectangle2_y(rectangle2_ys[2847]), .rectangle2_width(rectangle2_widths[2847]), .rectangle2_height(rectangle2_heights[2847]), .rectangle2_weight(rectangle2_weights[2847]), .rectangle3_x(rectangle3_xs[2847]), .rectangle3_y(rectangle3_ys[2847]), .rectangle3_width(rectangle3_widths[2847]), .rectangle3_height(rectangle3_heights[2847]), .rectangle3_weight(rectangle3_weights[2847]), .feature_threshold(feature_thresholds[2847]), .feature_above(feature_aboves[2847]), .feature_below(feature_belows[2847]), .scan_win_std_dev(scan_win_std_dev[2847]), .feature_accum(feature_accums[2847]));
  accum_calculator ac2848(.scan_win(scan_win2848), .rectangle1_x(rectangle1_xs[2848]), .rectangle1_y(rectangle1_ys[2848]), .rectangle1_width(rectangle1_widths[2848]), .rectangle1_height(rectangle1_heights[2848]), .rectangle1_weight(rectangle1_weights[2848]), .rectangle2_x(rectangle2_xs[2848]), .rectangle2_y(rectangle2_ys[2848]), .rectangle2_width(rectangle2_widths[2848]), .rectangle2_height(rectangle2_heights[2848]), .rectangle2_weight(rectangle2_weights[2848]), .rectangle3_x(rectangle3_xs[2848]), .rectangle3_y(rectangle3_ys[2848]), .rectangle3_width(rectangle3_widths[2848]), .rectangle3_height(rectangle3_heights[2848]), .rectangle3_weight(rectangle3_weights[2848]), .feature_threshold(feature_thresholds[2848]), .feature_above(feature_aboves[2848]), .feature_below(feature_belows[2848]), .scan_win_std_dev(scan_win_std_dev[2848]), .feature_accum(feature_accums[2848]));
  accum_calculator ac2849(.scan_win(scan_win2849), .rectangle1_x(rectangle1_xs[2849]), .rectangle1_y(rectangle1_ys[2849]), .rectangle1_width(rectangle1_widths[2849]), .rectangle1_height(rectangle1_heights[2849]), .rectangle1_weight(rectangle1_weights[2849]), .rectangle2_x(rectangle2_xs[2849]), .rectangle2_y(rectangle2_ys[2849]), .rectangle2_width(rectangle2_widths[2849]), .rectangle2_height(rectangle2_heights[2849]), .rectangle2_weight(rectangle2_weights[2849]), .rectangle3_x(rectangle3_xs[2849]), .rectangle3_y(rectangle3_ys[2849]), .rectangle3_width(rectangle3_widths[2849]), .rectangle3_height(rectangle3_heights[2849]), .rectangle3_weight(rectangle3_weights[2849]), .feature_threshold(feature_thresholds[2849]), .feature_above(feature_aboves[2849]), .feature_below(feature_belows[2849]), .scan_win_std_dev(scan_win_std_dev[2849]), .feature_accum(feature_accums[2849]));
  accum_calculator ac2850(.scan_win(scan_win2850), .rectangle1_x(rectangle1_xs[2850]), .rectangle1_y(rectangle1_ys[2850]), .rectangle1_width(rectangle1_widths[2850]), .rectangle1_height(rectangle1_heights[2850]), .rectangle1_weight(rectangle1_weights[2850]), .rectangle2_x(rectangle2_xs[2850]), .rectangle2_y(rectangle2_ys[2850]), .rectangle2_width(rectangle2_widths[2850]), .rectangle2_height(rectangle2_heights[2850]), .rectangle2_weight(rectangle2_weights[2850]), .rectangle3_x(rectangle3_xs[2850]), .rectangle3_y(rectangle3_ys[2850]), .rectangle3_width(rectangle3_widths[2850]), .rectangle3_height(rectangle3_heights[2850]), .rectangle3_weight(rectangle3_weights[2850]), .feature_threshold(feature_thresholds[2850]), .feature_above(feature_aboves[2850]), .feature_below(feature_belows[2850]), .scan_win_std_dev(scan_win_std_dev[2850]), .feature_accum(feature_accums[2850]));
  accum_calculator ac2851(.scan_win(scan_win2851), .rectangle1_x(rectangle1_xs[2851]), .rectangle1_y(rectangle1_ys[2851]), .rectangle1_width(rectangle1_widths[2851]), .rectangle1_height(rectangle1_heights[2851]), .rectangle1_weight(rectangle1_weights[2851]), .rectangle2_x(rectangle2_xs[2851]), .rectangle2_y(rectangle2_ys[2851]), .rectangle2_width(rectangle2_widths[2851]), .rectangle2_height(rectangle2_heights[2851]), .rectangle2_weight(rectangle2_weights[2851]), .rectangle3_x(rectangle3_xs[2851]), .rectangle3_y(rectangle3_ys[2851]), .rectangle3_width(rectangle3_widths[2851]), .rectangle3_height(rectangle3_heights[2851]), .rectangle3_weight(rectangle3_weights[2851]), .feature_threshold(feature_thresholds[2851]), .feature_above(feature_aboves[2851]), .feature_below(feature_belows[2851]), .scan_win_std_dev(scan_win_std_dev[2851]), .feature_accum(feature_accums[2851]));
  accum_calculator ac2852(.scan_win(scan_win2852), .rectangle1_x(rectangle1_xs[2852]), .rectangle1_y(rectangle1_ys[2852]), .rectangle1_width(rectangle1_widths[2852]), .rectangle1_height(rectangle1_heights[2852]), .rectangle1_weight(rectangle1_weights[2852]), .rectangle2_x(rectangle2_xs[2852]), .rectangle2_y(rectangle2_ys[2852]), .rectangle2_width(rectangle2_widths[2852]), .rectangle2_height(rectangle2_heights[2852]), .rectangle2_weight(rectangle2_weights[2852]), .rectangle3_x(rectangle3_xs[2852]), .rectangle3_y(rectangle3_ys[2852]), .rectangle3_width(rectangle3_widths[2852]), .rectangle3_height(rectangle3_heights[2852]), .rectangle3_weight(rectangle3_weights[2852]), .feature_threshold(feature_thresholds[2852]), .feature_above(feature_aboves[2852]), .feature_below(feature_belows[2852]), .scan_win_std_dev(scan_win_std_dev[2852]), .feature_accum(feature_accums[2852]));
  accum_calculator ac2853(.scan_win(scan_win2853), .rectangle1_x(rectangle1_xs[2853]), .rectangle1_y(rectangle1_ys[2853]), .rectangle1_width(rectangle1_widths[2853]), .rectangle1_height(rectangle1_heights[2853]), .rectangle1_weight(rectangle1_weights[2853]), .rectangle2_x(rectangle2_xs[2853]), .rectangle2_y(rectangle2_ys[2853]), .rectangle2_width(rectangle2_widths[2853]), .rectangle2_height(rectangle2_heights[2853]), .rectangle2_weight(rectangle2_weights[2853]), .rectangle3_x(rectangle3_xs[2853]), .rectangle3_y(rectangle3_ys[2853]), .rectangle3_width(rectangle3_widths[2853]), .rectangle3_height(rectangle3_heights[2853]), .rectangle3_weight(rectangle3_weights[2853]), .feature_threshold(feature_thresholds[2853]), .feature_above(feature_aboves[2853]), .feature_below(feature_belows[2853]), .scan_win_std_dev(scan_win_std_dev[2853]), .feature_accum(feature_accums[2853]));
  accum_calculator ac2854(.scan_win(scan_win2854), .rectangle1_x(rectangle1_xs[2854]), .rectangle1_y(rectangle1_ys[2854]), .rectangle1_width(rectangle1_widths[2854]), .rectangle1_height(rectangle1_heights[2854]), .rectangle1_weight(rectangle1_weights[2854]), .rectangle2_x(rectangle2_xs[2854]), .rectangle2_y(rectangle2_ys[2854]), .rectangle2_width(rectangle2_widths[2854]), .rectangle2_height(rectangle2_heights[2854]), .rectangle2_weight(rectangle2_weights[2854]), .rectangle3_x(rectangle3_xs[2854]), .rectangle3_y(rectangle3_ys[2854]), .rectangle3_width(rectangle3_widths[2854]), .rectangle3_height(rectangle3_heights[2854]), .rectangle3_weight(rectangle3_weights[2854]), .feature_threshold(feature_thresholds[2854]), .feature_above(feature_aboves[2854]), .feature_below(feature_belows[2854]), .scan_win_std_dev(scan_win_std_dev[2854]), .feature_accum(feature_accums[2854]));
  accum_calculator ac2855(.scan_win(scan_win2855), .rectangle1_x(rectangle1_xs[2855]), .rectangle1_y(rectangle1_ys[2855]), .rectangle1_width(rectangle1_widths[2855]), .rectangle1_height(rectangle1_heights[2855]), .rectangle1_weight(rectangle1_weights[2855]), .rectangle2_x(rectangle2_xs[2855]), .rectangle2_y(rectangle2_ys[2855]), .rectangle2_width(rectangle2_widths[2855]), .rectangle2_height(rectangle2_heights[2855]), .rectangle2_weight(rectangle2_weights[2855]), .rectangle3_x(rectangle3_xs[2855]), .rectangle3_y(rectangle3_ys[2855]), .rectangle3_width(rectangle3_widths[2855]), .rectangle3_height(rectangle3_heights[2855]), .rectangle3_weight(rectangle3_weights[2855]), .feature_threshold(feature_thresholds[2855]), .feature_above(feature_aboves[2855]), .feature_below(feature_belows[2855]), .scan_win_std_dev(scan_win_std_dev[2855]), .feature_accum(feature_accums[2855]));
  accum_calculator ac2856(.scan_win(scan_win2856), .rectangle1_x(rectangle1_xs[2856]), .rectangle1_y(rectangle1_ys[2856]), .rectangle1_width(rectangle1_widths[2856]), .rectangle1_height(rectangle1_heights[2856]), .rectangle1_weight(rectangle1_weights[2856]), .rectangle2_x(rectangle2_xs[2856]), .rectangle2_y(rectangle2_ys[2856]), .rectangle2_width(rectangle2_widths[2856]), .rectangle2_height(rectangle2_heights[2856]), .rectangle2_weight(rectangle2_weights[2856]), .rectangle3_x(rectangle3_xs[2856]), .rectangle3_y(rectangle3_ys[2856]), .rectangle3_width(rectangle3_widths[2856]), .rectangle3_height(rectangle3_heights[2856]), .rectangle3_weight(rectangle3_weights[2856]), .feature_threshold(feature_thresholds[2856]), .feature_above(feature_aboves[2856]), .feature_below(feature_belows[2856]), .scan_win_std_dev(scan_win_std_dev[2856]), .feature_accum(feature_accums[2856]));
  accum_calculator ac2857(.scan_win(scan_win2857), .rectangle1_x(rectangle1_xs[2857]), .rectangle1_y(rectangle1_ys[2857]), .rectangle1_width(rectangle1_widths[2857]), .rectangle1_height(rectangle1_heights[2857]), .rectangle1_weight(rectangle1_weights[2857]), .rectangle2_x(rectangle2_xs[2857]), .rectangle2_y(rectangle2_ys[2857]), .rectangle2_width(rectangle2_widths[2857]), .rectangle2_height(rectangle2_heights[2857]), .rectangle2_weight(rectangle2_weights[2857]), .rectangle3_x(rectangle3_xs[2857]), .rectangle3_y(rectangle3_ys[2857]), .rectangle3_width(rectangle3_widths[2857]), .rectangle3_height(rectangle3_heights[2857]), .rectangle3_weight(rectangle3_weights[2857]), .feature_threshold(feature_thresholds[2857]), .feature_above(feature_aboves[2857]), .feature_below(feature_belows[2857]), .scan_win_std_dev(scan_win_std_dev[2857]), .feature_accum(feature_accums[2857]));
  accum_calculator ac2858(.scan_win(scan_win2858), .rectangle1_x(rectangle1_xs[2858]), .rectangle1_y(rectangle1_ys[2858]), .rectangle1_width(rectangle1_widths[2858]), .rectangle1_height(rectangle1_heights[2858]), .rectangle1_weight(rectangle1_weights[2858]), .rectangle2_x(rectangle2_xs[2858]), .rectangle2_y(rectangle2_ys[2858]), .rectangle2_width(rectangle2_widths[2858]), .rectangle2_height(rectangle2_heights[2858]), .rectangle2_weight(rectangle2_weights[2858]), .rectangle3_x(rectangle3_xs[2858]), .rectangle3_y(rectangle3_ys[2858]), .rectangle3_width(rectangle3_widths[2858]), .rectangle3_height(rectangle3_heights[2858]), .rectangle3_weight(rectangle3_weights[2858]), .feature_threshold(feature_thresholds[2858]), .feature_above(feature_aboves[2858]), .feature_below(feature_belows[2858]), .scan_win_std_dev(scan_win_std_dev[2858]), .feature_accum(feature_accums[2858]));
  accum_calculator ac2859(.scan_win(scan_win2859), .rectangle1_x(rectangle1_xs[2859]), .rectangle1_y(rectangle1_ys[2859]), .rectangle1_width(rectangle1_widths[2859]), .rectangle1_height(rectangle1_heights[2859]), .rectangle1_weight(rectangle1_weights[2859]), .rectangle2_x(rectangle2_xs[2859]), .rectangle2_y(rectangle2_ys[2859]), .rectangle2_width(rectangle2_widths[2859]), .rectangle2_height(rectangle2_heights[2859]), .rectangle2_weight(rectangle2_weights[2859]), .rectangle3_x(rectangle3_xs[2859]), .rectangle3_y(rectangle3_ys[2859]), .rectangle3_width(rectangle3_widths[2859]), .rectangle3_height(rectangle3_heights[2859]), .rectangle3_weight(rectangle3_weights[2859]), .feature_threshold(feature_thresholds[2859]), .feature_above(feature_aboves[2859]), .feature_below(feature_belows[2859]), .scan_win_std_dev(scan_win_std_dev[2859]), .feature_accum(feature_accums[2859]));
  accum_calculator ac2860(.scan_win(scan_win2860), .rectangle1_x(rectangle1_xs[2860]), .rectangle1_y(rectangle1_ys[2860]), .rectangle1_width(rectangle1_widths[2860]), .rectangle1_height(rectangle1_heights[2860]), .rectangle1_weight(rectangle1_weights[2860]), .rectangle2_x(rectangle2_xs[2860]), .rectangle2_y(rectangle2_ys[2860]), .rectangle2_width(rectangle2_widths[2860]), .rectangle2_height(rectangle2_heights[2860]), .rectangle2_weight(rectangle2_weights[2860]), .rectangle3_x(rectangle3_xs[2860]), .rectangle3_y(rectangle3_ys[2860]), .rectangle3_width(rectangle3_widths[2860]), .rectangle3_height(rectangle3_heights[2860]), .rectangle3_weight(rectangle3_weights[2860]), .feature_threshold(feature_thresholds[2860]), .feature_above(feature_aboves[2860]), .feature_below(feature_belows[2860]), .scan_win_std_dev(scan_win_std_dev[2860]), .feature_accum(feature_accums[2860]));
  accum_calculator ac2861(.scan_win(scan_win2861), .rectangle1_x(rectangle1_xs[2861]), .rectangle1_y(rectangle1_ys[2861]), .rectangle1_width(rectangle1_widths[2861]), .rectangle1_height(rectangle1_heights[2861]), .rectangle1_weight(rectangle1_weights[2861]), .rectangle2_x(rectangle2_xs[2861]), .rectangle2_y(rectangle2_ys[2861]), .rectangle2_width(rectangle2_widths[2861]), .rectangle2_height(rectangle2_heights[2861]), .rectangle2_weight(rectangle2_weights[2861]), .rectangle3_x(rectangle3_xs[2861]), .rectangle3_y(rectangle3_ys[2861]), .rectangle3_width(rectangle3_widths[2861]), .rectangle3_height(rectangle3_heights[2861]), .rectangle3_weight(rectangle3_weights[2861]), .feature_threshold(feature_thresholds[2861]), .feature_above(feature_aboves[2861]), .feature_below(feature_belows[2861]), .scan_win_std_dev(scan_win_std_dev[2861]), .feature_accum(feature_accums[2861]));
  accum_calculator ac2862(.scan_win(scan_win2862), .rectangle1_x(rectangle1_xs[2862]), .rectangle1_y(rectangle1_ys[2862]), .rectangle1_width(rectangle1_widths[2862]), .rectangle1_height(rectangle1_heights[2862]), .rectangle1_weight(rectangle1_weights[2862]), .rectangle2_x(rectangle2_xs[2862]), .rectangle2_y(rectangle2_ys[2862]), .rectangle2_width(rectangle2_widths[2862]), .rectangle2_height(rectangle2_heights[2862]), .rectangle2_weight(rectangle2_weights[2862]), .rectangle3_x(rectangle3_xs[2862]), .rectangle3_y(rectangle3_ys[2862]), .rectangle3_width(rectangle3_widths[2862]), .rectangle3_height(rectangle3_heights[2862]), .rectangle3_weight(rectangle3_weights[2862]), .feature_threshold(feature_thresholds[2862]), .feature_above(feature_aboves[2862]), .feature_below(feature_belows[2862]), .scan_win_std_dev(scan_win_std_dev[2862]), .feature_accum(feature_accums[2862]));
  accum_calculator ac2863(.scan_win(scan_win2863), .rectangle1_x(rectangle1_xs[2863]), .rectangle1_y(rectangle1_ys[2863]), .rectangle1_width(rectangle1_widths[2863]), .rectangle1_height(rectangle1_heights[2863]), .rectangle1_weight(rectangle1_weights[2863]), .rectangle2_x(rectangle2_xs[2863]), .rectangle2_y(rectangle2_ys[2863]), .rectangle2_width(rectangle2_widths[2863]), .rectangle2_height(rectangle2_heights[2863]), .rectangle2_weight(rectangle2_weights[2863]), .rectangle3_x(rectangle3_xs[2863]), .rectangle3_y(rectangle3_ys[2863]), .rectangle3_width(rectangle3_widths[2863]), .rectangle3_height(rectangle3_heights[2863]), .rectangle3_weight(rectangle3_weights[2863]), .feature_threshold(feature_thresholds[2863]), .feature_above(feature_aboves[2863]), .feature_below(feature_belows[2863]), .scan_win_std_dev(scan_win_std_dev[2863]), .feature_accum(feature_accums[2863]));
  accum_calculator ac2864(.scan_win(scan_win2864), .rectangle1_x(rectangle1_xs[2864]), .rectangle1_y(rectangle1_ys[2864]), .rectangle1_width(rectangle1_widths[2864]), .rectangle1_height(rectangle1_heights[2864]), .rectangle1_weight(rectangle1_weights[2864]), .rectangle2_x(rectangle2_xs[2864]), .rectangle2_y(rectangle2_ys[2864]), .rectangle2_width(rectangle2_widths[2864]), .rectangle2_height(rectangle2_heights[2864]), .rectangle2_weight(rectangle2_weights[2864]), .rectangle3_x(rectangle3_xs[2864]), .rectangle3_y(rectangle3_ys[2864]), .rectangle3_width(rectangle3_widths[2864]), .rectangle3_height(rectangle3_heights[2864]), .rectangle3_weight(rectangle3_weights[2864]), .feature_threshold(feature_thresholds[2864]), .feature_above(feature_aboves[2864]), .feature_below(feature_belows[2864]), .scan_win_std_dev(scan_win_std_dev[2864]), .feature_accum(feature_accums[2864]));
  accum_calculator ac2865(.scan_win(scan_win2865), .rectangle1_x(rectangle1_xs[2865]), .rectangle1_y(rectangle1_ys[2865]), .rectangle1_width(rectangle1_widths[2865]), .rectangle1_height(rectangle1_heights[2865]), .rectangle1_weight(rectangle1_weights[2865]), .rectangle2_x(rectangle2_xs[2865]), .rectangle2_y(rectangle2_ys[2865]), .rectangle2_width(rectangle2_widths[2865]), .rectangle2_height(rectangle2_heights[2865]), .rectangle2_weight(rectangle2_weights[2865]), .rectangle3_x(rectangle3_xs[2865]), .rectangle3_y(rectangle3_ys[2865]), .rectangle3_width(rectangle3_widths[2865]), .rectangle3_height(rectangle3_heights[2865]), .rectangle3_weight(rectangle3_weights[2865]), .feature_threshold(feature_thresholds[2865]), .feature_above(feature_aboves[2865]), .feature_below(feature_belows[2865]), .scan_win_std_dev(scan_win_std_dev[2865]), .feature_accum(feature_accums[2865]));
  accum_calculator ac2866(.scan_win(scan_win2866), .rectangle1_x(rectangle1_xs[2866]), .rectangle1_y(rectangle1_ys[2866]), .rectangle1_width(rectangle1_widths[2866]), .rectangle1_height(rectangle1_heights[2866]), .rectangle1_weight(rectangle1_weights[2866]), .rectangle2_x(rectangle2_xs[2866]), .rectangle2_y(rectangle2_ys[2866]), .rectangle2_width(rectangle2_widths[2866]), .rectangle2_height(rectangle2_heights[2866]), .rectangle2_weight(rectangle2_weights[2866]), .rectangle3_x(rectangle3_xs[2866]), .rectangle3_y(rectangle3_ys[2866]), .rectangle3_width(rectangle3_widths[2866]), .rectangle3_height(rectangle3_heights[2866]), .rectangle3_weight(rectangle3_weights[2866]), .feature_threshold(feature_thresholds[2866]), .feature_above(feature_aboves[2866]), .feature_below(feature_belows[2866]), .scan_win_std_dev(scan_win_std_dev[2866]), .feature_accum(feature_accums[2866]));
  accum_calculator ac2867(.scan_win(scan_win2867), .rectangle1_x(rectangle1_xs[2867]), .rectangle1_y(rectangle1_ys[2867]), .rectangle1_width(rectangle1_widths[2867]), .rectangle1_height(rectangle1_heights[2867]), .rectangle1_weight(rectangle1_weights[2867]), .rectangle2_x(rectangle2_xs[2867]), .rectangle2_y(rectangle2_ys[2867]), .rectangle2_width(rectangle2_widths[2867]), .rectangle2_height(rectangle2_heights[2867]), .rectangle2_weight(rectangle2_weights[2867]), .rectangle3_x(rectangle3_xs[2867]), .rectangle3_y(rectangle3_ys[2867]), .rectangle3_width(rectangle3_widths[2867]), .rectangle3_height(rectangle3_heights[2867]), .rectangle3_weight(rectangle3_weights[2867]), .feature_threshold(feature_thresholds[2867]), .feature_above(feature_aboves[2867]), .feature_below(feature_belows[2867]), .scan_win_std_dev(scan_win_std_dev[2867]), .feature_accum(feature_accums[2867]));
  accum_calculator ac2868(.scan_win(scan_win2868), .rectangle1_x(rectangle1_xs[2868]), .rectangle1_y(rectangle1_ys[2868]), .rectangle1_width(rectangle1_widths[2868]), .rectangle1_height(rectangle1_heights[2868]), .rectangle1_weight(rectangle1_weights[2868]), .rectangle2_x(rectangle2_xs[2868]), .rectangle2_y(rectangle2_ys[2868]), .rectangle2_width(rectangle2_widths[2868]), .rectangle2_height(rectangle2_heights[2868]), .rectangle2_weight(rectangle2_weights[2868]), .rectangle3_x(rectangle3_xs[2868]), .rectangle3_y(rectangle3_ys[2868]), .rectangle3_width(rectangle3_widths[2868]), .rectangle3_height(rectangle3_heights[2868]), .rectangle3_weight(rectangle3_weights[2868]), .feature_threshold(feature_thresholds[2868]), .feature_above(feature_aboves[2868]), .feature_below(feature_belows[2868]), .scan_win_std_dev(scan_win_std_dev[2868]), .feature_accum(feature_accums[2868]));
  accum_calculator ac2869(.scan_win(scan_win2869), .rectangle1_x(rectangle1_xs[2869]), .rectangle1_y(rectangle1_ys[2869]), .rectangle1_width(rectangle1_widths[2869]), .rectangle1_height(rectangle1_heights[2869]), .rectangle1_weight(rectangle1_weights[2869]), .rectangle2_x(rectangle2_xs[2869]), .rectangle2_y(rectangle2_ys[2869]), .rectangle2_width(rectangle2_widths[2869]), .rectangle2_height(rectangle2_heights[2869]), .rectangle2_weight(rectangle2_weights[2869]), .rectangle3_x(rectangle3_xs[2869]), .rectangle3_y(rectangle3_ys[2869]), .rectangle3_width(rectangle3_widths[2869]), .rectangle3_height(rectangle3_heights[2869]), .rectangle3_weight(rectangle3_weights[2869]), .feature_threshold(feature_thresholds[2869]), .feature_above(feature_aboves[2869]), .feature_below(feature_belows[2869]), .scan_win_std_dev(scan_win_std_dev[2869]), .feature_accum(feature_accums[2869]));
  accum_calculator ac2870(.scan_win(scan_win2870), .rectangle1_x(rectangle1_xs[2870]), .rectangle1_y(rectangle1_ys[2870]), .rectangle1_width(rectangle1_widths[2870]), .rectangle1_height(rectangle1_heights[2870]), .rectangle1_weight(rectangle1_weights[2870]), .rectangle2_x(rectangle2_xs[2870]), .rectangle2_y(rectangle2_ys[2870]), .rectangle2_width(rectangle2_widths[2870]), .rectangle2_height(rectangle2_heights[2870]), .rectangle2_weight(rectangle2_weights[2870]), .rectangle3_x(rectangle3_xs[2870]), .rectangle3_y(rectangle3_ys[2870]), .rectangle3_width(rectangle3_widths[2870]), .rectangle3_height(rectangle3_heights[2870]), .rectangle3_weight(rectangle3_weights[2870]), .feature_threshold(feature_thresholds[2870]), .feature_above(feature_aboves[2870]), .feature_below(feature_belows[2870]), .scan_win_std_dev(scan_win_std_dev[2870]), .feature_accum(feature_accums[2870]));
  accum_calculator ac2871(.scan_win(scan_win2871), .rectangle1_x(rectangle1_xs[2871]), .rectangle1_y(rectangle1_ys[2871]), .rectangle1_width(rectangle1_widths[2871]), .rectangle1_height(rectangle1_heights[2871]), .rectangle1_weight(rectangle1_weights[2871]), .rectangle2_x(rectangle2_xs[2871]), .rectangle2_y(rectangle2_ys[2871]), .rectangle2_width(rectangle2_widths[2871]), .rectangle2_height(rectangle2_heights[2871]), .rectangle2_weight(rectangle2_weights[2871]), .rectangle3_x(rectangle3_xs[2871]), .rectangle3_y(rectangle3_ys[2871]), .rectangle3_width(rectangle3_widths[2871]), .rectangle3_height(rectangle3_heights[2871]), .rectangle3_weight(rectangle3_weights[2871]), .feature_threshold(feature_thresholds[2871]), .feature_above(feature_aboves[2871]), .feature_below(feature_belows[2871]), .scan_win_std_dev(scan_win_std_dev[2871]), .feature_accum(feature_accums[2871]));
  accum_calculator ac2872(.scan_win(scan_win2872), .rectangle1_x(rectangle1_xs[2872]), .rectangle1_y(rectangle1_ys[2872]), .rectangle1_width(rectangle1_widths[2872]), .rectangle1_height(rectangle1_heights[2872]), .rectangle1_weight(rectangle1_weights[2872]), .rectangle2_x(rectangle2_xs[2872]), .rectangle2_y(rectangle2_ys[2872]), .rectangle2_width(rectangle2_widths[2872]), .rectangle2_height(rectangle2_heights[2872]), .rectangle2_weight(rectangle2_weights[2872]), .rectangle3_x(rectangle3_xs[2872]), .rectangle3_y(rectangle3_ys[2872]), .rectangle3_width(rectangle3_widths[2872]), .rectangle3_height(rectangle3_heights[2872]), .rectangle3_weight(rectangle3_weights[2872]), .feature_threshold(feature_thresholds[2872]), .feature_above(feature_aboves[2872]), .feature_below(feature_belows[2872]), .scan_win_std_dev(scan_win_std_dev[2872]), .feature_accum(feature_accums[2872]));
  accum_calculator ac2873(.scan_win(scan_win2873), .rectangle1_x(rectangle1_xs[2873]), .rectangle1_y(rectangle1_ys[2873]), .rectangle1_width(rectangle1_widths[2873]), .rectangle1_height(rectangle1_heights[2873]), .rectangle1_weight(rectangle1_weights[2873]), .rectangle2_x(rectangle2_xs[2873]), .rectangle2_y(rectangle2_ys[2873]), .rectangle2_width(rectangle2_widths[2873]), .rectangle2_height(rectangle2_heights[2873]), .rectangle2_weight(rectangle2_weights[2873]), .rectangle3_x(rectangle3_xs[2873]), .rectangle3_y(rectangle3_ys[2873]), .rectangle3_width(rectangle3_widths[2873]), .rectangle3_height(rectangle3_heights[2873]), .rectangle3_weight(rectangle3_weights[2873]), .feature_threshold(feature_thresholds[2873]), .feature_above(feature_aboves[2873]), .feature_below(feature_belows[2873]), .scan_win_std_dev(scan_win_std_dev[2873]), .feature_accum(feature_accums[2873]));
  accum_calculator ac2874(.scan_win(scan_win2874), .rectangle1_x(rectangle1_xs[2874]), .rectangle1_y(rectangle1_ys[2874]), .rectangle1_width(rectangle1_widths[2874]), .rectangle1_height(rectangle1_heights[2874]), .rectangle1_weight(rectangle1_weights[2874]), .rectangle2_x(rectangle2_xs[2874]), .rectangle2_y(rectangle2_ys[2874]), .rectangle2_width(rectangle2_widths[2874]), .rectangle2_height(rectangle2_heights[2874]), .rectangle2_weight(rectangle2_weights[2874]), .rectangle3_x(rectangle3_xs[2874]), .rectangle3_y(rectangle3_ys[2874]), .rectangle3_width(rectangle3_widths[2874]), .rectangle3_height(rectangle3_heights[2874]), .rectangle3_weight(rectangle3_weights[2874]), .feature_threshold(feature_thresholds[2874]), .feature_above(feature_aboves[2874]), .feature_below(feature_belows[2874]), .scan_win_std_dev(scan_win_std_dev[2874]), .feature_accum(feature_accums[2874]));
  accum_calculator ac2875(.scan_win(scan_win2875), .rectangle1_x(rectangle1_xs[2875]), .rectangle1_y(rectangle1_ys[2875]), .rectangle1_width(rectangle1_widths[2875]), .rectangle1_height(rectangle1_heights[2875]), .rectangle1_weight(rectangle1_weights[2875]), .rectangle2_x(rectangle2_xs[2875]), .rectangle2_y(rectangle2_ys[2875]), .rectangle2_width(rectangle2_widths[2875]), .rectangle2_height(rectangle2_heights[2875]), .rectangle2_weight(rectangle2_weights[2875]), .rectangle3_x(rectangle3_xs[2875]), .rectangle3_y(rectangle3_ys[2875]), .rectangle3_width(rectangle3_widths[2875]), .rectangle3_height(rectangle3_heights[2875]), .rectangle3_weight(rectangle3_weights[2875]), .feature_threshold(feature_thresholds[2875]), .feature_above(feature_aboves[2875]), .feature_below(feature_belows[2875]), .scan_win_std_dev(scan_win_std_dev[2875]), .feature_accum(feature_accums[2875]));
  accum_calculator ac2876(.scan_win(scan_win2876), .rectangle1_x(rectangle1_xs[2876]), .rectangle1_y(rectangle1_ys[2876]), .rectangle1_width(rectangle1_widths[2876]), .rectangle1_height(rectangle1_heights[2876]), .rectangle1_weight(rectangle1_weights[2876]), .rectangle2_x(rectangle2_xs[2876]), .rectangle2_y(rectangle2_ys[2876]), .rectangle2_width(rectangle2_widths[2876]), .rectangle2_height(rectangle2_heights[2876]), .rectangle2_weight(rectangle2_weights[2876]), .rectangle3_x(rectangle3_xs[2876]), .rectangle3_y(rectangle3_ys[2876]), .rectangle3_width(rectangle3_widths[2876]), .rectangle3_height(rectangle3_heights[2876]), .rectangle3_weight(rectangle3_weights[2876]), .feature_threshold(feature_thresholds[2876]), .feature_above(feature_aboves[2876]), .feature_below(feature_belows[2876]), .scan_win_std_dev(scan_win_std_dev[2876]), .feature_accum(feature_accums[2876]));
  accum_calculator ac2877(.scan_win(scan_win2877), .rectangle1_x(rectangle1_xs[2877]), .rectangle1_y(rectangle1_ys[2877]), .rectangle1_width(rectangle1_widths[2877]), .rectangle1_height(rectangle1_heights[2877]), .rectangle1_weight(rectangle1_weights[2877]), .rectangle2_x(rectangle2_xs[2877]), .rectangle2_y(rectangle2_ys[2877]), .rectangle2_width(rectangle2_widths[2877]), .rectangle2_height(rectangle2_heights[2877]), .rectangle2_weight(rectangle2_weights[2877]), .rectangle3_x(rectangle3_xs[2877]), .rectangle3_y(rectangle3_ys[2877]), .rectangle3_width(rectangle3_widths[2877]), .rectangle3_height(rectangle3_heights[2877]), .rectangle3_weight(rectangle3_weights[2877]), .feature_threshold(feature_thresholds[2877]), .feature_above(feature_aboves[2877]), .feature_below(feature_belows[2877]), .scan_win_std_dev(scan_win_std_dev[2877]), .feature_accum(feature_accums[2877]));
  accum_calculator ac2878(.scan_win(scan_win2878), .rectangle1_x(rectangle1_xs[2878]), .rectangle1_y(rectangle1_ys[2878]), .rectangle1_width(rectangle1_widths[2878]), .rectangle1_height(rectangle1_heights[2878]), .rectangle1_weight(rectangle1_weights[2878]), .rectangle2_x(rectangle2_xs[2878]), .rectangle2_y(rectangle2_ys[2878]), .rectangle2_width(rectangle2_widths[2878]), .rectangle2_height(rectangle2_heights[2878]), .rectangle2_weight(rectangle2_weights[2878]), .rectangle3_x(rectangle3_xs[2878]), .rectangle3_y(rectangle3_ys[2878]), .rectangle3_width(rectangle3_widths[2878]), .rectangle3_height(rectangle3_heights[2878]), .rectangle3_weight(rectangle3_weights[2878]), .feature_threshold(feature_thresholds[2878]), .feature_above(feature_aboves[2878]), .feature_below(feature_belows[2878]), .scan_win_std_dev(scan_win_std_dev[2878]), .feature_accum(feature_accums[2878]));
  accum_calculator ac2879(.scan_win(scan_win2879), .rectangle1_x(rectangle1_xs[2879]), .rectangle1_y(rectangle1_ys[2879]), .rectangle1_width(rectangle1_widths[2879]), .rectangle1_height(rectangle1_heights[2879]), .rectangle1_weight(rectangle1_weights[2879]), .rectangle2_x(rectangle2_xs[2879]), .rectangle2_y(rectangle2_ys[2879]), .rectangle2_width(rectangle2_widths[2879]), .rectangle2_height(rectangle2_heights[2879]), .rectangle2_weight(rectangle2_weights[2879]), .rectangle3_x(rectangle3_xs[2879]), .rectangle3_y(rectangle3_ys[2879]), .rectangle3_width(rectangle3_widths[2879]), .rectangle3_height(rectangle3_heights[2879]), .rectangle3_weight(rectangle3_weights[2879]), .feature_threshold(feature_thresholds[2879]), .feature_above(feature_aboves[2879]), .feature_below(feature_belows[2879]), .scan_win_std_dev(scan_win_std_dev[2879]), .feature_accum(feature_accums[2879]));
  accum_calculator ac2880(.scan_win(scan_win2880), .rectangle1_x(rectangle1_xs[2880]), .rectangle1_y(rectangle1_ys[2880]), .rectangle1_width(rectangle1_widths[2880]), .rectangle1_height(rectangle1_heights[2880]), .rectangle1_weight(rectangle1_weights[2880]), .rectangle2_x(rectangle2_xs[2880]), .rectangle2_y(rectangle2_ys[2880]), .rectangle2_width(rectangle2_widths[2880]), .rectangle2_height(rectangle2_heights[2880]), .rectangle2_weight(rectangle2_weights[2880]), .rectangle3_x(rectangle3_xs[2880]), .rectangle3_y(rectangle3_ys[2880]), .rectangle3_width(rectangle3_widths[2880]), .rectangle3_height(rectangle3_heights[2880]), .rectangle3_weight(rectangle3_weights[2880]), .feature_threshold(feature_thresholds[2880]), .feature_above(feature_aboves[2880]), .feature_below(feature_belows[2880]), .scan_win_std_dev(scan_win_std_dev[2880]), .feature_accum(feature_accums[2880]));
  accum_calculator ac2881(.scan_win(scan_win2881), .rectangle1_x(rectangle1_xs[2881]), .rectangle1_y(rectangle1_ys[2881]), .rectangle1_width(rectangle1_widths[2881]), .rectangle1_height(rectangle1_heights[2881]), .rectangle1_weight(rectangle1_weights[2881]), .rectangle2_x(rectangle2_xs[2881]), .rectangle2_y(rectangle2_ys[2881]), .rectangle2_width(rectangle2_widths[2881]), .rectangle2_height(rectangle2_heights[2881]), .rectangle2_weight(rectangle2_weights[2881]), .rectangle3_x(rectangle3_xs[2881]), .rectangle3_y(rectangle3_ys[2881]), .rectangle3_width(rectangle3_widths[2881]), .rectangle3_height(rectangle3_heights[2881]), .rectangle3_weight(rectangle3_weights[2881]), .feature_threshold(feature_thresholds[2881]), .feature_above(feature_aboves[2881]), .feature_below(feature_belows[2881]), .scan_win_std_dev(scan_win_std_dev[2881]), .feature_accum(feature_accums[2881]));
  accum_calculator ac2882(.scan_win(scan_win2882), .rectangle1_x(rectangle1_xs[2882]), .rectangle1_y(rectangle1_ys[2882]), .rectangle1_width(rectangle1_widths[2882]), .rectangle1_height(rectangle1_heights[2882]), .rectangle1_weight(rectangle1_weights[2882]), .rectangle2_x(rectangle2_xs[2882]), .rectangle2_y(rectangle2_ys[2882]), .rectangle2_width(rectangle2_widths[2882]), .rectangle2_height(rectangle2_heights[2882]), .rectangle2_weight(rectangle2_weights[2882]), .rectangle3_x(rectangle3_xs[2882]), .rectangle3_y(rectangle3_ys[2882]), .rectangle3_width(rectangle3_widths[2882]), .rectangle3_height(rectangle3_heights[2882]), .rectangle3_weight(rectangle3_weights[2882]), .feature_threshold(feature_thresholds[2882]), .feature_above(feature_aboves[2882]), .feature_below(feature_belows[2882]), .scan_win_std_dev(scan_win_std_dev[2882]), .feature_accum(feature_accums[2882]));
  accum_calculator ac2883(.scan_win(scan_win2883), .rectangle1_x(rectangle1_xs[2883]), .rectangle1_y(rectangle1_ys[2883]), .rectangle1_width(rectangle1_widths[2883]), .rectangle1_height(rectangle1_heights[2883]), .rectangle1_weight(rectangle1_weights[2883]), .rectangle2_x(rectangle2_xs[2883]), .rectangle2_y(rectangle2_ys[2883]), .rectangle2_width(rectangle2_widths[2883]), .rectangle2_height(rectangle2_heights[2883]), .rectangle2_weight(rectangle2_weights[2883]), .rectangle3_x(rectangle3_xs[2883]), .rectangle3_y(rectangle3_ys[2883]), .rectangle3_width(rectangle3_widths[2883]), .rectangle3_height(rectangle3_heights[2883]), .rectangle3_weight(rectangle3_weights[2883]), .feature_threshold(feature_thresholds[2883]), .feature_above(feature_aboves[2883]), .feature_below(feature_belows[2883]), .scan_win_std_dev(scan_win_std_dev[2883]), .feature_accum(feature_accums[2883]));
  accum_calculator ac2884(.scan_win(scan_win2884), .rectangle1_x(rectangle1_xs[2884]), .rectangle1_y(rectangle1_ys[2884]), .rectangle1_width(rectangle1_widths[2884]), .rectangle1_height(rectangle1_heights[2884]), .rectangle1_weight(rectangle1_weights[2884]), .rectangle2_x(rectangle2_xs[2884]), .rectangle2_y(rectangle2_ys[2884]), .rectangle2_width(rectangle2_widths[2884]), .rectangle2_height(rectangle2_heights[2884]), .rectangle2_weight(rectangle2_weights[2884]), .rectangle3_x(rectangle3_xs[2884]), .rectangle3_y(rectangle3_ys[2884]), .rectangle3_width(rectangle3_widths[2884]), .rectangle3_height(rectangle3_heights[2884]), .rectangle3_weight(rectangle3_weights[2884]), .feature_threshold(feature_thresholds[2884]), .feature_above(feature_aboves[2884]), .feature_below(feature_belows[2884]), .scan_win_std_dev(scan_win_std_dev[2884]), .feature_accum(feature_accums[2884]));
  accum_calculator ac2885(.scan_win(scan_win2885), .rectangle1_x(rectangle1_xs[2885]), .rectangle1_y(rectangle1_ys[2885]), .rectangle1_width(rectangle1_widths[2885]), .rectangle1_height(rectangle1_heights[2885]), .rectangle1_weight(rectangle1_weights[2885]), .rectangle2_x(rectangle2_xs[2885]), .rectangle2_y(rectangle2_ys[2885]), .rectangle2_width(rectangle2_widths[2885]), .rectangle2_height(rectangle2_heights[2885]), .rectangle2_weight(rectangle2_weights[2885]), .rectangle3_x(rectangle3_xs[2885]), .rectangle3_y(rectangle3_ys[2885]), .rectangle3_width(rectangle3_widths[2885]), .rectangle3_height(rectangle3_heights[2885]), .rectangle3_weight(rectangle3_weights[2885]), .feature_threshold(feature_thresholds[2885]), .feature_above(feature_aboves[2885]), .feature_below(feature_belows[2885]), .scan_win_std_dev(scan_win_std_dev[2885]), .feature_accum(feature_accums[2885]));
  accum_calculator ac2886(.scan_win(scan_win2886), .rectangle1_x(rectangle1_xs[2886]), .rectangle1_y(rectangle1_ys[2886]), .rectangle1_width(rectangle1_widths[2886]), .rectangle1_height(rectangle1_heights[2886]), .rectangle1_weight(rectangle1_weights[2886]), .rectangle2_x(rectangle2_xs[2886]), .rectangle2_y(rectangle2_ys[2886]), .rectangle2_width(rectangle2_widths[2886]), .rectangle2_height(rectangle2_heights[2886]), .rectangle2_weight(rectangle2_weights[2886]), .rectangle3_x(rectangle3_xs[2886]), .rectangle3_y(rectangle3_ys[2886]), .rectangle3_width(rectangle3_widths[2886]), .rectangle3_height(rectangle3_heights[2886]), .rectangle3_weight(rectangle3_weights[2886]), .feature_threshold(feature_thresholds[2886]), .feature_above(feature_aboves[2886]), .feature_below(feature_belows[2886]), .scan_win_std_dev(scan_win_std_dev[2886]), .feature_accum(feature_accums[2886]));
  accum_calculator ac2887(.scan_win(scan_win2887), .rectangle1_x(rectangle1_xs[2887]), .rectangle1_y(rectangle1_ys[2887]), .rectangle1_width(rectangle1_widths[2887]), .rectangle1_height(rectangle1_heights[2887]), .rectangle1_weight(rectangle1_weights[2887]), .rectangle2_x(rectangle2_xs[2887]), .rectangle2_y(rectangle2_ys[2887]), .rectangle2_width(rectangle2_widths[2887]), .rectangle2_height(rectangle2_heights[2887]), .rectangle2_weight(rectangle2_weights[2887]), .rectangle3_x(rectangle3_xs[2887]), .rectangle3_y(rectangle3_ys[2887]), .rectangle3_width(rectangle3_widths[2887]), .rectangle3_height(rectangle3_heights[2887]), .rectangle3_weight(rectangle3_weights[2887]), .feature_threshold(feature_thresholds[2887]), .feature_above(feature_aboves[2887]), .feature_below(feature_belows[2887]), .scan_win_std_dev(scan_win_std_dev[2887]), .feature_accum(feature_accums[2887]));
  accum_calculator ac2888(.scan_win(scan_win2888), .rectangle1_x(rectangle1_xs[2888]), .rectangle1_y(rectangle1_ys[2888]), .rectangle1_width(rectangle1_widths[2888]), .rectangle1_height(rectangle1_heights[2888]), .rectangle1_weight(rectangle1_weights[2888]), .rectangle2_x(rectangle2_xs[2888]), .rectangle2_y(rectangle2_ys[2888]), .rectangle2_width(rectangle2_widths[2888]), .rectangle2_height(rectangle2_heights[2888]), .rectangle2_weight(rectangle2_weights[2888]), .rectangle3_x(rectangle3_xs[2888]), .rectangle3_y(rectangle3_ys[2888]), .rectangle3_width(rectangle3_widths[2888]), .rectangle3_height(rectangle3_heights[2888]), .rectangle3_weight(rectangle3_weights[2888]), .feature_threshold(feature_thresholds[2888]), .feature_above(feature_aboves[2888]), .feature_below(feature_belows[2888]), .scan_win_std_dev(scan_win_std_dev[2888]), .feature_accum(feature_accums[2888]));
  accum_calculator ac2889(.scan_win(scan_win2889), .rectangle1_x(rectangle1_xs[2889]), .rectangle1_y(rectangle1_ys[2889]), .rectangle1_width(rectangle1_widths[2889]), .rectangle1_height(rectangle1_heights[2889]), .rectangle1_weight(rectangle1_weights[2889]), .rectangle2_x(rectangle2_xs[2889]), .rectangle2_y(rectangle2_ys[2889]), .rectangle2_width(rectangle2_widths[2889]), .rectangle2_height(rectangle2_heights[2889]), .rectangle2_weight(rectangle2_weights[2889]), .rectangle3_x(rectangle3_xs[2889]), .rectangle3_y(rectangle3_ys[2889]), .rectangle3_width(rectangle3_widths[2889]), .rectangle3_height(rectangle3_heights[2889]), .rectangle3_weight(rectangle3_weights[2889]), .feature_threshold(feature_thresholds[2889]), .feature_above(feature_aboves[2889]), .feature_below(feature_belows[2889]), .scan_win_std_dev(scan_win_std_dev[2889]), .feature_accum(feature_accums[2889]));
  accum_calculator ac2890(.scan_win(scan_win2890), .rectangle1_x(rectangle1_xs[2890]), .rectangle1_y(rectangle1_ys[2890]), .rectangle1_width(rectangle1_widths[2890]), .rectangle1_height(rectangle1_heights[2890]), .rectangle1_weight(rectangle1_weights[2890]), .rectangle2_x(rectangle2_xs[2890]), .rectangle2_y(rectangle2_ys[2890]), .rectangle2_width(rectangle2_widths[2890]), .rectangle2_height(rectangle2_heights[2890]), .rectangle2_weight(rectangle2_weights[2890]), .rectangle3_x(rectangle3_xs[2890]), .rectangle3_y(rectangle3_ys[2890]), .rectangle3_width(rectangle3_widths[2890]), .rectangle3_height(rectangle3_heights[2890]), .rectangle3_weight(rectangle3_weights[2890]), .feature_threshold(feature_thresholds[2890]), .feature_above(feature_aboves[2890]), .feature_below(feature_belows[2890]), .scan_win_std_dev(scan_win_std_dev[2890]), .feature_accum(feature_accums[2890]));
  accum_calculator ac2891(.scan_win(scan_win2891), .rectangle1_x(rectangle1_xs[2891]), .rectangle1_y(rectangle1_ys[2891]), .rectangle1_width(rectangle1_widths[2891]), .rectangle1_height(rectangle1_heights[2891]), .rectangle1_weight(rectangle1_weights[2891]), .rectangle2_x(rectangle2_xs[2891]), .rectangle2_y(rectangle2_ys[2891]), .rectangle2_width(rectangle2_widths[2891]), .rectangle2_height(rectangle2_heights[2891]), .rectangle2_weight(rectangle2_weights[2891]), .rectangle3_x(rectangle3_xs[2891]), .rectangle3_y(rectangle3_ys[2891]), .rectangle3_width(rectangle3_widths[2891]), .rectangle3_height(rectangle3_heights[2891]), .rectangle3_weight(rectangle3_weights[2891]), .feature_threshold(feature_thresholds[2891]), .feature_above(feature_aboves[2891]), .feature_below(feature_belows[2891]), .scan_win_std_dev(scan_win_std_dev[2891]), .feature_accum(feature_accums[2891]));
  accum_calculator ac2892(.scan_win(scan_win2892), .rectangle1_x(rectangle1_xs[2892]), .rectangle1_y(rectangle1_ys[2892]), .rectangle1_width(rectangle1_widths[2892]), .rectangle1_height(rectangle1_heights[2892]), .rectangle1_weight(rectangle1_weights[2892]), .rectangle2_x(rectangle2_xs[2892]), .rectangle2_y(rectangle2_ys[2892]), .rectangle2_width(rectangle2_widths[2892]), .rectangle2_height(rectangle2_heights[2892]), .rectangle2_weight(rectangle2_weights[2892]), .rectangle3_x(rectangle3_xs[2892]), .rectangle3_y(rectangle3_ys[2892]), .rectangle3_width(rectangle3_widths[2892]), .rectangle3_height(rectangle3_heights[2892]), .rectangle3_weight(rectangle3_weights[2892]), .feature_threshold(feature_thresholds[2892]), .feature_above(feature_aboves[2892]), .feature_below(feature_belows[2892]), .scan_win_std_dev(scan_win_std_dev[2892]), .feature_accum(feature_accums[2892]));
  accum_calculator ac2893(.scan_win(scan_win2893), .rectangle1_x(rectangle1_xs[2893]), .rectangle1_y(rectangle1_ys[2893]), .rectangle1_width(rectangle1_widths[2893]), .rectangle1_height(rectangle1_heights[2893]), .rectangle1_weight(rectangle1_weights[2893]), .rectangle2_x(rectangle2_xs[2893]), .rectangle2_y(rectangle2_ys[2893]), .rectangle2_width(rectangle2_widths[2893]), .rectangle2_height(rectangle2_heights[2893]), .rectangle2_weight(rectangle2_weights[2893]), .rectangle3_x(rectangle3_xs[2893]), .rectangle3_y(rectangle3_ys[2893]), .rectangle3_width(rectangle3_widths[2893]), .rectangle3_height(rectangle3_heights[2893]), .rectangle3_weight(rectangle3_weights[2893]), .feature_threshold(feature_thresholds[2893]), .feature_above(feature_aboves[2893]), .feature_below(feature_belows[2893]), .scan_win_std_dev(scan_win_std_dev[2893]), .feature_accum(feature_accums[2893]));
  accum_calculator ac2894(.scan_win(scan_win2894), .rectangle1_x(rectangle1_xs[2894]), .rectangle1_y(rectangle1_ys[2894]), .rectangle1_width(rectangle1_widths[2894]), .rectangle1_height(rectangle1_heights[2894]), .rectangle1_weight(rectangle1_weights[2894]), .rectangle2_x(rectangle2_xs[2894]), .rectangle2_y(rectangle2_ys[2894]), .rectangle2_width(rectangle2_widths[2894]), .rectangle2_height(rectangle2_heights[2894]), .rectangle2_weight(rectangle2_weights[2894]), .rectangle3_x(rectangle3_xs[2894]), .rectangle3_y(rectangle3_ys[2894]), .rectangle3_width(rectangle3_widths[2894]), .rectangle3_height(rectangle3_heights[2894]), .rectangle3_weight(rectangle3_weights[2894]), .feature_threshold(feature_thresholds[2894]), .feature_above(feature_aboves[2894]), .feature_below(feature_belows[2894]), .scan_win_std_dev(scan_win_std_dev[2894]), .feature_accum(feature_accums[2894]));
  accum_calculator ac2895(.scan_win(scan_win2895), .rectangle1_x(rectangle1_xs[2895]), .rectangle1_y(rectangle1_ys[2895]), .rectangle1_width(rectangle1_widths[2895]), .rectangle1_height(rectangle1_heights[2895]), .rectangle1_weight(rectangle1_weights[2895]), .rectangle2_x(rectangle2_xs[2895]), .rectangle2_y(rectangle2_ys[2895]), .rectangle2_width(rectangle2_widths[2895]), .rectangle2_height(rectangle2_heights[2895]), .rectangle2_weight(rectangle2_weights[2895]), .rectangle3_x(rectangle3_xs[2895]), .rectangle3_y(rectangle3_ys[2895]), .rectangle3_width(rectangle3_widths[2895]), .rectangle3_height(rectangle3_heights[2895]), .rectangle3_weight(rectangle3_weights[2895]), .feature_threshold(feature_thresholds[2895]), .feature_above(feature_aboves[2895]), .feature_below(feature_belows[2895]), .scan_win_std_dev(scan_win_std_dev[2895]), .feature_accum(feature_accums[2895]));
  accum_calculator ac2896(.scan_win(scan_win2896), .rectangle1_x(rectangle1_xs[2896]), .rectangle1_y(rectangle1_ys[2896]), .rectangle1_width(rectangle1_widths[2896]), .rectangle1_height(rectangle1_heights[2896]), .rectangle1_weight(rectangle1_weights[2896]), .rectangle2_x(rectangle2_xs[2896]), .rectangle2_y(rectangle2_ys[2896]), .rectangle2_width(rectangle2_widths[2896]), .rectangle2_height(rectangle2_heights[2896]), .rectangle2_weight(rectangle2_weights[2896]), .rectangle3_x(rectangle3_xs[2896]), .rectangle3_y(rectangle3_ys[2896]), .rectangle3_width(rectangle3_widths[2896]), .rectangle3_height(rectangle3_heights[2896]), .rectangle3_weight(rectangle3_weights[2896]), .feature_threshold(feature_thresholds[2896]), .feature_above(feature_aboves[2896]), .feature_below(feature_belows[2896]), .scan_win_std_dev(scan_win_std_dev[2896]), .feature_accum(feature_accums[2896]));
  accum_calculator ac2897(.scan_win(scan_win2897), .rectangle1_x(rectangle1_xs[2897]), .rectangle1_y(rectangle1_ys[2897]), .rectangle1_width(rectangle1_widths[2897]), .rectangle1_height(rectangle1_heights[2897]), .rectangle1_weight(rectangle1_weights[2897]), .rectangle2_x(rectangle2_xs[2897]), .rectangle2_y(rectangle2_ys[2897]), .rectangle2_width(rectangle2_widths[2897]), .rectangle2_height(rectangle2_heights[2897]), .rectangle2_weight(rectangle2_weights[2897]), .rectangle3_x(rectangle3_xs[2897]), .rectangle3_y(rectangle3_ys[2897]), .rectangle3_width(rectangle3_widths[2897]), .rectangle3_height(rectangle3_heights[2897]), .rectangle3_weight(rectangle3_weights[2897]), .feature_threshold(feature_thresholds[2897]), .feature_above(feature_aboves[2897]), .feature_below(feature_belows[2897]), .scan_win_std_dev(scan_win_std_dev[2897]), .feature_accum(feature_accums[2897]));
  accum_calculator ac2898(.scan_win(scan_win2898), .rectangle1_x(rectangle1_xs[2898]), .rectangle1_y(rectangle1_ys[2898]), .rectangle1_width(rectangle1_widths[2898]), .rectangle1_height(rectangle1_heights[2898]), .rectangle1_weight(rectangle1_weights[2898]), .rectangle2_x(rectangle2_xs[2898]), .rectangle2_y(rectangle2_ys[2898]), .rectangle2_width(rectangle2_widths[2898]), .rectangle2_height(rectangle2_heights[2898]), .rectangle2_weight(rectangle2_weights[2898]), .rectangle3_x(rectangle3_xs[2898]), .rectangle3_y(rectangle3_ys[2898]), .rectangle3_width(rectangle3_widths[2898]), .rectangle3_height(rectangle3_heights[2898]), .rectangle3_weight(rectangle3_weights[2898]), .feature_threshold(feature_thresholds[2898]), .feature_above(feature_aboves[2898]), .feature_below(feature_belows[2898]), .scan_win_std_dev(scan_win_std_dev[2898]), .feature_accum(feature_accums[2898]));
  accum_calculator ac2899(.scan_win(scan_win2899), .rectangle1_x(rectangle1_xs[2899]), .rectangle1_y(rectangle1_ys[2899]), .rectangle1_width(rectangle1_widths[2899]), .rectangle1_height(rectangle1_heights[2899]), .rectangle1_weight(rectangle1_weights[2899]), .rectangle2_x(rectangle2_xs[2899]), .rectangle2_y(rectangle2_ys[2899]), .rectangle2_width(rectangle2_widths[2899]), .rectangle2_height(rectangle2_heights[2899]), .rectangle2_weight(rectangle2_weights[2899]), .rectangle3_x(rectangle3_xs[2899]), .rectangle3_y(rectangle3_ys[2899]), .rectangle3_width(rectangle3_widths[2899]), .rectangle3_height(rectangle3_heights[2899]), .rectangle3_weight(rectangle3_weights[2899]), .feature_threshold(feature_thresholds[2899]), .feature_above(feature_aboves[2899]), .feature_below(feature_belows[2899]), .scan_win_std_dev(scan_win_std_dev[2899]), .feature_accum(feature_accums[2899]));
  accum_calculator ac2900(.scan_win(scan_win2900), .rectangle1_x(rectangle1_xs[2900]), .rectangle1_y(rectangle1_ys[2900]), .rectangle1_width(rectangle1_widths[2900]), .rectangle1_height(rectangle1_heights[2900]), .rectangle1_weight(rectangle1_weights[2900]), .rectangle2_x(rectangle2_xs[2900]), .rectangle2_y(rectangle2_ys[2900]), .rectangle2_width(rectangle2_widths[2900]), .rectangle2_height(rectangle2_heights[2900]), .rectangle2_weight(rectangle2_weights[2900]), .rectangle3_x(rectangle3_xs[2900]), .rectangle3_y(rectangle3_ys[2900]), .rectangle3_width(rectangle3_widths[2900]), .rectangle3_height(rectangle3_heights[2900]), .rectangle3_weight(rectangle3_weights[2900]), .feature_threshold(feature_thresholds[2900]), .feature_above(feature_aboves[2900]), .feature_below(feature_belows[2900]), .scan_win_std_dev(scan_win_std_dev[2900]), .feature_accum(feature_accums[2900]));
  accum_calculator ac2901(.scan_win(scan_win2901), .rectangle1_x(rectangle1_xs[2901]), .rectangle1_y(rectangle1_ys[2901]), .rectangle1_width(rectangle1_widths[2901]), .rectangle1_height(rectangle1_heights[2901]), .rectangle1_weight(rectangle1_weights[2901]), .rectangle2_x(rectangle2_xs[2901]), .rectangle2_y(rectangle2_ys[2901]), .rectangle2_width(rectangle2_widths[2901]), .rectangle2_height(rectangle2_heights[2901]), .rectangle2_weight(rectangle2_weights[2901]), .rectangle3_x(rectangle3_xs[2901]), .rectangle3_y(rectangle3_ys[2901]), .rectangle3_width(rectangle3_widths[2901]), .rectangle3_height(rectangle3_heights[2901]), .rectangle3_weight(rectangle3_weights[2901]), .feature_threshold(feature_thresholds[2901]), .feature_above(feature_aboves[2901]), .feature_below(feature_belows[2901]), .scan_win_std_dev(scan_win_std_dev[2901]), .feature_accum(feature_accums[2901]));
  accum_calculator ac2902(.scan_win(scan_win2902), .rectangle1_x(rectangle1_xs[2902]), .rectangle1_y(rectangle1_ys[2902]), .rectangle1_width(rectangle1_widths[2902]), .rectangle1_height(rectangle1_heights[2902]), .rectangle1_weight(rectangle1_weights[2902]), .rectangle2_x(rectangle2_xs[2902]), .rectangle2_y(rectangle2_ys[2902]), .rectangle2_width(rectangle2_widths[2902]), .rectangle2_height(rectangle2_heights[2902]), .rectangle2_weight(rectangle2_weights[2902]), .rectangle3_x(rectangle3_xs[2902]), .rectangle3_y(rectangle3_ys[2902]), .rectangle3_width(rectangle3_widths[2902]), .rectangle3_height(rectangle3_heights[2902]), .rectangle3_weight(rectangle3_weights[2902]), .feature_threshold(feature_thresholds[2902]), .feature_above(feature_aboves[2902]), .feature_below(feature_belows[2902]), .scan_win_std_dev(scan_win_std_dev[2902]), .feature_accum(feature_accums[2902]));
  accum_calculator ac2903(.scan_win(scan_win2903), .rectangle1_x(rectangle1_xs[2903]), .rectangle1_y(rectangle1_ys[2903]), .rectangle1_width(rectangle1_widths[2903]), .rectangle1_height(rectangle1_heights[2903]), .rectangle1_weight(rectangle1_weights[2903]), .rectangle2_x(rectangle2_xs[2903]), .rectangle2_y(rectangle2_ys[2903]), .rectangle2_width(rectangle2_widths[2903]), .rectangle2_height(rectangle2_heights[2903]), .rectangle2_weight(rectangle2_weights[2903]), .rectangle3_x(rectangle3_xs[2903]), .rectangle3_y(rectangle3_ys[2903]), .rectangle3_width(rectangle3_widths[2903]), .rectangle3_height(rectangle3_heights[2903]), .rectangle3_weight(rectangle3_weights[2903]), .feature_threshold(feature_thresholds[2903]), .feature_above(feature_aboves[2903]), .feature_below(feature_belows[2903]), .scan_win_std_dev(scan_win_std_dev[2903]), .feature_accum(feature_accums[2903]));
  accum_calculator ac2904(.scan_win(scan_win2904), .rectangle1_x(rectangle1_xs[2904]), .rectangle1_y(rectangle1_ys[2904]), .rectangle1_width(rectangle1_widths[2904]), .rectangle1_height(rectangle1_heights[2904]), .rectangle1_weight(rectangle1_weights[2904]), .rectangle2_x(rectangle2_xs[2904]), .rectangle2_y(rectangle2_ys[2904]), .rectangle2_width(rectangle2_widths[2904]), .rectangle2_height(rectangle2_heights[2904]), .rectangle2_weight(rectangle2_weights[2904]), .rectangle3_x(rectangle3_xs[2904]), .rectangle3_y(rectangle3_ys[2904]), .rectangle3_width(rectangle3_widths[2904]), .rectangle3_height(rectangle3_heights[2904]), .rectangle3_weight(rectangle3_weights[2904]), .feature_threshold(feature_thresholds[2904]), .feature_above(feature_aboves[2904]), .feature_below(feature_belows[2904]), .scan_win_std_dev(scan_win_std_dev[2904]), .feature_accum(feature_accums[2904]));
  accum_calculator ac2905(.scan_win(scan_win2905), .rectangle1_x(rectangle1_xs[2905]), .rectangle1_y(rectangle1_ys[2905]), .rectangle1_width(rectangle1_widths[2905]), .rectangle1_height(rectangle1_heights[2905]), .rectangle1_weight(rectangle1_weights[2905]), .rectangle2_x(rectangle2_xs[2905]), .rectangle2_y(rectangle2_ys[2905]), .rectangle2_width(rectangle2_widths[2905]), .rectangle2_height(rectangle2_heights[2905]), .rectangle2_weight(rectangle2_weights[2905]), .rectangle3_x(rectangle3_xs[2905]), .rectangle3_y(rectangle3_ys[2905]), .rectangle3_width(rectangle3_widths[2905]), .rectangle3_height(rectangle3_heights[2905]), .rectangle3_weight(rectangle3_weights[2905]), .feature_threshold(feature_thresholds[2905]), .feature_above(feature_aboves[2905]), .feature_below(feature_belows[2905]), .scan_win_std_dev(scan_win_std_dev[2905]), .feature_accum(feature_accums[2905]));
  accum_calculator ac2906(.scan_win(scan_win2906), .rectangle1_x(rectangle1_xs[2906]), .rectangle1_y(rectangle1_ys[2906]), .rectangle1_width(rectangle1_widths[2906]), .rectangle1_height(rectangle1_heights[2906]), .rectangle1_weight(rectangle1_weights[2906]), .rectangle2_x(rectangle2_xs[2906]), .rectangle2_y(rectangle2_ys[2906]), .rectangle2_width(rectangle2_widths[2906]), .rectangle2_height(rectangle2_heights[2906]), .rectangle2_weight(rectangle2_weights[2906]), .rectangle3_x(rectangle3_xs[2906]), .rectangle3_y(rectangle3_ys[2906]), .rectangle3_width(rectangle3_widths[2906]), .rectangle3_height(rectangle3_heights[2906]), .rectangle3_weight(rectangle3_weights[2906]), .feature_threshold(feature_thresholds[2906]), .feature_above(feature_aboves[2906]), .feature_below(feature_belows[2906]), .scan_win_std_dev(scan_win_std_dev[2906]), .feature_accum(feature_accums[2906]));
  accum_calculator ac2907(.scan_win(scan_win2907), .rectangle1_x(rectangle1_xs[2907]), .rectangle1_y(rectangle1_ys[2907]), .rectangle1_width(rectangle1_widths[2907]), .rectangle1_height(rectangle1_heights[2907]), .rectangle1_weight(rectangle1_weights[2907]), .rectangle2_x(rectangle2_xs[2907]), .rectangle2_y(rectangle2_ys[2907]), .rectangle2_width(rectangle2_widths[2907]), .rectangle2_height(rectangle2_heights[2907]), .rectangle2_weight(rectangle2_weights[2907]), .rectangle3_x(rectangle3_xs[2907]), .rectangle3_y(rectangle3_ys[2907]), .rectangle3_width(rectangle3_widths[2907]), .rectangle3_height(rectangle3_heights[2907]), .rectangle3_weight(rectangle3_weights[2907]), .feature_threshold(feature_thresholds[2907]), .feature_above(feature_aboves[2907]), .feature_below(feature_belows[2907]), .scan_win_std_dev(scan_win_std_dev[2907]), .feature_accum(feature_accums[2907]));
  accum_calculator ac2908(.scan_win(scan_win2908), .rectangle1_x(rectangle1_xs[2908]), .rectangle1_y(rectangle1_ys[2908]), .rectangle1_width(rectangle1_widths[2908]), .rectangle1_height(rectangle1_heights[2908]), .rectangle1_weight(rectangle1_weights[2908]), .rectangle2_x(rectangle2_xs[2908]), .rectangle2_y(rectangle2_ys[2908]), .rectangle2_width(rectangle2_widths[2908]), .rectangle2_height(rectangle2_heights[2908]), .rectangle2_weight(rectangle2_weights[2908]), .rectangle3_x(rectangle3_xs[2908]), .rectangle3_y(rectangle3_ys[2908]), .rectangle3_width(rectangle3_widths[2908]), .rectangle3_height(rectangle3_heights[2908]), .rectangle3_weight(rectangle3_weights[2908]), .feature_threshold(feature_thresholds[2908]), .feature_above(feature_aboves[2908]), .feature_below(feature_belows[2908]), .scan_win_std_dev(scan_win_std_dev[2908]), .feature_accum(feature_accums[2908]));
  accum_calculator ac2909(.scan_win(scan_win2909), .rectangle1_x(rectangle1_xs[2909]), .rectangle1_y(rectangle1_ys[2909]), .rectangle1_width(rectangle1_widths[2909]), .rectangle1_height(rectangle1_heights[2909]), .rectangle1_weight(rectangle1_weights[2909]), .rectangle2_x(rectangle2_xs[2909]), .rectangle2_y(rectangle2_ys[2909]), .rectangle2_width(rectangle2_widths[2909]), .rectangle2_height(rectangle2_heights[2909]), .rectangle2_weight(rectangle2_weights[2909]), .rectangle3_x(rectangle3_xs[2909]), .rectangle3_y(rectangle3_ys[2909]), .rectangle3_width(rectangle3_widths[2909]), .rectangle3_height(rectangle3_heights[2909]), .rectangle3_weight(rectangle3_weights[2909]), .feature_threshold(feature_thresholds[2909]), .feature_above(feature_aboves[2909]), .feature_below(feature_belows[2909]), .scan_win_std_dev(scan_win_std_dev[2909]), .feature_accum(feature_accums[2909]));
  accum_calculator ac2910(.scan_win(scan_win2910), .rectangle1_x(rectangle1_xs[2910]), .rectangle1_y(rectangle1_ys[2910]), .rectangle1_width(rectangle1_widths[2910]), .rectangle1_height(rectangle1_heights[2910]), .rectangle1_weight(rectangle1_weights[2910]), .rectangle2_x(rectangle2_xs[2910]), .rectangle2_y(rectangle2_ys[2910]), .rectangle2_width(rectangle2_widths[2910]), .rectangle2_height(rectangle2_heights[2910]), .rectangle2_weight(rectangle2_weights[2910]), .rectangle3_x(rectangle3_xs[2910]), .rectangle3_y(rectangle3_ys[2910]), .rectangle3_width(rectangle3_widths[2910]), .rectangle3_height(rectangle3_heights[2910]), .rectangle3_weight(rectangle3_weights[2910]), .feature_threshold(feature_thresholds[2910]), .feature_above(feature_aboves[2910]), .feature_below(feature_belows[2910]), .scan_win_std_dev(scan_win_std_dev[2910]), .feature_accum(feature_accums[2910]));
  accum_calculator ac2911(.scan_win(scan_win2911), .rectangle1_x(rectangle1_xs[2911]), .rectangle1_y(rectangle1_ys[2911]), .rectangle1_width(rectangle1_widths[2911]), .rectangle1_height(rectangle1_heights[2911]), .rectangle1_weight(rectangle1_weights[2911]), .rectangle2_x(rectangle2_xs[2911]), .rectangle2_y(rectangle2_ys[2911]), .rectangle2_width(rectangle2_widths[2911]), .rectangle2_height(rectangle2_heights[2911]), .rectangle2_weight(rectangle2_weights[2911]), .rectangle3_x(rectangle3_xs[2911]), .rectangle3_y(rectangle3_ys[2911]), .rectangle3_width(rectangle3_widths[2911]), .rectangle3_height(rectangle3_heights[2911]), .rectangle3_weight(rectangle3_weights[2911]), .feature_threshold(feature_thresholds[2911]), .feature_above(feature_aboves[2911]), .feature_below(feature_belows[2911]), .scan_win_std_dev(scan_win_std_dev[2911]), .feature_accum(feature_accums[2911]));
  accum_calculator ac2912(.scan_win(scan_win2912), .rectangle1_x(rectangle1_xs[2912]), .rectangle1_y(rectangle1_ys[2912]), .rectangle1_width(rectangle1_widths[2912]), .rectangle1_height(rectangle1_heights[2912]), .rectangle1_weight(rectangle1_weights[2912]), .rectangle2_x(rectangle2_xs[2912]), .rectangle2_y(rectangle2_ys[2912]), .rectangle2_width(rectangle2_widths[2912]), .rectangle2_height(rectangle2_heights[2912]), .rectangle2_weight(rectangle2_weights[2912]), .rectangle3_x(rectangle3_xs[2912]), .rectangle3_y(rectangle3_ys[2912]), .rectangle3_width(rectangle3_widths[2912]), .rectangle3_height(rectangle3_heights[2912]), .rectangle3_weight(rectangle3_weights[2912]), .feature_threshold(feature_thresholds[2912]), .feature_above(feature_aboves[2912]), .feature_below(feature_belows[2912]), .scan_win_std_dev(scan_win_std_dev[2912]), .feature_accum(feature_accums[2912]));

endmodule

module accum_calculator(
  input  logic [`WINDOW_SIZE-1:0][`WINDOW_SIZE-1:0][31:0] scan_win,
  input  logic [31:0] rectangle1_x, rectangle1_y, rectangle1_width, rectangle1_height, rectangle1_weight,
                      rectangle2_x, rectangle2_y, rectangle2_width, rectangle2_height, rectangle2_weight,
                      rectangle3_x, rectangle3_y, rectangle3_width, rectangle3_height, rectangle3_weight, 
                      feature_threshold, feature_above, feature_below, scan_win_std_dev,
  output logic [31:0] feature_accum);

  logic [31:0] rectangle1_val, rectangle2_val, rectangle3_val, 
               rectangle1_product, rectangle2_product, rectangle3_product,
               feature_product, feature_sum;
  logic feature_comparison;

  assign rectangle1_val = scan_win[rectangle1_y + rectangle1_height][rectangle1_x + rectangle1_width] +
                          scan_win[rectangle1_y][rectangle1_x]-
                          scan_win[rectangle1_y][rectangle1_x + rectangle1_width] -
                          scan_win[rectangle1_y + rectangle1_height][rectangle1_x];
  assign rectangle2_val = scan_win[rectangle2_y + rectangle2_height][rectangle2_x + rectangle2_width] +
                          scan_win[rectangle2_y][rectangle2_x]-
                          scan_win[rectangle2_y][rectangle2_x + rectangle2_width] -
                          scan_win[rectangle2_y + rectangle2_height][rectangle2_x];
  assign rectangle3_val = scan_win[rectangle3_y + rectangle3_height][rectangle3_x + rectangle3_width] +
                          scan_win[rectangle3_y][rectangle3_x]-
                          scan_win[rectangle3_y][rectangle3_x + rectangle3_width] -
                          scan_win[rectangle3_y + rectangle3_height][rectangle3_x];
  multiplier m1(.out(rectangle1_product), .a(rectangle1_val), .b(rectangle1_weight));
  multiplier m2(.out(rectangle2_product), .a(rectangle2_val), .b(rectangle2_weight));
  multiplier m3(.out(rectangle3_product), .a(rectangle3_val), .b(rectangle3_weight));
  multiplier m4(.out(feature_product), .a(feature_threshold), .b(scan_win_std_dev));
  assign feature_sum = rectangle1_product + rectangle2_product + rectangle3_product;
  signed_comparator feature_c(.gt(feature_comparison), .A(feature_sum), .B(feature_product));
  assign feature_accum = (feature_comparison) ? feature_above : feature_below;

endmodule