/** @file vj_weights.vh
 *  @brief Viola-Jones weights data structure
 */

// assume we use haarcascade_frontalface_default.xml
`define NUM_STAGE 25
`define NUM_FEATURE 2913
`define WINDOW_SIZE 24
`define LAPTOP_WIDTH 320
`define LAPTOP_HEIGHT 240
`define PYRAMID_LEVELS 13

localparam int[13] pyramid_widths = {320, 266, 222, 185, 154, 128, 107, 89, 74, 62, 51, 43, 35};
localparam int[13] pyramid_heights = {240, 199, 166, 138, 115, 96, 80, 66, 55, 46, 38, 32, 26};
localparam logic [12:0][31:0] x_ratios = 
{32'd78841, 32'd78526, 32'd78644, 32'd78729, 32'd78849, 32'd78399, 32'd78791, 
 32'd78821, 32'd78221, 32'd79672, 32'd77729, 32'd80516};
localparam logic [12:0][31:0] y_ratios = 
{32'd79039, 32'd78565, 32'd78834, 32'd78644, 32'd78507, 32'd78644, 32'd79438, 
 32'd78644, 32'd78359, 32'd79334, 32'd77825, 32'd80660};

localparam logic [25:0][31:0] stage_num_feature = {32'sd0, 32'sd9, 32'sd25, 32'sd52, 32'sd84, 32'sd136, 32'sd189, 32'sd251, 32'sd323, 32'sd406, 32'sd497, 32'sd596, 32'sd711, 32'sd838, 32'sd973, 32'sd1109, 32'sd1246, 32'sd1405, 32'sd1560, 32'sd1729, 32'sd1925, 32'sd2122, 32'sd2303, 32'sd2502, 32'sd2713, 32'sd2913}

localparam logic [24:0][31:0] stage_threshold = {-32'sd258, -32'sd255, -32'sd238, -32'sd228, -32'sd225, -32'sd211, -32'sd206, -32'sd199, -32'sd197, -32'sd187, -32'sd198, -32'sd190, -32'sd183, -32'sd190, -32'sd175, -32'sd180, -32'sd184, -32'sd174, -32'sd166, -32'sd164, -32'sd168, -32'sd170, -32'sd167, -32'sd173, -32'sd153};

localparam logic [2912:0][31:0] rectangle1_xs = {32'sd6, 32'sd6, 32'sd3, 32'sd8, 32'sd3, 32'sd6, 32'sd5, 32'sd11, 32'sd4, 32'sd6, 32'sd6, 32'sd1, 32'sd0, 32'sd9, 32'sd5, 32'sd5, 32'sd13, 32'sd7, 32'sd10, 32'sd2, 32'sd18, 32'sd0, 32'sd9, 32'sd7, 32'sd5, 32'sd0, 32'sd5, 32'sd9, 32'sd9, 32'sd6, 32'sd3, 32'sd5, 32'sd18, 32'sd1, 32'sd0, 32'sd5, 32'sd2, 32'sd8, 32'sd2, 32'sd0, 32'sd20, 32'sd0, 32'sd18, 32'sd0, 32'sd12, 32'sd0, 32'sd12, 32'sd8, 32'sd5, 32'sd1, 32'sd17, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd4, 32'sd2, 32'sd19, 32'sd1, 32'sd0, 32'sd1, 32'sd14, 32'sd3, 32'sd6, 32'sd8, 32'sd15, 32'sd1, 32'sd4, 32'sd0, 32'sd3, 32'sd1, 32'sd5, 32'sd3, 32'sd14, 32'sd1, 32'sd11, 32'sd5, 32'sd6, 32'sd9, 32'sd9, 32'sd7, 32'sd10, 32'sd8, 32'sd3, 32'sd6, 32'sd0, 32'sd4, 32'sd11, 32'sd0, 32'sd11, 32'sd4, 32'sd11, 32'sd9, 32'sd9, 32'sd1, 32'sd10, 32'sd6, 32'sd7, 32'sd0, 32'sd6, 32'sd1, 32'sd6, 32'sd2, 32'sd20, 32'sd0, 32'sd2, 32'sd0, 32'sd12, 32'sd5, 32'sd11, 32'sd0, 32'sd12, 32'sd6, 32'sd8, 32'sd0, 32'sd10, 32'sd3, 32'sd2, 32'sd2, 32'sd3, 32'sd5, 32'sd9, 32'sd4, 32'sd4, 32'sd6, 32'sd3, 32'sd0, 32'sd6, 32'sd6, 32'sd3, 32'sd1, 32'sd8, 32'sd0, 32'sd12, 32'sd0, 32'sd19, 32'sd0, 32'sd6, 32'sd7, 32'sd9, 32'sd0, 32'sd4, 32'sd7, 32'sd18, 32'sd0, 32'sd18, 32'sd0, 32'sd16, 32'sd2, 32'sd9, 32'sd2, 32'sd14, 32'sd5, 32'sd15, 32'sd0, 32'sd8, 32'sd7, 32'sd0, 32'sd1, 32'sd14, 32'sd7, 32'sd10, 32'sd4, 32'sd10, 32'sd1, 32'sd10, 32'sd5, 32'sd8, 32'sd6, 32'sd7, 32'sd0, 32'sd1, 32'sd5, 32'sd12, 32'sd6, 32'sd7, 32'sd0, 32'sd2, 32'sd2, 32'sd14, 32'sd8, 32'sd14, 32'sd8, 32'sd17, 32'sd6, 32'sd13, 32'sd3, 32'sd9, 32'sd0, 32'sd0, 32'sd6, 32'sd7, 32'sd10, 32'sd1, 32'sd5, 32'sd9, 32'sd20, 32'sd2, 32'sd5, 32'sd0, 32'sd5, 32'sd0, 32'sd6, 32'sd0, 32'sd1, 32'sd2, 32'sd2, 32'sd0, 32'sd9, 32'sd7, 32'sd11, 32'sd6, 32'sd18, 32'sd3, 32'sd18, 32'sd1, 32'sd11, 32'sd0, 32'sd13, 32'sd7, 32'sd11, 32'sd8, 32'sd13, 32'sd2, 32'sd3, 32'sd0, 32'sd9, 32'sd4, 32'sd7, 32'sd0, 32'sd7, 32'sd7, 32'sd3, 32'sd0, 32'sd3, 32'sd4, 32'sd13, 32'sd9, 32'sd5, 32'sd1, 32'sd10, 32'sd0, 32'sd1, 32'sd4, 32'sd0, 32'sd2, 32'sd9, 32'sd5, 32'sd17, 32'sd1, 32'sd14, 32'sd3, 32'sd15, 32'sd9, 32'sd17, 32'sd3, 32'sd7, 32'sd1, 32'sd10, 32'sd0, 32'sd15, 32'sd3, 32'sd12, 32'sd6, 32'sd14, 32'sd1, 32'sd13, 32'sd7, 32'sd12, 32'sd6, 32'sd6, 32'sd7, 32'sd7, 32'sd8, 32'sd7, 32'sd0, 32'sd15, 32'sd0, 32'sd15, 32'sd7, 32'sd15, 32'sd0, 32'sd8, 32'sd0, 32'sd3, 32'sd0, 32'sd9, 32'sd10, 32'sd7, 32'sd5, 32'sd14, 32'sd2, 32'sd0, 32'sd4, 32'sd9, 32'sd0, 32'sd18, 32'sd0, 32'sd8, 32'sd8, 32'sd11, 32'sd7, 32'sd12, 32'sd6, 32'sd15, 32'sd5, 32'sd9, 32'sd7, 32'sd14, 32'sd2, 32'sd5, 32'sd9, 32'sd12, 32'sd9, 32'sd3, 32'sd6, 32'sd12, 32'sd1, 32'sd12, 32'sd1, 32'sd10, 32'sd3, 32'sd10, 32'sd0, 32'sd6, 32'sd6, 32'sd5, 32'sd4, 32'sd11, 32'sd7, 32'sd3, 32'sd2, 32'sd3, 32'sd8, 32'sd16, 32'sd7, 32'sd18, 32'sd0, 32'sd18, 32'sd3, 32'sd18, 32'sd0, 32'sd5, 32'sd6, 32'sd10, 32'sd8, 32'sd15, 32'sd3, 32'sd15, 32'sd2, 32'sd8, 32'sd8, 32'sd15, 32'sd4, 32'sd13, 32'sd7, 32'sd18, 32'sd1, 32'sd14, 32'sd1, 32'sd4, 32'sd1, 32'sd10, 32'sd0, 32'sd15, 32'sd3, 32'sd15, 32'sd3, 32'sd15, 32'sd0, 32'sd4, 32'sd2, 32'sd14, 32'sd6, 32'sd17, 32'sd1, 32'sd16, 32'sd7, 32'sd12, 32'sd4, 32'sd10, 32'sd2, 32'sd15, 32'sd0, 32'sd6, 32'sd1, 32'sd6, 32'sd0, 32'sd8, 32'sd9, 32'sd6, 32'sd0, 32'sd16, 32'sd0, 32'sd14, 32'sd1, 32'sd5, 32'sd4, 32'sd16, 32'sd0, 32'sd10, 32'sd9, 32'sd9, 32'sd3, 32'sd6, 32'sd8, 32'sd0, 32'sd14, 32'sd5, 32'sd9, 32'sd0, 32'sd3, 32'sd3, 32'sd20, 32'sd0, 32'sd8, 32'sd6, 32'sd9, 32'sd1, 32'sd9, 32'sd7, 32'sd13, 32'sd7, 32'sd14, 32'sd2, 32'sd18, 32'sd6, 32'sd18, 32'sd7, 32'sd18, 32'sd0, 32'sd9, 32'sd0, 32'sd17, 32'sd1, 32'sd14, 32'sd6, 32'sd3, 32'sd9, 32'sd12, 32'sd6, 32'sd6, 32'sd1, 32'sd10, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd1, 32'sd6, 32'sd4, 32'sd1, 32'sd5, 32'sd0, 32'sd3, 32'sd2, 32'sd6, 32'sd14, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd3, 32'sd6, 32'sd0, 32'sd13, 32'sd7, 32'sd9, 32'sd1, 32'sd13, 32'sd5, 32'sd16, 32'sd4, 32'sd0, 32'sd5, 32'sd12, 32'sd2, 32'sd15, 32'sd0, 32'sd12, 32'sd11, 32'sd9, 32'sd8, 32'sd12, 32'sd3, 32'sd6, 32'sd7, 32'sd12, 32'sd10, 32'sd16, 32'sd4, 32'sd2, 32'sd5, 32'sd10, 32'sd8, 32'sd6, 32'sd6, 32'sd0, 32'sd1, 32'sd3, 32'sd3, 32'sd0, 32'sd10, 32'sd8, 32'sd5, 32'sd0, 32'sd14, 32'sd9, 32'sd14, 32'sd1, 32'sd15, 32'sd0, 32'sd17, 32'sd2, 32'sd3, 32'sd9, 32'sd18, 32'sd0, 32'sd4, 32'sd2, 32'sd14, 32'sd0, 32'sd18, 32'sd5, 32'sd21, 32'sd6, 32'sd8, 32'sd7, 32'sd21, 32'sd10, 32'sd15, 32'sd0, 32'sd11, 32'sd7, 32'sd12, 32'sd6, 32'sd14, 32'sd6, 32'sd3, 32'sd3, 32'sd0, 32'sd10, 32'sd11, 32'sd6, 32'sd16, 32'sd3, 32'sd16, 32'sd0, 32'sd10, 32'sd0, 32'sd13, 32'sd7, 32'sd5, 32'sd0, 32'sd6, 32'sd3, 32'sd8, 32'sd2, 32'sd15, 32'sd3, 32'sd17, 32'sd1, 32'sd19, 32'sd1, 32'sd4, 32'sd6, 32'sd15, 32'sd0, 32'sd15, 32'sd3, 32'sd8, 32'sd6, 32'sd5, 32'sd10, 32'sd10, 32'sd0, 32'sd15, 32'sd0, 32'sd12, 32'sd9, 32'sd12, 32'sd6, 32'sd15, 32'sd0, 32'sd11, 32'sd6, 32'sd10, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd12, 32'sd2, 32'sd7, 32'sd0, 32'sd3, 32'sd6, 32'sd5, 32'sd11, 32'sd0, 32'sd18, 32'sd3, 32'sd9, 32'sd0, 32'sd13, 32'sd0, 32'sd13, 32'sd4, 32'sd13, 32'sd5, 32'sd7, 32'sd6, 32'sd14, 32'sd4, 32'sd11, 32'sd0, 32'sd13, 32'sd2, 32'sd10, 32'sd8, 32'sd14, 32'sd6, 32'sd8, 32'sd7, 32'sd8, 32'sd5, 32'sd3, 32'sd0, 32'sd5, 32'sd0, 32'sd3, 32'sd1, 32'sd5, 32'sd1, 32'sd1, 32'sd3, 32'sd6, 32'sd6, 32'sd14, 32'sd1, 32'sd11, 32'sd10, 32'sd11, 32'sd7, 32'sd12, 32'sd2, 32'sd14, 32'sd6, 32'sd14, 32'sd0, 32'sd5, 32'sd1, 32'sd13, 32'sd7, 32'sd12, 32'sd0, 32'sd7, 32'sd7, 32'sd8, 32'sd1, 32'sd13, 32'sd5, 32'sd14, 32'sd4, 32'sd12, 32'sd9, 32'sd11, 32'sd5, 32'sd8, 32'sd1, 32'sd9, 32'sd3, 32'sd12, 32'sd8, 32'sd2, 32'sd0, 32'sd14, 32'sd2, 32'sd2, 32'sd6, 32'sd5, 32'sd1, 32'sd7, 32'sd3, 32'sd9, 32'sd2, 32'sd18, 
                                                    32'sd3, 32'sd20, 32'sd2, 32'sd1, 32'sd0, 32'sd19, 32'sd0, 32'sd18, 32'sd0, 32'sd7, 32'sd0, 32'sd10, 32'sd8, 32'sd4, 32'sd2, 32'sd7, 32'sd3, 32'sd16, 32'sd5, 32'sd10, 32'sd4, 32'sd2, 32'sd6, 32'sd1, 32'sd12, 32'sd0, 32'sd15, 32'sd5, 32'sd8, 32'sd1, 32'sd17, 32'sd8, 32'sd17, 32'sd7, 32'sd15, 32'sd2, 32'sd10, 32'sd0, 32'sd20, 32'sd1, 32'sd15, 32'sd0, 32'sd16, 32'sd2, 32'sd10, 32'sd1, 32'sd11, 32'sd3, 32'sd3, 32'sd10, 32'sd3, 32'sd0, 32'sd12, 32'sd8, 32'sd10, 32'sd9, 32'sd4, 32'sd0, 32'sd9, 32'sd8, 32'sd13, 32'sd5, 32'sd0, 32'sd1, 32'sd19, 32'sd0, 32'sd16, 32'sd0, 32'sd12, 32'sd7, 32'sd9, 32'sd0, 32'sd1, 32'sd1, 32'sd13, 32'sd0, 32'sd12, 32'sd4, 32'sd15, 32'sd1, 32'sd3, 32'sd2, 32'sd13, 32'sd1, 32'sd3, 32'sd7, 32'sd12, 32'sd0, 32'sd13, 32'sd0, 32'sd15, 32'sd0, 32'sd13, 32'sd5, 32'sd0, 32'sd2, 32'sd0, 32'sd1, 32'sd15, 32'sd0, 32'sd6, 32'sd8, 32'sd10, 32'sd8, 32'sd12, 32'sd6, 32'sd13, 32'sd1, 32'sd15, 32'sd6, 32'sd13, 32'sd5, 32'sd6, 32'sd0, 32'sd11, 32'sd9, 32'sd10, 32'sd8, 32'sd3, 32'sd10, 32'sd4, 32'sd9, 32'sd5, 32'sd2, 32'sd13, 32'sd8, 32'sd12, 32'sd2, 32'sd7, 32'sd3, 32'sd11, 32'sd0, 32'sd3, 32'sd1, 32'sd11, 32'sd9, 32'sd9, 32'sd1, 32'sd6, 32'sd1, 32'sd8, 32'sd2, 32'sd11, 32'sd7, 32'sd11, 32'sd5, 32'sd11, 32'sd5, 32'sd4, 32'sd2, 32'sd7, 32'sd9, 32'sd2, 32'sd8, 32'sd3, 32'sd8, 32'sd0, 32'sd6, 32'sd0, 32'sd20, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd1, 32'sd5, 32'sd4, 32'sd8, 32'sd6, 32'sd2, 32'sd11, 32'sd2, 32'sd5, 32'sd9, 32'sd8, 32'sd6, 32'sd10, 32'sd0, 32'sd18, 32'sd2, 32'sd3, 32'sd2, 32'sd13, 32'sd6, 32'sd9, 32'sd7, 32'sd18, 32'sd9, 32'sd6, 32'sd0, 32'sd13, 32'sd0, 32'sd13, 32'sd5, 32'sd11, 32'sd4, 32'sd6, 32'sd0, 32'sd12, 32'sd0, 32'sd12, 32'sd5, 32'sd5, 32'sd5, 32'sd3, 32'sd7, 32'sd13, 32'sd2, 32'sd19, 32'sd1, 32'sd5, 32'sd0, 32'sd2, 32'sd5, 32'sd1, 32'sd3, 32'sd8, 32'sd6, 32'sd10, 32'sd1, 32'sd8, 32'sd3, 32'sd5, 32'sd4, 32'sd6, 32'sd7, 32'sd0, 32'sd0, 32'sd3, 32'sd2, 32'sd7, 32'sd5, 32'sd10, 32'sd9, 32'sd18, 32'sd4, 32'sd10, 32'sd9, 32'sd11, 32'sd7, 32'sd4, 32'sd2, 32'sd13, 32'sd7, 32'sd3, 32'sd1, 32'sd8, 32'sd3, 32'sd5, 32'sd8, 32'sd9, 32'sd0, 32'sd6, 32'sd0, 32'sd13, 32'sd5, 32'sd1, 32'sd9, 32'sd9, 32'sd5, 32'sd4, 32'sd0, 32'sd16, 32'sd9, 32'sd8, 32'sd8, 32'sd10, 32'sd7, 32'sd5, 32'sd2, 32'sd18, 32'sd1, 32'sd6, 32'sd9, 32'sd10, 32'sd6, 32'sd8, 32'sd1, 32'sd9, 32'sd6, 32'sd17, 32'sd2, 32'sd7, 32'sd1, 32'sd1, 32'sd9, 32'sd3, 32'sd16, 32'sd0, 32'sd16, 32'sd0, 32'sd8, 32'sd5, 32'sd4, 32'sd0, 32'sd6, 32'sd0, 32'sd20, 32'sd8, 32'sd6, 32'sd0, 32'sd6, 32'sd0, 32'sd20, 32'sd0, 32'sd15, 32'sd0, 32'sd13, 32'sd5, 32'sd5, 32'sd3, 32'sd6, 32'sd6, 32'sd10, 32'sd1, 32'sd11, 32'sd5, 32'sd12, 32'sd5, 32'sd13, 32'sd0, 32'sd8, 32'sd1, 32'sd2, 32'sd2, 32'sd17, 32'sd1, 32'sd7, 32'sd0, 32'sd15, 32'sd1, 32'sd9, 32'sd0, 32'sd16, 32'sd4, 32'sd7, 32'sd9, 32'sd12, 32'sd8, 32'sd15, 32'sd3, 32'sd15, 32'sd1, 32'sd15, 32'sd6, 32'sd10, 32'sd6, 32'sd11, 32'sd6, 32'sd11, 32'sd9, 32'sd3, 32'sd2, 32'sd3, 32'sd3, 32'sd4, 32'sd0, 32'sd10, 32'sd0, 32'sd5, 32'sd8, 32'sd11, 32'sd5, 32'sd5, 32'sd10, 32'sd10, 32'sd7, 32'sd1, 32'sd0, 32'sd12, 32'sd2, 32'sd12, 32'sd1, 32'sd12, 32'sd0, 32'sd5, 32'sd6, 32'sd14, 32'sd5, 32'sd9, 32'sd1, 32'sd8, 32'sd3, 32'sd12, 32'sd0, 32'sd8, 32'sd4, 32'sd12, 32'sd9, 32'sd9, 32'sd1, 32'sd8, 32'sd3, 32'sd7, 32'sd10, 32'sd10, 32'sd3, 32'sd12, 32'sd3, 32'sd10, 32'sd5, 32'sd7, 32'sd6, 32'sd12, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd1, 32'sd9, 32'sd2, 32'sd5, 32'sd4, 32'sd2, 32'sd7, 32'sd0, 32'sd2, 32'sd3, 32'sd6, 32'sd9, 32'sd15, 32'sd8, 32'sd3, 32'sd2, 32'sd19, 32'sd1, 32'sd14, 32'sd4, 32'sd14, 32'sd6, 32'sd14, 32'sd4, 32'sd0, 32'sd1, 32'sd20, 32'sd0, 32'sd8, 32'sd7, 32'sd16, 32'sd5, 32'sd11, 32'sd10, 32'sd10, 32'sd7, 32'sd14, 32'sd5, 32'sd12, 32'sd6, 32'sd11, 32'sd1, 32'sd15, 32'sd9, 32'sd10, 32'sd3, 32'sd16, 32'sd7, 32'sd15, 32'sd0, 32'sd13, 32'sd2, 32'sd5, 32'sd1, 32'sd5, 32'sd1, 32'sd14, 32'sd4, 32'sd14, 32'sd4, 32'sd18, 32'sd1, 32'sd2, 32'sd0, 32'sd12, 32'sd3, 32'sd16, 32'sd3, 32'sd9, 32'sd9, 32'sd15, 32'sd7, 32'sd17, 32'sd3, 32'sd3, 32'sd0, 32'sd2, 32'sd0, 32'sd13, 32'sd5, 32'sd5, 32'sd5, 32'sd18, 32'sd0, 32'sd3, 32'sd2, 32'sd2, 32'sd5, 32'sd6, 32'sd6, 32'sd13, 32'sd5, 32'sd6, 32'sd0, 32'sd18, 32'sd0, 32'sd12, 32'sd6, 32'sd0, 32'sd3, 32'sd9, 32'sd5, 32'sd4, 32'sd10, 32'sd8, 32'sd2, 32'sd8, 32'sd0, 32'sd18, 32'sd0, 32'sd9, 32'sd1, 32'sd2, 32'sd7, 32'sd8, 32'sd4, 32'sd10, 32'sd2, 32'sd15, 32'sd3, 32'sd15, 32'sd4, 32'sd15, 32'sd0, 32'sd15, 32'sd0, 32'sd10, 32'sd1, 32'sd7, 32'sd10, 32'sd8, 32'sd3, 32'sd7, 32'sd0, 32'sd10, 32'sd7, 32'sd5, 32'sd5, 32'sd6, 32'sd3, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd10, 32'sd4, 32'sd0, 32'sd9, 32'sd3, 32'sd6, 32'sd11, 32'sd5, 32'sd4, 32'sd2, 32'sd7, 32'sd1, 32'sd13, 32'sd5, 32'sd11, 32'sd6, 32'sd3, 32'sd0, 32'sd10, 32'sd6, 32'sd6, 32'sd0, 32'sd18, 32'sd0, 32'sd11, 32'sd0, 32'sd2, 32'sd1, 32'sd18, 32'sd0, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd7, 32'sd15, 32'sd3, 32'sd15, 32'sd0, 32'sd15, 32'sd0, 32'sd5, 32'sd0, 32'sd9, 32'sd3, 32'sd9, 32'sd5, 32'sd9, 32'sd8, 32'sd10, 32'sd5, 32'sd9, 32'sd7, 32'sd11, 32'sd9, 32'sd6, 32'sd1, 32'sd16, 32'sd0, 32'sd8, 32'sd0, 32'sd3, 32'sd0, 32'sd6, 32'sd0, 32'sd14, 32'sd1, 32'sd13, 32'sd4, 32'sd12, 32'sd2, 32'sd16, 32'sd3, 32'sd14, 32'sd8, 32'sd9, 32'sd0, 32'sd4, 32'sd5, 32'sd15, 32'sd0, 32'sd8, 32'sd1, 32'sd14, 32'sd4, 32'sd16, 32'sd3, 32'sd18, 32'sd1, 32'sd11, 32'sd0, 32'sd15, 32'sd7, 32'sd22, 32'sd0, 32'sd18, 32'sd0, 32'sd3, 32'sd6, 32'sd7, 32'sd2, 32'sd4, 32'sd9, 32'sd4, 32'sd3, 32'sd18, 32'sd2, 32'sd4, 32'sd7, 32'sd7, 32'sd6, 32'sd12, 32'sd0, 32'sd8, 32'sd2, 32'sd13, 32'sd5, 32'sd9, 32'sd5, 32'sd3, 32'sd2, 32'sd11, 32'sd3, 32'sd9, 32'sd1, 32'sd15, 32'sd1, 32'sd9, 32'sd6, 32'sd10, 32'sd7, 32'sd10, 32'sd4, 32'sd0, 
                                                    32'sd3, 32'sd19, 32'sd0, 32'sd17, 32'sd1, 32'sd18, 32'sd0, 32'sd3, 32'sd2, 32'sd9, 32'sd5, 32'sd10, 32'sd8, 32'sd7, 32'sd9, 32'sd5, 32'sd8, 32'sd8, 32'sd6, 32'sd14, 32'sd6, 32'sd8, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd7, 32'sd6, 32'sd14, 32'sd4, 32'sd2, 32'sd6, 32'sd9, 32'sd7, 32'sd6, 32'sd5, 32'sd18, 32'sd0, 32'sd18, 32'sd2, 32'sd5, 32'sd11, 32'sd15, 32'sd7, 32'sd7, 32'sd10, 32'sd10, 32'sd2, 32'sd14, 32'sd8, 32'sd14, 32'sd3, 32'sd14, 32'sd1, 32'sd3, 32'sd1, 32'sd18, 32'sd0, 32'sd5, 32'sd6, 32'sd14, 32'sd4, 32'sd15, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd1, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd10, 32'sd10, 32'sd6, 32'sd11, 32'sd9, 32'sd2, 32'sd1, 32'sd13, 32'sd6, 32'sd10, 32'sd6, 32'sd14, 32'sd6, 32'sd9, 32'sd8, 32'sd17, 32'sd1, 32'sd14, 32'sd7, 32'sd3, 32'sd1, 32'sd14, 32'sd0, 32'sd12, 32'sd0, 32'sd10, 32'sd1, 32'sd15, 32'sd6, 32'sd6, 32'sd8, 32'sd14, 32'sd0, 32'sd10, 32'sd6, 32'sd7, 32'sd9, 32'sd10, 32'sd8, 32'sd7, 32'sd4, 32'sd17, 32'sd3, 32'sd10, 32'sd2, 32'sd3, 32'sd4, 32'sd15, 32'sd7, 32'sd15, 32'sd1, 32'sd11, 32'sd5, 32'sd10, 32'sd4, 32'sd0, 32'sd4, 32'sd10, 32'sd0, 32'sd6, 32'sd1, 32'sd18, 32'sd4, 32'sd6, 32'sd1, 32'sd1, 32'sd2, 32'sd12, 32'sd0, 32'sd10, 32'sd7, 32'sd9, 32'sd4, 32'sd6, 32'sd5, 32'sd10, 32'sd8, 32'sd9, 32'sd3, 32'sd4, 32'sd6, 32'sd8, 32'sd0, 32'sd11, 32'sd2, 32'sd8, 32'sd0, 32'sd0, 32'sd2, 32'sd4, 32'sd10, 32'sd7, 32'sd9, 32'sd17, 32'sd0, 32'sd16, 32'sd1, 32'sd12, 32'sd3, 32'sd12, 32'sd3, 32'sd12, 32'sd8, 32'sd10, 32'sd6, 32'sd13, 32'sd1, 32'sd7, 32'sd2, 32'sd0, 32'sd9, 32'sd0, 32'sd9, 32'sd2, 32'sd13, 32'sd4, 32'sd20, 32'sd8, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd13, 32'sd5, 32'sd13, 32'sd2, 32'sd9, 32'sd8, 32'sd12, 32'sd8, 32'sd8, 32'sd11, 32'sd9, 32'sd0, 32'sd9, 32'sd1, 32'sd12, 32'sd6, 32'sd13, 32'sd1, 32'sd9, 32'sd2, 32'sd15, 32'sd0, 32'sd9, 32'sd2, 32'sd15, 32'sd4, 32'sd17, 32'sd0, 32'sd15, 32'sd0, 32'sd9, 32'sd3, 32'sd16, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd5, 32'sd8, 32'sd4, 32'sd10, 32'sd8, 32'sd11, 32'sd4, 32'sd14, 32'sd2, 32'sd4, 32'sd8, 32'sd1, 32'sd7, 32'sd13, 32'sd8, 32'sd4, 32'sd3, 32'sd14, 32'sd8, 32'sd3, 32'sd4, 32'sd3, 32'sd9, 32'sd9, 32'sd7, 32'sd12, 32'sd6, 32'sd18, 32'sd3, 32'sd18, 32'sd0, 32'sd13, 32'sd5, 32'sd11, 32'sd3, 32'sd16, 32'sd5, 32'sd7, 32'sd1, 32'sd2, 32'sd3, 32'sd17, 32'sd5, 32'sd13, 32'sd0, 32'sd15, 32'sd1, 32'sd12, 32'sd1, 32'sd3, 32'sd6, 32'sd5, 32'sd9, 32'sd11, 32'sd4, 32'sd6, 32'sd5, 32'sd11, 32'sd5, 32'sd1, 32'sd7, 32'sd6, 32'sd6, 32'sd11, 32'sd5, 32'sd6, 32'sd0, 32'sd2, 32'sd0, 32'sd9, 32'sd9, 32'sd12, 32'sd0, 32'sd1, 32'sd3, 32'sd2, 32'sd5, 32'sd10, 32'sd8, 32'sd5, 32'sd6, 32'sd7, 32'sd5, 32'sd4, 32'sd0, 32'sd9, 32'sd9, 32'sd6, 32'sd9, 32'sd10, 32'sd5, 32'sd14, 32'sd5, 32'sd14, 32'sd0, 32'sd16, 32'sd4, 32'sd8, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd6, 32'sd10, 32'sd1, 32'sd0, 32'sd2, 32'sd2, 32'sd1, 32'sd10, 32'sd7, 32'sd9, 32'sd7, 32'sd3, 32'sd7, 32'sd3, 32'sd8, 32'sd3, 32'sd6, 32'sd1, 32'sd5, 32'sd8, 32'sd3, 32'sd0, 32'sd2, 32'sd4, 32'sd9, 32'sd9, 32'sd14, 32'sd7, 32'sd14, 32'sd4, 32'sd17, 32'sd1, 32'sd14, 32'sd0, 32'sd9, 32'sd3, 32'sd14, 32'sd4, 32'sd7, 32'sd7, 32'sd14, 32'sd10, 32'sd14, 32'sd5, 32'sd4, 32'sd9, 32'sd3, 32'sd4, 32'sd16, 32'sd4, 32'sd6, 32'sd10, 32'sd9, 32'sd6, 32'sd5, 32'sd3, 32'sd6, 32'sd0, 32'sd6, 32'sd0, 32'sd4, 32'sd0, 32'sd15, 32'sd0, 32'sd6, 32'sd3, 32'sd12, 32'sd6, 32'sd6, 32'sd9, 32'sd10, 32'sd7, 32'sd14, 32'sd2, 32'sd11, 32'sd1, 32'sd15, 32'sd1, 32'sd10, 32'sd4, 32'sd7, 32'sd10, 32'sd13, 32'sd3, 32'sd13, 32'sd5, 32'sd10, 32'sd7, 32'sd15, 32'sd5, 32'sd8, 32'sd7, 32'sd12, 32'sd6, 32'sd7, 32'sd6, 32'sd5, 32'sd3, 32'sd3, 32'sd0, 32'sd14, 32'sd0, 32'sd1, 32'sd1, 32'sd7, 32'sd9, 32'sd10, 32'sd2, 32'sd8, 32'sd0, 32'sd5, 32'sd2, 32'sd14, 32'sd3, 32'sd9, 32'sd4, 32'sd0, 32'sd7, 32'sd11, 32'sd0, 32'sd14, 32'sd2, 32'sd11, 32'sd7, 32'sd6, 32'sd4, 32'sd14, 32'sd4, 32'sd13, 32'sd8, 32'sd17, 32'sd4, 32'sd15, 32'sd3, 32'sd12, 32'sd0, 32'sd16, 32'sd2, 32'sd15, 32'sd0, 32'sd18, 32'sd0, 32'sd16, 32'sd5, 32'sd12, 32'sd0, 32'sd5, 32'sd0, 32'sd8, 32'sd5, 32'sd10, 32'sd6, 32'sd6, 32'sd3, 32'sd12, 32'sd0, 32'sd0, 32'sd5, 32'sd10, 32'sd9, 32'sd8, 32'sd0, 32'sd16, 32'sd3, 32'sd6, 32'sd0, 32'sd14, 32'sd0, 32'sd2, 32'sd4, 32'sd12, 32'sd0, 32'sd6, 32'sd1, 32'sd11, 32'sd3, 32'sd15, 32'sd6, 32'sd9, 32'sd4, 32'sd7, 32'sd5, 32'sd11, 32'sd7, 32'sd8, 32'sd0, 32'sd10, 32'sd0, 32'sd20, 32'sd0, 32'sd12, 32'sd1, 32'sd5, 32'sd1, 32'sd6, 32'sd5, 32'sd11, 32'sd1, 32'sd11, 32'sd0, 32'sd3, 32'sd1, 32'sd0, 32'sd1, 32'sd11, 32'sd4, 32'sd12, 32'sd4, 32'sd13, 32'sd1, 32'sd9, 32'sd0, 32'sd6, 32'sd6, 32'sd10, 32'sd6, 32'sd13, 32'sd2, 32'sd11, 32'sd1, 32'sd1, 32'sd0, 32'sd13, 32'sd5, 32'sd18, 32'sd0, 32'sd11, 32'sd0, 32'sd12, 32'sd1, 32'sd7, 32'sd8, 32'sd6, 32'sd2, 32'sd14, 32'sd3, 32'sd15, 32'sd5, 32'sd11, 32'sd7, 32'sd11, 32'sd9, 32'sd4, 32'sd9, 32'sd17, 32'sd1, 32'sd7, 32'sd6, 32'sd9, 32'sd1, 32'sd19, 32'sd0, 32'sd3, 32'sd1, 32'sd2, 32'sd4, 32'sd6, 32'sd4, 32'sd15, 32'sd3, 32'sd8, 32'sd3, 32'sd15, 32'sd3, 32'sd5, 32'sd1, 32'sd14, 32'sd0, 32'sd15, 32'sd3, 32'sd9, 32'sd1, 32'sd13, 32'sd1, 32'sd6, 32'sd8, 32'sd0, 32'sd0, 32'sd4, 32'sd1, 32'sd14, 32'sd1, 32'sd10, 32'sd6, 32'sd10, 32'sd7, 32'sd14, 32'sd6, 32'sd8, 32'sd3, 32'sd5, 32'sd0, 32'sd9, 32'sd4, 32'sd10, 32'sd8, 32'sd7, 32'sd8, 32'sd11, 32'sd7, 32'sd4, 32'sd0, 32'sd7, 32'sd1, 32'sd11, 32'sd6, 32'sd7, 32'sd7, 32'sd9, 32'sd0, 32'sd7, 32'sd1, 32'sd9, 32'sd0, 32'sd1, 32'sd1, 32'sd9, 32'sd3, 32'sd9, 32'sd9, 32'sd16, 32'sd2, 32'sd13, 32'sd1, 32'sd14, 32'sd3, 32'sd13, 32'sd7, 32'sd4, 32'sd9, 32'sd7, 32'sd0, 32'sd15, 32'sd1, 32'sd14, 32'sd4, 32'sd15, 32'sd3, 32'sd0, 32'sd7, 32'sd1, 32'sd1, 32'sd6, 32'sd1, 32'sd15, 32'sd3, 32'sd4, 32'sd0, 32'sd6, 32'sd4, 32'sd6, 32'sd0, 32'sd3, 32'sd4, 32'sd20, 32'sd0, 
                                                    32'sd11, 32'sd6, 32'sd11, 32'sd1, 32'sd11, 32'sd1, 32'sd11, 32'sd0, 32'sd3, 32'sd7, 32'sd17, 32'sd5, 32'sd16, 32'sd0, 32'sd6, 32'sd0, 32'sd3, 32'sd2, 32'sd10, 32'sd10, 32'sd11, 32'sd9, 32'sd5, 32'sd6, 32'sd10, 32'sd0, 32'sd6, 32'sd4, 32'sd14, 32'sd0, 32'sd1, 32'sd8, 32'sd13, 32'sd10, 32'sd7, 32'sd8, 32'sd7, 32'sd2, 32'sd11, 32'sd7, 32'sd13, 32'sd0, 32'sd12, 32'sd8, 32'sd12, 32'sd6, 32'sd14, 32'sd0, 32'sd14, 32'sd0, 32'sd4, 32'sd1, 32'sd4, 32'sd0, 32'sd3, 32'sd9, 32'sd0, 32'sd6, 32'sd2, 32'sd18, 32'sd0, 32'sd11, 32'sd9, 32'sd7, 32'sd1, 32'sd18, 32'sd5, 32'sd18, 32'sd0, 32'sd9, 32'sd2, 32'sd10, 32'sd5, 32'sd9, 32'sd7, 32'sd10, 32'sd4, 32'sd6, 32'sd0, 32'sd3, 32'sd9, 32'sd6, 32'sd2, 32'sd19, 32'sd0, 32'sd5, 32'sd5, 32'sd1, 32'sd8, 32'sd6, 32'sd9, 32'sd2, 32'sd5, 32'sd8, 32'sd9, 32'sd14, 32'sd2, 32'sd10, 32'sd1, 32'sd11, 32'sd4, 32'sd6, 32'sd5, 32'sd9, 32'sd7, 32'sd7, 32'sd2, 32'sd5, 32'sd7, 32'sd0, 32'sd0, 32'sd16, 32'sd5, 32'sd5, 32'sd0, 32'sd11, 32'sd0, 32'sd4, 32'sd2, 32'sd3, 32'sd2, 32'sd6, 32'sd0, 32'sd3, 32'sd0, 32'sd5, 32'sd1, 32'sd19, 32'sd3, 32'sd19, 32'sd7, 32'sd9, 32'sd0, 32'sd15, 32'sd1, 32'sd9, 32'sd7, 32'sd9, 32'sd7, 32'sd9, 32'sd7, 32'sd9, 32'sd10, 32'sd5, 32'sd0, 32'sd9, 32'sd2, 32'sd15, 32'sd1, 32'sd6, 32'sd0, 32'sd6, 32'sd0, 32'sd13, 32'sd2, 32'sd13, 32'sd5, 32'sd11, 32'sd7, 32'sd10, 32'sd3, 32'sd14, 32'sd4, 32'sd4, 32'sd5, 32'sd7, 32'sd2, 32'sd10, 32'sd3, 32'sd16, 32'sd0, 32'sd0, 32'sd4, 32'sd10, 32'sd7, 32'sd13, 32'sd3, 32'sd16, 32'sd2, 32'sd3, 32'sd4, 32'sd4, 32'sd3, 32'sd8, 32'sd2, 32'sd14, 32'sd7, 32'sd4, 32'sd0, 32'sd10, 32'sd5, 32'sd0, 32'sd0, 32'sd3, 32'sd9, 32'sd0, 32'sd6, 32'sd8, 32'sd2, 32'sd12, 32'sd5, 32'sd14, 32'sd5, 32'sd6, 32'sd7, 32'sd11, 32'sd7, 32'sd13, 32'sd0, 32'sd1, 32'sd6, 32'sd10, 32'sd3, 32'sd0, 32'sd0, 32'sd3, 32'sd7, 32'sd10, 32'sd8, 32'sd12, 32'sd6, 32'sd16, 32'sd2, 32'sd10, 32'sd8, 32'sd14, 32'sd0, 32'sd11, 32'sd3, 32'sd10, 32'sd0, 32'sd19, 32'sd4, 32'sd4, 32'sd0, 32'sd6, 32'sd19, 32'sd0, 32'sd18, 32'sd0, 32'sd5, 32'sd10, 32'sd9, 32'sd0, 32'sd7, 32'sd1, 32'sd8, 32'sd0, 32'sd13, 32'sd10, 32'sd13, 32'sd7, 32'sd4, 32'sd0, 32'sd0, 32'sd6, 32'sd7, 32'sd0, 32'sd13, 32'sd3, 32'sd12, 32'sd2, 32'sd9, 32'sd6, 32'sd14, 32'sd5, 32'sd10, 32'sd6, 32'sd14, 32'sd4, 32'sd14, 32'sd0, 32'sd13, 32'sd2, 32'sd6, 32'sd0, 32'sd19, 32'sd1, 32'sd15, 32'sd3, 32'sd11, 32'sd7, 32'sd14, 32'sd3, 32'sd20, 32'sd7, 32'sd7, 32'sd2, 32'sd15, 32'sd7, 32'sd13, 32'sd5, 32'sd3, 32'sd5, 32'sd9, 32'sd3, 32'sd19, 32'sd0, 32'sd20, 32'sd0, 32'sd7, 32'sd4, 32'sd10, 32'sd0, 32'sd7, 32'sd0, 32'sd13, 32'sd1, 32'sd7, 32'sd0, 32'sd6, 32'sd8, 32'sd7, 32'sd1, 32'sd16, 32'sd5, 32'sd7, 32'sd4, 32'sd6, 32'sd9, 32'sd15, 32'sd6, 32'sd12, 32'sd7, 32'sd6, 32'sd10, 32'sd10, 32'sd3, 32'sd4, 32'sd2, 32'sd13, 32'sd7, 32'sd1, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd3, 32'sd13, 32'sd2, 32'sd10, 32'sd6, 32'sd2, 32'sd2, 32'sd10, 32'sd8, 32'sd13, 32'sd3, 32'sd3, 32'sd2, 32'sd14, 32'sd3, 32'sd5, 32'sd2, 32'sd17, 32'sd2, 32'sd0, 32'sd7, 32'sd15, 32'sd5, 32'sd11, 32'sd6, 32'sd11, 32'sd5, 32'sd15, 32'sd4, 32'sd12, 32'sd6, 32'sd5, 32'sd9, 32'sd12, 32'sd4, 32'sd4, 32'sd5, 32'sd14, 32'sd9, 32'sd9, 32'sd9, 32'sd1, 32'sd2, 32'sd12, 32'sd6, 32'sd12, 32'sd8, 32'sd7, 32'sd0, 32'sd4, 32'sd2, 32'sd15, 32'sd0, 32'sd6, 32'sd6, 32'sd8, 32'sd1, 32'sd6, 32'sd7, 32'sd10, 32'sd3, 32'sd15, 32'sd1, 32'sd15, 32'sd10, 32'sd15, 32'sd6, 32'sd15, 32'sd6, 32'sd16, 32'sd2, 32'sd2, 32'sd6, 32'sd9, 32'sd2, 32'sd16, 32'sd0, 32'sd15, 32'sd8, 32'sd15, 32'sd0, 32'sd12, 32'sd3, 32'sd13, 32'sd0, 32'sd10, 32'sd7, 32'sd4, 32'sd0, 32'sd6, 32'sd3, 32'sd9, 32'sd5, 32'sd5, 32'sd3, 32'sd5, 32'sd6, 32'sd0, 32'sd2, 32'sd8, 32'sd18, 32'sd0, 32'sd4, 32'sd6, 32'sd4, 32'sd4, 32'sd7, 32'sd0, 32'sd13, 32'sd5, 32'sd3, 32'sd0, 32'sd14, 32'sd0, 32'sd14, 32'sd0, 32'sd6, 32'sd0, 32'sd14, 32'sd6, 32'sd15, 32'sd8, 32'sd4, 32'sd5, 32'sd7, 32'sd10, 32'sd5, 32'sd1, 32'sd18, 32'sd0, 32'sd13, 32'sd0, 32'sd12, 32'sd7, 32'sd14, 32'sd0, 32'sd14, 32'sd2, 32'sd14, 32'sd1, 32'sd3, 32'sd5, 32'sd5, 32'sd8, 32'sd9, 32'sd6, 32'sd5, 32'sd8, 32'sd6, 32'sd3, 32'sd13, 32'sd3, 32'sd12, 32'sd7, 32'sd13, 32'sd7, 32'sd11, 32'sd7, 32'sd5, 32'sd8, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd3, 32'sd12, 32'sd8, 32'sd10, 32'sd5, 32'sd2, 32'sd6, 32'sd8, 32'sd9, 32'sd15, 32'sd1, 32'sd11, 32'sd5, 32'sd6, 32'sd1, 32'sd2, 32'sd7, 32'sd10, 32'sd3, 32'sd7, 32'sd7, 32'sd9, 32'sd1, 32'sd13, 32'sd3, 32'sd8, 32'sd6, 32'sd4, 32'sd0, 32'sd3, 32'sd2, 32'sd16, 32'sd4, 32'sd16, 32'sd1, 32'sd15, 32'sd3, 32'sd18, 32'sd0, 32'sd4, 32'sd2, 32'sd17, 32'sd1, 32'sd8, 32'sd0, 32'sd11, 32'sd0, 32'sd19, 32'sd2, 32'sd3, 32'sd4, 32'sd7, 32'sd3, 32'sd8, 32'sd4, 32'sd10, 32'sd3, 32'sd15, 32'sd0, 32'sd6, 32'sd9, 32'sd12, 32'sd8, 32'sd16, 32'sd8, 32'sd6, 32'sd0, 32'sd17, 32'sd0, 32'sd9, 32'sd1, 32'sd7, 32'sd7, 32'sd7, 32'sd3, 32'sd9, 32'sd3, 32'sd6, 32'sd1, 32'sd16, 32'sd0, 32'sd0, 32'sd3, 32'sd4, 32'sd0, 32'sd20, 32'sd1, 32'sd18, 32'sd0, 32'sd8, 32'sd4, 32'sd7, 32'sd6, 32'sd7, 32'sd9, 32'sd8, 32'sd8, 32'sd8, 32'sd4, 32'sd7, 32'sd0, 32'sd12, 32'sd4, 32'sd8, 32'sd9, 32'sd14, 32'sd7, 32'sd4, 32'sd10, 32'sd12, 32'sd0, 32'sd16, 32'sd5, 32'sd10, 32'sd2, 32'sd2, 32'sd7, 32'sd3, 32'sd2, 32'sd15, 32'sd2, 32'sd10, 32'sd4, 32'sd15, 32'sd0, 32'sd18, 32'sd0, 32'sd15, 32'sd3, 32'sd12, 32'sd0, 32'sd11, 32'sd9, 32'sd12, 32'sd3, 32'sd5, 32'sd0, 32'sd8, 32'sd6, 32'sd14, 32'sd9, 32'sd6, 32'sd6, 32'sd1, 32'sd12, 32'sd3, 32'sd9, 32'sd4, 32'sd11, 32'sd3, 32'sd5, 32'sd4, 32'sd9, 32'sd8, 32'sd16, 32'sd3, 32'sd6, 32'sd8, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd2, 32'sd9, 32'sd9, 32'sd9, 32'sd5, 32'sd2, 32'sd6, 32'sd5, 32'sd18, 32'sd0, 32'sd10, 32'sd6, 32'sd3, 32'sd5, 32'sd17, 32'sd0, 32'sd9, 32'sd5, 32'sd11, 32'sd0, 32'sd6, 32'sd4, 32'sd9, 32'sd5, 32'sd6, 32'sd7, 32'sd11, 
                                                    32'sd1, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd19, 32'sd4, 32'sd19, 32'sd1, 32'sd3, 32'sd0, 32'sd12, 32'sd7, 32'sd12, 32'sd2, 32'sd14, 32'sd0, 32'sd15, 32'sd0, 32'sd14, 32'sd0, 32'sd5, 32'sd0, 32'sd3, 32'sd5, 32'sd4, 32'sd3, 32'sd4, 32'sd4, 32'sd16, 32'sd6, 32'sd13, 32'sd3, 32'sd12, 32'sd5, 32'sd10, 32'sd6, 32'sd6, 32'sd0, 32'sd12, 32'sd0, 32'sd12, 32'sd9, 32'sd6, 32'sd0, 32'sd2, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd4, 32'sd12, 32'sd6, 32'sd15, 32'sd3, 32'sd6, 32'sd5, 32'sd12, 32'sd0, 32'sd11, 32'sd10, 32'sd9, 32'sd1, 32'sd6, 32'sd1, 32'sd7, 32'sd0, 32'sd10, 32'sd9, 32'sd10, 32'sd8, 32'sd9, 32'sd1, 32'sd0, 32'sd6, 32'sd8, 32'sd5, 32'sd4, 32'sd4, 32'sd8, 32'sd1, 32'sd10, 32'sd1, 32'sd0, 32'sd1, 32'sd5, 32'sd0, 32'sd9, 32'sd1, 32'sd8, 32'sd8, 32'sd5, 32'sd9, 32'sd6, 32'sd2, 32'sd10, 32'sd7, 32'sd14, 32'sd8, 32'sd9, 32'sd3, 32'sd5, 32'sd4, 32'sd6, 32'sd9, 32'sd12, 32'sd6, 32'sd9, 32'sd5, 32'sd5, 32'sd9, 32'sd11, 32'sd2, 32'sd15, 32'sd3, 32'sd3, 32'sd5, 32'sd16, 32'sd0, 32'sd13, 32'sd1, 32'sd15, 32'sd5, 32'sd6, 32'sd2, 32'sd14, 32'sd10, 32'sd13, 32'sd3, 32'sd13, 32'sd3, 32'sd11, 32'sd0, 32'sd0, 32'sd6, 32'sd18, 32'sd0, 32'sd15, 32'sd1, 32'sd15, 32'sd0, 32'sd3, 32'sd0, 32'sd15, 32'sd0, 32'sd12, 32'sd3, 32'sd16, 32'sd0, 32'sd9}

localparam logic [2912:0][31:0] rectangle1_ys = {32'sd4, 32'sd4, 32'sd9, 32'sd18, 32'sd5, 32'sd5, 32'sd8, 32'sd14, 32'sd0, 32'sd6, 32'sd4, 32'sd8, 32'sd2, 32'sd9, 32'sd6, 32'sd0, 32'sd11, 32'sd5, 32'sd8, 32'sd5, 32'sd0, 32'sd6, 32'sd6, 32'sd18, 32'sd7, 32'sd3, 32'sd8, 32'sd6, 32'sd5, 32'sd6, 32'sd21, 32'sd6, 32'sd1, 32'sd1, 32'sd8, 32'sd6, 32'sd12, 32'sd1, 32'sd13, 32'sd1, 32'sd2, 32'sd5, 32'sd4, 32'sd3, 32'sd1, 32'sd6, 32'sd1, 32'sd1, 32'sd5, 32'sd10, 32'sd13, 32'sd4, 32'sd4, 32'sd5, 32'sd1, 32'sd10, 32'sd17, 32'sd3, 32'sd3, 32'sd1, 32'sd7, 32'sd7, 32'sd12, 32'sd6, 32'sd7, 32'sd15, 32'sd17, 32'sd4, 32'sd1, 32'sd0, 32'sd5, 32'sd8, 32'sd14, 32'sd15, 32'sd15, 32'sd6, 32'sd5, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd6, 32'sd6, 32'sd8, 32'sd0, 32'sd0, 32'sd7, 32'sd6, 32'sd20, 32'sd6, 32'sd13, 32'sd6, 32'sd6, 32'sd12, 32'sd22, 32'sd7, 32'sd7, 32'sd6, 32'sd14, 32'sd18, 32'sd1, 32'sd16, 32'sd4, 32'sd4, 32'sd4, 32'sd16, 32'sd12, 32'sd0, 32'sd10, 32'sd8, 32'sd8, 32'sd0, 32'sd0, 32'sd14, 32'sd16, 32'sd8, 32'sd19, 32'sd10, 32'sd9, 32'sd0, 32'sd6, 32'sd5, 32'sd5, 32'sd14, 32'sd13, 32'sd16, 32'sd0, 32'sd6, 32'sd1, 32'sd2, 32'sd8, 32'sd9, 32'sd12, 32'sd16, 32'sd16, 32'sd1, 32'sd2, 32'sd8, 32'sd5, 32'sd17, 32'sd7, 32'sd1, 32'sd5, 32'sd1, 32'sd1, 32'sd0, 32'sd0, 32'sd7, 32'sd10, 32'sd9, 32'sd15, 32'sd7, 32'sd6, 32'sd8, 32'sd8, 32'sd6, 32'sd7, 32'sd14, 32'sd10, 32'sd12, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd18, 32'sd3, 32'sd3, 32'sd10, 32'sd10, 32'sd11, 32'sd11, 32'sd11, 32'sd10, 32'sd13, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd1, 32'sd1, 32'sd6, 32'sd14, 32'sd14, 32'sd18, 32'sd4, 32'sd17, 32'sd2, 32'sd8, 32'sd5, 32'sd5, 32'sd4, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd22, 32'sd0, 32'sd6, 32'sd1, 32'sd5, 32'sd1, 32'sd2, 32'sd8, 32'sd12, 32'sd12, 32'sd7, 32'sd1, 32'sd2, 32'sd4, 32'sd1, 32'sd15, 32'sd5, 32'sd5, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd6, 32'sd7, 32'sd17, 32'sd18, 32'sd18, 32'sd20, 32'sd15, 32'sd4, 32'sd6, 32'sd14, 32'sd9, 32'sd6, 32'sd6, 32'sd10, 32'sd16, 32'sd6, 32'sd0, 32'sd0, 32'sd7, 32'sd20, 32'sd5, 32'sd2, 32'sd1, 32'sd0, 32'sd0, 32'sd21, 32'sd7, 32'sd7, 32'sd8, 32'sd15, 32'sd15, 32'sd0, 32'sd6, 32'sd1, 32'sd2, 32'sd14, 32'sd6, 32'sd2, 32'sd4, 32'sd17, 32'sd7, 32'sd1, 32'sd13, 32'sd13, 32'sd6, 32'sd12, 32'sd1, 32'sd0, 32'sd2, 32'sd2, 32'sd18, 32'sd6, 32'sd7, 32'sd3, 32'sd4, 32'sd1, 32'sd2, 32'sd3, 32'sd3, 32'sd0, 32'sd8, 32'sd8, 32'sd14, 32'sd14, 32'sd10, 32'sd0, 32'sd1, 32'sd6, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd9, 32'sd8, 32'sd12, 32'sd12, 32'sd12, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd2, 32'sd10, 32'sd14, 32'sd13, 32'sd5, 32'sd17, 32'sd18, 32'sd0, 32'sd4, 32'sd4, 32'sd3, 32'sd1, 32'sd16, 32'sd3, 32'sd5, 32'sd2, 32'sd14, 32'sd21, 32'sd14, 32'sd2, 32'sd4, 32'sd6, 32'sd8, 32'sd14, 32'sd6, 32'sd6, 32'sd7, 32'sd3, 32'sd12, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd2, 32'sd18, 32'sd2, 32'sd2, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd6, 32'sd12, 32'sd5, 32'sd8, 32'sd6, 32'sd12, 32'sd12, 32'sd1, 32'sd1, 32'sd9, 32'sd21, 32'sd13, 32'sd13, 32'sd6, 32'sd0, 32'sd7, 32'sd4, 32'sd0, 32'sd0, 32'sd12, 32'sd12, 32'sd12, 32'sd12, 32'sd14, 32'sd13, 32'sd15, 32'sd0, 32'sd1, 32'sd1, 32'sd14, 32'sd3, 32'sd1, 32'sd0, 32'sd6, 32'sd10, 32'sd15, 32'sd1, 32'sd9, 32'sd0, 32'sd15, 32'sd15, 32'sd7, 32'sd12, 32'sd8, 32'sd14, 32'sd10, 32'sd3, 32'sd17, 32'sd13, 32'sd0, 32'sd3, 32'sd5, 32'sd7, 32'sd6, 32'sd8, 32'sd15, 32'sd1, 32'sd8, 32'sd5, 32'sd2, 32'sd7, 32'sd7, 32'sd6, 32'sd1, 32'sd1, 32'sd18, 32'sd4, 32'sd16, 32'sd7, 32'sd7, 32'sd2, 32'sd20, 32'sd12, 32'sd2, 32'sd0, 32'sd0, 32'sd15, 32'sd8, 32'sd3, 32'sd5, 32'sd4, 32'sd6, 32'sd4, 32'sd4, 32'sd4, 32'sd22, 32'sd14, 32'sd14, 32'sd11, 32'sd11, 32'sd9, 32'sd12, 32'sd0, 32'sd0, 32'sd17, 32'sd17, 32'sd6, 32'sd6, 32'sd4, 32'sd0, 32'sd0, 32'sd15, 32'sd8, 32'sd12, 32'sd2, 32'sd20, 32'sd0, 32'sd13, 32'sd10, 32'sd3, 32'sd5, 32'sd7, 32'sd0, 32'sd0, 32'sd1, 32'sd17, 32'sd15, 32'sd15, 32'sd16, 32'sd13, 32'sd0, 32'sd4, 32'sd5, 32'sd4, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd5, 32'sd13, 32'sd0, 32'sd7, 32'sd2, 32'sd2, 32'sd2, 32'sd6, 32'sd5, 32'sd6, 32'sd0, 32'sd3, 32'sd7, 32'sd7, 32'sd7, 32'sd6, 32'sd14, 32'sd0, 32'sd2, 32'sd4, 32'sd3, 32'sd4, 32'sd0, 32'sd6, 32'sd0, 32'sd10, 32'sd21, 32'sd6, 32'sd5, 32'sd2, 32'sd7, 32'sd7, 32'sd17, 32'sd18, 32'sd6, 32'sd18, 32'sd18, 32'sd9, 32'sd9, 32'sd3, 32'sd17, 32'sd15, 32'sd17, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd11, 32'sd0, 32'sd0, 32'sd8, 32'sd12, 32'sd0, 32'sd6, 32'sd0, 32'sd2, 32'sd7, 32'sd6, 32'sd1, 32'sd4, 32'sd3, 32'sd1, 32'sd0, 32'sd0, 32'sd13, 32'sd5, 32'sd1, 32'sd2, 32'sd10, 32'sd4, 32'sd10, 32'sd10, 32'sd14, 32'sd7, 32'sd1, 32'sd1, 32'sd5, 32'sd9, 32'sd16, 32'sd12, 32'sd14, 32'sd13, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd1, 32'sd1, 32'sd15, 32'sd9, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd17, 32'sd5, 32'sd2, 32'sd2, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd6, 32'sd7, 32'sd6, 32'sd6, 32'sd3, 32'sd0, 32'sd9, 32'sd7, 32'sd6, 32'sd0, 32'sd14, 32'sd14, 32'sd12, 32'sd2, 32'sd16, 32'sd16, 32'sd0, 32'sd0, 32'sd8, 32'sd5, 32'sd13, 32'sd14, 32'sd6, 32'sd0, 32'sd1, 32'sd6, 32'sd0, 32'sd11, 32'sd20, 32'sd11, 32'sd12, 32'sd11, 32'sd11, 32'sd4, 32'sd15, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd18, 32'sd7, 32'sd14, 32'sd2, 32'sd3, 32'sd6, 32'sd8, 32'sd4, 32'sd8, 32'sd2, 32'sd16, 32'sd0, 32'sd2, 32'sd11, 32'sd3, 32'sd16, 32'sd17, 32'sd13, 32'sd9, 32'sd7, 32'sd8, 32'sd2, 32'sd17, 32'sd18, 32'sd3, 32'sd6, 32'sd0, 32'sd0, 32'sd10, 32'sd11, 32'sd5, 32'sd6, 32'sd5, 32'sd3, 32'sd21, 32'sd10, 32'sd4, 32'sd8, 32'sd9, 32'sd6, 32'sd6, 32'sd5, 32'sd4, 32'sd4, 32'sd10, 32'sd10, 32'sd2, 32'sd2, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd18, 32'sd18, 32'sd2, 32'sd2, 32'sd5, 32'sd8, 32'sd7, 32'sd5, 32'sd14, 32'sd14, 32'sd11, 32'sd9, 32'sd6, 32'sd19, 32'sd5, 32'sd5, 32'sd4, 
                                                    32'sd6, 32'sd10, 32'sd7, 32'sd2, 32'sd18, 32'sd9, 32'sd2, 32'sd0, 32'sd3, 32'sd2, 32'sd5, 32'sd0, 32'sd3, 32'sd14, 32'sd9, 32'sd11, 32'sd5, 32'sd6, 32'sd6, 32'sd5, 32'sd5, 32'sd10, 32'sd10, 32'sd0, 32'sd3, 32'sd1, 32'sd7, 32'sd12, 32'sd6, 32'sd7, 32'sd18, 32'sd2, 32'sd3, 32'sd2, 32'sd0, 32'sd0, 32'sd5, 32'sd22, 32'sd10, 32'sd1, 32'sd0, 32'sd3, 32'sd15, 32'sd13, 32'sd8, 32'sd8, 32'sd2, 32'sd5, 32'sd8, 32'sd8, 32'sd6, 32'sd0, 32'sd9, 32'sd0, 32'sd5, 32'sd5, 32'sd5, 32'sd4, 32'sd16, 32'sd16, 32'sd9, 32'sd13, 32'sd10, 32'sd9, 32'sd0, 32'sd11, 32'sd5, 32'sd5, 32'sd6, 32'sd6, 32'sd5, 32'sd6, 32'sd13, 32'sd5, 32'sd2, 32'sd15, 32'sd17, 32'sd13, 32'sd10, 32'sd6, 32'sd14, 32'sd12, 32'sd10, 32'sd0, 32'sd11, 32'sd2, 32'sd4, 32'sd0, 32'sd17, 32'sd6, 32'sd10, 32'sd16, 32'sd16, 32'sd16, 32'sd11, 32'sd11, 32'sd3, 32'sd4, 32'sd0, 32'sd16, 32'sd15, 32'sd15, 32'sd17, 32'sd8, 32'sd6, 32'sd8, 32'sd8, 32'sd5, 32'sd6, 32'sd7, 32'sd5, 32'sd9, 32'sd8, 32'sd8, 32'sd11, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd3, 32'sd10, 32'sd0, 32'sd3, 32'sd4, 32'sd0, 32'sd5, 32'sd0, 32'sd4, 32'sd10, 32'sd10, 32'sd11, 32'sd10, 32'sd12, 32'sd21, 32'sd20, 32'sd15, 32'sd17, 32'sd12, 32'sd6, 32'sd13, 32'sd16, 32'sd5, 32'sd1, 32'sd19, 32'sd1, 32'sd2, 32'sd10, 32'sd11, 32'sd9, 32'sd10, 32'sd7, 32'sd0, 32'sd6, 32'sd0, 32'sd2, 32'sd17, 32'sd0, 32'sd0, 32'sd17, 32'sd7, 32'sd3, 32'sd2, 32'sd2, 32'sd1, 32'sd16, 32'sd13, 32'sd15, 32'sd5, 32'sd13, 32'sd2, 32'sd14, 32'sd12, 32'sd13, 32'sd8, 32'sd12, 32'sd16, 32'sd1, 32'sd2, 32'sd6, 32'sd7, 32'sd0, 32'sd8, 32'sd12, 32'sd21, 32'sd0, 32'sd6, 32'sd4, 32'sd7, 32'sd8, 32'sd8, 32'sd14, 32'sd11, 32'sd12, 32'sd0, 32'sd10, 32'sd2, 32'sd0, 32'sd6, 32'sd6, 32'sd11, 32'sd11, 32'sd16, 32'sd6, 32'sd16, 32'sd7, 32'sd10, 32'sd4, 32'sd18, 32'sd0, 32'sd3, 32'sd0, 32'sd1, 32'sd1, 32'sd16, 32'sd3, 32'sd16, 32'sd3, 32'sd9, 32'sd4, 32'sd7, 32'sd7, 32'sd4, 32'sd12, 32'sd3, 32'sd6, 32'sd6, 32'sd3, 32'sd3, 32'sd6, 32'sd1, 32'sd17, 32'sd18, 32'sd5, 32'sd6, 32'sd2, 32'sd7, 32'sd0, 32'sd8, 32'sd7, 32'sd5, 32'sd9, 32'sd14, 32'sd14, 32'sd8, 32'sd11, 32'sd0, 32'sd0, 32'sd1, 32'sd11, 32'sd18, 32'sd9, 32'sd10, 32'sd6, 32'sd14, 32'sd7, 32'sd4, 32'sd16, 32'sd13, 32'sd8, 32'sd16, 32'sd0, 32'sd5, 32'sd5, 32'sd6, 32'sd7, 32'sd10, 32'sd12, 32'sd10, 32'sd0, 32'sd4, 32'sd10, 32'sd6, 32'sd11, 32'sd8, 32'sd11, 32'sd9, 32'sd12, 32'sd4, 32'sd4, 32'sd9, 32'sd5, 32'sd9, 32'sd0, 32'sd9, 32'sd9, 32'sd4, 32'sd3, 32'sd1, 32'sd6, 32'sd18, 32'sd8, 32'sd19, 32'sd8, 32'sd8, 32'sd12, 32'sd7, 32'sd1, 32'sd12, 32'sd0, 32'sd0, 32'sd3, 32'sd6, 32'sd11, 32'sd8, 32'sd17, 32'sd14, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd11, 32'sd20, 32'sd6, 32'sd0, 32'sd3, 32'sd5, 32'sd12, 32'sd0, 32'sd0, 32'sd5, 32'sd12, 32'sd13, 32'sd1, 32'sd0, 32'sd2, 32'sd2, 32'sd10, 32'sd10, 32'sd6, 32'sd12, 32'sd14, 32'sd1, 32'sd11, 32'sd15, 32'sd14, 32'sd3, 32'sd6, 32'sd6, 32'sd1, 32'sd1, 32'sd15, 32'sd15, 32'sd1, 32'sd3, 32'sd0, 32'sd3, 32'sd5, 32'sd0, 32'sd1, 32'sd7, 32'sd3, 32'sd3, 32'sd7, 32'sd7, 32'sd13, 32'sd5, 32'sd1, 32'sd1, 32'sd15, 32'sd2, 32'sd5, 32'sd15, 32'sd12, 32'sd12, 32'sd0, 32'sd2, 32'sd7, 32'sd9, 32'sd5, 32'sd5, 32'sd17, 32'sd18, 32'sd17, 32'sd17, 32'sd17, 32'sd0, 32'sd0, 32'sd14, 32'sd13, 32'sd20, 32'sd9, 32'sd10, 32'sd8, 32'sd10, 32'sd10, 32'sd15, 32'sd5, 32'sd13, 32'sd17, 32'sd12, 32'sd9, 32'sd9, 32'sd7, 32'sd4, 32'sd8, 32'sd7, 32'sd15, 32'sd8, 32'sd17, 32'sd17, 32'sd1, 32'sd7, 32'sd5, 32'sd4, 32'sd16, 32'sd16, 32'sd0, 32'sd6, 32'sd4, 32'sd0, 32'sd1, 32'sd6, 32'sd9, 32'sd2, 32'sd2, 32'sd3, 32'sd1, 32'sd9, 32'sd10, 32'sd0, 32'sd4, 32'sd1, 32'sd8, 32'sd0, 32'sd22, 32'sd15, 32'sd0, 32'sd7, 32'sd14, 32'sd14, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd2, 32'sd2, 32'sd0, 32'sd4, 32'sd16, 32'sd0, 32'sd12, 32'sd21, 32'sd5, 32'sd5, 32'sd6, 32'sd5, 32'sd14, 32'sd5, 32'sd8, 32'sd6, 32'sd13, 32'sd10, 32'sd13, 32'sd0, 32'sd1, 32'sd4, 32'sd3, 32'sd13, 32'sd13, 32'sd13, 32'sd16, 32'sd16, 32'sd16, 32'sd16, 32'sd0, 32'sd1, 32'sd2, 32'sd15, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd0, 32'sd12, 32'sd2, 32'sd10, 32'sd3, 32'sd7, 32'sd11, 32'sd8, 32'sd0, 32'sd0, 32'sd3, 32'sd18, 32'sd18, 32'sd3, 32'sd7, 32'sd3, 32'sd17, 32'sd5, 32'sd6, 32'sd16, 32'sd2, 32'sd2, 32'sd4, 32'sd13, 32'sd1, 32'sd12, 32'sd7, 32'sd5, 32'sd11, 32'sd11, 32'sd4, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd13, 32'sd7, 32'sd8, 32'sd14, 32'sd0, 32'sd15, 32'sd9, 32'sd4, 32'sd10, 32'sd5, 32'sd18, 32'sd18, 32'sd20, 32'sd8, 32'sd8, 32'sd5, 32'sd5, 32'sd6, 32'sd0, 32'sd4, 32'sd4, 32'sd12, 32'sd0, 32'sd12, 32'sd12, 32'sd15, 32'sd15, 32'sd0, 32'sd0, 32'sd6, 32'sd12, 32'sd4, 32'sd22, 32'sd7, 32'sd0, 32'sd1, 32'sd16, 32'sd7, 32'sd10, 32'sd2, 32'sd9, 32'sd2, 32'sd2, 32'sd3, 32'sd13, 32'sd14, 32'sd2, 32'sd4, 32'sd1, 32'sd6, 32'sd21, 32'sd5, 32'sd6, 32'sd6, 32'sd3, 32'sd10, 32'sd15, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd10, 32'sd2, 32'sd5, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd2, 32'sd10, 32'sd7, 32'sd0, 32'sd3, 32'sd7, 32'sd6, 32'sd2, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd17, 32'sd14, 32'sd15, 32'sd15, 32'sd14, 32'sd8, 32'sd7, 32'sd8, 32'sd0, 32'sd8, 32'sd5, 32'sd6, 32'sd7, 32'sd8, 32'sd8, 32'sd10, 32'sd5, 32'sd12, 32'sd9, 32'sd14, 32'sd9, 32'sd18, 32'sd6, 32'sd6, 32'sd16, 32'sd16, 32'sd11, 32'sd6, 32'sd7, 32'sd6, 32'sd7, 32'sd10, 32'sd12, 32'sd14, 32'sd12, 32'sd13, 32'sd0, 32'sd1, 32'sd16, 32'sd17, 32'sd2, 32'sd0, 32'sd0, 32'sd2, 32'sd1, 32'sd8, 32'sd8, 32'sd5, 32'sd5, 32'sd4, 32'sd7, 32'sd15, 32'sd2, 32'sd1, 32'sd1, 32'sd1, 32'sd1, 32'sd11, 32'sd11, 32'sd6, 32'sd10, 32'sd9, 32'sd18, 32'sd21, 32'sd12, 32'sd6, 32'sd6, 32'sd4, 32'sd12, 32'sd14, 32'sd7, 32'sd13, 32'sd7, 32'sd12, 32'sd2, 32'sd0, 32'sd9, 32'sd10, 32'sd10, 32'sd15, 32'sd16, 32'sd2, 32'sd5, 32'sd0, 32'sd16, 32'sd12, 32'sd15, 
                                                    32'sd10, 32'sd9, 32'sd11, 32'sd7, 32'sd15, 32'sd8, 32'sd4, 32'sd6, 32'sd6, 32'sd7, 32'sd8, 32'sd8, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd11, 32'sd11, 32'sd8, 32'sd6, 32'sd18, 32'sd4, 32'sd1, 32'sd11, 32'sd12, 32'sd12, 32'sd0, 32'sd12, 32'sd20, 32'sd4, 32'sd2, 32'sd8, 32'sd7, 32'sd0, 32'sd11, 32'sd0, 32'sd7, 32'sd17, 32'sd10, 32'sd5, 32'sd11, 32'sd4, 32'sd0, 32'sd4, 32'sd4, 32'sd18, 32'sd0, 32'sd4, 32'sd4, 32'sd11, 32'sd6, 32'sd0, 32'sd9, 32'sd15, 32'sd7, 32'sd15, 32'sd12, 32'sd12, 32'sd12, 32'sd7, 32'sd7, 32'sd4, 32'sd4, 32'sd11, 32'sd16, 32'sd15, 32'sd15, 32'sd1, 32'sd21, 32'sd20, 32'sd1, 32'sd17, 32'sd16, 32'sd16, 32'sd16, 32'sd10, 32'sd18, 32'sd5, 32'sd2, 32'sd7, 32'sd6, 32'sd0, 32'sd7, 32'sd1, 32'sd18, 32'sd2, 32'sd7, 32'sd1, 32'sd0, 32'sd3, 32'sd15, 32'sd10, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd17, 32'sd20, 32'sd3, 32'sd3, 32'sd6, 32'sd6, 32'sd9, 32'sd18, 32'sd0, 32'sd1, 32'sd0, 32'sd10, 32'sd16, 32'sd16, 32'sd12, 32'sd16, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd4, 32'sd8, 32'sd3, 32'sd3, 32'sd1, 32'sd5, 32'sd6, 32'sd10, 32'sd4, 32'sd2, 32'sd4, 32'sd4, 32'sd8, 32'sd8, 32'sd13, 32'sd13, 32'sd13, 32'sd2, 32'sd2, 32'sd2, 32'sd0, 32'sd2, 32'sd5, 32'sd3, 32'sd21, 32'sd10, 32'sd10, 32'sd8, 32'sd8, 32'sd8, 32'sd15, 32'sd13, 32'sd8, 32'sd13, 32'sd15, 32'sd4, 32'sd15, 32'sd15, 32'sd11, 32'sd6, 32'sd2, 32'sd2, 32'sd1, 32'sd7, 32'sd6, 32'sd11, 32'sd16, 32'sd0, 32'sd11, 32'sd9, 32'sd5, 32'sd2, 32'sd3, 32'sd15, 32'sd0, 32'sd0, 32'sd1, 32'sd0, 32'sd2, 32'sd2, 32'sd2, 32'sd4, 32'sd1, 32'sd1, 32'sd5, 32'sd4, 32'sd5, 32'sd5, 32'sd5, 32'sd0, 32'sd8, 32'sd6, 32'sd3, 32'sd18, 32'sd8, 32'sd2, 32'sd5, 32'sd4, 32'sd6, 32'sd1, 32'sd4, 32'sd6, 32'sd17, 32'sd6, 32'sd6, 32'sd5, 32'sd2, 32'sd2, 32'sd6, 32'sd3, 32'sd3, 32'sd3, 32'sd1, 32'sd2, 32'sd2, 32'sd14, 32'sd8, 32'sd0, 32'sd0, 32'sd6, 32'sd5, 32'sd7, 32'sd16, 32'sd17, 32'sd8, 32'sd13, 32'sd17, 32'sd17, 32'sd0, 32'sd2, 32'sd3, 32'sd17, 32'sd17, 32'sd18, 32'sd15, 32'sd13, 32'sd14, 32'sd18, 32'sd13, 32'sd14, 32'sd2, 32'sd9, 32'sd3, 32'sd2, 32'sd4, 32'sd5, 32'sd5, 32'sd6, 32'sd4, 32'sd4, 32'sd7, 32'sd9, 32'sd0, 32'sd3, 32'sd1, 32'sd22, 32'sd10, 32'sd0, 32'sd0, 32'sd2, 32'sd13, 32'sd21, 32'sd1, 32'sd7, 32'sd0, 32'sd1, 32'sd1, 32'sd2, 32'sd5, 32'sd2, 32'sd2, 32'sd11, 32'sd7, 32'sd9, 32'sd9, 32'sd4, 32'sd6, 32'sd21, 32'sd21, 32'sd5, 32'sd10, 32'sd0, 32'sd2, 32'sd0, 32'sd12, 32'sd13, 32'sd0, 32'sd1, 32'sd13, 32'sd21, 32'sd3, 32'sd10, 32'sd3, 32'sd2, 32'sd1, 32'sd0, 32'sd1, 32'sd18, 32'sd15, 32'sd10, 32'sd9, 32'sd11, 32'sd7, 32'sd2, 32'sd2, 32'sd4, 32'sd5, 32'sd7, 32'sd4, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd1, 32'sd0, 32'sd5, 32'sd0, 32'sd14, 32'sd14, 32'sd18, 32'sd0, 32'sd4, 32'sd2, 32'sd1, 32'sd8, 32'sd15, 32'sd10, 32'sd17, 32'sd4, 32'sd0, 32'sd6, 32'sd9, 32'sd9, 32'sd11, 32'sd2, 32'sd0, 32'sd15, 32'sd18, 32'sd17, 32'sd11, 32'sd11, 32'sd9, 32'sd16, 32'sd16, 32'sd1, 32'sd2, 32'sd15, 32'sd11, 32'sd18, 32'sd14, 32'sd7, 32'sd8, 32'sd1, 32'sd14, 32'sd7, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd8, 32'sd21, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd1, 32'sd1, 32'sd13, 32'sd0, 32'sd5, 32'sd10, 32'sd7, 32'sd10, 32'sd6, 32'sd2, 32'sd13, 32'sd6, 32'sd13, 32'sd20, 32'sd4, 32'sd6, 32'sd0, 32'sd13, 32'sd16, 32'sd0, 32'sd6, 32'sd5, 32'sd15, 32'sd7, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd18, 32'sd15, 32'sd3, 32'sd3, 32'sd14, 32'sd14, 32'sd15, 32'sd17, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd7, 32'sd8, 32'sd9, 32'sd0, 32'sd1, 32'sd4, 32'sd1, 32'sd2, 32'sd1, 32'sd0, 32'sd17, 32'sd14, 32'sd15, 32'sd21, 32'sd15, 32'sd15, 32'sd6, 32'sd3, 32'sd1, 32'sd4, 32'sd1, 32'sd2, 32'sd2, 32'sd2, 32'sd7, 32'sd3, 32'sd6, 32'sd1, 32'sd8, 32'sd0, 32'sd16, 32'sd16, 32'sd19, 32'sd16, 32'sd8, 32'sd15, 32'sd18, 32'sd18, 32'sd3, 32'sd5, 32'sd5, 32'sd6, 32'sd2, 32'sd6, 32'sd2, 32'sd8, 32'sd5, 32'sd8, 32'sd0, 32'sd12, 32'sd12, 32'sd7, 32'sd14, 32'sd6, 32'sd6, 32'sd13, 32'sd10, 32'sd10, 32'sd9, 32'sd3, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd1, 32'sd1, 32'sd0, 32'sd10, 32'sd9, 32'sd9, 32'sd7, 32'sd15, 32'sd10, 32'sd4, 32'sd2, 32'sd0, 32'sd9, 32'sd2, 32'sd0, 32'sd15, 32'sd14, 32'sd1, 32'sd0, 32'sd3, 32'sd2, 32'sd4, 32'sd16, 32'sd16, 32'sd18, 32'sd0, 32'sd3, 32'sd12, 32'sd3, 32'sd3, 32'sd8, 32'sd15, 32'sd13, 32'sd6, 32'sd9, 32'sd0, 32'sd3, 32'sd3, 32'sd5, 32'sd4, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd1, 32'sd2, 32'sd13, 32'sd13, 32'sd2, 32'sd9, 32'sd6, 32'sd8, 32'sd7, 32'sd12, 32'sd10, 32'sd6, 32'sd12, 32'sd15, 32'sd14, 32'sd8, 32'sd10, 32'sd10, 32'sd9, 32'sd12, 32'sd12, 32'sd12, 32'sd12, 32'sd12, 32'sd10, 32'sd15, 32'sd10, 32'sd1, 32'sd4, 32'sd5, 32'sd10, 32'sd12, 32'sd0, 32'sd10, 32'sd2, 32'sd20, 32'sd10, 32'sd17, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd7, 32'sd1, 32'sd14, 32'sd13, 32'sd6, 32'sd2, 32'sd6, 32'sd19, 32'sd15, 32'sd5, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd1, 32'sd13, 32'sd1, 32'sd17, 32'sd13, 32'sd18, 32'sd14, 32'sd1, 32'sd4, 32'sd0, 32'sd5, 32'sd5, 32'sd1, 32'sd1, 32'sd0, 32'sd4, 32'sd6, 32'sd18, 32'sd18, 32'sd15, 32'sd7, 32'sd7, 32'sd9, 32'sd13, 32'sd15, 32'sd15, 32'sd13, 32'sd13, 32'sd5, 32'sd18, 32'sd19, 32'sd19, 32'sd19, 32'sd14, 32'sd0, 32'sd1, 32'sd9, 32'sd15, 32'sd0, 32'sd10, 32'sd10, 32'sd8, 32'sd5, 32'sd5, 32'sd4, 32'sd4, 32'sd7, 32'sd6, 32'sd4, 32'sd0, 32'sd1, 32'sd1, 32'sd14, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd7, 32'sd22, 32'sd16, 32'sd3, 32'sd10, 32'sd16, 32'sd0, 32'sd5, 32'sd8, 32'sd1, 32'sd6, 32'sd3, 32'sd13, 32'sd12, 32'sd5, 32'sd5, 32'sd6, 32'sd1, 32'sd19, 32'sd14, 32'sd6, 32'sd0, 32'sd0, 32'sd1, 32'sd8, 32'sd7, 32'sd12, 32'sd1, 32'sd1, 32'sd7, 32'sd10, 32'sd7, 32'sd3, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd2, 32'sd1, 32'sd0, 32'sd17, 
                                                    32'sd18, 32'sd17, 32'sd15, 32'sd15, 32'sd14, 32'sd10, 32'sd18, 32'sd12, 32'sd10, 32'sd10, 32'sd2, 32'sd6, 32'sd14, 32'sd14, 32'sd1, 32'sd21, 32'sd1, 32'sd16, 32'sd1, 32'sd0, 32'sd1, 32'sd1, 32'sd7, 32'sd14, 32'sd1, 32'sd0, 32'sd1, 32'sd1, 32'sd0, 32'sd14, 32'sd7, 32'sd11, 32'sd5, 32'sd6, 32'sd1, 32'sd1, 32'sd9, 32'sd4, 32'sd16, 32'sd0, 32'sd5, 32'sd3, 32'sd12, 32'sd11, 32'sd10, 32'sd9, 32'sd2, 32'sd6, 32'sd8, 32'sd1, 32'sd1, 32'sd14, 32'sd16, 32'sd16, 32'sd4, 32'sd19, 32'sd8, 32'sd1, 32'sd8, 32'sd8, 32'sd5, 32'sd6, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd0, 32'sd1, 32'sd6, 32'sd6, 32'sd17, 32'sd22, 32'sd12, 32'sd12, 32'sd12, 32'sd14, 32'sd6, 32'sd7, 32'sd3, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd12, 32'sd2, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd6, 32'sd1, 32'sd7, 32'sd7, 32'sd20, 32'sd6, 32'sd2, 32'sd3, 32'sd4, 32'sd1, 32'sd0, 32'sd2, 32'sd2, 32'sd15, 32'sd17, 32'sd6, 32'sd0, 32'sd4, 32'sd6, 32'sd12, 32'sd14, 32'sd14, 32'sd18, 32'sd3, 32'sd3, 32'sd6, 32'sd5, 32'sd4, 32'sd16, 32'sd8, 32'sd6, 32'sd5, 32'sd1, 32'sd1, 32'sd10, 32'sd2, 32'sd0, 32'sd1, 32'sd6, 32'sd1, 32'sd4, 32'sd0, 32'sd16, 32'sd16, 32'sd0, 32'sd3, 32'sd7, 32'sd9, 32'sd14, 32'sd14, 32'sd21, 32'sd21, 32'sd4, 32'sd7, 32'sd4, 32'sd15, 32'sd13, 32'sd6, 32'sd16, 32'sd5, 32'sd8, 32'sd8, 32'sd8, 32'sd8, 32'sd8, 32'sd6, 32'sd8, 32'sd5, 32'sd5, 32'sd1, 32'sd10, 32'sd17, 32'sd16, 32'sd10, 32'sd4, 32'sd18, 32'sd18, 32'sd16, 32'sd15, 32'sd15, 32'sd1, 32'sd1, 32'sd5, 32'sd5, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd5, 32'sd6, 32'sd2, 32'sd2, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd8, 32'sd0, 32'sd10, 32'sd0, 32'sd1, 32'sd1, 32'sd6, 32'sd12, 32'sd9, 32'sd10, 32'sd18, 32'sd16, 32'sd14, 32'sd14, 32'sd10, 32'sd13, 32'sd13, 32'sd0, 32'sd8, 32'sd5, 32'sd0, 32'sd11, 32'sd5, 32'sd18, 32'sd8, 32'sd7, 32'sd0, 32'sd0, 32'sd2, 32'sd8, 32'sd9, 32'sd7, 32'sd2, 32'sd0, 32'sd14, 32'sd12, 32'sd12, 32'sd6, 32'sd0, 32'sd8, 32'sd6, 32'sd11, 32'sd3, 32'sd12, 32'sd16, 32'sd6, 32'sd10, 32'sd10, 32'sd12, 32'sd12, 32'sd15, 32'sd15, 32'sd20, 32'sd20, 32'sd17, 32'sd2, 32'sd1, 32'sd15, 32'sd2, 32'sd12, 32'sd7, 32'sd1, 32'sd8, 32'sd3, 32'sd6, 32'sd0, 32'sd0, 32'sd15, 32'sd7, 32'sd6, 32'sd21, 32'sd3, 32'sd7, 32'sd2, 32'sd10, 32'sd9, 32'sd5, 32'sd9, 32'sd11, 32'sd13, 32'sd0, 32'sd18, 32'sd4, 32'sd8, 32'sd3, 32'sd15, 32'sd18, 32'sd14, 32'sd15, 32'sd6, 32'sd6, 32'sd6, 32'sd14, 32'sd8, 32'sd6, 32'sd9, 32'sd9, 32'sd15, 32'sd20, 32'sd18, 32'sd18, 32'sd16, 32'sd16, 32'sd2, 32'sd2, 32'sd0, 32'sd20, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd12, 32'sd12, 32'sd5, 32'sd6, 32'sd5, 32'sd16, 32'sd8, 32'sd8, 32'sd4, 32'sd4, 32'sd7, 32'sd19, 32'sd11, 32'sd1, 32'sd2, 32'sd13, 32'sd0, 32'sd11, 32'sd1, 32'sd10, 32'sd19, 32'sd10, 32'sd1, 32'sd1, 32'sd4, 32'sd4, 32'sd6, 32'sd9, 32'sd5, 32'sd2, 32'sd0, 32'sd0, 32'sd7, 32'sd2, 32'sd0, 32'sd6, 32'sd8, 32'sd18, 32'sd14, 32'sd15, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd2, 32'sd6, 32'sd1, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd2, 32'sd11, 32'sd8, 32'sd8, 32'sd8, 32'sd11, 32'sd9, 32'sd4, 32'sd17, 32'sd21, 32'sd4, 32'sd15, 32'sd8, 32'sd12, 32'sd17, 32'sd16, 32'sd1, 32'sd1, 32'sd13, 32'sd1, 32'sd4, 32'sd8, 32'sd7, 32'sd7, 32'sd6, 32'sd6, 32'sd9, 32'sd1, 32'sd6, 32'sd5, 32'sd6, 32'sd4, 32'sd8, 32'sd10, 32'sd5, 32'sd4, 32'sd4, 32'sd7, 32'sd6, 32'sd5, 32'sd7, 32'sd7, 32'sd2, 32'sd1, 32'sd13, 32'sd13, 32'sd15, 32'sd15, 32'sd0, 32'sd6, 32'sd7, 32'sd9, 32'sd6, 32'sd7, 32'sd12, 32'sd14, 32'sd17, 32'sd12, 32'sd17, 32'sd3, 32'sd17, 32'sd1, 32'sd17, 32'sd5, 32'sd7, 32'sd4, 32'sd1, 32'sd5, 32'sd0, 32'sd11, 32'sd7, 32'sd7, 32'sd17, 32'sd6, 32'sd15, 32'sd15, 32'sd10, 32'sd10, 32'sd15, 32'sd1, 32'sd0, 32'sd0, 32'sd1, 32'sd21, 32'sd9, 32'sd4, 32'sd1, 32'sd9, 32'sd1, 32'sd0, 32'sd0, 32'sd6, 32'sd1, 32'sd12, 32'sd17, 32'sd1, 32'sd0, 32'sd6, 32'sd0, 32'sd7, 32'sd12, 32'sd9, 32'sd1, 32'sd11, 32'sd11, 32'sd10, 32'sd2, 32'sd16, 32'sd16, 32'sd13, 32'sd16, 32'sd16, 32'sd18, 32'sd13, 32'sd2, 32'sd8, 32'sd13, 32'sd20, 32'sd8, 32'sd7, 32'sd6, 32'sd20, 32'sd20, 32'sd1, 32'sd1, 32'sd3, 32'sd2, 32'sd9, 32'sd3, 32'sd0, 32'sd9, 32'sd4, 32'sd4, 32'sd13, 32'sd13, 32'sd15, 32'sd13, 32'sd0, 32'sd2, 32'sd1, 32'sd1, 32'sd6, 32'sd2, 32'sd11, 32'sd1, 32'sd0, 32'sd3, 32'sd1, 32'sd7, 32'sd0, 32'sd0, 32'sd9, 32'sd15, 32'sd7, 32'sd9, 32'sd17, 32'sd3, 32'sd1, 32'sd15, 32'sd0, 32'sd3, 32'sd1, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd11, 32'sd7, 32'sd6, 32'sd14, 32'sd14, 32'sd0, 32'sd0, 32'sd1, 32'sd12, 32'sd8, 32'sd6, 32'sd5, 32'sd9, 32'sd8, 32'sd12, 32'sd19, 32'sd0, 32'sd4, 32'sd16, 32'sd7, 32'sd7, 32'sd6, 32'sd17, 32'sd17, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd12, 32'sd9, 32'sd5, 32'sd5, 32'sd7, 32'sd1, 32'sd0, 32'sd6, 32'sd8, 32'sd6, 32'sd12, 32'sd4, 32'sd1, 32'sd1, 32'sd10, 32'sd4, 32'sd13, 32'sd13, 32'sd15, 32'sd14, 32'sd14, 32'sd8, 32'sd10, 32'sd10, 32'sd7, 32'sd10, 32'sd1, 32'sd15, 32'sd6, 32'sd1, 32'sd6, 32'sd18, 32'sd0, 32'sd13, 32'sd6, 32'sd6, 32'sd6, 32'sd7, 32'sd8, 32'sd8, 32'sd8, 32'sd2, 32'sd10, 32'sd10, 32'sd7, 32'sd7, 32'sd9, 32'sd2, 32'sd2, 32'sd1, 32'sd2, 32'sd3, 32'sd8, 32'sd8, 32'sd18, 32'sd6, 32'sd6, 32'sd3, 32'sd6, 32'sd8, 32'sd2, 32'sd14, 32'sd2, 32'sd3, 32'sd6, 32'sd2, 32'sd17, 32'sd7, 32'sd11, 32'sd1, 32'sd0, 32'sd0, 32'sd7, 32'sd2, 32'sd1, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd18, 32'sd8, 32'sd6, 32'sd2, 32'sd7, 32'sd6, 32'sd2, 32'sd9, 32'sd4, 32'sd8, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd6, 32'sd0, 32'sd1, 32'sd4, 32'sd5, 32'sd13, 32'sd14, 32'sd2, 32'sd1, 32'sd1, 32'sd4, 32'sd5, 32'sd1, 32'sd12, 32'sd12, 32'sd18, 32'sd13, 32'sd3, 32'sd9, 32'sd3, 32'sd2, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd16, 32'sd20, 32'sd10, 32'sd6, 32'sd1, 32'sd13, 32'sd15, 32'sd12, 32'sd11, 32'sd6, 32'sd0, 32'sd0, 
                                                    32'sd3, 32'sd3, 32'sd5, 32'sd5, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd6, 32'sd16, 32'sd16, 32'sd6, 32'sd7, 32'sd6, 32'sd1, 32'sd9, 32'sd5, 32'sd11, 32'sd8, 32'sd8, 32'sd6, 32'sd5, 32'sd7, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd6, 32'sd21, 32'sd19, 32'sd18, 32'sd18, 32'sd16, 32'sd16, 32'sd0, 32'sd0, 32'sd14, 32'sd14, 32'sd14, 32'sd14, 32'sd18, 32'sd18, 32'sd5, 32'sd3, 32'sd0, 32'sd0, 32'sd12, 32'sd3, 32'sd4, 32'sd4, 32'sd14, 32'sd14, 32'sd6, 32'sd11, 32'sd5, 32'sd4, 32'sd8, 32'sd8, 32'sd6, 32'sd14, 32'sd6, 32'sd6, 32'sd14, 32'sd5, 32'sd5, 32'sd0, 32'sd3, 32'sd3, 32'sd12, 32'sd10, 32'sd8, 32'sd14, 32'sd10, 32'sd10, 32'sd12, 32'sd8, 32'sd11, 32'sd11, 32'sd2, 32'sd2, 32'sd12, 32'sd10, 32'sd9, 32'sd8, 32'sd7, 32'sd0, 32'sd0, 32'sd5, 32'sd6, 32'sd0, 32'sd1, 32'sd0, 32'sd3, 32'sd14, 32'sd9, 32'sd2, 32'sd4, 32'sd4, 32'sd5, 32'sd7, 32'sd5, 32'sd5, 32'sd4, 32'sd14, 32'sd17, 32'sd16, 32'sd17, 32'sd20, 32'sd14, 32'sd6, 32'sd4, 32'sd3, 32'sd8, 32'sd6, 32'sd6, 32'sd5, 32'sd5, 32'sd5, 32'sd2, 32'sd1, 32'sd2, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd1, 32'sd9, 32'sd8, 32'sd9, 32'sd9, 32'sd0, 32'sd1, 32'sd1, 32'sd20, 32'sd0, 32'sd8, 32'sd8, 32'sd13, 32'sd13, 32'sd8, 32'sd8, 32'sd11, 32'sd11, 32'sd12, 32'sd1, 32'sd11, 32'sd10, 32'sd8, 32'sd8, 32'sd14, 32'sd18, 32'sd16, 32'sd20, 32'sd12, 32'sd12, 32'sd17, 32'sd6, 32'sd17, 32'sd18, 32'sd15, 32'sd13, 32'sd17, 32'sd17, 32'sd17, 32'sd17, 32'sd2, 32'sd13, 32'sd1}

localparam logic [2912:0][31:0] rectangle1_widths = {32'sd12, 32'sd12, 32'sd18, 32'sd9, 32'sd4, 32'sd12, 32'sd12, 32'sd4, 32'sd7, 32'sd12, 32'sd12, 32'sd19, 32'sd24, 32'sd6, 32'sd14, 32'sd14, 32'sd9, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd24, 32'sd6, 32'sd10, 32'sd14, 32'sd24, 32'sd15, 32'sd5, 32'sd6, 32'sd3, 32'sd18, 32'sd13, 32'sd6, 32'sd6, 32'sd24, 32'sd14, 32'sd21, 32'sd4, 32'sd20, 32'sd6, 32'sd4, 32'sd22, 32'sd6, 32'sd6, 32'sd4, 32'sd19, 32'sd4, 32'sd4, 32'sd14, 32'sd18, 32'sd4, 32'sd6, 32'sd12, 32'sd12, 32'sd24, 32'sd18, 32'sd12, 32'sd4, 32'sd4, 32'sd24, 32'sd8, 32'sd3, 32'sd16, 32'sd12, 32'sd6, 32'sd9, 32'sd18, 32'sd16, 32'sd4, 32'sd18, 32'sd20, 32'sd14, 32'sd7, 32'sd9, 32'sd9, 32'sd8, 32'sd14, 32'sd12, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd12, 32'sd24, 32'sd16, 32'sd6, 32'sd24, 32'sd4, 32'sd15, 32'sd4, 32'sd4, 32'sd6, 32'sd18, 32'sd4, 32'sd8, 32'sd10, 32'sd10, 32'sd18, 32'sd22, 32'sd18, 32'sd6, 32'sd4, 32'sd4, 32'sd20, 32'sd8, 32'sd6, 32'sd6, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd12, 32'sd20, 32'sd18, 32'sd18, 32'sd14, 32'sd10, 32'sd12, 32'sd18, 32'sd8, 32'sd18, 32'sd6, 32'sd12, 32'sd4, 32'sd19, 32'sd22, 32'sd11, 32'sd15, 32'sd12, 32'sd12, 32'sd5, 32'sd24, 32'sd12, 32'sd9, 32'sd6, 32'sd22, 32'sd17, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd8, 32'sd19, 32'sd6, 32'sd17, 32'sd3, 32'sd8, 32'sd9, 32'sd9, 32'sd10, 32'sd3, 32'sd24, 32'sd18, 32'sd6, 32'sd10, 32'sd9, 32'sd16, 32'sd9, 32'sd20, 32'sd9, 32'sd9, 32'sd10, 32'sd6, 32'sd12, 32'sd18, 32'sd22, 32'sd8, 32'sd6, 32'sd6, 32'sd11, 32'sd24, 32'sd22, 32'sd20, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd9, 32'sd9, 32'sd18, 32'sd8, 32'sd18, 32'sd12, 32'sd14, 32'sd6, 32'sd6, 32'sd9, 32'sd18, 32'sd5, 32'sd4, 32'sd18, 32'sd19, 32'sd4, 32'sd19, 32'sd6, 32'sd14, 32'sd20, 32'sd22, 32'sd7, 32'sd22, 32'sd22, 32'sd6, 32'sd9, 32'sd4, 32'sd12, 32'sd6, 32'sd18, 32'sd6, 32'sd16, 32'sd6, 32'sd24, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd9, 32'sd14, 32'sd18, 32'sd15, 32'sd15, 32'sd16, 32'sd10, 32'sd15, 32'sd10, 32'sd6, 32'sd18, 32'sd18, 32'sd18, 32'sd14, 32'sd2, 32'sd2, 32'sd15, 32'sd21, 32'sd5, 32'sd24, 32'sd22, 32'sd15, 32'sd24, 32'sd18, 32'sd10, 32'sd10, 32'sd6, 32'sd20, 32'sd10, 32'sd16, 32'sd7, 32'sd6, 32'sd6, 32'sd12, 32'sd10, 32'sd6, 32'sd5, 32'sd24, 32'sd5, 32'sd6, 32'sd6, 32'sd6, 32'sd3, 32'sd13, 32'sd4, 32'sd9, 32'sd6, 32'sd6, 32'sd12, 32'sd6, 32'sd12, 32'sd8, 32'sd10, 32'sd6, 32'sd2, 32'sd6, 32'sd2, 32'sd2, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd18, 32'sd24, 32'sd8, 32'sd4, 32'sd10, 32'sd3, 32'sd6, 32'sd6, 32'sd24, 32'sd13, 32'sd6, 32'sd16, 32'sd6, 32'sd6, 32'sd10, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd5, 32'sd3, 32'sd18, 32'sd19, 32'sd6, 32'sd3, 32'sd3, 32'sd18, 32'sd6, 32'sd9, 32'sd20, 32'sd6, 32'sd22, 32'sd5, 32'sd18, 32'sd6, 32'sd24, 32'sd12, 32'sd12, 32'sd14, 32'sd8, 32'sd5, 32'sd3, 32'sd18, 32'sd20, 32'sd19, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd15, 32'sd6, 32'sd6, 32'sd18, 32'sd12, 32'sd6, 32'sd6, 32'sd9, 32'sd13, 32'sd9, 32'sd6, 32'sd9, 32'sd3, 32'sd9, 32'sd10, 32'sd4, 32'sd4, 32'sd6, 32'sd18, 32'sd10, 32'sd22, 32'sd16, 32'sd18, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd19, 32'sd19, 32'sd10, 32'sd10, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd4, 32'sd14, 32'sd6, 32'sd18, 32'sd9, 32'sd21, 32'sd17, 32'sd11, 32'sd13, 32'sd9, 32'sd15, 32'sd6, 32'sd18, 32'sd24, 32'sd3, 32'sd24, 32'sd10, 32'sd18, 32'sd18, 32'sd16, 32'sd3, 32'sd18, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd12, 32'sd6, 32'sd24, 32'sd5, 32'sd5, 32'sd6, 32'sd6, 32'sd19, 32'sd12, 32'sd4, 32'sd10, 32'sd10, 32'sd10, 32'sd9, 32'sd21, 32'sd9, 32'sd9, 32'sd4, 32'sd4, 32'sd9, 32'sd18, 32'sd6, 32'sd11, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd19, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd18, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd18, 32'sd11, 32'sd14, 32'sd15, 32'sd22, 32'sd24, 32'sd18, 32'sd12, 32'sd7, 32'sd22, 32'sd14, 32'sd24, 32'sd18, 32'sd22, 32'sd11, 32'sd6, 32'sd24, 32'sd10, 32'sd10, 32'sd24, 32'sd18, 32'sd16, 32'sd16, 32'sd18, 32'sd21, 32'sd6, 32'sd6, 32'sd9, 32'sd2, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd24, 32'sd10, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd10, 32'sd2, 32'sd15, 32'sd6, 32'sd6, 32'sd9, 32'sd14, 32'sd8, 32'sd7, 32'sd4, 32'sd6, 32'sd6, 32'sd21, 32'sd5, 32'sd4, 32'sd5, 32'sd11, 32'sd12, 32'sd24, 32'sd23, 32'sd18, 32'sd21, 32'sd6, 32'sd4, 32'sd8, 32'sd15, 32'sd10, 32'sd9, 32'sd6, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd18, 32'sd21, 32'sd6, 32'sd6, 32'sd6, 32'sd16, 32'sd10, 32'sd10, 32'sd10, 32'sd6, 32'sd12, 32'sd3, 32'sd6, 32'sd9, 32'sd8, 32'sd3, 32'sd4, 32'sd9, 32'sd24, 32'sd6, 32'sd6, 32'sd6, 32'sd12, 32'sd2, 32'sd12, 32'sd18, 32'sd18, 32'sd24, 32'sd4, 32'sd6, 32'sd6, 32'sd8, 32'sd16, 32'sd8, 32'sd8, 32'sd11, 32'sd24, 32'sd4, 32'sd4, 32'sd16, 32'sd6, 32'sd18, 32'sd6, 32'sd9, 32'sd8, 32'sd3, 32'sd18, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd18, 32'sd12, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd3, 32'sd14, 32'sd3, 32'sd14, 32'sd14, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd8, 32'sd9, 32'sd8, 32'sd10, 32'sd4, 32'sd6, 32'sd18, 32'sd8, 32'sd24, 32'sd3, 32'sd10, 32'sd10, 32'sd10, 32'sd24, 32'sd15, 32'sd12, 32'sd14, 32'sd4, 32'sd6, 32'sd6, 32'sd18, 32'sd14, 32'sd6, 32'sd6, 32'sd24, 32'sd6, 32'sd10, 32'sd6, 32'sd6, 32'sd11, 32'sd10, 32'sd6, 32'sd6, 32'sd4, 32'sd20, 32'sd10, 32'sd6, 32'sd10, 32'sd4, 32'sd10, 32'sd12, 32'sd8, 32'sd4, 32'sd9, 32'sd14, 32'sd19, 32'sd10, 32'sd16, 32'sd24, 32'sd18, 32'sd18, 32'sd18, 32'sd9, 32'sd23, 32'sd18, 32'sd12, 32'sd3, 32'sd10, 32'sd10, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd3, 32'sd9, 32'sd3, 32'sd6, 32'sd18, 32'sd18, 32'sd8, 32'sd9, 32'sd9, 32'sd5, 32'sd14, 32'sd3, 32'sd15, 32'sd15, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd8, 32'sd8, 32'sd10, 32'sd21, 32'sd12, 32'sd12, 
                                                    32'sd12, 32'sd6, 32'sd20, 32'sd12, 32'sd8, 32'sd8, 32'sd20, 32'sd12, 32'sd16, 32'sd9, 32'sd12, 32'sd14, 32'sd9, 32'sd19, 32'sd6, 32'sd18, 32'sd4, 32'sd20, 32'sd22, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd10, 32'sd12, 32'sd24, 32'sd4, 32'sd4, 32'sd17, 32'sd18, 32'sd14, 32'sd14, 32'sd3, 32'sd3, 32'sd14, 32'sd9, 32'sd18, 32'sd12, 32'sd8, 32'sd7, 32'sd22, 32'sd4, 32'sd7, 32'sd9, 32'sd22, 32'sd6, 32'sd8, 32'sd6, 32'sd6, 32'sd9, 32'sd18, 32'sd12, 32'sd4, 32'sd4, 32'sd6, 32'sd9, 32'sd8, 32'sd6, 32'sd6, 32'sd4, 32'sd19, 32'sd9, 32'sd12, 32'sd18, 32'sd4, 32'sd18, 32'sd4, 32'sd4, 32'sd4, 32'sd6, 32'sd4, 32'sd18, 32'sd20, 32'sd6, 32'sd8, 32'sd3, 32'sd14, 32'sd24, 32'sd18, 32'sd5, 32'sd5, 32'sd8, 32'sd8, 32'sd12, 32'sd6, 32'sd6, 32'sd12, 32'sd23, 32'sd19, 32'sd11, 32'sd8, 32'sd10, 32'sd9, 32'sd9, 32'sd9, 32'sd20, 32'sd9, 32'sd9, 32'sd8, 32'sd21, 32'sd10, 32'sd12, 32'sd23, 32'sd8, 32'sd18, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd24, 32'sd18, 32'sd24, 32'sd18, 32'sd9, 32'sd9, 32'sd18, 32'sd6, 32'sd6, 32'sd5, 32'sd6, 32'sd6, 32'sd8, 32'sd21, 32'sd3, 32'sd11, 32'sd10, 32'sd12, 32'sd18, 32'sd22, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd3, 32'sd16, 32'sd6, 32'sd16, 32'sd18, 32'sd6, 32'sd8, 32'sd10, 32'sd10, 32'sd12, 32'sd8, 32'sd9, 32'sd24, 32'sd18, 32'sd9, 32'sd10, 32'sd4, 32'sd9, 32'sd6, 32'sd12, 32'sd20, 32'sd9, 32'sd9, 32'sd4, 32'sd8, 32'sd9, 32'sd12, 32'sd9, 32'sd6, 32'sd5, 32'sd21, 32'sd10, 32'sd6, 32'sd18, 32'sd8, 32'sd18, 32'sd9, 32'sd18, 32'sd12, 32'sd6, 32'sd4, 32'sd4, 32'sd24, 32'sd9, 32'sd9, 32'sd19, 32'sd22, 32'sd6, 32'sd20, 32'sd6, 32'sd16, 32'sd8, 32'sd6, 32'sd16, 32'sd16, 32'sd4, 32'sd8, 32'sd12, 32'sd6, 32'sd8, 32'sd6, 32'sd6, 32'sd21, 32'sd16, 32'sd7, 32'sd4, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd12, 32'sd23, 32'sd6, 32'sd12, 32'sd10, 32'sd6, 32'sd9, 32'sd9, 32'sd18, 32'sd18, 32'sd12, 32'sd21, 32'sd12, 32'sd6, 32'sd19, 32'sd14, 32'sd18, 32'sd4, 32'sd11, 32'sd9, 32'sd4, 32'sd4, 32'sd18, 32'sd11, 32'sd20, 32'sd13, 32'sd22, 32'sd14, 32'sd10, 32'sd10, 32'sd6, 32'sd9, 32'sd8, 32'sd16, 32'sd14, 32'sd9, 32'sd18, 32'sd9, 32'sd24, 32'sd10, 32'sd18, 32'sd6, 32'sd11, 32'sd12, 32'sd4, 32'sd4, 32'sd6, 32'sd15, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd16, 32'sd20, 32'sd4, 32'sd4, 32'sd18, 32'sd6, 32'sd9, 32'sd15, 32'sd19, 32'sd7, 32'sd9, 32'sd8, 32'sd18, 32'sd12, 32'sd9, 32'sd14, 32'sd22, 32'sd6, 32'sd10, 32'sd10, 32'sd16, 32'sd6, 32'sd8, 32'sd6, 32'sd8, 32'sd4, 32'sd8, 32'sd10, 32'sd14, 32'sd20, 32'sd4, 32'sd12, 32'sd12, 32'sd6, 32'sd8, 32'sd8, 32'sd9, 32'sd16, 32'sd6, 32'sd3, 32'sd5, 32'sd5, 32'sd10, 32'sd23, 32'sd21, 32'sd6, 32'sd12, 32'sd8, 32'sd24, 32'sd8, 32'sd8, 32'sd8, 32'sd5, 32'sd19, 32'sd24, 32'sd13, 32'sd24, 32'sd4, 32'sd6, 32'sd12, 32'sd12, 32'sd18, 32'sd9, 32'sd4, 32'sd4, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd19, 32'sd18, 32'sd16, 32'sd9, 32'sd4, 32'sd15, 32'sd8, 32'sd6, 32'sd6, 32'sd12, 32'sd11, 32'sd21, 32'sd8, 32'sd6, 32'sd21, 32'sd19, 32'sd6, 32'sd6, 32'sd14, 32'sd9, 32'sd8, 32'sd22, 32'sd9, 32'sd18, 32'sd7, 32'sd16, 32'sd12, 32'sd4, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd3, 32'sd6, 32'sd3, 32'sd12, 32'sd4, 32'sd3, 32'sd3, 32'sd10, 32'sd3, 32'sd6, 32'sd19, 32'sd18, 32'sd18, 32'sd6, 32'sd20, 32'sd20, 32'sd6, 32'sd24, 32'sd18, 32'sd6, 32'sd8, 32'sd8, 32'sd14, 32'sd4, 32'sd5, 32'sd8, 32'sd22, 32'sd6, 32'sd9, 32'sd19, 32'sd9, 32'sd18, 32'sd9, 32'sd24, 32'sd14, 32'sd9, 32'sd6, 32'sd13, 32'sd6, 32'sd21, 32'sd9, 32'sd9, 32'sd10, 32'sd24, 32'sd9, 32'sd6, 32'sd9, 32'sd6, 32'sd14, 32'sd14, 32'sd9, 32'sd6, 32'sd10, 32'sd4, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd9, 32'sd4, 32'sd12, 32'sd9, 32'sd10, 32'sd10, 32'sd24, 32'sd9, 32'sd24, 32'sd11, 32'sd22, 32'sd6, 32'sd20, 32'sd14, 32'sd16, 32'sd19, 32'sd10, 32'sd4, 32'sd21, 32'sd6, 32'sd14, 32'sd6, 32'sd9, 32'sd4, 32'sd19, 32'sd20, 32'sd4, 32'sd8, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd24, 32'sd6, 32'sd4, 32'sd4, 32'sd9, 32'sd6, 32'sd7, 32'sd14, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd10, 32'sd14, 32'sd12, 32'sd12, 32'sd6, 32'sd20, 32'sd9, 32'sd6, 32'sd5, 32'sd16, 32'sd8, 32'sd6, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd18, 32'sd18, 32'sd18, 32'sd19, 32'sd6, 32'sd15, 32'sd6, 32'sd6, 32'sd6, 32'sd22, 32'sd21, 32'sd18, 32'sd6, 32'sd18, 32'sd8, 32'sd18, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd7, 32'sd9, 32'sd21, 32'sd7, 32'sd22, 32'sd24, 32'sd9, 32'sd12, 32'sd14, 32'sd14, 32'sd6, 32'sd6, 32'sd20, 32'sd9, 32'sd21, 32'sd14, 32'sd12, 32'sd9, 32'sd6, 32'sd6, 32'sd18, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd24, 32'sd18, 32'sd10, 32'sd12, 32'sd19, 32'sd4, 32'sd9, 32'sd15, 32'sd12, 32'sd6, 32'sd6, 32'sd16, 32'sd14, 32'sd20, 32'sd20, 32'sd6, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd15, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd8, 32'sd4, 32'sd10, 32'sd4, 32'sd10, 32'sd18, 32'sd11, 32'sd12, 32'sd12, 32'sd9, 32'sd15, 32'sd12, 32'sd12, 32'sd12, 32'sd8, 32'sd8, 32'sd24, 32'sd8, 32'sd4, 32'sd4, 32'sd15, 32'sd24, 32'sd5, 32'sd18, 32'sd3, 32'sd4, 32'sd9, 32'sd20, 32'sd18, 32'sd10, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd18, 32'sd20, 32'sd4, 32'sd6, 32'sd18, 32'sd18, 32'sd6, 32'sd6, 32'sd6, 32'sd20, 32'sd20, 32'sd18, 32'sd6, 32'sd22, 32'sd6, 32'sd6, 32'sd24, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd18, 32'sd9, 32'sd23, 32'sd18, 32'sd9, 32'sd8, 32'sd15, 32'sd8, 32'sd6, 32'sd8, 32'sd6, 32'sd4, 32'sd12, 32'sd8, 32'sd8, 32'sd6, 32'sd6, 32'sd12, 32'sd18, 32'sd8, 32'sd22, 32'sd12, 32'sd20, 32'sd20, 32'sd10, 32'sd18, 32'sd19, 32'sd6, 32'sd22, 32'sd7, 32'sd11, 32'sd10, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd18, 32'sd13, 32'sd8, 32'sd8, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd5, 32'sd5, 32'sd6, 32'sd6, 32'sd12, 32'sd24, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd18, 32'sd7, 32'sd12, 32'sd18, 32'sd20, 32'sd6, 32'sd18, 32'sd18, 
                                                    32'sd6, 32'sd9, 32'sd18, 32'sd6, 32'sd12, 32'sd12, 32'sd6, 32'sd4, 32'sd9, 32'sd12, 32'sd6, 32'sd6, 32'sd9, 32'sd12, 32'sd20, 32'sd12, 32'sd3, 32'sd15, 32'sd6, 32'sd12, 32'sd8, 32'sd8, 32'sd9, 32'sd12, 32'sd6, 32'sd9, 32'sd8, 32'sd6, 32'sd24, 32'sd6, 32'sd5, 32'sd5, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd9, 32'sd10, 32'sd10, 32'sd6, 32'sd6, 32'sd10, 32'sd6, 32'sd18, 32'sd6, 32'sd9, 32'sd6, 32'sd4, 32'sd4, 32'sd12, 32'sd10, 32'sd22, 32'sd2, 32'sd24, 32'sd10, 32'sd8, 32'sd6, 32'sd5, 32'sd20, 32'sd12, 32'sd6, 32'sd10, 32'sd12, 32'sd6, 32'sd4, 32'sd6, 32'sd4, 32'sd4, 32'sd19, 32'sd2, 32'sd2, 32'sd2, 32'sd10, 32'sd4, 32'sd6, 32'sd16, 32'sd6, 32'sd6, 32'sd6, 32'sd12, 32'sd9, 32'sd9, 32'sd18, 32'sd22, 32'sd6, 32'sd6, 32'sd16, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd24, 32'sd24, 32'sd6, 32'sd18, 32'sd18, 32'sd22, 32'sd9, 32'sd21, 32'sd12, 32'sd24, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd20, 32'sd12, 32'sd4, 32'sd12, 32'sd4, 32'sd3, 32'sd10, 32'sd12, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd18, 32'sd22, 32'sd10, 32'sd10, 32'sd12, 32'sd12, 32'sd5, 32'sd21, 32'sd9, 32'sd12, 32'sd12, 32'sd8, 32'sd10, 32'sd10, 32'sd12, 32'sd10, 32'sd12, 32'sd4, 32'sd6, 32'sd6, 32'sd11, 32'sd6, 32'sd4, 32'sd4, 32'sd8, 32'sd16, 32'sd18, 32'sd16, 32'sd8, 32'sd9, 32'sd8, 32'sd8, 32'sd8, 32'sd8, 32'sd5, 32'sd7, 32'sd24, 32'sd8, 32'sd8, 32'sd24, 32'sd12, 32'sd12, 32'sd6, 32'sd8, 32'sd18, 32'sd18, 32'sd22, 32'sd12, 32'sd12, 32'sd12, 32'sd6, 32'sd9, 32'sd7, 32'sd9, 32'sd18, 32'sd4, 32'sd6, 32'sd6, 32'sd12, 32'sd14, 32'sd17, 32'sd12, 32'sd9, 32'sd24, 32'sd9, 32'sd18, 32'sd9, 32'sd9, 32'sd24, 32'sd20, 32'sd16, 32'sd4, 32'sd10, 32'sd6, 32'sd7, 32'sd7, 32'sd6, 32'sd19, 32'sd9, 32'sd9, 32'sd10, 32'sd18, 32'sd4, 32'sd4, 32'sd8, 32'sd12, 32'sd6, 32'sd12, 32'sd10, 32'sd21, 32'sd9, 32'sd6, 32'sd6, 32'sd12, 32'sd20, 32'sd10, 32'sd5, 32'sd4, 32'sd8, 32'sd24, 32'sd4, 32'sd18, 32'sd16, 32'sd6, 32'sd14, 32'sd8, 32'sd20, 32'sd9, 32'sd6, 32'sd4, 32'sd4, 32'sd8, 32'sd2, 32'sd9, 32'sd19, 32'sd9, 32'sd18, 32'sd6, 32'sd6, 32'sd4, 32'sd18, 32'sd14, 32'sd18, 32'sd9, 32'sd12, 32'sd7, 32'sd20, 32'sd9, 32'sd15, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd12, 32'sd6, 32'sd8, 32'sd24, 32'sd6, 32'sd8, 32'sd24, 32'sd12, 32'sd9, 32'sd16, 32'sd4, 32'sd5, 32'sd9, 32'sd9, 32'sd6, 32'sd20, 32'sd17, 32'sd7, 32'sd23, 32'sd6, 32'sd4, 32'sd6, 32'sd18, 32'sd9, 32'sd2, 32'sd2, 32'sd18, 32'sd15, 32'sd18, 32'sd4, 32'sd10, 32'sd10, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd6, 32'sd6, 32'sd11, 32'sd10, 32'sd10, 32'sd10, 32'sd6, 32'sd10, 32'sd16, 32'sd16, 32'sd22, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd7, 32'sd8, 32'sd6, 32'sd3, 32'sd8, 32'sd19, 32'sd4, 32'sd18, 32'sd5, 32'sd4, 32'sd16, 32'sd18, 32'sd10, 32'sd12, 32'sd12, 32'sd22, 32'sd9, 32'sd12, 32'sd10, 32'sd8, 32'sd8, 32'sd18, 32'sd10, 32'sd21, 32'sd22, 32'sd6, 32'sd3, 32'sd12, 32'sd12, 32'sd22, 32'sd18, 32'sd22, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd6, 32'sd12, 32'sd12, 32'sd18, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd6, 32'sd6, 32'sd10, 32'sd5, 32'sd5, 32'sd9, 32'sd23, 32'sd8, 32'sd6, 32'sd9, 32'sd18, 32'sd11, 32'sd11, 32'sd24, 32'sd8, 32'sd14, 32'sd21, 32'sd24, 32'sd8, 32'sd21, 32'sd12, 32'sd4, 32'sd4, 32'sd6, 32'sd9, 32'sd19, 32'sd10, 32'sd18, 32'sd6, 32'sd17, 32'sd12, 32'sd6, 32'sd16, 32'sd5, 32'sd18, 32'sd6, 32'sd20, 32'sd15, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd3, 32'sd14, 32'sd12, 32'sd4, 32'sd6, 32'sd4, 32'sd6, 32'sd14, 32'sd16, 32'sd6, 32'sd21, 32'sd6, 32'sd5, 32'sd16, 32'sd14, 32'sd4, 32'sd12, 32'sd12, 32'sd14, 32'sd18, 32'sd18, 32'sd24, 32'sd18, 32'sd9, 32'sd19, 32'sd24, 32'sd9, 32'sd9, 32'sd18, 32'sd18, 32'sd3, 32'sd8, 32'sd18, 32'sd3, 32'sd4, 32'sd10, 32'sd6, 32'sd10, 32'sd5, 32'sd12, 32'sd9, 32'sd8, 32'sd5, 32'sd14, 32'sd10, 32'sd4, 32'sd6, 32'sd18, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd9, 32'sd14, 32'sd15, 32'sd8, 32'sd6, 32'sd6, 32'sd12, 32'sd12, 32'sd16, 32'sd18, 32'sd18, 32'sd24, 32'sd9, 32'sd24, 32'sd22, 32'sd9, 32'sd10, 32'sd6, 32'sd12, 32'sd12, 32'sd16, 32'sd10, 32'sd18, 32'sd9, 32'sd10, 32'sd18, 32'sd15, 32'sd15, 32'sd24, 32'sd6, 32'sd6, 32'sd6, 32'sd10, 32'sd18, 32'sd10, 32'sd10, 32'sd14, 32'sd9, 32'sd6, 32'sd6, 32'sd8, 32'sd4, 32'sd3, 32'sd16, 32'sd6, 32'sd6, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd4, 32'sd12, 32'sd12, 32'sd12, 32'sd14, 32'sd20, 32'sd8, 32'sd13, 32'sd6, 32'sd6, 32'sd12, 32'sd15, 32'sd12, 32'sd18, 32'sd24, 32'sd3, 32'sd4, 32'sd4, 32'sd12, 32'sd17, 32'sd5, 32'sd5, 32'sd18, 32'sd12, 32'sd6, 32'sd6, 32'sd21, 32'sd6, 32'sd12, 32'sd16, 32'sd18, 32'sd15, 32'sd9, 32'sd15, 32'sd3, 32'sd3, 32'sd10, 32'sd16, 32'sd12, 32'sd9, 32'sd6, 32'sd6, 32'sd10, 32'sd18, 32'sd14, 32'sd14, 32'sd3, 32'sd5, 32'sd12, 32'sd20, 32'sd19, 32'sd9, 32'sd14, 32'sd14, 32'sd9, 32'sd18, 32'sd6, 32'sd18, 32'sd20, 32'sd20, 32'sd24, 32'sd20, 32'sd9, 32'sd9, 32'sd8, 32'sd8, 32'sd4, 32'sd20, 32'sd6, 32'sd21, 32'sd13, 32'sd12, 32'sd10, 32'sd5, 32'sd6, 32'sd18, 32'sd9, 32'sd21, 32'sd22, 32'sd18, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd9, 32'sd9, 32'sd15, 32'sd3, 32'sd12, 32'sd20, 32'sd6, 32'sd18, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd16, 32'sd6, 32'sd6, 32'sd18, 32'sd10, 32'sd10, 32'sd9, 32'sd6, 32'sd5, 32'sd8, 32'sd19, 32'sd12, 32'sd21, 32'sd16, 32'sd18, 32'sd10, 32'sd4, 32'sd18, 32'sd12, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd12, 32'sd10, 32'sd10, 32'sd6, 32'sd6, 32'sd8, 32'sd12, 32'sd10, 32'sd10, 32'sd18, 32'sd4, 32'sd24, 32'sd6, 32'sd20, 32'sd19, 32'sd10, 32'sd21, 32'sd8, 32'sd10, 32'sd4, 32'sd6, 32'sd4, 32'sd4, 32'sd9, 32'sd16, 32'sd16, 32'sd24, 32'sd9, 32'sd14, 32'sd7, 32'sd8, 32'sd12, 32'sd4, 32'sd3, 32'sd9, 32'sd20, 32'sd24, 32'sd12, 32'sd8, 32'sd6, 32'sd10, 32'sd14, 32'sd10, 32'sd9, 32'sd24, 
                                                    32'sd12, 32'sd22, 32'sd12, 32'sd9, 32'sd23, 32'sd19, 32'sd6, 32'sd18, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd4, 32'sd8, 32'sd7, 32'sd18, 32'sd4, 32'sd4, 32'sd20, 32'sd6, 32'sd10, 32'sd4, 32'sd8, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd24, 32'sd10, 32'sd23, 32'sd19, 32'sd18, 32'sd9, 32'sd6, 32'sd6, 32'sd20, 32'sd6, 32'sd18, 32'sd9, 32'sd18, 32'sd18, 32'sd18, 32'sd10, 32'sd4, 32'sd4, 32'sd4, 32'sd12, 32'sd4, 32'sd10, 32'sd4, 32'sd3, 32'sd4, 32'sd6, 32'sd19, 32'sd9, 32'sd7, 32'sd14, 32'sd8, 32'sd8, 32'sd18, 32'sd9, 32'sd18, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd4, 32'sd18, 32'sd6, 32'sd8, 32'sd18, 32'sd14, 32'sd15, 32'sd10, 32'sd4, 32'sd22, 32'sd6, 32'sd6, 32'sd4, 32'sd10, 32'sd8, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd4, 32'sd19, 32'sd6, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd24, 32'sd10, 32'sd10, 32'sd19, 32'sd19, 32'sd16, 32'sd24, 32'sd6, 32'sd6, 32'sd18, 32'sd18, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd10, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd15, 32'sd20, 32'sd4, 32'sd12, 32'sd6, 32'sd9, 32'sd6, 32'sd12, 32'sd18, 32'sd18, 32'sd18, 32'sd6, 32'sd12, 32'sd18, 32'sd4, 32'sd19, 32'sd15, 32'sd14, 32'sd22, 32'sd6, 32'sd18, 32'sd3, 32'sd20, 32'sd5, 32'sd12, 32'sd6, 32'sd8, 32'sd8, 32'sd12, 32'sd6, 32'sd3, 32'sd14, 32'sd12, 32'sd4, 32'sd15, 32'sd6, 32'sd10, 32'sd18, 32'sd15, 32'sd8, 32'sd24, 32'sd6, 32'sd8, 32'sd10, 32'sd18, 32'sd24, 32'sd6, 32'sd8, 32'sd18, 32'sd18, 32'sd18, 32'sd20, 32'sd14, 32'sd12, 32'sd21, 32'sd21, 32'sd18, 32'sd18, 32'sd4, 32'sd18, 32'sd4, 32'sd10, 32'sd11, 32'sd4, 32'sd9, 32'sd4, 32'sd8, 32'sd8, 32'sd12, 32'sd9, 32'sd12, 32'sd9, 32'sd12, 32'sd4, 32'sd14, 32'sd11, 32'sd6, 32'sd11, 32'sd9, 32'sd18, 32'sd12, 32'sd18, 32'sd18, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd18, 32'sd6, 32'sd15, 32'sd15, 32'sd4, 32'sd6, 32'sd8, 32'sd8, 32'sd24, 32'sd14, 32'sd8, 32'sd10, 32'sd8, 32'sd4, 32'sd6, 32'sd6, 32'sd18, 32'sd16, 32'sd16, 32'sd8, 32'sd16, 32'sd12, 32'sd9, 32'sd9, 32'sd16, 32'sd19, 32'sd9, 32'sd3, 32'sd24, 32'sd5, 32'sd19, 32'sd6, 32'sd24, 32'sd9, 32'sd10, 32'sd20, 32'sd7, 32'sd7, 32'sd2, 32'sd10, 32'sd12, 32'sd3, 32'sd12, 32'sd6, 32'sd9, 32'sd22, 32'sd22, 32'sd9, 32'sd4, 32'sd18, 32'sd24, 32'sd24, 32'sd18, 32'sd4, 32'sd10, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd10, 32'sd10, 32'sd9, 32'sd14, 32'sd10, 32'sd10, 32'sd3, 32'sd9, 32'sd5, 32'sd24, 32'sd12, 32'sd4, 32'sd9, 32'sd6, 32'sd6, 32'sd19, 32'sd4, 32'sd6, 32'sd18, 32'sd10, 32'sd18, 32'sd9, 32'sd24, 32'sd8, 32'sd4, 32'sd8, 32'sd10, 32'sd18, 32'sd19, 32'sd24, 32'sd8, 32'sd10, 32'sd6, 32'sd7, 32'sd12, 32'sd6, 32'sd15, 32'sd6, 32'sd7, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd9, 32'sd18, 32'sd9, 32'sd9, 32'sd18, 32'sd18, 32'sd4, 32'sd4, 32'sd2, 32'sd16, 32'sd4, 32'sd10, 32'sd6, 32'sd7, 32'sd4, 32'sd6, 32'sd10, 32'sd18, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd18, 32'sd9, 32'sd9, 32'sd10, 32'sd5, 32'sd5, 32'sd4, 32'sd4, 32'sd10, 32'sd14, 32'sd12, 32'sd24, 32'sd14, 32'sd6, 32'sd4, 32'sd14, 32'sd16, 32'sd21, 32'sd15, 32'sd6, 32'sd16, 32'sd16, 32'sd3, 32'sd3, 32'sd10, 32'sd6, 32'sd12, 32'sd5, 32'sd9, 32'sd11, 32'sd4, 32'sd9, 32'sd13, 32'sd4, 32'sd6, 32'sd10, 32'sd20, 32'sd9, 32'sd4, 32'sd4, 32'sd22, 32'sd9, 32'sd24, 32'sd16, 32'sd18, 32'sd6, 32'sd9, 32'sd9, 32'sd4, 32'sd7, 32'sd20, 32'sd19, 32'sd6, 32'sd6, 32'sd4, 32'sd9, 32'sd18, 32'sd2, 32'sd8, 32'sd18, 32'sd15, 32'sd12, 32'sd6, 32'sd20, 32'sd24, 32'sd9, 32'sd4, 32'sd4, 32'sd8, 32'sd6, 32'sd3, 32'sd12, 32'sd5, 32'sd5, 32'sd6, 32'sd6, 32'sd14, 32'sd3, 32'sd6, 32'sd4, 32'sd16, 32'sd7, 32'sd8, 32'sd6, 32'sd9, 32'sd3, 32'sd22, 32'sd18, 32'sd6, 32'sd9, 32'sd4, 32'sd4, 32'sd10, 32'sd3, 32'sd18, 32'sd18, 32'sd9, 32'sd9, 32'sd18, 32'sd6, 32'sd10, 32'sd18, 32'sd18, 32'sd9, 32'sd6, 32'sd18, 32'sd9, 32'sd10, 32'sd9, 32'sd3, 32'sd9, 32'sd11, 32'sd9, 32'sd11, 32'sd8, 32'sd20, 32'sd21, 32'sd12, 32'sd6, 32'sd8, 32'sd8, 32'sd8, 32'sd9, 32'sd8, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd10, 32'sd6, 32'sd6, 32'sd10, 32'sd16, 32'sd19, 32'sd18, 32'sd9, 32'sd6, 32'sd6, 32'sd14, 32'sd8, 32'sd7, 32'sd12, 32'sd8, 32'sd22, 32'sd6, 32'sd6, 32'sd6, 32'sd17, 32'sd12, 32'sd18, 32'sd10, 32'sd10, 32'sd24, 32'sd6, 32'sd6, 32'sd19, 32'sd6, 32'sd10, 32'sd10, 32'sd9, 32'sd18, 32'sd18, 32'sd9, 32'sd9, 32'sd6, 32'sd4, 32'sd8, 32'sd18, 32'sd4, 32'sd12, 32'sd4, 32'sd18, 32'sd18, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd12, 32'sd4, 32'sd6, 32'sd12, 32'sd8, 32'sd8, 32'sd9, 32'sd9, 32'sd18, 32'sd9, 32'sd18, 32'sd6, 32'sd9, 32'sd9, 32'sd14, 32'sd6, 32'sd12, 32'sd18, 32'sd6, 32'sd16, 32'sd3, 32'sd6, 32'sd4, 32'sd4, 32'sd5, 32'sd9, 32'sd18, 32'sd5, 32'sd17, 32'sd18, 32'sd24, 32'sd18, 32'sd6, 32'sd14, 32'sd3, 32'sd6, 32'sd6, 32'sd6, 32'sd21, 32'sd12, 32'sd9, 32'sd6, 32'sd8, 32'sd8, 32'sd8, 32'sd8, 32'sd12, 32'sd18, 32'sd20, 32'sd9, 32'sd8, 32'sd16, 32'sd10, 32'sd10, 32'sd15, 32'sd18, 32'sd10, 32'sd18, 32'sd10, 32'sd10, 32'sd18, 32'sd18, 32'sd18, 32'sd6, 32'sd8, 32'sd8, 32'sd8, 32'sd18, 32'sd9, 32'sd18, 32'sd6, 32'sd6, 32'sd18, 32'sd12, 32'sd6, 32'sd2, 32'sd10, 32'sd20, 32'sd12, 32'sd3, 32'sd3, 32'sd3, 32'sd18, 32'sd10, 32'sd14, 32'sd14, 32'sd9, 32'sd8, 32'sd4, 32'sd5, 32'sd9, 32'sd9, 32'sd12, 32'sd5, 32'sd3, 32'sd6, 32'sd7, 32'sd4, 32'sd14, 32'sd19, 32'sd6, 32'sd15, 32'sd10, 32'sd8, 32'sd12, 32'sd9, 32'sd14, 32'sd14, 32'sd13, 32'sd6, 32'sd17, 32'sd17, 32'sd8, 32'sd8, 32'sd24, 32'sd15, 32'sd18, 32'sd18, 32'sd3, 32'sd3, 32'sd6, 32'sd6, 32'sd11, 32'sd12, 32'sd12, 32'sd9, 32'sd12, 32'sd6, 32'sd9, 32'sd6, 32'sd9, 32'sd16, 32'sd10, 32'sd7, 32'sd11, 32'sd12, 32'sd8, 32'sd4, 32'sd3, 32'sd3, 32'sd18, 32'sd4, 32'sd3, 32'sd18, 32'sd3, 32'sd3, 32'sd5, 32'sd18, 32'sd20, 32'sd9, 32'sd19, 32'sd19, 32'sd9, 32'sd18, 32'sd14, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 
                                                    32'sd6, 32'sd12, 32'sd12, 32'sd4, 32'sd6, 32'sd3, 32'sd18, 32'sd16, 32'sd10, 32'sd9, 32'sd9, 32'sd10, 32'sd3, 32'sd12, 32'sd12, 32'sd8, 32'sd6, 32'sd12, 32'sd12, 32'sd6, 32'sd7, 32'sd18, 32'sd19, 32'sd12, 32'sd6, 32'sd6, 32'sd5, 32'sd5, 32'sd14, 32'sd3, 32'sd24, 32'sd20, 32'sd18, 32'sd6, 32'sd20, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd15, 32'sd18, 32'sd3, 32'sd6, 32'sd6, 32'sd8, 32'sd8, 32'sd20, 32'sd13, 32'sd7, 32'sd7, 32'sd10, 32'sd10, 32'sd3, 32'sd18, 32'sd18, 32'sd9, 32'sd15, 32'sd12, 32'sd12, 32'sd6, 32'sd13, 32'sd22, 32'sd6, 32'sd6, 32'sd24, 32'sd10, 32'sd18, 32'sd10, 32'sd3, 32'sd12, 32'sd4, 32'sd4, 32'sd18, 32'sd9, 32'sd12, 32'sd9, 32'sd10, 32'sd10, 32'sd10, 32'sd10, 32'sd9, 32'sd9, 32'sd10, 32'sd10, 32'sd18, 32'sd18, 32'sd18, 32'sd7, 32'sd19, 32'sd16, 32'sd16, 32'sd12, 32'sd2, 32'sd2, 32'sd8, 32'sd8, 32'sd3, 32'sd12, 32'sd8, 32'sd12, 32'sd18, 32'sd18, 32'sd3, 32'sd18, 32'sd3, 32'sd3, 32'sd18, 32'sd18, 32'sd22, 32'sd21, 32'sd18, 32'sd18, 32'sd24, 32'sd16, 32'sd6, 32'sd8, 32'sd6, 32'sd6, 32'sd18, 32'sd10, 32'sd9, 32'sd9, 32'sd3, 32'sd3, 32'sd6, 32'sd6, 32'sd16, 32'sd9, 32'sd16, 32'sd18, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd18, 32'sd24, 32'sd9, 32'sd8, 32'sd13, 32'sd16, 32'sd14, 32'sd9, 32'sd16, 32'sd13, 32'sd13, 32'sd24, 32'sd10, 32'sd18, 32'sd18, 32'sd9, 32'sd22, 32'sd8, 32'sd8, 32'sd18, 32'sd5, 32'sd12, 32'sd18, 32'sd4, 32'sd6, 32'sd2, 32'sd2, 32'sd10, 32'sd18, 32'sd17, 32'sd12, 32'sd16, 32'sd5, 32'sd6, 32'sd6, 32'sd6, 32'sd13, 32'sd19, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd4, 32'sd8, 32'sd8, 32'sd10, 32'sd10, 32'sd4, 32'sd4, 32'sd16, 32'sd16, 32'sd7, 32'sd3, 32'sd9, 32'sd17, 32'sd8, 32'sd8, 32'sd10, 32'sd22, 32'sd24, 32'sd12, 32'sd6, 32'sd6, 32'sd9, 32'sd22, 32'sd9, 32'sd18, 32'sd19, 32'sd18, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd3, 32'sd24, 32'sd6}

localparam logic [2912:0][31:0] rectangle1_heights = {32'sd9, 32'sd7, 32'sd9, 32'sd6, 32'sd19, 32'sd16, 32'sd6, 32'sd10, 32'sd6, 32'sd6, 32'sd7, 32'sd12, 32'sd3, 32'sd15, 32'sd10, 32'sd9, 32'sd6, 32'sd10, 32'sd10, 32'sd9, 32'sd11, 32'sd13, 32'sd9, 32'sd6, 32'sd12, 32'sd3, 32'sd6, 32'sd14, 32'sd10, 32'sd12, 32'sd3, 32'sd6, 32'sd15, 32'sd15, 32'sd15, 32'sd12, 32'sd12, 32'sd10, 32'sd10, 32'sd13, 32'sd13, 32'sd19, 32'sd9, 32'sd11, 32'sd9, 32'sd3, 32'sd9, 32'sd9, 32'sd14, 32'sd2, 32'sd11, 32'sd9, 32'sd9, 32'sd6, 32'sd5, 32'sd6, 32'sd6, 32'sd13, 32'sd13, 32'sd23, 32'sd12, 32'sd14, 32'sd6, 32'sd6, 32'sd12, 32'sd6, 32'sd3, 32'sd12, 32'sd20, 32'sd2, 32'sd14, 32'sd12, 32'sd9, 32'sd6, 32'sd6, 32'sd10, 32'sd14, 32'sd5, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd4, 32'sd9, 32'sd6, 32'sd12, 32'sd6, 32'sd3, 32'sd9, 32'sd4, 32'sd9, 32'sd9, 32'sd12, 32'sd2, 32'sd10, 32'sd10, 32'sd6, 32'sd4, 32'sd2, 32'sd3, 32'sd3, 32'sd15, 32'sd10, 32'sd10, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd10, 32'sd3, 32'sd2, 32'sd12, 32'sd24, 32'sd10, 32'sd12, 32'sd12, 32'sd3, 32'sd8, 32'sd6, 32'sd6, 32'sd18, 32'sd14, 32'sd2, 32'sd13, 32'sd4, 32'sd10, 32'sd6, 32'sd6, 32'sd12, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd15, 32'sd9, 32'sd10, 32'sd8, 32'sd7, 32'sd22, 32'sd22, 32'sd16, 32'sd6, 32'sd12, 32'sd6, 32'sd14, 32'sd10, 32'sd11, 32'sd11, 32'sd18, 32'sd14, 32'sd8, 32'sd14, 32'sd6, 32'sd16, 32'sd6, 32'sd4, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd3, 32'sd3, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd12, 32'sd17, 32'sd24, 32'sd24, 32'sd22, 32'sd22, 32'sd18, 32'sd6, 32'sd4, 32'sd3, 32'sd18, 32'sd3, 32'sd4, 32'sd6, 32'sd6, 32'sd16, 32'sd16, 32'sd9, 32'sd8, 32'sd9, 32'sd3, 32'sd2, 32'sd9, 32'sd18, 32'sd9, 32'sd12, 32'sd2, 32'sd3, 32'sd9, 32'sd4, 32'sd4, 32'sd11, 32'sd6, 32'sd10, 32'sd12, 32'sd15, 32'sd3, 32'sd9, 32'sd6, 32'sd9, 32'sd14, 32'sd13, 32'sd13, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd9, 32'sd4, 32'sd6, 32'sd10, 32'sd14, 32'sd9, 32'sd3, 32'sd3, 32'sd4, 32'sd6, 32'sd18, 32'sd18, 32'sd10, 32'sd4, 32'sd18, 32'sd6, 32'sd8, 32'sd9, 32'sd19, 32'sd3, 32'sd4, 32'sd4, 32'sd16, 32'sd4, 32'sd6, 32'sd9, 32'sd15, 32'sd13, 32'sd14, 32'sd10, 32'sd6, 32'sd14, 32'sd12, 32'sd5, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd16, 32'sd6, 32'sd9, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd9, 32'sd3, 32'sd21, 32'sd12, 32'sd9, 32'sd20, 32'sd9, 32'sd21, 32'sd23, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd4, 32'sd19, 32'sd12, 32'sd10, 32'sd12, 32'sd19, 32'sd10, 32'sd12, 32'sd2, 32'sd4, 32'sd9, 32'sd4, 32'sd9, 32'sd9, 32'sd4, 32'sd9, 32'sd9, 32'sd9, 32'sd15, 32'sd15, 32'sd4, 32'sd7, 32'sd10, 32'sd8, 32'sd16, 32'sd3, 32'sd3, 32'sd9, 32'sd18, 32'sd18, 32'sd9, 32'sd14, 32'sd6, 32'sd16, 32'sd12, 32'sd16, 32'sd10, 32'sd3, 32'sd10, 32'sd4, 32'sd9, 32'sd5, 32'sd12, 32'sd10, 32'sd14, 32'sd16, 32'sd8, 32'sd2, 32'sd6, 32'sd9, 32'sd14, 32'sd12, 32'sd18, 32'sd18, 32'sd9, 32'sd6, 32'sd9, 32'sd9, 32'sd2, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd15, 32'sd6, 32'sd14, 32'sd6, 32'sd4, 32'sd19, 32'sd19, 32'sd9, 32'sd3, 32'sd9, 32'sd4, 32'sd6, 32'sd22, 32'sd14, 32'sd20, 32'sd9, 32'sd9, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd3, 32'sd3, 32'sd6, 32'sd12, 32'sd12, 32'sd12, 32'sd9, 32'sd12, 32'sd12, 32'sd8, 32'sd9, 32'sd3, 32'sd6, 32'sd23, 32'sd4, 32'sd18, 32'sd6, 32'sd6, 32'sd4, 32'sd9, 32'sd3, 32'sd4, 32'sd12, 32'sd3, 32'sd6, 32'sd3, 32'sd9, 32'sd9, 32'sd12, 32'sd4, 32'sd9, 32'sd10, 32'sd9, 32'sd21, 32'sd7, 32'sd9, 32'sd4, 32'sd12, 32'sd12, 32'sd9, 32'sd17, 32'sd9, 32'sd6, 32'sd19, 32'sd7, 32'sd12, 32'sd12, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd14, 32'sd14, 32'sd6, 32'sd5, 32'sd11, 32'sd14, 32'sd9, 32'sd6, 32'sd9, 32'sd9, 32'sd4, 32'sd2, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd7, 32'sd10, 32'sd9, 32'sd9, 32'sd3, 32'sd3, 32'sd12, 32'sd6, 32'sd4, 32'sd2, 32'sd24, 32'sd4, 32'sd9, 32'sd12, 32'sd6, 32'sd3, 32'sd16, 32'sd4, 32'sd2, 32'sd8, 32'sd6, 32'sd6, 32'sd10, 32'sd10, 32'sd4, 32'sd3, 32'sd6, 32'sd6, 32'sd3, 32'sd10, 32'sd24, 32'sd11, 32'sd6, 32'sd20, 32'sd24, 32'sd24, 32'sd14, 32'sd12, 32'sd14, 32'sd6, 32'sd9, 32'sd14, 32'sd15, 32'sd9, 32'sd14, 32'sd18, 32'sd6, 32'sd10, 32'sd9, 32'sd7, 32'sd3, 32'sd6, 32'sd12, 32'sd18, 32'sd9, 32'sd13, 32'sd3, 32'sd12, 32'sd10, 32'sd8, 32'sd9, 32'sd5, 32'sd5, 32'sd6, 32'sd3, 32'sd6, 32'sd12, 32'sd15, 32'sd10, 32'sd12, 32'sd6, 32'sd6, 32'sd16, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd3, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd10, 32'sd16, 32'sd5, 32'sd5, 32'sd10, 32'sd6, 32'sd18, 32'sd9, 32'sd7, 32'sd10, 32'sd18, 32'sd9, 32'sd6, 32'sd3, 32'sd9, 32'sd10, 32'sd12, 32'sd12, 32'sd21, 32'sd8, 32'sd8, 32'sd3, 32'sd4, 32'sd9, 32'sd9, 32'sd22, 32'sd14, 32'sd15, 32'sd14, 32'sd14, 32'sd6, 32'sd9, 32'sd16, 32'sd16, 32'sd8, 32'sd9, 32'sd3, 32'sd9, 32'sd6, 32'sd10, 32'sd18, 32'sd3, 32'sd11, 32'sd11, 32'sd9, 32'sd9, 32'sd9, 32'sd4, 32'sd6, 32'sd6, 32'sd17, 32'sd17, 32'sd4, 32'sd18, 32'sd12, 32'sd12, 32'sd15, 32'sd15, 32'sd6, 32'sd6, 32'sd14, 32'sd9, 32'sd15, 32'sd15, 32'sd9, 32'sd21, 32'sd12, 32'sd12, 32'sd18, 32'sd9, 32'sd3, 32'sd10, 32'sd4, 32'sd20, 32'sd8, 32'sd8, 32'sd9, 32'sd3, 32'sd4, 32'sd6, 32'sd6, 32'sd10, 32'sd7, 32'sd6, 32'sd3, 32'sd18, 32'sd6, 32'sd6, 32'sd3, 32'sd7, 32'sd6, 32'sd6, 32'sd7, 32'sd12, 32'sd4, 32'sd9, 32'sd9, 32'sd15, 32'sd3, 32'sd6, 32'sd11, 32'sd9, 32'sd9, 32'sd4, 32'sd6, 32'sd10, 32'sd16, 32'sd4, 32'sd9, 32'sd8, 32'sd8, 32'sd18, 32'sd11, 32'sd5, 32'sd3, 32'sd3, 32'sd6, 32'sd10, 32'sd3, 32'sd3, 32'sd22, 32'sd6, 32'sd6, 32'sd12, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd9, 32'sd19, 32'sd6, 32'sd19, 32'sd9, 32'sd3, 32'sd4, 32'sd10, 32'sd6, 32'sd8, 32'sd12, 32'sd6, 32'sd19, 32'sd20, 32'sd20, 32'sd6, 32'sd6, 32'sd14, 32'sd14, 32'sd7, 32'sd9, 32'sd10, 32'sd10, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd10, 
                                                    32'sd10, 32'sd13, 32'sd5, 32'sd6, 32'sd4, 32'sd5, 32'sd12, 32'sd6, 32'sd3, 32'sd9, 32'sd2, 32'sd18, 32'sd3, 32'sd3, 32'sd18, 32'sd23, 32'sd19, 32'sd9, 32'sd6, 32'sd12, 32'sd6, 32'sd10, 32'sd15, 32'sd6, 32'sd8, 32'sd6, 32'sd6, 32'sd18, 32'sd18, 32'sd4, 32'sd4, 32'sd9, 32'sd8, 32'sd5, 32'sd8, 32'sd4, 32'sd15, 32'sd8, 32'sd4, 32'sd4, 32'sd17, 32'sd18, 32'sd12, 32'sd9, 32'sd12, 32'sd2, 32'sd6, 32'sd11, 32'sd10, 32'sd17, 32'sd6, 32'sd9, 32'sd12, 32'sd12, 32'sd15, 32'sd3, 32'sd7, 32'sd9, 32'sd3, 32'sd12, 32'sd14, 32'sd9, 32'sd18, 32'sd18, 32'sd10, 32'sd11, 32'sd3, 32'sd3, 32'sd12, 32'sd8, 32'sd12, 32'sd14, 32'sd10, 32'sd2, 32'sd12, 32'sd12, 32'sd18, 32'sd18, 32'sd12, 32'sd9, 32'sd11, 32'sd12, 32'sd3, 32'sd3, 32'sd4, 32'sd5, 32'sd4, 32'sd9, 32'sd6, 32'sd6, 32'sd8, 32'sd18, 32'sd10, 32'sd5, 32'sd6, 32'sd14, 32'sd4, 32'sd4, 32'sd10, 32'sd3, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd3, 32'sd4, 32'sd3, 32'sd6, 32'sd6, 32'sd3, 32'sd10, 32'sd9, 32'sd8, 32'sd8, 32'sd11, 32'sd9, 32'sd6, 32'sd12, 32'sd12, 32'sd8, 32'sd3, 32'sd4, 32'sd22, 32'sd8, 32'sd9, 32'sd9, 32'sd14, 32'sd8, 32'sd14, 32'sd20, 32'sd10, 32'sd4, 32'sd4, 32'sd9, 32'sd5, 32'sd4, 32'sd4, 32'sd5, 32'sd10, 32'sd8, 32'sd3, 32'sd4, 32'sd6, 32'sd4, 32'sd12, 32'sd6, 32'sd9, 32'sd4, 32'sd3, 32'sd9, 32'sd4, 32'sd18, 32'sd12, 32'sd8, 32'sd5, 32'sd6, 32'sd9, 32'sd12, 32'sd6, 32'sd6, 32'sd15, 32'sd2, 32'sd6, 32'sd2, 32'sd6, 32'sd3, 32'sd5, 32'sd9, 32'sd9, 32'sd9, 32'sd4, 32'sd6, 32'sd6, 32'sd3, 32'sd12, 32'sd6, 32'sd3, 32'sd10, 32'sd6, 32'sd9, 32'sd14, 32'sd6, 32'sd8, 32'sd12, 32'sd10, 32'sd6, 32'sd9, 32'sd12, 32'sd9, 32'sd6, 32'sd3, 32'sd6, 32'sd6, 32'sd14, 32'sd9, 32'sd14, 32'sd16, 32'sd10, 32'sd5, 32'sd3, 32'sd12, 32'sd5, 32'sd4, 32'sd12, 32'sd6, 32'sd6, 32'sd13, 32'sd13, 32'sd6, 32'sd3, 32'sd6, 32'sd14, 32'sd2, 32'sd4, 32'sd4, 32'sd9, 32'sd4, 32'sd6, 32'sd23, 32'sd23, 32'sd3, 32'sd4, 32'sd3, 32'sd4, 32'sd15, 32'sd3, 32'sd4, 32'sd4, 32'sd9, 32'sd6, 32'sd10, 32'sd6, 32'sd6, 32'sd6, 32'sd2, 32'sd6, 32'sd3, 32'sd6, 32'sd3, 32'sd16, 32'sd6, 32'sd22, 32'sd10, 32'sd18, 32'sd9, 32'sd10, 32'sd9, 32'sd10, 32'sd10, 32'sd10, 32'sd9, 32'sd3, 32'sd13, 32'sd13, 32'sd7, 32'sd9, 32'sd6, 32'sd6, 32'sd2, 32'sd16, 32'sd6, 32'sd12, 32'sd3, 32'sd6, 32'sd4, 32'sd14, 32'sd6, 32'sd9, 32'sd10, 32'sd10, 32'sd6, 32'sd9, 32'sd14, 32'sd12, 32'sd12, 32'sd9, 32'sd16, 32'sd6, 32'sd14, 32'sd2, 32'sd16, 32'sd10, 32'sd4, 32'sd7, 32'sd16, 32'sd16, 32'sd6, 32'sd12, 32'sd8, 32'sd18, 32'sd14, 32'sd14, 32'sd6, 32'sd18, 32'sd3, 32'sd9, 32'sd6, 32'sd16, 32'sd4, 32'sd16, 32'sd16, 32'sd10, 32'sd8, 32'sd2, 32'sd9, 32'sd8, 32'sd3, 32'sd11, 32'sd9, 32'sd8, 32'sd6, 32'sd3, 32'sd6, 32'sd9, 32'sd9, 32'sd19, 32'sd19, 32'sd8, 32'sd8, 32'sd3, 32'sd4, 32'sd6, 32'sd6, 32'sd14, 32'sd12, 32'sd5, 32'sd9, 32'sd9, 32'sd8, 32'sd6, 32'sd3, 32'sd12, 32'sd12, 32'sd2, 32'sd3, 32'sd14, 32'sd14, 32'sd14, 32'sd6, 32'sd9, 32'sd4, 32'sd6, 32'sd3, 32'sd9, 32'sd4, 32'sd5, 32'sd9, 32'sd10, 32'sd10, 32'sd9, 32'sd9, 32'sd19, 32'sd9, 32'sd19, 32'sd4, 32'sd9, 32'sd19, 32'sd12, 32'sd5, 32'sd18, 32'sd12, 32'sd3, 32'sd3, 32'sd4, 32'sd9, 32'sd4, 32'sd4, 32'sd6, 32'sd8, 32'sd3, 32'sd6, 32'sd5, 32'sd5, 32'sd6, 32'sd15, 32'sd12, 32'sd14, 32'sd6, 32'sd6, 32'sd4, 32'sd3, 32'sd4, 32'sd3, 32'sd4, 32'sd3, 32'sd4, 32'sd6, 32'sd9, 32'sd4, 32'sd12, 32'sd3, 32'sd6, 32'sd7, 32'sd8, 32'sd3, 32'sd6, 32'sd9, 32'sd4, 32'sd6, 32'sd10, 32'sd10, 32'sd17, 32'sd20, 32'sd4, 32'sd9, 32'sd9, 32'sd16, 32'sd4, 32'sd4, 32'sd6, 32'sd10, 32'sd6, 32'sd8, 32'sd8, 32'sd8, 32'sd4, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd18, 32'sd4, 32'sd14, 32'sd6, 32'sd3, 32'sd4, 32'sd15, 32'sd3, 32'sd6, 32'sd9, 32'sd9, 32'sd9, 32'sd21, 32'sd2, 32'sd3, 32'sd13, 32'sd8, 32'sd9, 32'sd9, 32'sd10, 32'sd10, 32'sd6, 32'sd6, 32'sd21, 32'sd13, 32'sd21, 32'sd20, 32'sd6, 32'sd9, 32'sd9, 32'sd3, 32'sd9, 32'sd10, 32'sd9, 32'sd9, 32'sd4, 32'sd14, 32'sd6, 32'sd12, 32'sd10, 32'sd8, 32'sd6, 32'sd9, 32'sd14, 32'sd6, 32'sd9, 32'sd10, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd11, 32'sd6, 32'sd11, 32'sd11, 32'sd9, 32'sd4, 32'sd12, 32'sd3, 32'sd9, 32'sd3, 32'sd9, 32'sd3, 32'sd9, 32'sd9, 32'sd18, 32'sd18, 32'sd9, 32'sd6, 32'sd3, 32'sd9, 32'sd3, 32'sd16, 32'sd4, 32'sd8, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd10, 32'sd8, 32'sd15, 32'sd8, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd2, 32'sd11, 32'sd15, 32'sd13, 32'sd9, 32'sd9, 32'sd4, 32'sd4, 32'sd4, 32'sd3, 32'sd3, 32'sd20, 32'sd6, 32'sd4, 32'sd7, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd9, 32'sd8, 32'sd8, 32'sd9, 32'sd16, 32'sd12, 32'sd12, 32'sd6, 32'sd22, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd10, 32'sd16, 32'sd6, 32'sd10, 32'sd6, 32'sd2, 32'sd6, 32'sd10, 32'sd6, 32'sd4, 32'sd16, 32'sd13, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd11, 32'sd10, 32'sd10, 32'sd21, 32'sd9, 32'sd6, 32'sd16, 32'sd3, 32'sd12, 32'sd9, 32'sd8, 32'sd2, 32'sd3, 32'sd6, 32'sd18, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd2, 32'sd4, 32'sd12, 32'sd12, 32'sd22, 32'sd22, 32'sd11, 32'sd11, 32'sd9, 32'sd3, 32'sd2, 32'sd2, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd10, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd3, 32'sd6, 32'sd6, 32'sd3, 32'sd6, 32'sd10, 32'sd6, 32'sd10, 32'sd12, 32'sd10, 32'sd9, 32'sd18, 32'sd4, 32'sd10, 32'sd10, 32'sd14, 32'sd19, 32'sd6, 32'sd6, 32'sd10, 32'sd8, 32'sd6, 32'sd18, 32'sd12, 32'sd8, 32'sd3, 32'sd3, 32'sd9, 32'sd4, 32'sd12, 32'sd9, 32'sd8, 32'sd7, 32'sd9, 32'sd12, 32'sd6, 32'sd9, 32'sd23, 32'sd6, 32'sd3, 32'sd14, 32'sd12, 32'sd12, 32'sd7, 32'sd9, 32'sd12, 32'sd12, 32'sd15, 32'sd15, 32'sd9, 32'sd15, 32'sd8, 32'sd4, 32'sd19, 32'sd19, 32'sd20, 32'sd20, 32'sd12, 32'sd12, 32'sd14, 32'sd8, 32'sd12, 32'sd5, 32'sd3, 32'sd12, 32'sd3, 32'sd3, 32'sd9, 32'sd6, 32'sd4, 32'sd14, 32'sd6, 32'sd9, 32'sd6, 32'sd10, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 
                                                    32'sd6, 32'sd3, 32'sd6, 32'sd24, 32'sd4, 32'sd12, 32'sd8, 32'sd14, 32'sd14, 32'sd10, 32'sd6, 32'sd9, 32'sd7, 32'sd10, 32'sd9, 32'sd12, 32'sd14, 32'sd8, 32'sd8, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd8, 32'sd8, 32'sd12, 32'sd11, 32'sd4, 32'sd7, 32'sd3, 32'sd9, 32'sd7, 32'sd6, 32'sd11, 32'sd11, 32'sd18, 32'sd5, 32'sd3, 32'sd20, 32'sd4, 32'sd4, 32'sd10, 32'sd14, 32'sd8, 32'sd9, 32'sd8, 32'sd6, 32'sd4, 32'sd9, 32'sd8, 32'sd17, 32'sd6, 32'sd17, 32'sd17, 32'sd3, 32'sd18, 32'sd18, 32'sd18, 32'sd8, 32'sd9, 32'sd9, 32'sd8, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd3, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd9, 32'sd9, 32'sd23, 32'sd3, 32'sd4, 32'sd23, 32'sd3, 32'sd3, 32'sd4, 32'sd6, 32'sd3, 32'sd6, 32'sd4, 32'sd15, 32'sd12, 32'sd9, 32'sd9, 32'sd9, 32'sd3, 32'sd6, 32'sd13, 32'sd4, 32'sd13, 32'sd18, 32'sd5, 32'sd8, 32'sd9, 32'sd9, 32'sd14, 32'sd14, 32'sd16, 32'sd10, 32'sd6, 32'sd4, 32'sd5, 32'sd5, 32'sd16, 32'sd16, 32'sd15, 32'sd2, 32'sd6, 32'sd4, 32'sd12, 32'sd12, 32'sd8, 32'sd8, 32'sd5, 32'sd8, 32'sd6, 32'sd18, 32'sd14, 32'sd14, 32'sd12, 32'sd16, 32'sd21, 32'sd21, 32'sd18, 32'sd8, 32'sd12, 32'sd12, 32'sd20, 32'sd6, 32'sd20, 32'sd20, 32'sd14, 32'sd14, 32'sd8, 32'sd9, 32'sd10, 32'sd11, 32'sd16, 32'sd6, 32'sd9, 32'sd12, 32'sd9, 32'sd10, 32'sd3, 32'sd2, 32'sd3, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd12, 32'sd6, 32'sd4, 32'sd16, 32'sd9, 32'sd9, 32'sd10, 32'sd6, 32'sd8, 32'sd21, 32'sd9, 32'sd3, 32'sd10, 32'sd3, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd12, 32'sd15, 32'sd4, 32'sd8, 32'sd10, 32'sd10, 32'sd12, 32'sd8, 32'sd4, 32'sd4, 32'sd6, 32'sd2, 32'sd9, 32'sd9, 32'sd10, 32'sd13, 32'sd6, 32'sd3, 32'sd6, 32'sd5, 32'sd9, 32'sd9, 32'sd7, 32'sd6, 32'sd6, 32'sd4, 32'sd18, 32'sd9, 32'sd14, 32'sd6, 32'sd9, 32'sd3, 32'sd6, 32'sd9, 32'sd6, 32'sd10, 32'sd3, 32'sd6, 32'sd9, 32'sd11, 32'sd11, 32'sd10, 32'sd18, 32'sd6, 32'sd3, 32'sd6, 32'sd5, 32'sd9, 32'sd9, 32'sd15, 32'sd3, 32'sd6, 32'sd3, 32'sd6, 32'sd6, 32'sd8, 32'sd3, 32'sd6, 32'sd4, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd10, 32'sd4, 32'sd6, 32'sd10, 32'sd6, 32'sd8, 32'sd6, 32'sd4, 32'sd10, 32'sd8, 32'sd12, 32'sd12, 32'sd9, 32'sd12, 32'sd16, 32'sd6, 32'sd2, 32'sd9, 32'sd9, 32'sd13, 32'sd2, 32'sd6, 32'sd24, 32'sd24, 32'sd10, 32'sd6, 32'sd3, 32'sd11, 32'sd4, 32'sd18, 32'sd16, 32'sd16, 32'sd6, 32'sd2, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd7, 32'sd7, 32'sd6, 32'sd8, 32'sd3, 32'sd3, 32'sd14, 32'sd10, 32'sd12, 32'sd18, 32'sd9, 32'sd9, 32'sd10, 32'sd12, 32'sd12, 32'sd10, 32'sd2, 32'sd13, 32'sd3, 32'sd12, 32'sd15, 32'sd4, 32'sd3, 32'sd8, 32'sd6, 32'sd3, 32'sd4, 32'sd6, 32'sd5, 32'sd7, 32'sd10, 32'sd10, 32'sd6, 32'sd9, 32'sd6, 32'sd16, 32'sd22, 32'sd12, 32'sd18, 32'sd18, 32'sd4, 32'sd4, 32'sd6, 32'sd9, 32'sd9, 32'sd9, 32'sd3, 32'sd13, 32'sd4, 32'sd6, 32'sd3, 32'sd12, 32'sd9, 32'sd13, 32'sd2, 32'sd9, 32'sd9, 32'sd8, 32'sd8, 32'sd8, 32'sd6, 32'sd15, 32'sd12, 32'sd9, 32'sd4, 32'sd3, 32'sd6, 32'sd6, 32'sd6, 32'sd8, 32'sd6, 32'sd3, 32'sd3, 32'sd5, 32'sd3, 32'sd6, 32'sd10, 32'sd10, 32'sd12, 32'sd6, 32'sd2, 32'sd10, 32'sd12, 32'sd12, 32'sd9, 32'sd11, 32'sd13, 32'sd6, 32'sd12, 32'sd3, 32'sd6, 32'sd3, 32'sd10, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd9, 32'sd9, 32'sd16, 32'sd16, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd16, 32'sd12, 32'sd6, 32'sd20, 32'sd9, 32'sd9, 32'sd9, 32'sd4, 32'sd12, 32'sd9, 32'sd4, 32'sd9, 32'sd8, 32'sd16, 32'sd6, 32'sd15, 32'sd8, 32'sd4, 32'sd6, 32'sd10, 32'sd21, 32'sd21, 32'sd3, 32'sd6, 32'sd2, 32'sd2, 32'sd4, 32'sd4, 32'sd2, 32'sd3, 32'sd23, 32'sd6, 32'sd3, 32'sd23, 32'sd10, 32'sd12, 32'sd14, 32'sd9, 32'sd12, 32'sd10, 32'sd4, 32'sd10, 32'sd12, 32'sd24, 32'sd4, 32'sd10, 32'sd9, 32'sd3, 32'sd9, 32'sd9, 32'sd18, 32'sd11, 32'sd4, 32'sd8, 32'sd9, 32'sd10, 32'sd12, 32'sd12, 32'sd4, 32'sd10, 32'sd6, 32'sd9, 32'sd5, 32'sd22, 32'sd6, 32'sd8, 32'sd4, 32'sd6, 32'sd4, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd3, 32'sd6, 32'sd9, 32'sd3, 32'sd6, 32'sd6, 32'sd4, 32'sd12, 32'sd9, 32'sd12, 32'sd6, 32'sd9, 32'sd9, 32'sd8, 32'sd6, 32'sd7, 32'sd12, 32'sd12, 32'sd6, 32'sd14, 32'sd18, 32'sd12, 32'sd14, 32'sd14, 32'sd20, 32'sd20, 32'sd17, 32'sd17, 32'sd6, 32'sd6, 32'sd13, 32'sd13, 32'sd9, 32'sd7, 32'sd6, 32'sd6, 32'sd9, 32'sd3, 32'sd10, 32'sd9, 32'sd18, 32'sd9, 32'sd4, 32'sd12, 32'sd5, 32'sd3, 32'sd5, 32'sd18, 32'sd14, 32'sd9, 32'sd6, 32'sd4, 32'sd8, 32'sd8, 32'sd2, 32'sd5, 32'sd12, 32'sd12, 32'sd3, 32'sd12, 32'sd6, 32'sd9, 32'sd5, 32'sd6, 32'sd6, 32'sd11, 32'sd18, 32'sd18, 32'sd8, 32'sd8, 32'sd3, 32'sd13, 32'sd9, 32'sd9, 32'sd9, 32'sd2, 32'sd6, 32'sd6, 32'sd21, 32'sd12, 32'sd6, 32'sd3, 32'sd3, 32'sd6, 32'sd12, 32'sd18, 32'sd7, 32'sd4, 32'sd9, 32'sd4, 32'sd6, 32'sd6, 32'sd2, 32'sd8, 32'sd7, 32'sd7, 32'sd5, 32'sd5, 32'sd10, 32'sd2, 32'sd6, 32'sd3, 32'sd9, 32'sd5, 32'sd6, 32'sd8, 32'sd9, 32'sd6, 32'sd4, 32'sd3, 32'sd2, 32'sd3, 32'sd9, 32'sd9, 32'sd20, 32'sd20, 32'sd14, 32'sd9, 32'sd4, 32'sd4, 32'sd6, 32'sd18, 32'sd6, 32'sd4, 32'sd9, 32'sd14, 32'sd18, 32'sd18, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd11, 32'sd12, 32'sd3, 32'sd8, 32'sd6, 32'sd4, 32'sd12, 32'sd12, 32'sd8, 32'sd3, 32'sd6, 32'sd8, 32'sd8, 32'sd3, 32'sd14, 32'sd10, 32'sd3, 32'sd6, 32'sd9, 32'sd8, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd8, 32'sd6, 32'sd4, 32'sd4, 32'sd3, 32'sd10, 32'sd6, 32'sd9, 32'sd6, 32'sd8, 32'sd6, 32'sd14, 32'sd8, 32'sd4, 32'sd9, 32'sd10, 32'sd13, 32'sd13, 32'sd6, 32'sd6, 32'sd14, 32'sd4, 32'sd6, 32'sd4, 32'sd9, 32'sd10, 32'sd5, 32'sd13, 32'sd19, 32'sd6, 32'sd2, 32'sd4, 32'sd5, 32'sd14, 32'sd6, 32'sd24, 32'sd14, 32'sd8, 32'sd6, 32'sd3, 32'sd5, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd12, 32'sd21, 32'sd3, 32'sd9, 32'sd12, 32'sd9, 32'sd9, 32'sd22, 32'sd12, 32'sd9, 32'sd4, 32'sd22, 32'sd22, 32'sd4, 32'sd7, 32'sd4, 32'sd15, 32'sd12, 32'sd12, 32'sd16, 
                                                    32'sd16, 32'sd16, 32'sd16, 32'sd3, 32'sd4, 32'sd8, 32'sd3, 32'sd2, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd14, 32'sd3, 32'sd7, 32'sd5, 32'sd5, 32'sd9, 32'sd10, 32'sd9, 32'sd9, 32'sd20, 32'sd3, 32'sd20, 32'sd8, 32'sd20, 32'sd19, 32'sd20, 32'sd9, 32'sd4, 32'sd6, 32'sd6, 32'sd8, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd8, 32'sd9, 32'sd9, 32'sd18, 32'sd20, 32'sd20, 32'sd6, 32'sd9, 32'sd6, 32'sd8, 32'sd12, 32'sd7, 32'sd6, 32'sd10, 32'sd3, 32'sd10, 32'sd12, 32'sd18, 32'sd16, 32'sd12, 32'sd14, 32'sd6, 32'sd6, 32'sd6, 32'sd10, 32'sd3, 32'sd8, 32'sd22, 32'sd8, 32'sd8, 32'sd9, 32'sd4, 32'sd6, 32'sd6, 32'sd3, 32'sd3, 32'sd9, 32'sd5, 32'sd15, 32'sd9, 32'sd3, 32'sd2, 32'sd9, 32'sd9, 32'sd9, 32'sd10, 32'sd16, 32'sd10, 32'sd13, 32'sd13, 32'sd9, 32'sd11, 32'sd11, 32'sd6, 32'sd3, 32'sd9, 32'sd14, 32'sd9, 32'sd6, 32'sd9, 32'sd20, 32'sd3, 32'sd3, 32'sd3, 32'sd9, 32'sd15, 32'sd3, 32'sd18, 32'sd3, 32'sd4, 32'sd5, 32'sd14, 32'sd9, 32'sd3, 32'sd18, 32'sd3, 32'sd12, 32'sd5, 32'sd12, 32'sd10, 32'sd10, 32'sd6, 32'sd9, 32'sd20, 32'sd6, 32'sd13, 32'sd15, 32'sd4, 32'sd14, 32'sd6, 32'sd3, 32'sd8, 32'sd18, 32'sd3, 32'sd13, 32'sd10, 32'sd9, 32'sd3, 32'sd3, 32'sd11, 32'sd10, 32'sd3, 32'sd3, 32'sd10, 32'sd21, 32'sd3, 32'sd6, 32'sd4, 32'sd4, 32'sd3, 32'sd3, 32'sd18, 32'sd3, 32'sd18, 32'sd6, 32'sd9, 32'sd10, 32'sd6, 32'sd18, 32'sd10, 32'sd10, 32'sd5, 32'sd7, 32'sd5, 32'sd7, 32'sd5, 32'sd18, 32'sd12, 32'sd4, 32'sd10, 32'sd6, 32'sd6, 32'sd2, 32'sd13, 32'sd3, 32'sd3, 32'sd6, 32'sd6, 32'sd6, 32'sd16, 32'sd16, 32'sd10, 32'sd10, 32'sd24, 32'sd20, 32'sd9, 32'sd9, 32'sd5, 32'sd9, 32'sd8, 32'sd8, 32'sd9, 32'sd12, 32'sd18, 32'sd18, 32'sd6, 32'sd3, 32'sd15, 32'sd14, 32'sd10, 32'sd9, 32'sd8, 32'sd8, 32'sd12, 32'sd4, 32'sd15, 32'sd10, 32'sd6, 32'sd5, 32'sd4, 32'sd6, 32'sd12, 32'sd6, 32'sd6, 32'sd23, 32'sd6, 32'sd12, 32'sd18, 32'sd12, 32'sd8, 32'sd4, 32'sd6, 32'sd3, 32'sd20, 32'sd20, 32'sd18, 32'sd12, 32'sd8, 32'sd14, 32'sd16, 32'sd9, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd9, 32'sd7, 32'sd6, 32'sd10, 32'sd21, 32'sd10, 32'sd8, 32'sd9, 32'sd12, 32'sd12, 32'sd12, 32'sd12, 32'sd9, 32'sd9, 32'sd4, 32'sd4, 32'sd6, 32'sd4, 32'sd4, 32'sd4, 32'sd19, 32'sd8, 32'sd12, 32'sd3, 32'sd4, 32'sd10, 32'sd6, 32'sd22, 32'sd22, 32'sd3, 32'sd15, 32'sd9, 32'sd3, 32'sd15, 32'sd3, 32'sd6, 32'sd14, 32'sd10, 32'sd9, 32'sd10, 32'sd10, 32'sd4, 32'sd2, 32'sd6, 32'sd16, 32'sd4, 32'sd9, 32'sd9, 32'sd6, 32'sd9, 32'sd8, 32'sd16, 32'sd12, 32'sd9, 32'sd9, 32'sd9, 32'sd18, 32'sd12, 32'sd12, 32'sd6, 32'sd4, 32'sd6, 32'sd6, 32'sd3, 32'sd3, 32'sd22, 32'sd22, 32'sd24, 32'sd4, 32'sd18, 32'sd14, 32'sd9, 32'sd9, 32'sd20, 32'sd9, 32'sd14, 32'sd6, 32'sd24, 32'sd24, 32'sd7, 32'sd7, 32'sd19, 32'sd6, 32'sd6, 32'sd8, 32'sd15, 32'sd15, 32'sd20, 32'sd20, 32'sd4, 32'sd4, 32'sd3, 32'sd3, 32'sd20, 32'sd9, 32'sd19, 32'sd3, 32'sd20, 32'sd9, 32'sd5, 32'sd6, 32'sd20, 32'sd20, 32'sd12, 32'sd12, 32'sd8, 32'sd6, 32'sd4, 32'sd15, 32'sd6, 32'sd10, 32'sd12, 32'sd4, 32'sd6, 32'sd18, 32'sd9, 32'sd6, 32'sd3, 32'sd6, 32'sd19, 32'sd19, 32'sd2, 32'sd6, 32'sd18, 32'sd8, 32'sd6, 32'sd10, 32'sd6, 32'sd6, 32'sd15, 32'sd10, 32'sd4, 32'sd3, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd5, 32'sd20, 32'sd6, 32'sd2, 32'sd6, 32'sd6, 32'sd9, 32'sd4, 32'sd6, 32'sd4, 32'sd22, 32'sd22, 32'sd9, 32'sd9, 32'sd18, 32'sd6, 32'sd8, 32'sd8, 32'sd12, 32'sd12, 32'sd8, 32'sd14, 32'sd12, 32'sd18, 32'sd18, 32'sd20, 32'sd12, 32'sd14, 32'sd6, 32'sd18, 32'sd14, 32'sd2, 32'sd12, 32'sd7, 32'sd12, 32'sd12, 32'sd22, 32'sd20, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd24, 32'sd12, 32'sd4, 32'sd6, 32'sd3, 32'sd8, 32'sd12, 32'sd3, 32'sd7, 32'sd6, 32'sd7, 32'sd19, 32'sd7, 32'sd9, 32'sd7, 32'sd6, 32'sd5, 32'sd19, 32'sd6, 32'sd14, 32'sd9, 32'sd5, 32'sd5, 32'sd5, 32'sd7, 32'sd10, 32'sd9, 32'sd9, 32'sd7, 32'sd7, 32'sd8, 32'sd12, 32'sd12, 32'sd12, 32'sd8, 32'sd3, 32'sd4, 32'sd6, 32'sd15, 32'sd6, 32'sd9, 32'sd20, 32'sd9, 32'sd5, 32'sd14, 32'sd4, 32'sd6, 32'sd7, 32'sd6, 32'sd18, 32'sd6, 32'sd4, 32'sd6, 32'sd12, 32'sd3, 32'sd6, 32'sd6, 32'sd3, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd3, 32'sd3, 32'sd6, 32'sd6, 32'sd9, 32'sd12, 32'sd8, 32'sd3, 32'sd12, 32'sd3, 32'sd9, 32'sd3, 32'sd3, 32'sd20, 32'sd20, 32'sd18, 32'sd12, 32'sd6, 32'sd18, 32'sd9, 32'sd6, 32'sd20, 32'sd20, 32'sd6, 32'sd6, 32'sd3, 32'sd6, 32'sd3, 32'sd7, 32'sd6, 32'sd6, 32'sd6, 32'sd13, 32'sd6, 32'sd15, 32'sd7, 32'sd6, 32'sd12, 32'sd9, 32'sd24, 32'sd24, 32'sd12, 32'sd6, 32'sd6, 32'sd12, 32'sd6, 32'sd14, 32'sd2, 32'sd3, 32'sd9, 32'sd12, 32'sd12, 32'sd9, 32'sd10, 32'sd9, 32'sd7, 32'sd5, 32'sd8, 32'sd18, 32'sd10, 32'sd10, 32'sd10, 32'sd10, 32'sd5, 32'sd2, 32'sd6, 32'sd7, 32'sd16, 32'sd8, 32'sd4, 32'sd8, 32'sd4, 32'sd9, 32'sd8, 32'sd4, 32'sd12, 32'sd12, 32'sd7, 32'sd3, 32'sd3, 32'sd10, 32'sd24, 32'sd15, 32'sd24, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd4, 32'sd20, 32'sd23, 32'sd18, 32'sd6, 32'sd6, 32'sd5, 32'sd19, 32'sd18, 32'sd18, 32'sd3, 32'sd9, 32'sd7, 32'sd7, 32'sd6, 32'sd10, 32'sd10, 32'sd16, 32'sd6, 32'sd6, 32'sd9, 32'sd8, 32'sd12, 32'sd9, 32'sd6, 32'sd22, 32'sd3, 32'sd3, 32'sd24, 32'sd6, 32'sd14, 32'sd10, 32'sd5, 32'sd6, 32'sd14, 32'sd14, 32'sd4, 32'sd12, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd10, 32'sd8, 32'sd8, 32'sd4, 32'sd18, 32'sd19, 32'sd16, 32'sd16, 32'sd6, 32'sd5, 32'sd5, 32'sd6, 32'sd5, 32'sd7, 32'sd6, 32'sd9, 32'sd6, 32'sd20, 32'sd12, 32'sd12, 32'sd6, 32'sd8, 32'sd10, 32'sd9, 32'sd22, 32'sd22, 32'sd4, 32'sd15, 32'sd12, 32'sd13, 32'sd24, 32'sd24, 32'sd8, 32'sd2, 32'sd3, 32'sd6, 32'sd10, 32'sd3, 32'sd4, 32'sd8, 32'sd4, 32'sd16, 32'sd16, 32'sd16, 32'sd14, 32'sd14, 32'sd22, 32'sd22, 32'sd20, 32'sd20, 32'sd9, 32'sd16, 32'sd12, 32'sd6, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd8, 32'sd12, 32'sd9, 32'sd6, 32'sd5, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd3, 32'sd2, 32'sd6, 32'sd9, 32'sd9, 32'sd15, 32'sd15, 32'sd6, 
                                                    32'sd14, 32'sd5, 32'sd3, 32'sd2, 32'sd10, 32'sd3, 32'sd11, 32'sd8, 32'sd9, 32'sd2, 32'sd6, 32'sd3, 32'sd18, 32'sd10, 32'sd10, 32'sd9, 32'sd9, 32'sd3, 32'sd4, 32'sd14, 32'sd14, 32'sd6, 32'sd6, 32'sd18, 32'sd3, 32'sd3, 32'sd10, 32'sd4, 32'sd6, 32'sd9, 32'sd12, 32'sd6, 32'sd13, 32'sd6, 32'sd6, 32'sd3, 32'sd6, 32'sd3, 32'sd6, 32'sd19, 32'sd16, 32'sd18, 32'sd18, 32'sd3, 32'sd4, 32'sd6, 32'sd4, 32'sd8, 32'sd8, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd2, 32'sd3, 32'sd12, 32'sd9, 32'sd15, 32'sd4, 32'sd12, 32'sd15, 32'sd19, 32'sd19, 32'sd10, 32'sd10, 32'sd18, 32'sd6, 32'sd10, 32'sd10, 32'sd10, 32'sd10, 32'sd18, 32'sd3, 32'sd18, 32'sd18, 32'sd3, 32'sd3, 32'sd3, 32'sd10, 32'sd17, 32'sd17, 32'sd11, 32'sd6, 32'sd8, 32'sd7, 32'sd14, 32'sd14, 32'sd2, 32'sd6, 32'sd4, 32'sd6, 32'sd18, 32'sd18, 32'sd10, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd3, 32'sd9, 32'sd6, 32'sd18, 32'sd9, 32'sd9, 32'sd9, 32'sd3, 32'sd4, 32'sd10, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd9, 32'sd3, 32'sd3, 32'sd6, 32'sd4, 32'sd6, 32'sd15, 32'sd3, 32'sd10, 32'sd3, 32'sd6, 32'sd18, 32'sd6, 32'sd18, 32'sd18, 32'sd6, 32'sd12, 32'sd22, 32'sd6, 32'sd6, 32'sd18, 32'sd9, 32'sd9, 32'sd12, 32'sd4, 32'sd3, 32'sd8, 32'sd15, 32'sd14, 32'sd14, 32'sd14, 32'sd4, 32'sd20, 32'sd12, 32'sd12, 32'sd8, 32'sd8, 32'sd15, 32'sd15, 32'sd12, 32'sd12, 32'sd9, 32'sd21, 32'sd4, 32'sd9, 32'sd15, 32'sd15, 32'sd8, 32'sd6, 32'sd4, 32'sd3, 32'sd12, 32'sd12, 32'sd6, 32'sd10, 32'sd6, 32'sd2, 32'sd3, 32'sd3, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd20, 32'sd8, 32'sd22}

localparam logic [2912:0][31:0] rectangle1_weights = {-32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, 
                                                    -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, 
                                                    -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, 
                                                    -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, 
                                                    -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, 
                                                    -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128, -32'sd128};

localparam logic [2912:0][31:0] rectangle2_xs = {32'sd6, 32'sd10, 32'sd3, 32'sd8, 32'sd5, 32'sd6, 32'sd5, 32'sd11, 32'sd4, 32'sd6, 32'sd10, 32'sd1, 32'sd8, 32'sd9, 32'sd5, 32'sd5, 32'sd16, 32'sd9, 32'sd12, 32'sd4, 32'sd20, 32'sd8, 32'sd11, 32'sd7, 32'sd5, 32'sd8, 32'sd5, 32'sd9, 32'sd11, 32'sd6, 32'sd9, 32'sd5, 32'sd18, 32'sd4, 32'sd8, 32'sd5, 32'sd2, 32'sd10, 32'sd2, 32'sd2, 32'sd20, 32'sd11, 32'sd20, 32'sd2, 32'sd12, 32'sd0, 32'sd12, 32'sd10, 32'sd12, 32'sd1, 32'sd17, 32'sd0, 32'sd6, 32'sd10, 32'sd8, 32'sd4, 32'sd2, 32'sd19, 32'sd3, 32'sd8, 32'sd1, 32'sd14, 32'sd3, 32'sd6, 32'sd8, 32'sd15, 32'sd1, 32'sd4, 32'sd2, 32'sd3, 32'sd1, 32'sd5, 32'sd3, 32'sd14, 32'sd1, 32'sd15, 32'sd5, 32'sd10, 32'sd9, 32'sd11, 32'sd9, 32'sd12, 32'sd10, 32'sd9, 32'sd6, 32'sd8, 32'sd4, 32'sd11, 32'sd8, 32'sd11, 32'sd9, 32'sd11, 32'sd11, 32'sd9, 32'sd1, 32'sd10, 32'sd6, 32'sd7, 32'sd0, 32'sd6, 32'sd1, 32'sd6, 32'sd5, 32'sd20, 32'sd2, 32'sd12, 32'sd4, 32'sd14, 32'sd8, 32'sd17, 32'sd0, 32'sd14, 32'sd8, 32'sd8, 32'sd0, 32'sd12, 32'sd9, 32'sd2, 32'sd2, 32'sd3, 32'sd5, 32'sd14, 32'sd4, 32'sd4, 32'sd6, 32'sd3, 32'sd3, 32'sd10, 32'sd8, 32'sd3, 32'sd12, 32'sd8, 32'sd5, 32'sd16, 32'sd4, 32'sd19, 32'sd8, 32'sd6, 32'sd10, 32'sd9, 32'sd0, 32'sd4, 32'sd9, 32'sd18, 32'sd3, 32'sd18, 32'sd3, 32'sd16, 32'sd2, 32'sd9, 32'sd2, 32'sd14, 32'sd5, 32'sd18, 32'sd3, 32'sd8, 32'sd7, 32'sd8, 32'sd10, 32'sd14, 32'sd7, 32'sd13, 32'sd12, 32'sd13, 32'sd1, 32'sd13, 32'sd8, 32'sd8, 32'sd8, 32'sd7, 32'sd0, 32'sd1, 32'sd9, 32'sd12, 32'sd9, 32'sd7, 32'sd0, 32'sd13, 32'sd12, 32'sd14, 32'sd9, 32'sd14, 32'sd9, 32'sd18, 32'sd6, 32'sd13, 32'sd3, 32'sd13, 32'sd0, 32'sd6, 32'sd6, 32'sd10, 32'sd10, 32'sd4, 32'sd5, 32'sd9, 32'sd20, 32'sd2, 32'sd5, 32'sd2, 32'sd5, 32'sd2, 32'sd13, 32'sd0, 32'sd1, 32'sd2, 32'sd13, 32'sd0, 32'sd11, 32'sd10, 32'sd11, 32'sd6, 32'sd18, 32'sd3, 32'sd18, 32'sd1, 32'sd13, 32'sd0, 32'sd13, 32'sd9, 32'sd13, 32'sd10, 32'sd13, 32'sd2, 32'sd12, 32'sd5, 32'sd14, 32'sd4, 32'sd7, 32'sd5, 32'sd12, 32'sd9, 32'sd3, 32'sd0, 32'sd12, 32'sd4, 32'sd13, 32'sd10, 32'sd10, 32'sd8, 32'sd10, 32'sd0, 32'sd12, 32'sd4, 32'sd8, 32'sd11, 32'sd9, 32'sd10, 32'sd20, 32'sd1, 32'sd14, 32'sd3, 32'sd15, 32'sd11, 32'sd17, 32'sd3, 32'sd7, 32'sd4, 32'sd10, 32'sd8, 32'sd15, 32'sd3, 32'sd12, 32'sd6, 32'sd14, 32'sd1, 32'sd13, 32'sd10, 32'sd12, 32'sd9, 32'sd6, 32'sd9, 32'sd7, 32'sd8, 32'sd7, 32'sd0, 32'sd15, 32'sd0, 32'sd15, 32'sd8, 32'sd15, 32'sd0, 32'sd8, 32'sd0, 32'sd9, 32'sd8, 32'sd9, 32'sd12, 32'sd12, 32'sd6, 32'sd16, 32'sd2, 32'sd0, 32'sd4, 32'sd9, 32'sd0, 32'sd18, 32'sd0, 32'sd8, 32'sd10, 32'sd13, 32'sd9, 32'sd14, 32'sd8, 32'sd15, 32'sd8, 32'sd9, 32'sd7, 32'sd14, 32'sd2, 32'sd5, 32'sd11, 32'sd13, 32'sd10, 32'sd9, 32'sd8, 32'sd12, 32'sd1, 32'sd15, 32'sd1, 32'sd10, 32'sd3, 32'sd12, 32'sd8, 32'sd6, 32'sd10, 32'sd5, 32'sd4, 32'sd11, 32'sd7, 32'sd9, 32'sd2, 32'sd3, 32'sd10, 32'sd16, 32'sd9, 32'sd21, 32'sd0, 32'sd18, 32'sd3, 32'sd18, 32'sd0, 32'sd5, 32'sd6, 32'sd12, 32'sd10, 32'sd15, 32'sd3, 32'sd15, 32'sd5, 32'sd11, 32'sd8, 32'sd15, 32'sd9, 32'sd13, 32'sd9, 32'sd18, 32'sd1, 32'sd14, 32'sd1, 32'sd12, 32'sd1, 32'sd14, 32'sd0, 32'sd17, 32'sd5, 32'sd18, 32'sd3, 32'sd15, 32'sd0, 32'sd4, 32'sd2, 32'sd14, 32'sd6, 32'sd20, 32'sd1, 32'sd16, 32'sd7, 32'sd12, 32'sd4, 32'sd12, 32'sd8, 32'sd15, 32'sd7, 32'sd6, 32'sd1, 32'sd6, 32'sd0, 32'sd13, 32'sd9, 32'sd12, 32'sd8, 32'sd16, 32'sd0, 32'sd14, 32'sd7, 32'sd5, 32'sd4, 32'sd16, 32'sd6, 32'sd12, 32'sd11, 32'sd11, 32'sd12, 32'sd6, 32'sd10, 32'sd8, 32'sd14, 32'sd5, 32'sd11, 32'sd3, 32'sd3, 32'sd3, 32'sd20, 32'sd5, 32'sd13, 32'sd6, 32'sd12, 32'sd8, 32'sd9, 32'sd10, 32'sd13, 32'sd9, 32'sd14, 32'sd8, 32'sd20, 32'sd6, 32'sd18, 32'sd7, 32'sd18, 32'sd0, 32'sd9, 32'sd0, 32'sd17, 32'sd1, 32'sd14, 32'sd8, 32'sd9, 32'sd9, 32'sd14, 32'sd8, 32'sd6, 32'sd1, 32'sd10, 32'sd5, 32'sd5, 32'sd0, 32'sd8, 32'sd10, 32'sd6, 32'sd4, 32'sd12, 32'sd12, 32'sd12, 32'sd3, 32'sd2, 32'sd6, 32'sd14, 32'sd0, 32'sd19, 32'sd0, 32'sd12, 32'sd0, 32'sd13, 32'sd3, 32'sd6, 32'sd0, 32'sd15, 32'sd9, 32'sd12, 32'sd1, 32'sd15, 32'sd7, 32'sd19, 32'sd6, 32'sd8, 32'sd5, 32'sd14, 32'sd2, 32'sd18, 32'sd2, 32'sd17, 32'sd12, 32'sd14, 32'sd10, 32'sd14, 32'sd6, 32'sd6, 32'sd11, 32'sd12, 32'sd10, 32'sd16, 32'sd6, 32'sd9, 32'sd5, 32'sd10, 32'sd8, 32'sd6, 32'sd10, 32'sd8, 32'sd1, 32'sd9, 32'sd3, 32'sd2, 32'sd10, 32'sd8, 32'sd10, 32'sd0, 32'sd14, 32'sd9, 32'sd14, 32'sd1, 32'sd15, 32'sd0, 32'sd19, 32'sd2, 32'sd3, 32'sd9, 32'sd18, 32'sd0, 32'sd12, 32'sd2, 32'sd14, 32'sd5, 32'sd18, 32'sd5, 32'sd22, 32'sd8, 32'sd11, 32'sd7, 32'sd22, 32'sd12, 32'sd15, 32'sd0, 32'sd13, 32'sd9, 32'sd14, 32'sd6, 32'sd14, 32'sd6, 32'sd3, 32'sd3, 32'sd12, 32'sd12, 32'sd13, 32'sd8, 32'sd20, 32'sd3, 32'sd20, 32'sd0, 32'sd10, 32'sd8, 32'sd13, 32'sd9, 32'sd13, 32'sd0, 32'sd6, 32'sd3, 32'sd8, 32'sd2, 32'sd15, 32'sd3, 32'sd19, 32'sd3, 32'sd19, 32'sd3, 32'sd4, 32'sd6, 32'sd15, 32'sd0, 32'sd17, 32'sd5, 32'sd8, 32'sd6, 32'sd5, 32'sd10, 32'sd10, 32'sd0, 32'sd15, 32'sd0, 32'sd14, 32'sd11, 32'sd14, 32'sd8, 32'sd15, 32'sd3, 32'sd11, 32'sd6, 32'sd12, 32'sd0, 32'sd3, 32'sd3, 32'sd12, 32'sd1, 32'sd17, 32'sd2, 32'sd7, 32'sd8, 32'sd3, 32'sd10, 32'sd5, 32'sd11, 32'sd3, 32'sd18, 32'sd3, 32'sd9, 32'sd3, 32'sd13, 32'sd8, 32'sd13, 32'sd4, 32'sd13, 32'sd8, 32'sd7, 32'sd6, 32'sd16, 32'sd6, 32'sd11, 32'sd0, 32'sd13, 32'sd5, 32'sd10, 32'sd10, 32'sd14, 32'sd6, 32'sd12, 32'sd7, 32'sd8, 32'sd5, 32'sd3, 32'sd5, 32'sd5, 32'sd8, 32'sd3, 32'sd1, 32'sd5, 32'sd1, 32'sd1, 32'sd3, 32'sd6, 32'sd7, 32'sd14, 32'sd1, 32'sd13, 32'sd12, 32'sd13, 32'sd9, 32'sd15, 32'sd5, 32'sd15, 32'sd6, 32'sd15, 32'sd0, 32'sd5, 32'sd7, 32'sd17, 32'sd10, 32'sd15, 32'sd0, 32'sd14, 32'sd8, 32'sd13, 32'sd6, 32'sd13, 32'sd8, 32'sd17, 32'sd4, 32'sd12, 32'sd11, 32'sd11, 32'sd9, 32'sd8, 32'sd1, 32'sd9, 32'sd9, 32'sd18, 32'sd8, 32'sd2, 32'sd0, 
                                                    32'sd18, 32'sd2, 32'sd2, 32'sd12, 32'sd13, 32'sd1, 32'sd11, 32'sd3, 32'sd12, 32'sd2, 32'sd18, 32'sd3, 32'sd22, 32'sd2, 32'sd1, 32'sd0, 32'sd19, 32'sd3, 32'sd20, 32'sd0, 32'sd13, 32'sd0, 32'sd10, 32'sd8, 32'sd4, 32'sd2, 32'sd14, 32'sd3, 32'sd17, 32'sd6, 32'sd10, 32'sd4, 32'sd2, 32'sd10, 32'sd5, 32'sd12, 32'sd0, 32'sd15, 32'sd5, 32'sd8, 32'sd1, 32'sd19, 32'sd8, 32'sd20, 32'sd9, 32'sd15, 32'sd2, 32'sd16, 32'sd2, 32'sd20, 32'sd3, 32'sd15, 32'sd0, 32'sd16, 32'sd2, 32'sd10, 32'sd1, 32'sd14, 32'sd3, 32'sd3, 32'sd10, 32'sd3, 32'sd2, 32'sd12, 32'sd10, 32'sd12, 32'sd11, 32'sd4, 32'sd0, 32'sd9, 32'sd8, 32'sd13, 32'sd5, 32'sd12, 32'sd1, 32'sd19, 32'sd0, 32'sd20, 32'sd0, 32'sd18, 32'sd9, 32'sd11, 32'sd0, 32'sd1, 32'sd1, 32'sd13, 32'sd4, 32'sd12, 32'sd4, 32'sd15, 32'sd1, 32'sd13, 32'sd5, 32'sd16, 32'sd5, 32'sd10, 32'sd7, 32'sd12, 32'sd0, 32'sd17, 32'sd0, 32'sd15, 32'sd0, 32'sd13, 32'sd8, 32'sd12, 32'sd2, 32'sd12, 32'sd1, 32'sd15, 32'sd0, 32'sd6, 32'sd10, 32'sd12, 32'sd8, 32'sd12, 32'sd8, 32'sd13, 32'sd1, 32'sd15, 32'sd6, 32'sd18, 32'sd11, 32'sd12, 32'sd0, 32'sd11, 32'sd11, 32'sd12, 32'sd8, 32'sd9, 32'sd10, 32'sd4, 32'sd11, 32'sd5, 32'sd8, 32'sd15, 32'sd12, 32'sd12, 32'sd7, 32'sd11, 32'sd3, 32'sd14, 32'sd8, 32'sd9, 32'sd1, 32'sd11, 32'sd9, 32'sd12, 32'sd1, 32'sd6, 32'sd1, 32'sd8, 32'sd2, 32'sd11, 32'sd7, 32'sd14, 32'sd9, 32'sd14, 32'sd7, 32'sd4, 32'sd9, 32'sd7, 32'sd11, 32'sd2, 32'sd8, 32'sd3, 32'sd11, 32'sd0, 32'sd10, 32'sd2, 32'sd20, 32'sd2, 32'sd12, 32'sd0, 32'sd14, 32'sd0, 32'sd12, 32'sd8, 32'sd4, 32'sd10, 32'sd14, 32'sd2, 32'sd14, 32'sd2, 32'sd5, 32'sd9, 32'sd12, 32'sd6, 32'sd12, 32'sd0, 32'sd18, 32'sd5, 32'sd10, 32'sd2, 32'sd13, 32'sd6, 32'sd11, 32'sd7, 32'sd18, 32'sd11, 32'sd10, 32'sd0, 32'sd15, 32'sd4, 32'sd13, 32'sd7, 32'sd14, 32'sd7, 32'sd12, 32'sd6, 32'sd16, 32'sd0, 32'sd16, 32'sd5, 32'sd5, 32'sd5, 32'sd9, 32'sd9, 32'sd13, 32'sd5, 32'sd19, 32'sd3, 32'sd5, 32'sd0, 32'sd2, 32'sd5, 32'sd1, 32'sd10, 32'sd8, 32'sd11, 32'sd12, 32'sd4, 32'sd12, 32'sd3, 32'sd5, 32'sd4, 32'sd6, 32'sd10, 32'sd0, 32'sd0, 32'sd3, 32'sd2, 32'sd7, 32'sd5, 32'sd10, 32'sd9, 32'sd18, 32'sd9, 32'sd12, 32'sd11, 32'sd13, 32'sd9, 32'sd4, 32'sd2, 32'sd13, 32'sd9, 32'sd9, 32'sd1, 32'sd8, 32'sd3, 32'sd5, 32'sd8, 32'sd9, 32'sd0, 32'sd6, 32'sd4, 32'sd13, 32'sd5, 32'sd12, 32'sd11, 32'sd14, 32'sd5, 32'sd12, 32'sd0, 32'sd20, 32'sd9, 32'sd12, 32'sd10, 32'sd14, 32'sd7, 32'sd12, 32'sd2, 32'sd18, 32'sd1, 32'sd6, 32'sd12, 32'sd14, 32'sd6, 32'sd11, 32'sd1, 32'sd9, 32'sd7, 32'sd17, 32'sd2, 32'sd7, 32'sd1, 32'sd8, 32'sd11, 32'sd3, 32'sd20, 32'sd8, 32'sd20, 32'sd0, 32'sd8, 32'sd5, 32'sd4, 32'sd8, 32'sd6, 32'sd0, 32'sd20, 32'sd10, 32'sd12, 32'sd0, 32'sd6, 32'sd0, 32'sd20, 32'sd2, 32'sd18, 32'sd3, 32'sd13, 32'sd8, 32'sd5, 32'sd9, 32'sd6, 32'sd9, 32'sd10, 32'sd1, 32'sd11, 32'sd7, 32'sd14, 32'sd5, 32'sd13, 32'sd0, 32'sd12, 32'sd1, 32'sd2, 32'sd2, 32'sd20, 32'sd1, 32'sd14, 32'sd0, 32'sd15, 32'sd1, 32'sd9, 32'sd0, 32'sd16, 32'sd12, 32'sd7, 32'sd11, 32'sd12, 32'sd10, 32'sd15, 32'sd3, 32'sd16, 32'sd3, 32'sd16, 32'sd12, 32'sd10, 32'sd7, 32'sd11, 32'sd11, 32'sd12, 32'sd11, 32'sd3, 32'sd2, 32'sd12, 32'sd5, 32'sd14, 32'sd0, 32'sd10, 32'sd8, 32'sd5, 32'sd11, 32'sd11, 32'sd9, 32'sd5, 32'sd10, 32'sd10, 32'sd7, 32'sd12, 32'sd0, 32'sd12, 32'sd2, 32'sd12, 32'sd1, 32'sd12, 32'sd0, 32'sd5, 32'sd6, 32'sd14, 32'sd5, 32'sd9, 32'sd8, 32'sd11, 32'sd6, 32'sd17, 32'sd8, 32'sd8, 32'sd4, 32'sd12, 32'sd9, 32'sd16, 32'sd1, 32'sd11, 32'sd3, 32'sd7, 32'sd12, 32'sd12, 32'sd3, 32'sd12, 32'sd3, 32'sd13, 32'sd5, 32'sd11, 32'sd9, 32'sd17, 32'sd2, 32'sd12, 32'sd0, 32'sd12, 32'sd5, 32'sd12, 32'sd9, 32'sd2, 32'sd5, 32'sd4, 32'sd2, 32'sd7, 32'sd0, 32'sd2, 32'sd6, 32'sd6, 32'sd11, 32'sd15, 32'sd8, 32'sd3, 32'sd2, 32'sd19, 32'sd1, 32'sd14, 32'sd4, 32'sd14, 32'sd8, 32'sd14, 32'sd4, 32'sd8, 32'sd3, 32'sd20, 32'sd2, 32'sd8, 32'sd9, 32'sd16, 32'sd12, 32'sd11, 32'sd12, 32'sd12, 32'sd10, 32'sd14, 32'sd5, 32'sd18, 32'sd6, 32'sd13, 32'sd1, 32'sd15, 32'sd9, 32'sd10, 32'sd3, 32'sd16, 32'sd9, 32'sd15, 32'sd0, 32'sd13, 32'sd2, 32'sd5, 32'sd1, 32'sd5, 32'sd1, 32'sd16, 32'sd9, 32'sd16, 32'sd6, 32'sd18, 32'sd1, 32'sd9, 32'sd0, 32'sd14, 32'sd3, 32'sd16, 32'sd3, 32'sd11, 32'sd11, 32'sd15, 32'sd8, 32'sd17, 32'sd3, 32'sd3, 32'sd0, 32'sd2, 32'sd0, 32'sd13, 32'sd5, 32'sd12, 32'sd5, 32'sd18, 32'sd0, 32'sd13, 32'sd5, 32'sd9, 32'sd12, 32'sd6, 32'sd9, 32'sd13, 32'sd8, 32'sd6, 32'sd2, 32'sd20, 32'sd2, 32'sd14, 32'sd8, 32'sd8, 32'sd12, 32'sd9, 32'sd11, 32'sd4, 32'sd10, 32'sd8, 32'sd7, 32'sd12, 32'sd0, 32'sd18, 32'sd0, 32'sd16, 32'sd1, 32'sd12, 32'sd9, 32'sd12, 32'sd8, 32'sd12, 32'sd4, 32'sd15, 32'sd3, 32'sd15, 32'sd4, 32'sd15, 32'sd0, 32'sd15, 32'sd0, 32'sd14, 32'sd3, 32'sd7, 32'sd10, 32'sd8, 32'sd12, 32'sd7, 32'sd0, 32'sd16, 32'sd7, 32'sd10, 32'sd11, 32'sd12, 32'sd3, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd10, 32'sd4, 32'sd8, 32'sd9, 32'sd9, 32'sd6, 32'sd11, 32'sd8, 32'sd4, 32'sd8, 32'sd7, 32'sd1, 32'sd15, 32'sd7, 32'sd13, 32'sd9, 32'sd3, 32'sd0, 32'sd10, 32'sd6, 32'sd15, 32'sd0, 32'sd20, 32'sd2, 32'sd13, 32'sd0, 32'sd2, 32'sd1, 32'sd18, 32'sd0, 32'sd17, 32'sd0, 32'sd0, 32'sd2, 32'sd12, 32'sd9, 32'sd17, 32'sd5, 32'sd15, 32'sd0, 32'sd15, 32'sd0, 32'sd5, 32'sd0, 32'sd13, 32'sd8, 32'sd13, 32'sd8, 32'sd13, 32'sd10, 32'sd12, 32'sd11, 32'sd13, 32'sd7, 32'sd14, 32'sd12, 32'sd12, 32'sd1, 32'sd20, 32'sd0, 32'sd14, 32'sd0, 32'sd13, 32'sd0, 32'sd6, 32'sd0, 32'sd14, 32'sd1, 32'sd13, 32'sd4, 32'sd17, 32'sd5, 32'sd16, 32'sd3, 32'sd14, 32'sd10, 32'sd11, 32'sd0, 32'sd4, 32'sd5, 32'sd19, 32'sd0, 32'sd8, 32'sd3, 32'sd17, 32'sd4, 32'sd16, 32'sd3, 32'sd18, 32'sd1, 32'sd17, 32'sd0, 32'sd15, 32'sd8, 32'sd22, 32'sd1, 32'sd20, 32'sd2, 32'sd3, 32'sd6, 32'sd7, 32'sd11, 32'sd4, 32'sd9, 32'sd4, 32'sd3, 32'sd18, 32'sd2, 32'sd13, 32'sd7, 
                                                    32'sd13, 32'sd10, 32'sd12, 32'sd0, 32'sd11, 32'sd2, 32'sd13, 32'sd5, 32'sd9, 32'sd5, 32'sd3, 32'sd6, 32'sd12, 32'sd8, 32'sd9, 32'sd1, 32'sd19, 32'sd1, 32'sd9, 32'sd6, 32'sd12, 32'sd10, 32'sd14, 32'sd4, 32'sd8, 32'sd6, 32'sd19, 32'sd0, 32'sd17, 32'sd1, 32'sd18, 32'sd0, 32'sd3, 32'sd2, 32'sd14, 32'sd5, 32'sd10, 32'sd11, 32'sd7, 32'sd12, 32'sd5, 32'sd10, 32'sd11, 32'sd9, 32'sd14, 32'sd8, 32'sd12, 32'sd7, 32'sd2, 32'sd1, 32'sd8, 32'sd7, 32'sd6, 32'sd17, 32'sd4, 32'sd2, 32'sd6, 32'sd9, 32'sd7, 32'sd10, 32'sd8, 32'sd18, 32'sd3, 32'sd18, 32'sd4, 32'sd5, 32'sd11, 32'sd15, 32'sd7, 32'sd12, 32'sd12, 32'sd12, 32'sd2, 32'sd14, 32'sd10, 32'sd14, 32'sd3, 32'sd14, 32'sd1, 32'sd3, 32'sd1, 32'sd18, 32'sd0, 32'sd5, 32'sd6, 32'sd14, 32'sd4, 32'sd17, 32'sd8, 32'sd8, 32'sd5, 32'sd3, 32'sd0, 32'sd12, 32'sd0, 32'sd9, 32'sd2, 32'sd0, 32'sd10, 32'sd10, 32'sd8, 32'sd13, 32'sd11, 32'sd2, 32'sd1, 32'sd13, 32'sd12, 32'sd10, 32'sd7, 32'sd14, 32'sd10, 32'sd11, 32'sd10, 32'sd20, 32'sd1, 32'sd17, 32'sd9, 32'sd12, 32'sd12, 32'sd14, 32'sd5, 32'sd16, 32'sd4, 32'sd10, 32'sd1, 32'sd15, 32'sd12, 32'sd12, 32'sd8, 32'sd19, 32'sd0, 32'sd14, 32'sd6, 32'sd13, 32'sd9, 32'sd13, 32'sd8, 32'sd7, 32'sd4, 32'sd17, 32'sd3, 32'sd14, 32'sd2, 32'sd3, 32'sd4, 32'sd19, 32'sd10, 32'sd19, 32'sd1, 32'sd15, 32'sd5, 32'sd10, 32'sd4, 32'sd0, 32'sd8, 32'sd14, 32'sd0, 32'sd6, 32'sd1, 32'sd18, 32'sd4, 32'sd6, 32'sd1, 32'sd1, 32'sd2, 32'sd18, 32'sd0, 32'sd12, 32'sd7, 32'sd9, 32'sd7, 32'sd12, 32'sd7, 32'sd12, 32'sd10, 32'sd15, 32'sd3, 32'sd4, 32'sd6, 32'sd8, 32'sd12, 32'sd11, 32'sd2, 32'sd8, 32'sd0, 32'sd0, 32'sd2, 32'sd12, 32'sd10, 32'sd7, 32'sd9, 32'sd17, 32'sd0, 32'sd19, 32'sd1, 32'sd12, 32'sd3, 32'sd12, 32'sd12, 32'sd12, 32'sd10, 32'sd14, 32'sd10, 32'sd13, 32'sd7, 32'sd7, 32'sd9, 32'sd0, 32'sd11, 32'sd3, 32'sd15, 32'sd2, 32'sd13, 32'sd4, 32'sd20, 32'sd8, 32'sd12, 32'sd2, 32'sd3, 32'sd3, 32'sd13, 32'sd5, 32'sd17, 32'sd2, 32'sd12, 32'sd10, 32'sd12, 32'sd10, 32'sd12, 32'sd12, 32'sd12, 32'sd0, 32'sd9, 32'sd7, 32'sd14, 32'sd8, 32'sd13, 32'sd1, 32'sd9, 32'sd2, 32'sd15, 32'sd0, 32'sd9, 32'sd2, 32'sd15, 32'sd4, 32'sd17, 32'sd0, 32'sd15, 32'sd0, 32'sd15, 32'sd3, 32'sd20, 32'sd8, 32'sd13, 32'sd0, 32'sd0, 32'sd5, 32'sd11, 32'sd4, 32'sd10, 32'sd8, 32'sd11, 32'sd4, 32'sd14, 32'sd2, 32'sd4, 32'sd8, 32'sd1, 32'sd9, 32'sd13, 32'sd10, 32'sd4, 32'sd6, 32'sd14, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd11, 32'sd9, 32'sd12, 32'sd14, 32'sd8, 32'sd18, 32'sd3, 32'sd18, 32'sd0, 32'sd13, 32'sd10, 32'sd11, 32'sd8, 32'sd16, 32'sd5, 32'sd7, 32'sd9, 32'sd13, 32'sd3, 32'sd20, 32'sd7, 32'sd15, 32'sd0, 32'sd19, 32'sd1, 32'sd12, 32'sd1, 32'sd3, 32'sd8, 32'sd5, 32'sd9, 32'sd11, 32'sd4, 32'sd6, 32'sd5, 32'sd17, 32'sd11, 32'sd1, 32'sd10, 32'sd10, 32'sd11, 32'sd11, 32'sd9, 32'sd15, 32'sd0, 32'sd2, 32'sd0, 32'sd9, 32'sd9, 32'sd18, 32'sd0, 32'sd12, 32'sd3, 32'sd2, 32'sd5, 32'sd12, 32'sd10, 32'sd5, 32'sd9, 32'sd7, 32'sd9, 32'sd4, 32'sd0, 32'sd11, 32'sd11, 32'sd6, 32'sd11, 32'sd12, 32'sd5, 32'sd14, 32'sd5, 32'sd14, 32'sd0, 32'sd16, 32'sd4, 32'sd8, 32'sd0, 32'sd13, 32'sd0, 32'sd12, 32'sd6, 32'sd10, 32'sd1, 32'sd0, 32'sd6, 32'sd9, 32'sd1, 32'sd10, 32'sd7, 32'sd9, 32'sd10, 32'sd3, 32'sd7, 32'sd3, 32'sd10, 32'sd3, 32'sd10, 32'sd4, 32'sd5, 32'sd8, 32'sd9, 32'sd3, 32'sd2, 32'sd9, 32'sd11, 32'sd11, 32'sd16, 32'sd7, 32'sd16, 32'sd6, 32'sd19, 32'sd3, 32'sd14, 32'sd0, 32'sd9, 32'sd6, 32'sd14, 32'sd4, 32'sd7, 32'sd9, 32'sd14, 32'sd12, 32'sd14, 32'sd5, 32'sd4, 32'sd11, 32'sd3, 32'sd4, 32'sd16, 32'sd4, 32'sd13, 32'sd10, 32'sd15, 32'sd12, 32'sd12, 32'sd3, 32'sd12, 32'sd8, 32'sd6, 32'sd0, 32'sd4, 32'sd0, 32'sd15, 32'sd0, 32'sd6, 32'sd3, 32'sd13, 32'sd6, 32'sd6, 32'sd10, 32'sd10, 32'sd7, 32'sd17, 32'sd2, 32'sd11, 32'sd1, 32'sd15, 32'sd1, 32'sd10, 32'sd11, 32'sd7, 32'sd10, 32'sd15, 32'sd3, 32'sd15, 32'sd7, 32'sd12, 32'sd9, 32'sd15, 32'sd5, 32'sd8, 32'sd7, 32'sd12, 32'sd9, 32'sd7, 32'sd10, 32'sd13, 32'sd9, 32'sd9, 32'sd0, 32'sd14, 32'sd0, 32'sd12, 32'sd1, 32'sd7, 32'sd11, 32'sd16, 32'sd2, 32'sd8, 32'sd0, 32'sd5, 32'sd2, 32'sd14, 32'sd3, 32'sd9, 32'sd4, 32'sd12, 32'sd9, 32'sd13, 32'sd0, 32'sd14, 32'sd2, 32'sd11, 32'sd7, 32'sd13, 32'sd7, 32'sd17, 32'sd4, 32'sd13, 32'sd10, 32'sd18, 32'sd12, 32'sd17, 32'sd5, 32'sd16, 32'sd4, 32'sd18, 32'sd4, 32'sd15, 32'sd0, 32'sd20, 32'sd2, 32'sd16, 32'sd9, 32'sd12, 32'sd0, 32'sd5, 32'sd0, 32'sd12, 32'sd5, 32'sd10, 32'sd8, 32'sd6, 32'sd3, 32'sd16, 32'sd6, 32'sd8, 32'sd6, 32'sd10, 32'sd11, 32'sd14, 32'sd0, 32'sd16, 32'sd3, 32'sd6, 32'sd4, 32'sd17, 32'sd2, 32'sd2, 32'sd4, 32'sd18, 32'sd8, 32'sd6, 32'sd6, 32'sd14, 32'sd8, 32'sd15, 32'sd6, 32'sd14, 32'sd4, 32'sd7, 32'sd8, 32'sd13, 32'sd9, 32'sd8, 32'sd0, 32'sd17, 32'sd0, 32'sd21, 32'sd0, 32'sd12, 32'sd1, 32'sd5, 32'sd1, 32'sd6, 32'sd5, 32'sd14, 32'sd1, 32'sd11, 32'sd0, 32'sd13, 32'sd1, 32'sd0, 32'sd1, 32'sd14, 32'sd7, 32'sd12, 32'sd8, 32'sd13, 32'sd11, 32'sd9, 32'sd7, 32'sd6, 32'sd10, 32'sd10, 32'sd6, 32'sd15, 32'sd8, 32'sd11, 32'sd8, 32'sd1, 32'sd0, 32'sd15, 32'sd7, 32'sd20, 32'sd2, 32'sd14, 32'sd2, 32'sd12, 32'sd1, 32'sd7, 32'sd8, 32'sd12, 32'sd2, 32'sd14, 32'sd3, 32'sd17, 32'sd5, 32'sd13, 32'sd9, 32'sd13, 32'sd12, 32'sd12, 32'sd11, 32'sd20, 32'sd1, 32'sd7, 32'sd6, 32'sd9, 32'sd1, 32'sd19, 32'sd4, 32'sd3, 32'sd1, 32'sd9, 32'sd4, 32'sd6, 32'sd4, 32'sd15, 32'sd9, 32'sd12, 32'sd6, 32'sd15, 32'sd3, 32'sd14, 32'sd1, 32'sd14, 32'sd0, 32'sd15, 32'sd3, 32'sd9, 32'sd1, 32'sd13, 32'sd1, 32'sd6, 32'sd8, 32'sd0, 32'sd0, 32'sd14, 32'sd1, 32'sd14, 32'sd8, 32'sd10, 32'sd11, 32'sd10, 32'sd9, 32'sd14, 32'sd8, 32'sd11, 32'sd3, 32'sd13, 32'sd0, 32'sd12, 32'sd11, 32'sd10, 32'sd8, 32'sd11, 32'sd10, 32'sd12, 32'sd10, 32'sd4, 32'sd0, 32'sd11, 32'sd1, 32'sd11, 32'sd6, 32'sd14, 32'sd7, 32'sd12, 32'sd12, 32'sd11, 32'sd1, 32'sd9, 32'sd0, 32'sd1, 32'sd1, 32'sd9, 32'sd9, 
                                                    32'sd11, 32'sd11, 32'sd18, 32'sd4, 32'sd15, 32'sd1, 32'sd14, 32'sd3, 32'sd15, 32'sd7, 32'sd14, 32'sd12, 32'sd7, 32'sd0, 32'sd19, 32'sd1, 32'sd16, 32'sd6, 32'sd17, 32'sd5, 32'sd0, 32'sd7, 32'sd1, 32'sd1, 32'sd6, 32'sd1, 32'sd15, 32'sd3, 32'sd4, 32'sd0, 32'sd6, 32'sd7, 32'sd12, 32'sd6, 32'sd9, 32'sd4, 32'sd20, 32'sd2, 32'sd13, 32'sd12, 32'sd13, 32'sd1, 32'sd13, 32'sd2, 32'sd13, 32'sd2, 32'sd3, 32'sd7, 32'sd17, 32'sd5, 32'sd16, 32'sd0, 32'sd15, 32'sd0, 32'sd9, 32'sd4, 32'sd12, 32'sd10, 32'sd13, 32'sd9, 32'sd14, 32'sd8, 32'sd10, 32'sd0, 32'sd13, 32'sd9, 32'sd14, 32'sd0, 32'sd1, 32'sd10, 32'sd16, 32'sd10, 32'sd12, 32'sd8, 32'sd13, 32'sd2, 32'sd11, 32'sd7, 32'sd13, 32'sd0, 32'sd12, 32'sd8, 32'sd12, 32'sd6, 32'sd14, 32'sd0, 32'sd14, 32'sd0, 32'sd4, 32'sd1, 32'sd4, 32'sd8, 32'sd3, 32'sd11, 32'sd0, 32'sd6, 32'sd2, 32'sd18, 32'sd0, 32'sd11, 32'sd9, 32'sd7, 32'sd3, 32'sd18, 32'sd7, 32'sd18, 32'sd3, 32'sd9, 32'sd2, 32'sd10, 32'sd5, 32'sd11, 32'sd10, 32'sd12, 32'sd4, 32'sd6, 32'sd9, 32'sd9, 32'sd11, 32'sd10, 32'sd2, 32'sd21, 32'sd0, 32'sd5, 32'sd12, 32'sd1, 32'sd10, 32'sd6, 32'sd9, 32'sd2, 32'sd5, 32'sd12, 32'sd9, 32'sd18, 32'sd2, 32'sd16, 32'sd1, 32'sd12, 32'sd4, 32'sd10, 32'sd5, 32'sd14, 32'sd7, 32'sd7, 32'sd2, 32'sd5, 32'sd7, 32'sd0, 32'sd2, 32'sd20, 32'sd5, 32'sd5, 32'sd0, 32'sd13, 32'sd0, 32'sd4, 32'sd2, 32'sd12, 32'sd12, 32'sd6, 32'sd0, 32'sd10, 32'sd7, 32'sd11, 32'sd7, 32'sd21, 32'sd3, 32'sd21, 32'sd7, 32'sd9, 32'sd0, 32'sd15, 32'sd1, 32'sd13, 32'sd7, 32'sd13, 32'sd10, 32'sd13, 32'sd10, 32'sd13, 32'sd10, 32'sd5, 32'sd0, 32'sd11, 32'sd2, 32'sd15, 32'sd1, 32'sd10, 32'sd0, 32'sd6, 32'sd0, 32'sd13, 32'sd2, 32'sd13, 32'sd8, 32'sd13, 32'sd9, 32'sd12, 32'sd3, 32'sd16, 32'sd6, 32'sd10, 32'sd7, 32'sd12, 32'sd7, 32'sd10, 32'sd3, 32'sd16, 32'sd4, 32'sd0, 32'sd11, 32'sd10, 32'sd12, 32'sd17, 32'sd5, 32'sd16, 32'sd5, 32'sd3, 32'sd4, 32'sd4, 32'sd3, 32'sd16, 32'sd6, 32'sd14, 32'sd7, 32'sd4, 32'sd0, 32'sd10, 32'sd6, 32'sd0, 32'sd0, 32'sd3, 32'sd9, 32'sd12, 32'sd6, 32'sd8, 32'sd2, 32'sd12, 32'sd5, 32'sd14, 32'sd10, 32'sd12, 32'sd7, 32'sd17, 32'sd9, 32'sd13, 32'sd0, 32'sd12, 32'sd9, 32'sd10, 32'sd9, 32'sd0, 32'sd8, 32'sd9, 32'sd9, 32'sd15, 32'sd10, 32'sd15, 32'sd6, 32'sd19, 32'sd2, 32'sd12, 32'sd10, 32'sd14, 32'sd5, 32'sd11, 32'sd3, 32'sd10, 32'sd5, 32'sd20, 32'sd7, 32'sd4, 32'sd8, 32'sd6, 32'sd19, 32'sd3, 32'sd20, 32'sd2, 32'sd5, 32'sd10, 32'sd11, 32'sd0, 32'sd7, 32'sd1, 32'sd11, 32'sd0, 32'sd17, 32'sd12, 32'sd17, 32'sd7, 32'sd13, 32'sd0, 32'sd8, 32'sd6, 32'sd7, 32'sd0, 32'sd13, 32'sd3, 32'sd12, 32'sd2, 32'sd9, 32'sd6, 32'sd14, 32'sd5, 32'sd12, 32'sd6, 32'sd17, 32'sd4, 32'sd14, 32'sd0, 32'sd13, 32'sd2, 32'sd6, 32'sd0, 32'sd21, 32'sd1, 32'sd15, 32'sd11, 32'sd13, 32'sd7, 32'sd14, 32'sd3, 32'sd22, 32'sd7, 32'sd12, 32'sd11, 32'sd15, 32'sd8, 32'sd13, 32'sd8, 32'sd9, 32'sd8, 32'sd12, 32'sd3, 32'sd19, 32'sd0, 32'sd22, 32'sd0, 32'sd7, 32'sd11, 32'sd10, 32'sd0, 32'sd14, 32'sd2, 32'sd13, 32'sd8, 32'sd15, 32'sd7, 32'sd11, 32'sd11, 32'sd15, 32'sd1, 32'sd16, 32'sd5, 32'sd12, 32'sd4, 32'sd6, 32'sd9, 32'sd15, 32'sd6, 32'sd12, 32'sd7, 32'sd6, 32'sd10, 32'sd12, 32'sd3, 32'sd4, 32'sd2, 32'sd13, 32'sd9, 32'sd1, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd5, 32'sd16, 32'sd5, 32'sd10, 32'sd6, 32'sd12, 32'sd2, 32'sd12, 32'sd10, 32'sd13, 32'sd6, 32'sd9, 32'sd2, 32'sd14, 32'sd3, 32'sd10, 32'sd2, 32'sd17, 32'sd2, 32'sd0, 32'sd7, 32'sd17, 32'sd5, 32'sd11, 32'sd8, 32'sd11, 32'sd5, 32'sd15, 32'sd4, 32'sd15, 32'sd6, 32'sd12, 32'sd9, 32'sd12, 32'sd4, 32'sd4, 32'sd5, 32'sd14, 32'sd9, 32'sd12, 32'sd10, 32'sd12, 32'sd2, 32'sd12, 32'sd9, 32'sd12, 32'sd8, 32'sd7, 32'sd1, 32'sd13, 32'sd2, 32'sd15, 32'sd0, 32'sd15, 32'sd6, 32'sd8, 32'sd1, 32'sd6, 32'sd10, 32'sd12, 32'sd3, 32'sd18, 32'sd1, 32'sd18, 32'sd11, 32'sd18, 32'sd6, 32'sd18, 32'sd6, 32'sd16, 32'sd12, 32'sd9, 32'sd6, 32'sd11, 32'sd6, 32'sd16, 32'sd4, 32'sd18, 32'sd8, 32'sd18, 32'sd3, 32'sd15, 32'sd6, 32'sd18, 32'sd0, 32'sd13, 32'sd7, 32'sd4, 32'sd0, 32'sd15, 32'sd3, 32'sd9, 32'sd8, 32'sd5, 32'sd3, 32'sd5, 32'sd10, 32'sd4, 32'sd2, 32'sd8, 32'sd18, 32'sd3, 32'sd4, 32'sd6, 32'sd13, 32'sd4, 32'sd12, 32'sd8, 32'sd13, 32'sd8, 32'sd3, 32'sd0, 32'sd14, 32'sd0, 32'sd14, 32'sd0, 32'sd6, 32'sd0, 32'sd14, 32'sd8, 32'sd15, 32'sd8, 32'sd10, 32'sd7, 32'sd7, 32'sd12, 32'sd11, 32'sd7, 32'sd21, 32'sd0, 32'sd15, 32'sd0, 32'sd18, 32'sd7, 32'sd16, 32'sd0, 32'sd18, 32'sd2, 32'sd14, 32'sd1, 32'sd9, 32'sd5, 32'sd5, 32'sd11, 32'sd12, 32'sd9, 32'sd12, 32'sd10, 32'sd12, 32'sd9, 32'sd13, 32'sd3, 32'sd12, 32'sd9, 32'sd13, 32'sd9, 32'sd11, 32'sd7, 32'sd5, 32'sd8, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd3, 32'sd12, 32'sd10, 32'sd12, 32'sd7, 32'sd9, 32'sd10, 32'sd11, 32'sd9, 32'sd19, 32'sd1, 32'sd15, 32'sd5, 32'sd6, 32'sd10, 32'sd12, 32'sd10, 32'sd14, 32'sd3, 32'sd7, 32'sd7, 32'sd14, 32'sd7, 32'sd18, 32'sd9, 32'sd13, 32'sd6, 32'sd10, 32'sd0, 32'sd3, 32'sd4, 32'sd16, 32'sd8, 32'sd16, 32'sd7, 32'sd15, 32'sd3, 32'sd18, 32'sd0, 32'sd13, 32'sd2, 32'sd17, 32'sd1, 32'sd8, 32'sd0, 32'sd15, 32'sd1, 32'sd20, 32'sd3, 32'sd9, 32'sd9, 32'sd7, 32'sd10, 32'sd11, 32'sd4, 32'sd10, 32'sd3, 32'sd15, 32'sd0, 32'sd6, 32'sd9, 32'sd12, 32'sd10, 32'sd16, 32'sd10, 32'sd6, 32'sd0, 32'sd17, 32'sd5, 32'sd14, 32'sd1, 32'sd7, 32'sd10, 32'sd14, 32'sd3, 32'sd9, 32'sd3, 32'sd6, 32'sd1, 32'sd16, 32'sd0, 32'sd12, 32'sd8, 32'sd10, 32'sd0, 32'sd21, 32'sd2, 32'sd20, 32'sd2, 32'sd8, 32'sd8, 32'sd11, 32'sd9, 32'sd7, 32'sd12, 32'sd11, 32'sd8, 32'sd11, 32'sd4, 32'sd12, 32'sd0, 32'sd12, 32'sd4, 32'sd12, 32'sd11, 32'sd15, 32'sd8, 32'sd13, 32'sd10, 32'sd12, 32'sd9, 32'sd17, 32'sd6, 32'sd10, 32'sd2, 32'sd2, 32'sd7, 32'sd3, 32'sd2, 32'sd15, 32'sd8, 32'sd10, 32'sd7, 32'sd18, 32'sd3, 32'sd20, 32'sd2, 32'sd17, 32'sd5, 32'sd16, 32'sd4, 32'sd11, 32'sd12, 32'sd12, 32'sd3, 32'sd13, 
                                                    32'sd0, 32'sd8, 32'sd9, 32'sd19, 32'sd9, 32'sd6, 32'sd10, 32'sd5, 32'sd12, 32'sd3, 32'sd15, 32'sd4, 32'sd11, 32'sd9, 32'sd5, 32'sd4, 32'sd11, 32'sd10, 32'sd16, 32'sd3, 32'sd13, 32'sd8, 32'sd8, 32'sd10, 32'sd5, 32'sd2, 32'sd2, 32'sd11, 32'sd9, 32'sd9, 32'sd5, 32'sd2, 32'sd6, 32'sd6, 32'sd20, 32'sd2, 32'sd10, 32'sd10, 32'sd3, 32'sd5, 32'sd17, 32'sd0, 32'sd9, 32'sd10, 32'sd11, 32'sd0, 32'sd6, 32'sd4, 32'sd9, 32'sd5, 32'sd6, 32'sd7, 32'sd11, 32'sd12, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd20, 32'sd4, 32'sd21, 32'sd1, 32'sd3, 32'sd0, 32'sd18, 32'sd7, 32'sd17, 32'sd2, 32'sd19, 32'sd0, 32'sd15, 32'sd0, 32'sd14, 32'sd0, 32'sd5, 32'sd0, 32'sd12, 32'sd5, 32'sd4, 32'sd3, 32'sd4, 32'sd10, 32'sd16, 32'sd7, 32'sd17, 32'sd3, 32'sd12, 32'sd5, 32'sd14, 32'sd6, 32'sd15, 32'sd0, 32'sd12, 32'sd0, 32'sd12, 32'sd9, 32'sd6, 32'sd0, 32'sd2, 32'sd7, 32'sd12, 32'sd6, 32'sd8, 32'sd4, 32'sd12, 32'sd10, 32'sd18, 32'sd3, 32'sd6, 32'sd5, 32'sd12, 32'sd0, 32'sd12, 32'sd11, 32'sd11, 32'sd1, 32'sd14, 32'sd1, 32'sd7, 32'sd0, 32'sd12, 32'sd12, 32'sd12, 32'sd10, 32'sd9, 32'sd1, 32'sd0, 32'sd6, 32'sd12, 32'sd5, 32'sd4, 32'sd4, 32'sd8, 32'sd1, 32'sd10, 32'sd1, 32'sd12, 32'sd1, 32'sd5, 32'sd0, 32'sd9, 32'sd1, 32'sd8, 32'sd8, 32'sd5, 32'sd9, 32'sd6, 32'sd2, 32'sd12, 32'sd10, 32'sd14, 32'sd8, 32'sd9, 32'sd12, 32'sd5, 32'sd4, 32'sd14, 32'sd9, 32'sd14, 32'sd8, 32'sd11, 32'sd5, 32'sd5, 32'sd9, 32'sd11, 32'sd2, 32'sd18, 32'sd3, 32'sd12, 32'sd5, 32'sd20, 32'sd0, 32'sd18, 32'sd1, 32'sd15, 32'sd5, 32'sd6, 32'sd2, 32'sd14, 32'sd10, 32'sd13, 32'sd3, 32'sd13, 32'sd3, 32'sd16, 32'sd0, 32'sd0, 32'sd12, 32'sd21, 32'sd0, 32'sd15, 32'sd1, 32'sd15, 32'sd0, 32'sd3, 32'sd0, 32'sd15, 32'sd0, 32'sd12, 32'sd3, 32'sd17, 32'sd0, 32'sd12}

localparam logic [2912:0][31:0] rectangle2_ys = {32'sd7, 32'sd4, 32'sd12, 32'sd20, 32'sd5, 32'sd13, 32'sd11, 32'sd19, 32'sd3, 32'sd8, 32'sd4, 32'sd12, 32'sd2, 32'sd14, 32'sd11, 32'sd3, 32'sd11, 32'sd5, 32'sd8, 32'sd5, 32'sd0, 32'sd6, 32'sd6, 32'sd20, 32'sd13, 32'sd3, 32'sd11, 32'sd13, 32'sd5, 32'sd12, 32'sd21, 32'sd8, 32'sd1, 32'sd1, 32'sd8, 32'sd6, 32'sd16, 32'sd1, 32'sd13, 32'sd1, 32'sd2, 32'sd5, 32'sd4, 32'sd3, 32'sd1, 32'sd7, 32'sd1, 32'sd1, 32'sd5, 32'sd11, 32'sd13, 32'sd7, 32'sd7, 32'sd5, 32'sd1, 32'sd12, 32'sd17, 32'sd3, 32'sd3, 32'sd1, 32'sd11, 32'sd14, 32'sd12, 32'sd8, 32'sd13, 32'sd17, 32'sd18, 32'sd10, 32'sd1, 32'sd1, 32'sd5, 32'sd12, 32'sd17, 32'sd17, 32'sd17, 32'sd6, 32'sd5, 32'sd0, 32'sd3, 32'sd6, 32'sd0, 32'sd6, 32'sd6, 32'sd8, 32'sd3, 32'sd0, 32'sd11, 32'sd6, 32'sd20, 32'sd6, 32'sd13, 32'sd6, 32'sd6, 32'sd18, 32'sd23, 32'sd12, 32'sd12, 32'sd8, 32'sd16, 32'sd19, 32'sd2, 32'sd17, 32'sd4, 32'sd4, 32'sd4, 32'sd16, 32'sd12, 32'sd0, 32'sd10, 32'sd8, 32'sd8, 32'sd0, 32'sd0, 32'sd16, 32'sd18, 32'sd8, 32'sd19, 32'sd11, 32'sd9, 32'sd0, 32'sd6, 32'sd5, 32'sd5, 32'sd15, 32'sd17, 32'sd19, 32'sd0, 32'sd6, 32'sd1, 32'sd3, 32'sd8, 32'sd11, 32'sd12, 32'sd16, 32'sd16, 32'sd5, 32'sd2, 32'sd10, 32'sd5, 32'sd20, 32'sd12, 32'sd4, 32'sd5, 32'sd1, 32'sd1, 32'sd0, 32'sd0, 32'sd7, 32'sd12, 32'sd13, 32'sd17, 32'sd14, 32'sd6, 32'sd8, 32'sd8, 32'sd15, 32'sd14, 32'sd14, 32'sd10, 32'sd15, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd20, 32'sd3, 32'sd5, 32'sd11, 32'sd11, 32'sd11, 32'sd11, 32'sd11, 32'sd12, 32'sd13, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd1, 32'sd1, 32'sd6, 32'sd16, 32'sd16, 32'sd19, 32'sd4, 32'sd18, 32'sd2, 32'sd11, 32'sd5, 32'sd13, 32'sd4, 32'sd3, 32'sd19, 32'sd0, 32'sd1, 32'sd23, 32'sd0, 32'sd12, 32'sd1, 32'sd5, 32'sd2, 32'sd3, 32'sd11, 32'sd12, 32'sd12, 32'sd7, 32'sd1, 32'sd7, 32'sd10, 32'sd6, 32'sd16, 32'sd8, 32'sd5, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd6, 32'sd7, 32'sd19, 32'sd18, 32'sd18, 32'sd20, 32'sd15, 32'sd6, 32'sd8, 32'sd14, 32'sd9, 32'sd6, 32'sd7, 32'sd11, 32'sd16, 32'sd6, 32'sd0, 32'sd0, 32'sd7, 32'sd20, 32'sd14, 32'sd2, 32'sd1, 32'sd3, 32'sd0, 32'sd21, 32'sd7, 32'sd7, 32'sd8, 32'sd15, 32'sd17, 32'sd3, 32'sd11, 32'sd1, 32'sd2, 32'sd14, 32'sd8, 32'sd2, 32'sd8, 32'sd17, 32'sd11, 32'sd1, 32'sd16, 32'sd16, 32'sd14, 32'sd14, 32'sd1, 32'sd0, 32'sd2, 32'sd2, 32'sd20, 32'sd6, 32'sd7, 32'sd10, 32'sd8, 32'sd4, 32'sd2, 32'sd6, 32'sd3, 32'sd0, 32'sd10, 32'sd10, 32'sd16, 32'sd16, 32'sd10, 32'sd0, 32'sd7, 32'sd6, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd11, 32'sd11, 32'sd14, 32'sd15, 32'sd15, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd4, 32'sd10, 32'sd19, 32'sd17, 32'sd13, 32'sd18, 32'sd19, 32'sd0, 32'sd4, 32'sd4, 32'sd3, 32'sd1, 32'sd19, 32'sd3, 32'sd5, 32'sd2, 32'sd19, 32'sd22, 32'sd14, 32'sd2, 32'sd7, 32'sd6, 32'sd12, 32'sd14, 32'sd13, 32'sd14, 32'sd7, 32'sd4, 32'sd14, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd5, 32'sd20, 32'sd5, 32'sd5, 32'sd11, 32'sd2, 32'sd0, 32'sd0, 32'sd14, 32'sd8, 32'sd14, 32'sd5, 32'sd8, 32'sd13, 32'sd14, 32'sd12, 32'sd1, 32'sd1, 32'sd12, 32'sd22, 32'sd16, 32'sd13, 32'sd6, 32'sd0, 32'sd7, 32'sd4, 32'sd0, 32'sd0, 32'sd12, 32'sd12, 32'sd14, 32'sd14, 32'sd15, 32'sd14, 32'sd17, 32'sd0, 32'sd1, 32'sd1, 32'sd17, 32'sd9, 32'sd7, 32'sd4, 32'sd6, 32'sd10, 32'sd17, 32'sd1, 32'sd11, 32'sd6, 32'sd17, 32'sd17, 32'sd7, 32'sd15, 32'sd8, 32'sd14, 32'sd16, 32'sd4, 32'sd19, 32'sd13, 32'sd3, 32'sd6, 32'sd11, 32'sd7, 32'sd6, 32'sd8, 32'sd15, 32'sd1, 32'sd8, 32'sd5, 32'sd2, 32'sd11, 32'sd11, 32'sd6, 32'sd1, 32'sd4, 32'sd18, 32'sd4, 32'sd16, 32'sd7, 32'sd7, 32'sd2, 32'sd20, 32'sd14, 32'sd2, 32'sd0, 32'sd0, 32'sd17, 32'sd8, 32'sd3, 32'sd12, 32'sd7, 32'sd8, 32'sd7, 32'sd7, 32'sd6, 32'sd23, 32'sd17, 32'sd17, 32'sd11, 32'sd11, 32'sd9, 32'sd17, 32'sd0, 32'sd0, 32'sd18, 32'sd18, 32'sd12, 32'sd6, 32'sd6, 32'sd1, 32'sd0, 32'sd15, 32'sd11, 32'sd16, 32'sd2, 32'sd20, 32'sd0, 32'sd13, 32'sd11, 32'sd7, 32'sd8, 32'sd9, 32'sd0, 32'sd0, 32'sd1, 32'sd18, 32'sd15, 32'sd15, 32'sd17, 32'sd18, 32'sd0, 32'sd4, 32'sd5, 32'sd14, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd5, 32'sd15, 32'sd0, 32'sd7, 32'sd2, 32'sd2, 32'sd2, 32'sd6, 32'sd5, 32'sd6, 32'sd0, 32'sd3, 32'sd7, 32'sd7, 32'sd13, 32'sd6, 32'sd17, 32'sd0, 32'sd2, 32'sd8, 32'sd8, 32'sd8, 32'sd3, 32'sd6, 32'sd0, 32'sd12, 32'sd21, 32'sd8, 32'sd5, 32'sd7, 32'sd12, 32'sd7, 32'sd19, 32'sd20, 32'sd14, 32'sd20, 32'sd20, 32'sd11, 32'sd11, 32'sd3, 32'sd18, 32'sd17, 32'sd20, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd11, 32'sd0, 32'sd0, 32'sd8, 32'sd12, 32'sd0, 32'sd6, 32'sd2, 32'sd3, 32'sd7, 32'sd6, 32'sd1, 32'sd10, 32'sd3, 32'sd5, 32'sd4, 32'sd1, 32'sd13, 32'sd5, 32'sd1, 32'sd2, 32'sd10, 32'sd9, 32'sd10, 32'sd10, 32'sd17, 32'sd7, 32'sd1, 32'sd1, 32'sd5, 32'sd12, 32'sd17, 32'sd15, 32'sd16, 32'sd13, 32'sd11, 32'sd6, 32'sd5, 32'sd5, 32'sd1, 32'sd1, 32'sd15, 32'sd11, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd19, 32'sd11, 32'sd8, 32'sd8, 32'sd12, 32'sd12, 32'sd2, 32'sd2, 32'sd6, 32'sd7, 32'sd6, 32'sd6, 32'sd3, 32'sd0, 32'sd13, 32'sd7, 32'sd6, 32'sd3, 32'sd15, 32'sd14, 32'sd12, 32'sd2, 32'sd16, 32'sd16, 32'sd3, 32'sd0, 32'sd10, 32'sd5, 32'sd16, 32'sd19, 32'sd6, 32'sd0, 32'sd2, 32'sd12, 32'sd0, 32'sd11, 32'sd20, 32'sd11, 32'sd14, 32'sd11, 32'sd11, 32'sd8, 32'sd17, 32'sd0, 32'sd0, 32'sd7, 32'sd1, 32'sd20, 32'sd7, 32'sd17, 32'sd2, 32'sd3, 32'sd6, 32'sd8, 32'sd12, 32'sd10, 32'sd5, 32'sd20, 32'sd0, 32'sd2, 32'sd11, 32'sd3, 32'sd17, 32'sd18, 32'sd15, 32'sd14, 32'sd8, 32'sd8, 32'sd2, 32'sd19, 32'sd20, 32'sd3, 32'sd6, 32'sd0, 32'sd0, 32'sd10, 32'sd11, 32'sd5, 32'sd8, 32'sd5, 32'sd6, 32'sd22, 32'sd10, 32'sd4, 32'sd8, 32'sd9, 32'sd10, 32'sd6, 32'sd5, 32'sd4, 32'sd4, 32'sd10, 32'sd10, 32'sd2, 32'sd2, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd20, 32'sd20, 32'sd2, 32'sd2, 32'sd5, 32'sd11, 32'sd9, 32'sd5, 
                                                    32'sd14, 32'sd14, 32'sd11, 32'sd9, 32'sd6, 32'sd21, 32'sd5, 32'sd5, 32'sd4, 32'sd7, 32'sd13, 32'sd8, 32'sd2, 32'sd19, 32'sd10, 32'sd2, 32'sd0, 32'sd3, 32'sd2, 32'sd7, 32'sd0, 32'sd3, 32'sd19, 32'sd14, 32'sd14, 32'sd5, 32'sd6, 32'sd6, 32'sd5, 32'sd5, 32'sd12, 32'sd12, 32'sd3, 32'sd3, 32'sd1, 32'sd11, 32'sd14, 32'sd11, 32'sd11, 32'sd20, 32'sd4, 32'sd3, 32'sd11, 32'sd0, 32'sd0, 32'sd11, 32'sd23, 32'sd10, 32'sd1, 32'sd0, 32'sd3, 32'sd17, 32'sd16, 32'sd12, 32'sd12, 32'sd7, 32'sd6, 32'sd8, 32'sd11, 32'sd7, 32'sd6, 32'sd9, 32'sd0, 32'sd5, 32'sd5, 32'sd5, 32'sd4, 32'sd17, 32'sd17, 32'sd13, 32'sd17, 32'sd16, 32'sd9, 32'sd0, 32'sd12, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd5, 32'sd6, 32'sd13, 32'sd5, 32'sd3, 32'sd16, 32'sd19, 32'sd13, 32'sd10, 32'sd9, 32'sd16, 32'sd14, 32'sd10, 32'sd0, 32'sd11, 32'sd2, 32'sd4, 32'sd0, 32'sd19, 32'sd8, 32'sd10, 32'sd17, 32'sd18, 32'sd18, 32'sd11, 32'sd11, 32'sd3, 32'sd5, 32'sd0, 32'sd17, 32'sd17, 32'sd17, 32'sd18, 32'sd8, 32'sd6, 32'sd12, 32'sd12, 32'sd5, 32'sd9, 32'sd9, 32'sd11, 32'sd13, 32'sd8, 32'sd8, 32'sd11, 32'sd11, 32'sd6, 32'sd0, 32'sd0, 32'sd3, 32'sd10, 32'sd7, 32'sd13, 32'sd4, 32'sd2, 32'sd5, 32'sd0, 32'sd4, 32'sd10, 32'sd10, 32'sd11, 32'sd10, 32'sd12, 32'sd21, 32'sd20, 32'sd17, 32'sd19, 32'sd18, 32'sd6, 32'sd16, 32'sd18, 32'sd6, 32'sd4, 32'sd21, 32'sd7, 32'sd2, 32'sd10, 32'sd11, 32'sd9, 32'sd10, 32'sd11, 32'sd0, 32'sd8, 32'sd0, 32'sd3, 32'sd20, 32'sd1, 32'sd0, 32'sd18, 32'sd7, 32'sd3, 32'sd2, 32'sd2, 32'sd1, 32'sd18, 32'sd15, 32'sd16, 32'sd5, 32'sd13, 32'sd3, 32'sd14, 32'sd12, 32'sd16, 32'sd8, 32'sd12, 32'sd20, 32'sd7, 32'sd2, 32'sd6, 32'sd7, 32'sd0, 32'sd11, 32'sd12, 32'sd21, 32'sd3, 32'sd9, 32'sd11, 32'sd7, 32'sd8, 32'sd16, 32'sd14, 32'sd11, 32'sd13, 32'sd0, 32'sd10, 32'sd4, 32'sd0, 32'sd6, 32'sd6, 32'sd11, 32'sd11, 32'sd16, 32'sd7, 32'sd16, 32'sd14, 32'sd11, 32'sd6, 32'sd18, 32'sd0, 32'sd5, 32'sd0, 32'sd1, 32'sd1, 32'sd17, 32'sd5, 32'sd17, 32'sd5, 32'sd9, 32'sd4, 32'sd7, 32'sd7, 32'sd4, 32'sd12, 32'sd3, 32'sd6, 32'sd9, 32'sd5, 32'sd4, 32'sd6, 32'sd2, 32'sd19, 32'sd19, 32'sd5, 32'sd8, 32'sd13, 32'sd12, 32'sd6, 32'sd11, 32'sd7, 32'sd5, 32'sd9, 32'sd14, 32'sd14, 32'sd11, 32'sd12, 32'sd0, 32'sd0, 32'sd1, 32'sd14, 32'sd20, 32'sd11, 32'sd11, 32'sd14, 32'sd16, 32'sd11, 32'sd5, 32'sd16, 32'sd15, 32'sd8, 32'sd16, 32'sd0, 32'sd5, 32'sd5, 32'sd6, 32'sd10, 32'sd10, 32'sd18, 32'sd10, 32'sd0, 32'sd4, 32'sd12, 32'sd6, 32'sd12, 32'sd16, 32'sd11, 32'sd11, 32'sd12, 32'sd4, 32'sd4, 32'sd9, 32'sd5, 32'sd9, 32'sd0, 32'sd16, 32'sd16, 32'sd7, 32'sd9, 32'sd1, 32'sd6, 32'sd18, 32'sd8, 32'sd19, 32'sd8, 32'sd8, 32'sd17, 32'sd11, 32'sd2, 32'sd12, 32'sd4, 32'sd1, 32'sd3, 32'sd6, 32'sd11, 32'sd8, 32'sd18, 32'sd16, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd12, 32'sd20, 32'sd8, 32'sd0, 32'sd10, 32'sd11, 32'sd12, 32'sd0, 32'sd0, 32'sd5, 32'sd14, 32'sd14, 32'sd1, 32'sd0, 32'sd3, 32'sd3, 32'sd10, 32'sd10, 32'sd6, 32'sd14, 32'sd17, 32'sd1, 32'sd13, 32'sd16, 32'sd17, 32'sd3, 32'sd6, 32'sd6, 32'sd1, 32'sd1, 32'sd18, 32'sd18, 32'sd1, 32'sd3, 32'sd0, 32'sd3, 32'sd5, 32'sd0, 32'sd7, 32'sd7, 32'sd3, 32'sd3, 32'sd8, 32'sd8, 32'sd13, 32'sd5, 32'sd1, 32'sd1, 32'sd15, 32'sd2, 32'sd6, 32'sd15, 32'sd12, 32'sd12, 32'sd2, 32'sd7, 32'sd11, 32'sd9, 32'sd5, 32'sd8, 32'sd19, 32'sd19, 32'sd19, 32'sd18, 32'sd19, 32'sd1, 32'sd2, 32'sd16, 32'sd16, 32'sd22, 32'sd13, 32'sd10, 32'sd8, 32'sd10, 32'sd10, 32'sd15, 32'sd7, 32'sd16, 32'sd19, 32'sd15, 32'sd9, 32'sd9, 32'sd7, 32'sd4, 32'sd8, 32'sd7, 32'sd15, 32'sd8, 32'sd19, 32'sd19, 32'sd1, 32'sd12, 32'sd5, 32'sd4, 32'sd16, 32'sd16, 32'sd0, 32'sd8, 32'sd4, 32'sd2, 32'sd1, 32'sd15, 32'sd11, 32'sd9, 32'sd5, 32'sd4, 32'sd3, 32'sd14, 32'sd11, 32'sd0, 32'sd7, 32'sd1, 32'sd11, 32'sd7, 32'sd23, 32'sd16, 32'sd0, 32'sd11, 32'sd17, 32'sd17, 32'sd5, 32'sd5, 32'sd8, 32'sd8, 32'sd2, 32'sd2, 32'sd0, 32'sd4, 32'sd18, 32'sd0, 32'sd15, 32'sd21, 32'sd5, 32'sd5, 32'sd6, 32'sd5, 32'sd16, 32'sd5, 32'sd8, 32'sd6, 32'sd13, 32'sd10, 32'sd15, 32'sd3, 32'sd8, 32'sd6, 32'sd6, 32'sd13, 32'sd15, 32'sd15, 32'sd18, 32'sd18, 32'sd17, 32'sd17, 32'sd1, 32'sd2, 32'sd2, 32'sd15, 32'sd2, 32'sd2, 32'sd5, 32'sd2, 32'sd0, 32'sd13, 32'sd2, 32'sd11, 32'sd6, 32'sd8, 32'sd11, 32'sd8, 32'sd0, 32'sd0, 32'sd6, 32'sd20, 32'sd19, 32'sd6, 32'sd8, 32'sd3, 32'sd19, 32'sd5, 32'sd6, 32'sd16, 32'sd5, 32'sd5, 32'sd4, 32'sd13, 32'sd1, 32'sd12, 32'sd7, 32'sd5, 32'sd11, 32'sd11, 32'sd5, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd13, 32'sd7, 32'sd8, 32'sd15, 32'sd10, 32'sd17, 32'sd9, 32'sd4, 32'sd13, 32'sd8, 32'sd18, 32'sd18, 32'sd20, 32'sd8, 32'sd8, 32'sd5, 32'sd5, 32'sd6, 32'sd0, 32'sd8, 32'sd8, 32'sd14, 32'sd11, 32'sd14, 32'sd14, 32'sd17, 32'sd17, 32'sd0, 32'sd0, 32'sd8, 32'sd17, 32'sd6, 32'sd22, 32'sd9, 32'sd0, 32'sd1, 32'sd18, 32'sd7, 32'sd10, 32'sd2, 32'sd12, 32'sd5, 32'sd5, 32'sd3, 32'sd13, 32'sd19, 32'sd9, 32'sd7, 32'sd1, 32'sd14, 32'sd21, 32'sd11, 32'sd6, 32'sd6, 32'sd4, 32'sd10, 32'sd17, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd1, 32'sd10, 32'sd8, 32'sd5, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd1, 32'sd3, 32'sd11, 32'sd10, 32'sd3, 32'sd6, 32'sd10, 32'sd8, 32'sd2, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd18, 32'sd16, 32'sd17, 32'sd16, 32'sd16, 32'sd8, 32'sd7, 32'sd8, 32'sd0, 32'sd8, 32'sd5, 32'sd6, 32'sd7, 32'sd8, 32'sd8, 32'sd10, 32'sd5, 32'sd12, 32'sd9, 32'sd14, 32'sd9, 32'sd18, 32'sd6, 32'sd6, 32'sd16, 32'sd17, 32'sd12, 32'sd9, 32'sd7, 32'sd10, 32'sd10, 32'sd10, 32'sd12, 32'sd17, 32'sd16, 32'sd16, 32'sd0, 32'sd1, 32'sd18, 32'sd18, 32'sd9, 32'sd0, 32'sd0, 32'sd2, 32'sd1, 32'sd8, 32'sd8, 32'sd10, 32'sd10, 32'sd7, 32'sd12, 32'sd15, 32'sd2, 32'sd1, 32'sd1, 32'sd1, 32'sd1, 32'sd11, 32'sd11, 32'sd13, 32'sd14, 32'sd13, 32'sd18, 32'sd22, 32'sd12, 32'sd7, 32'sd7, 32'sd7, 32'sd14, 32'sd14, 32'sd7, 
                                                    32'sd13, 32'sd7, 32'sd12, 32'sd7, 32'sd0, 32'sd12, 32'sd13, 32'sd13, 32'sd17, 32'sd19, 32'sd3, 32'sd5, 32'sd0, 32'sd16, 32'sd18, 32'sd15, 32'sd10, 32'sd9, 32'sd16, 32'sd9, 32'sd15, 32'sd8, 32'sd4, 32'sd9, 32'sd6, 32'sd7, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd3, 32'sd3, 32'sd11, 32'sd11, 32'sd8, 32'sd6, 32'sd19, 32'sd4, 32'sd1, 32'sd11, 32'sd12, 32'sd12, 32'sd0, 32'sd12, 32'sd21, 32'sd4, 32'sd2, 32'sd10, 32'sd7, 32'sd0, 32'sd15, 32'sd3, 32'sd7, 32'sd20, 32'sd12, 32'sd5, 32'sd11, 32'sd4, 32'sd0, 32'sd4, 32'sd4, 32'sd19, 32'sd9, 32'sd13, 32'sd13, 32'sd11, 32'sd6, 32'sd0, 32'sd9, 32'sd18, 32'sd7, 32'sd18, 32'sd14, 32'sd14, 32'sd14, 32'sd8, 32'sd9, 32'sd7, 32'sd7, 32'sd14, 32'sd18, 32'sd18, 32'sd18, 32'sd1, 32'sd21, 32'sd20, 32'sd1, 32'sd18, 32'sd17, 32'sd16, 32'sd18, 32'sd10, 32'sd18, 32'sd7, 32'sd7, 32'sd13, 32'sd6, 32'sd0, 32'sd7, 32'sd2, 32'sd18, 32'sd2, 32'sd7, 32'sd1, 32'sd0, 32'sd3, 32'sd15, 32'sd10, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd17, 32'sd20, 32'sd3, 32'sd3, 32'sd6, 32'sd6, 32'sd14, 32'sd19, 32'sd2, 32'sd1, 32'sd0, 32'sd10, 32'sd16, 32'sd16, 32'sd12, 32'sd16, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd10, 32'sd8, 32'sd10, 32'sd10, 32'sd1, 32'sd5, 32'sd10, 32'sd14, 32'sd4, 32'sd2, 32'sd4, 32'sd4, 32'sd8, 32'sd8, 32'sd17, 32'sd16, 32'sd18, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd2, 32'sd8, 32'sd3, 32'sd22, 32'sd11, 32'sd11, 32'sd11, 32'sd8, 32'sd8, 32'sd15, 32'sd15, 32'sd14, 32'sd13, 32'sd15, 32'sd4, 32'sd15, 32'sd15, 32'sd11, 32'sd8, 32'sd6, 32'sd9, 32'sd4, 32'sd7, 32'sd11, 32'sd12, 32'sd18, 32'sd2, 32'sd13, 32'sd12, 32'sd5, 32'sd7, 32'sd5, 32'sd19, 32'sd5, 32'sd5, 32'sd1, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd1, 32'sd1, 32'sd5, 32'sd4, 32'sd5, 32'sd5, 32'sd7, 32'sd0, 32'sd11, 32'sd6, 32'sd3, 32'sd18, 32'sd8, 32'sd4, 32'sd11, 32'sd4, 32'sd13, 32'sd1, 32'sd4, 32'sd7, 32'sd19, 32'sd9, 32'sd6, 32'sd5, 32'sd3, 32'sd2, 32'sd6, 32'sd3, 32'sd3, 32'sd3, 32'sd1, 32'sd2, 32'sd3, 32'sd16, 32'sd8, 32'sd0, 32'sd0, 32'sd11, 32'sd6, 32'sd9, 32'sd17, 32'sd19, 32'sd8, 32'sd17, 32'sd18, 32'sd19, 32'sd2, 32'sd5, 32'sd6, 32'sd19, 32'sd19, 32'sd18, 32'sd18, 32'sd13, 32'sd14, 32'sd18, 32'sd13, 32'sd17, 32'sd2, 32'sd9, 32'sd5, 32'sd7, 32'sd8, 32'sd9, 32'sd9, 32'sd9, 32'sd8, 32'sd12, 32'sd10, 32'sd10, 32'sd0, 32'sd3, 32'sd1, 32'sd23, 32'sd10, 32'sd0, 32'sd0, 32'sd2, 32'sd13, 32'sd21, 32'sd1, 32'sd7, 32'sd0, 32'sd1, 32'sd1, 32'sd5, 32'sd6, 32'sd5, 32'sd5, 32'sd13, 32'sd7, 32'sd9, 32'sd9, 32'sd4, 32'sd6, 32'sd21, 32'sd21, 32'sd5, 32'sd10, 32'sd0, 32'sd2, 32'sd0, 32'sd15, 32'sd13, 32'sd0, 32'sd7, 32'sd13, 32'sd22, 32'sd3, 32'sd11, 32'sd7, 32'sd7, 32'sd3, 32'sd1, 32'sd1, 32'sd18, 32'sd15, 32'sd10, 32'sd9, 32'sd11, 32'sd7, 32'sd2, 32'sd2, 32'sd4, 32'sd8, 32'sd9, 32'sd4, 32'sd11, 32'sd7, 32'sd0, 32'sd0, 32'sd1, 32'sd2, 32'sd7, 32'sd3, 32'sd14, 32'sd14, 32'sd19, 32'sd0, 32'sd4, 32'sd2, 32'sd2, 32'sd12, 32'sd15, 32'sd10, 32'sd18, 32'sd4, 32'sd0, 32'sd6, 32'sd13, 32'sd13, 32'sd13, 32'sd7, 32'sd6, 32'sd18, 32'sd20, 32'sd18, 32'sd13, 32'sd13, 32'sd9, 32'sd20, 32'sd18, 32'sd2, 32'sd2, 32'sd15, 32'sd11, 32'sd18, 32'sd19, 32'sd12, 32'sd12, 32'sd1, 32'sd15, 32'sd7, 32'sd12, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd11, 32'sd14, 32'sd21, 32'sd0, 32'sd1, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd18, 32'sd0, 32'sd0, 32'sd1, 32'sd1, 32'sd16, 32'sd3, 32'sd5, 32'sd10, 32'sd15, 32'sd10, 32'sd8, 32'sd2, 32'sd16, 32'sd6, 32'sd16, 32'sd22, 32'sd10, 32'sd6, 32'sd2, 32'sd16, 32'sd20, 32'sd0, 32'sd6, 32'sd10, 32'sd15, 32'sd7, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd19, 32'sd17, 32'sd4, 32'sd4, 32'sd16, 32'sd16, 32'sd16, 32'sd18, 32'sd0, 32'sd3, 32'sd17, 32'sd0, 32'sd12, 32'sd12, 32'sd9, 32'sd3, 32'sd7, 32'sd4, 32'sd3, 32'sd2, 32'sd5, 32'sd0, 32'sd19, 32'sd19, 32'sd15, 32'sd22, 32'sd15, 32'sd15, 32'sd6, 32'sd3, 32'sd3, 32'sd8, 32'sd4, 32'sd2, 32'sd2, 32'sd2, 32'sd7, 32'sd3, 32'sd6, 32'sd1, 32'sd8, 32'sd0, 32'sd18, 32'sd20, 32'sd19, 32'sd18, 32'sd8, 32'sd15, 32'sd18, 32'sd18, 32'sd6, 32'sd7, 32'sd6, 32'sd9, 32'sd5, 32'sd7, 32'sd4, 32'sd10, 32'sd5, 32'sd8, 32'sd0, 32'sd12, 32'sd14, 32'sd10, 32'sd17, 32'sd6, 32'sd6, 32'sd13, 32'sd10, 32'sd10, 32'sd9, 32'sd3, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd8, 32'sd8, 32'sd1, 32'sd1, 32'sd0, 32'sd10, 32'sd11, 32'sd11, 32'sd10, 32'sd16, 32'sd10, 32'sd7, 32'sd8, 32'sd0, 32'sd11, 32'sd6, 32'sd0, 32'sd15, 32'sd14, 32'sd1, 32'sd0, 32'sd3, 32'sd2, 32'sd6, 32'sd20, 32'sd20, 32'sd19, 32'sd0, 32'sd3, 32'sd12, 32'sd4, 32'sd3, 32'sd8, 32'sd15, 32'sd13, 32'sd6, 32'sd9, 32'sd0, 32'sd9, 32'sd9, 32'sd5, 32'sd4, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd3, 32'sd13, 32'sd13, 32'sd2, 32'sd13, 32'sd8, 32'sd9, 32'sd8, 32'sd14, 32'sd14, 32'sd12, 32'sd12, 32'sd17, 32'sd17, 32'sd8, 32'sd10, 32'sd10, 32'sd9, 32'sd12, 32'sd12, 32'sd12, 32'sd12, 32'sd12, 32'sd10, 32'sd15, 32'sd10, 32'sd1, 32'sd7, 32'sd5, 32'sd12, 32'sd16, 32'sd0, 32'sd10, 32'sd4, 32'sd20, 32'sd11, 32'sd18, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd7, 32'sd1, 32'sd16, 32'sd15, 32'sd8, 32'sd8, 32'sd6, 32'sd19, 32'sd18, 32'sd5, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd1, 32'sd13, 32'sd1, 32'sd18, 32'sd17, 32'sd20, 32'sd16, 32'sd1, 32'sd8, 32'sd0, 32'sd6, 32'sd5, 32'sd1, 32'sd5, 32'sd1, 32'sd11, 32'sd11, 32'sd18, 32'sd18, 32'sd15, 32'sd11, 32'sd11, 32'sd9, 32'sd15, 32'sd17, 32'sd17, 32'sd16, 32'sd16, 32'sd5, 32'sd18, 32'sd21, 32'sd21, 32'sd20, 32'sd19, 32'sd2, 32'sd4, 32'sd9, 32'sd19, 32'sd2, 32'sd10, 32'sd10, 32'sd8, 32'sd5, 32'sd5, 32'sd4, 32'sd4, 32'sd7, 32'sd6, 32'sd4, 32'sd0, 32'sd1, 32'sd1, 32'sd17, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd7, 32'sd22, 32'sd16, 32'sd3, 32'sd10, 32'sd19, 32'sd0, 32'sd5, 32'sd8, 32'sd1, 32'sd6, 32'sd3, 32'sd13, 32'sd14, 32'sd7, 32'sd7, 32'sd10, 32'sd8, 32'sd19, 32'sd14, 
                                                    32'sd6, 32'sd0, 32'sd0, 32'sd1, 32'sd14, 32'sd10, 32'sd12, 32'sd1, 32'sd1, 32'sd7, 32'sd10, 32'sd7, 32'sd8, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd4, 32'sd18, 32'sd19, 32'sd19, 32'sd18, 32'sd18, 32'sd17, 32'sd10, 32'sd19, 32'sd12, 32'sd10, 32'sd10, 32'sd2, 32'sd6, 32'sd14, 32'sd14, 32'sd1, 32'sd21, 32'sd1, 32'sd16, 32'sd1, 32'sd0, 32'sd1, 32'sd1, 32'sd9, 32'sd16, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd0, 32'sd16, 32'sd7, 32'sd11, 32'sd5, 32'sd6, 32'sd1, 32'sd1, 32'sd9, 32'sd4, 32'sd16, 32'sd0, 32'sd5, 32'sd3, 32'sd14, 32'sd16, 32'sd11, 32'sd9, 32'sd2, 32'sd6, 32'sd8, 32'sd1, 32'sd1, 32'sd16, 32'sd19, 32'sd19, 32'sd4, 32'sd20, 32'sd12, 32'sd12, 32'sd12, 32'sd12, 32'sd8, 32'sd8, 32'sd14, 32'sd14, 32'sd7, 32'sd7, 32'sd3, 32'sd1, 32'sd11, 32'sd6, 32'sd18, 32'sd23, 32'sd15, 32'sd15, 32'sd15, 32'sd19, 32'sd14, 32'sd12, 32'sd3, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd14, 32'sd3, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd6, 32'sd1, 32'sd7, 32'sd7, 32'sd20, 32'sd6, 32'sd2, 32'sd4, 32'sd4, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd15, 32'sd18, 32'sd12, 32'sd1, 32'sd8, 32'sd6, 32'sd12, 32'sd14, 32'sd14, 32'sd18, 32'sd6, 32'sd3, 32'sd6, 32'sd5, 32'sd9, 32'sd16, 32'sd8, 32'sd8, 32'sd6, 32'sd5, 32'sd10, 32'sd11, 32'sd2, 32'sd0, 32'sd4, 32'sd7, 32'sd2, 32'sd4, 32'sd0, 32'sd17, 32'sd17, 32'sd0, 32'sd3, 32'sd7, 32'sd9, 32'sd14, 32'sd14, 32'sd21, 32'sd21, 32'sd4, 32'sd8, 32'sd4, 32'sd17, 32'sd16, 32'sd11, 32'sd18, 32'sd5, 32'sd8, 32'sd8, 32'sd8, 32'sd8, 32'sd8, 32'sd6, 32'sd8, 32'sd11, 32'sd11, 32'sd3, 32'sd10, 32'sd19, 32'sd18, 32'sd11, 32'sd4, 32'sd19, 32'sd19, 32'sd18, 32'sd17, 32'sd17, 32'sd1, 32'sd1, 32'sd5, 32'sd5, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd5, 32'sd6, 32'sd2, 32'sd2, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd9, 32'sd7, 32'sd8, 32'sd0, 32'sd10, 32'sd0, 32'sd1, 32'sd1, 32'sd10, 32'sd14, 32'sd14, 32'sd10, 32'sd18, 32'sd16, 32'sd16, 32'sd16, 32'sd14, 32'sd15, 32'sd15, 32'sd0, 32'sd10, 32'sd9, 32'sd9, 32'sd11, 32'sd5, 32'sd20, 32'sd10, 32'sd8, 32'sd10, 32'sd10, 32'sd11, 32'sd8, 32'sd9, 32'sd14, 32'sd2, 32'sd0, 32'sd16, 32'sd12, 32'sd12, 32'sd6, 32'sd0, 32'sd8, 32'sd8, 32'sd11, 32'sd3, 32'sd12, 32'sd16, 32'sd6, 32'sd10, 32'sd10, 32'sd12, 32'sd12, 32'sd15, 32'sd15, 32'sd20, 32'sd20, 32'sd19, 32'sd4, 32'sd3, 32'sd15, 32'sd2, 32'sd12, 32'sd11, 32'sd1, 32'sd10, 32'sd3, 32'sd6, 32'sd0, 32'sd0, 32'sd16, 32'sd12, 32'sd6, 32'sd22, 32'sd8, 32'sd8, 32'sd2, 32'sd17, 32'sd9, 32'sd5, 32'sd9, 32'sd11, 32'sd13, 32'sd1, 32'sd18, 32'sd12, 32'sd10, 32'sd6, 32'sd18, 32'sd18, 32'sd17, 32'sd19, 32'sd14, 32'sd10, 32'sd9, 32'sd17, 32'sd8, 32'sd6, 32'sd9, 32'sd9, 32'sd17, 32'sd20, 32'sd20, 32'sd20, 32'sd17, 32'sd17, 32'sd2, 32'sd2, 32'sd0, 32'sd20, 32'sd6, 32'sd9, 32'sd9, 32'sd9, 32'sd4, 32'sd9, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd12, 32'sd12, 32'sd5, 32'sd6, 32'sd5, 32'sd16, 32'sd13, 32'sd13, 32'sd4, 32'sd4, 32'sd7, 32'sd19, 32'sd11, 32'sd2, 32'sd2, 32'sd13, 32'sd0, 32'sd11, 32'sd1, 32'sd10, 32'sd19, 32'sd10, 32'sd1, 32'sd1, 32'sd10, 32'sd10, 32'sd6, 32'sd12, 32'sd7, 32'sd7, 32'sd2, 32'sd5, 32'sd13, 32'sd4, 32'sd2, 32'sd6, 32'sd8, 32'sd20, 32'sd15, 32'sd17, 32'sd0, 32'sd0, 32'sd5, 32'sd2, 32'sd9, 32'sd6, 32'sd8, 32'sd1, 32'sd0, 32'sd0, 32'sd7, 32'sd5, 32'sd2, 32'sd12, 32'sd8, 32'sd8, 32'sd8, 32'sd11, 32'sd9, 32'sd14, 32'sd20, 32'sd22, 32'sd4, 32'sd17, 32'sd11, 32'sd12, 32'sd19, 32'sd18, 32'sd1, 32'sd1, 32'sd16, 32'sd1, 32'sd10, 32'sd8, 32'sd11, 32'sd11, 32'sd6, 32'sd6, 32'sd9, 32'sd8, 32'sd10, 32'sd5, 32'sd12, 32'sd14, 32'sd14, 32'sd10, 32'sd5, 32'sd4, 32'sd4, 32'sd8, 32'sd10, 32'sd5, 32'sd13, 32'sd13, 32'sd13, 32'sd1, 32'sd13, 32'sd13, 32'sd17, 32'sd17, 32'sd0, 32'sd10, 32'sd9, 32'sd9, 32'sd7, 32'sd7, 32'sd12, 32'sd15, 32'sd17, 32'sd14, 32'sd17, 32'sd3, 32'sd17, 32'sd4, 32'sd17, 32'sd8, 32'sd7, 32'sd4, 32'sd1, 32'sd5, 32'sd0, 32'sd11, 32'sd7, 32'sd7, 32'sd17, 32'sd6, 32'sd15, 32'sd15, 32'sd10, 32'sd10, 32'sd15, 32'sd1, 32'sd0, 32'sd0, 32'sd1, 32'sd22, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd4, 32'sd0, 32'sd3, 32'sd6, 32'sd1, 32'sd14, 32'sd20, 32'sd1, 32'sd0, 32'sd12, 32'sd0, 32'sd7, 32'sd14, 32'sd9, 32'sd1, 32'sd11, 32'sd11, 32'sd11, 32'sd5, 32'sd18, 32'sd18, 32'sd15, 32'sd17, 32'sd17, 32'sd20, 32'sd15, 32'sd2, 32'sd8, 32'sd17, 32'sd20, 32'sd8, 32'sd7, 32'sd6, 32'sd20, 32'sd20, 32'sd1, 32'sd1, 32'sd3, 32'sd6, 32'sd9, 32'sd3, 32'sd0, 32'sd9, 32'sd4, 32'sd4, 32'sd15, 32'sd15, 32'sd15, 32'sd15, 32'sd1, 32'sd2, 32'sd1, 32'sd1, 32'sd6, 32'sd2, 32'sd11, 32'sd1, 32'sd0, 32'sd6, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd13, 32'sd17, 32'sd9, 32'sd13, 32'sd19, 32'sd3, 32'sd2, 32'sd16, 32'sd0, 32'sd9, 32'sd7, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd11, 32'sd7, 32'sd6, 32'sd14, 32'sd14, 32'sd0, 32'sd0, 32'sd1, 32'sd12, 32'sd8, 32'sd6, 32'sd5, 32'sd9, 32'sd8, 32'sd12, 32'sd19, 32'sd0, 32'sd4, 32'sd16, 32'sd7, 32'sd7, 32'sd6, 32'sd18, 32'sd18, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd14, 32'sd9, 32'sd8, 32'sd8, 32'sd7, 32'sd1, 32'sd0, 32'sd15, 32'sd10, 32'sd6, 32'sd12, 32'sd4, 32'sd1, 32'sd1, 32'sd10, 32'sd4, 32'sd13, 32'sd13, 32'sd15, 32'sd14, 32'sd19, 32'sd16, 32'sd12, 32'sd12, 32'sd10, 32'sd14, 32'sd7, 32'sd15, 32'sd9, 32'sd1, 32'sd6, 32'sd19, 32'sd0, 32'sd13, 32'sd6, 32'sd6, 32'sd6, 32'sd7, 32'sd8, 32'sd8, 32'sd10, 32'sd2, 32'sd13, 32'sd13, 32'sd10, 32'sd10, 32'sd9, 32'sd2, 32'sd2, 32'sd1, 32'sd2, 32'sd3, 32'sd8, 32'sd8, 32'sd20, 32'sd6, 32'sd6, 32'sd3, 32'sd6, 32'sd8, 32'sd2, 32'sd17, 32'sd2, 32'sd3, 32'sd6, 32'sd6, 32'sd19, 32'sd7, 32'sd11, 32'sd1, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd19, 32'sd9, 32'sd8, 32'sd7, 32'sd8, 32'sd8, 32'sd2, 32'sd9, 32'sd4, 32'sd8, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd6, 32'sd0, 32'sd7, 32'sd4, 32'sd5, 32'sd15, 32'sd16, 32'sd2, 32'sd1, 
                                                    32'sd7, 32'sd7, 32'sd5, 32'sd1, 32'sd16, 32'sd14, 32'sd18, 32'sd16, 32'sd12, 32'sd9, 32'sd4, 32'sd2, 32'sd6, 32'sd6, 32'sd14, 32'sd14, 32'sd6, 32'sd13, 32'sd16, 32'sd20, 32'sd11, 32'sd6, 32'sd2, 32'sd13, 32'sd19, 32'sd15, 32'sd12, 32'sd8, 32'sd1, 32'sd0, 32'sd3, 32'sd3, 32'sd5, 32'sd5, 32'sd3, 32'sd4, 32'sd7, 32'sd7, 32'sd11, 32'sd11, 32'sd12, 32'sd17, 32'sd17, 32'sd11, 32'sd9, 32'sd6, 32'sd4, 32'sd9, 32'sd7, 32'sd11, 32'sd11, 32'sd11, 32'sd7, 32'sd7, 32'sd8, 32'sd2, 32'sd0, 32'sd6, 32'sd6, 32'sd6, 32'sd22, 32'sd21, 32'sd18, 32'sd20, 32'sd16, 32'sd16, 32'sd0, 32'sd0, 32'sd16, 32'sd16, 32'sd16, 32'sd16, 32'sd19, 32'sd19, 32'sd5, 32'sd6, 32'sd5, 32'sd2, 32'sd12, 32'sd3, 32'sd4, 32'sd4, 32'sd14, 32'sd14, 32'sd12, 32'sd11, 32'sd5, 32'sd4, 32'sd8, 32'sd8, 32'sd12, 32'sd15, 32'sd12, 32'sd12, 32'sd15, 32'sd6, 32'sd6, 32'sd0, 32'sd3, 32'sd3, 32'sd12, 32'sd13, 32'sd12, 32'sd14, 32'sd10, 32'sd10, 32'sd13, 32'sd10, 32'sd13, 32'sd13, 32'sd2, 32'sd2, 32'sd12, 32'sd13, 32'sd9, 32'sd10, 32'sd9, 32'sd1, 32'sd0, 32'sd5, 32'sd6, 32'sd0, 32'sd4, 32'sd3, 32'sd4, 32'sd16, 32'sd9, 32'sd5, 32'sd7, 32'sd7, 32'sd7, 32'sd9, 32'sd8, 32'sd8, 32'sd4, 32'sd17, 32'sd18, 32'sd17, 32'sd19, 32'sd20, 32'sd17, 32'sd11, 32'sd5, 32'sd8, 32'sd8, 32'sd6, 32'sd6, 32'sd5, 32'sd14, 32'sd14, 32'sd2, 32'sd1, 32'sd13, 32'sd2, 32'sd9, 32'sd9, 32'sd0, 32'sd0, 32'sd1, 32'sd11, 32'sd9, 32'sd13, 32'sd14, 32'sd0, 32'sd1, 32'sd1, 32'sd20, 32'sd0, 32'sd8, 32'sd8, 32'sd13, 32'sd13, 32'sd13, 32'sd13, 32'sd15, 32'sd15, 32'sd15, 32'sd8, 32'sd13, 32'sd13, 32'sd13, 32'sd13, 32'sd14, 32'sd18, 32'sd16, 32'sd20, 32'sd12, 32'sd12, 32'sd19, 32'sd6, 32'sd19, 32'sd19, 32'sd16, 32'sd14, 32'sd19, 32'sd19, 32'sd19, 32'sd19, 32'sd2, 32'sd17, 32'sd1}

localparam logic [2912:0][31:0] rectangle2_widths = {32'sd12, 32'sd4, 32'sd18, 32'sd9, 32'sd2, 32'sd12, 32'sd12, 32'sd4, 32'sd7, 32'sd12, 32'sd4, 32'sd19, 32'sd8, 32'sd6, 32'sd14, 32'sd14, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd8, 32'sd2, 32'sd10, 32'sd14, 32'sd8, 32'sd15, 32'sd5, 32'sd2, 32'sd3, 32'sd6, 32'sd13, 32'sd3, 32'sd3, 32'sd8, 32'sd7, 32'sd21, 32'sd2, 32'sd10, 32'sd2, 32'sd2, 32'sd11, 32'sd2, 32'sd2, 32'sd2, 32'sd19, 32'sd2, 32'sd2, 32'sd7, 32'sd18, 32'sd2, 32'sd6, 32'sd12, 32'sd4, 32'sd8, 32'sd18, 32'sd6, 32'sd2, 32'sd2, 32'sd8, 32'sd8, 32'sd3, 32'sd8, 32'sd12, 32'sd6, 32'sd9, 32'sd18, 32'sd16, 32'sd2, 32'sd18, 32'sd10, 32'sd14, 32'sd7, 32'sd9, 32'sd9, 32'sd4, 32'sd7, 32'sd4, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd6, 32'sd12, 32'sd8, 32'sd16, 32'sd3, 32'sd8, 32'sd2, 32'sd5, 32'sd2, 32'sd2, 32'sd6, 32'sd18, 32'sd4, 32'sd8, 32'sd10, 32'sd10, 32'sd18, 32'sd22, 32'sd18, 32'sd3, 32'sd2, 32'sd2, 32'sd10, 32'sd4, 32'sd2, 32'sd3, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd9, 32'sd9, 32'sd2, 32'sd6, 32'sd20, 32'sd9, 32'sd9, 32'sd7, 32'sd5, 32'sd6, 32'sd18, 32'sd8, 32'sd18, 32'sd3, 32'sd4, 32'sd2, 32'sd19, 32'sd11, 32'sd11, 32'sd5, 32'sd4, 32'sd4, 32'sd5, 32'sd8, 32'sd12, 32'sd3, 32'sd6, 32'sd22, 32'sd17, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd4, 32'sd19, 32'sd6, 32'sd17, 32'sd3, 32'sd4, 32'sd3, 32'sd3, 32'sd10, 32'sd3, 32'sd8, 32'sd9, 32'sd6, 32'sd5, 32'sd3, 32'sd8, 32'sd3, 32'sd10, 32'sd3, 32'sd3, 32'sd10, 32'sd2, 32'sd12, 32'sd18, 32'sd22, 32'sd4, 32'sd3, 32'sd3, 32'sd11, 32'sd12, 32'sd11, 32'sd10, 32'sd1, 32'sd1, 32'sd1, 32'sd1, 32'sd1, 32'sd9, 32'sd9, 32'sd18, 32'sd4, 32'sd18, 32'sd6, 32'sd14, 32'sd3, 32'sd6, 32'sd3, 32'sd18, 32'sd5, 32'sd2, 32'sd18, 32'sd19, 32'sd2, 32'sd19, 32'sd2, 32'sd7, 32'sd20, 32'sd22, 32'sd7, 32'sd11, 32'sd11, 32'sd2, 32'sd3, 32'sd4, 32'sd12, 32'sd6, 32'sd18, 32'sd6, 32'sd8, 32'sd2, 32'sd12, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd7, 32'sd9, 32'sd5, 32'sd5, 32'sd16, 32'sd10, 32'sd5, 32'sd5, 32'sd2, 32'sd18, 32'sd18, 32'sd9, 32'sd7, 32'sd1, 32'sd1, 32'sd5, 32'sd7, 32'sd5, 32'sd12, 32'sd11, 32'sd15, 32'sd8, 32'sd9, 32'sd5, 32'sd5, 32'sd3, 32'sd10, 32'sd10, 32'sd16, 32'sd7, 32'sd2, 32'sd3, 32'sd6, 32'sd10, 32'sd3, 32'sd5, 32'sd8, 32'sd5, 32'sd3, 32'sd6, 32'sd6, 32'sd3, 32'sd13, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd12, 32'sd2, 32'sd6, 32'sd8, 32'sd10, 32'sd6, 32'sd1, 32'sd6, 32'sd1, 32'sd1, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd8, 32'sd8, 32'sd2, 32'sd5, 32'sd1, 32'sd2, 32'sd3, 32'sd24, 32'sd13, 32'sd6, 32'sd16, 32'sd6, 32'sd6, 32'sd5, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd3, 32'sd6, 32'sd5, 32'sd3, 32'sd18, 32'sd19, 32'sd2, 32'sd1, 32'sd1, 32'sd6, 32'sd2, 32'sd9, 32'sd10, 32'sd3, 32'sd11, 32'sd5, 32'sd18, 32'sd2, 32'sd8, 32'sd12, 32'sd4, 32'sd14, 32'sd4, 32'sd5, 32'sd3, 32'sd6, 32'sd20, 32'sd19, 32'sd2, 32'sd3, 32'sd2, 32'sd3, 32'sd3, 32'sd6, 32'sd15, 32'sd6, 32'sd6, 32'sd18, 32'sd12, 32'sd2, 32'sd2, 32'sd9, 32'sd13, 32'sd9, 32'sd3, 32'sd3, 32'sd3, 32'sd9, 32'sd5, 32'sd2, 32'sd2, 32'sd6, 32'sd18, 32'sd10, 32'sd11, 32'sd8, 32'sd9, 32'sd4, 32'sd3, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd9, 32'sd9, 32'sd19, 32'sd19, 32'sd10, 32'sd5, 32'sd3, 32'sd3, 32'sd6, 32'sd9, 32'sd4, 32'sd14, 32'sd2, 32'sd6, 32'sd9, 32'sd7, 32'sd17, 32'sd11, 32'sd13, 32'sd9, 32'sd5, 32'sd6, 32'sd6, 32'sd8, 32'sd3, 32'sd24, 32'sd10, 32'sd6, 32'sd18, 32'sd16, 32'sd3, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd6, 32'sd2, 32'sd8, 32'sd5, 32'sd5, 32'sd2, 32'sd3, 32'sd19, 32'sd6, 32'sd2, 32'sd5, 32'sd5, 32'sd5, 32'sd3, 32'sd7, 32'sd9, 32'sd3, 32'sd2, 32'sd2, 32'sd9, 32'sd6, 32'sd2, 32'sd11, 32'sd6, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd19, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd18, 32'sd18, 32'sd11, 32'sd7, 32'sd15, 32'sd22, 32'sd8, 32'sd9, 32'sd12, 32'sd7, 32'sd11, 32'sd7, 32'sd12, 32'sd9, 32'sd22, 32'sd11, 32'sd6, 32'sd24, 32'sd5, 32'sd5, 32'sd12, 32'sd18, 32'sd8, 32'sd8, 32'sd18, 32'sd21, 32'sd2, 32'sd2, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd2, 32'sd8, 32'sd10, 32'sd2, 32'sd3, 32'sd3, 32'sd2, 32'sd5, 32'sd1, 32'sd5, 32'sd2, 32'sd2, 32'sd3, 32'sd7, 32'sd4, 32'sd7, 32'sd2, 32'sd6, 32'sd2, 32'sd7, 32'sd5, 32'sd4, 32'sd5, 32'sd11, 32'sd4, 32'sd8, 32'sd23, 32'sd6, 32'sd21, 32'sd2, 32'sd4, 32'sd8, 32'sd5, 32'sd10, 32'sd9, 32'sd6, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd2, 32'sd18, 32'sd21, 32'sd6, 32'sd6, 32'sd6, 32'sd8, 32'sd5, 32'sd5, 32'sd5, 32'sd3, 32'sd6, 32'sd1, 32'sd2, 32'sd3, 32'sd4, 32'sd1, 32'sd2, 32'sd9, 32'sd24, 32'sd2, 32'sd2, 32'sd2, 32'sd12, 32'sd1, 32'sd12, 32'sd18, 32'sd18, 32'sd12, 32'sd2, 32'sd2, 32'sd2, 32'sd4, 32'sd16, 32'sd4, 32'sd4, 32'sd11, 32'sd8, 32'sd2, 32'sd2, 32'sd8, 32'sd6, 32'sd18, 32'sd6, 32'sd9, 32'sd4, 32'sd3, 32'sd18, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd12, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd9, 32'sd3, 32'sd14, 32'sd3, 32'sd14, 32'sd14, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd4, 32'sd3, 32'sd8, 32'sd5, 32'sd2, 32'sd6, 32'sd18, 32'sd4, 32'sd12, 32'sd1, 32'sd5, 32'sd5, 32'sd10, 32'sd8, 32'sd15, 32'sd4, 32'sd14, 32'sd4, 32'sd3, 32'sd3, 32'sd18, 32'sd14, 32'sd3, 32'sd3, 32'sd8, 32'sd3, 32'sd10, 32'sd3, 32'sd3, 32'sd11, 32'sd10, 32'sd2, 32'sd2, 32'sd4, 32'sd20, 32'sd10, 32'sd3, 32'sd10, 32'sd2, 32'sd5, 32'sd6, 32'sd4, 32'sd4, 32'sd9, 32'sd14, 32'sd19, 32'sd5, 32'sd8, 32'sd8, 32'sd9, 32'sd18, 32'sd18, 32'sd9, 32'sd23, 32'sd18, 32'sd6, 32'sd1, 32'sd10, 32'sd10, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd1, 32'sd9, 32'sd1, 32'sd6, 32'sd18, 32'sd6, 32'sd4, 32'sd3, 32'sd3, 32'sd5, 32'sd7, 32'sd1, 32'sd5, 32'sd5, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd4, 32'sd4, 32'sd10, 32'sd21, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd20, 32'sd6, 32'sd4, 32'sd4, 32'sd10, 32'sd6, 32'sd8, 32'sd9, 32'sd4, 32'sd7, 32'sd3, 32'sd19, 32'sd6, 
                                                    32'sd18, 32'sd2, 32'sd20, 32'sd22, 32'sd2, 32'sd2, 32'sd3, 32'sd2, 32'sd10, 32'sd6, 32'sd12, 32'sd4, 32'sd4, 32'sd17, 32'sd9, 32'sd7, 32'sd7, 32'sd1, 32'sd1, 32'sd14, 32'sd9, 32'sd18, 32'sd4, 32'sd4, 32'sd7, 32'sd22, 32'sd4, 32'sd7, 32'sd9, 32'sd22, 32'sd2, 32'sd8, 32'sd3, 32'sd2, 32'sd9, 32'sd18, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd8, 32'sd6, 32'sd6, 32'sd4, 32'sd19, 32'sd3, 32'sd12, 32'sd18, 32'sd4, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd18, 32'sd20, 32'sd6, 32'sd8, 32'sd3, 32'sd7, 32'sd12, 32'sd18, 32'sd5, 32'sd5, 32'sd4, 32'sd4, 32'sd6, 32'sd2, 32'sd2, 32'sd6, 32'sd23, 32'sd19, 32'sd11, 32'sd4, 32'sd5, 32'sd9, 32'sd9, 32'sd9, 32'sd10, 32'sd3, 32'sd3, 32'sd4, 32'sd7, 32'sd5, 32'sd12, 32'sd23, 32'sd4, 32'sd18, 32'sd9, 32'sd9, 32'sd3, 32'sd3, 32'sd12, 32'sd18, 32'sd12, 32'sd18, 32'sd9, 32'sd9, 32'sd18, 32'sd2, 32'sd2, 32'sd5, 32'sd6, 32'sd2, 32'sd8, 32'sd21, 32'sd3, 32'sd11, 32'sd5, 32'sd6, 32'sd6, 32'sd22, 32'sd6, 32'sd2, 32'sd2, 32'sd3, 32'sd6, 32'sd3, 32'sd16, 32'sd2, 32'sd16, 32'sd6, 32'sd2, 32'sd4, 32'sd5, 32'sd5, 32'sd4, 32'sd4, 32'sd3, 32'sd8, 32'sd6, 32'sd9, 32'sd10, 32'sd4, 32'sd3, 32'sd6, 32'sd12, 32'sd20, 32'sd9, 32'sd9, 32'sd4, 32'sd4, 32'sd3, 32'sd4, 32'sd3, 32'sd2, 32'sd5, 32'sd7, 32'sd10, 32'sd2, 32'sd18, 32'sd8, 32'sd18, 32'sd3, 32'sd18, 32'sd4, 32'sd2, 32'sd2, 32'sd2, 32'sd12, 32'sd9, 32'sd9, 32'sd19, 32'sd11, 32'sd3, 32'sd20, 32'sd2, 32'sd8, 32'sd8, 32'sd3, 32'sd8, 32'sd16, 32'sd4, 32'sd4, 32'sd6, 32'sd2, 32'sd4, 32'sd6, 32'sd3, 32'sd7, 32'sd16, 32'sd7, 32'sd4, 32'sd2, 32'sd3, 32'sd4, 32'sd2, 32'sd4, 32'sd23, 32'sd2, 32'sd4, 32'sd10, 32'sd2, 32'sd3, 32'sd3, 32'sd6, 32'sd6, 32'sd4, 32'sd21, 32'sd4, 32'sd6, 32'sd19, 32'sd14, 32'sd6, 32'sd2, 32'sd11, 32'sd3, 32'sd2, 32'sd2, 32'sd18, 32'sd11, 32'sd20, 32'sd13, 32'sd11, 32'sd7, 32'sd5, 32'sd5, 32'sd2, 32'sd3, 32'sd4, 32'sd8, 32'sd14, 32'sd9, 32'sd18, 32'sd3, 32'sd24, 32'sd10, 32'sd18, 32'sd3, 32'sd11, 32'sd12, 32'sd4, 32'sd4, 32'sd6, 32'sd5, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd16, 32'sd20, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd9, 32'sd15, 32'sd19, 32'sd7, 32'sd9, 32'sd8, 32'sd18, 32'sd4, 32'sd9, 32'sd7, 32'sd11, 32'sd2, 32'sd5, 32'sd5, 32'sd8, 32'sd6, 32'sd4, 32'sd6, 32'sd4, 32'sd2, 32'sd4, 32'sd10, 32'sd7, 32'sd20, 32'sd4, 32'sd6, 32'sd12, 32'sd3, 32'sd4, 32'sd4, 32'sd3, 32'sd8, 32'sd3, 32'sd1, 32'sd5, 32'sd5, 32'sd10, 32'sd23, 32'sd7, 32'sd2, 32'sd6, 32'sd4, 32'sd8, 32'sd4, 32'sd4, 32'sd8, 32'sd5, 32'sd19, 32'sd8, 32'sd13, 32'sd24, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd18, 32'sd9, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd19, 32'sd6, 32'sd16, 32'sd3, 32'sd4, 32'sd15, 32'sd4, 32'sd2, 32'sd2, 32'sd6, 32'sd11, 32'sd21, 32'sd4, 32'sd3, 32'sd21, 32'sd19, 32'sd3, 32'sd3, 32'sd7, 32'sd9, 32'sd8, 32'sd11, 32'sd9, 32'sd18, 32'sd7, 32'sd8, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd1, 32'sd2, 32'sd1, 32'sd6, 32'sd2, 32'sd1, 32'sd3, 32'sd5, 32'sd1, 32'sd2, 32'sd19, 32'sd18, 32'sd9, 32'sd2, 32'sd10, 32'sd10, 32'sd3, 32'sd8, 32'sd18, 32'sd3, 32'sd4, 32'sd4, 32'sd14, 32'sd4, 32'sd5, 32'sd4, 32'sd11, 32'sd6, 32'sd9, 32'sd19, 32'sd9, 32'sd18, 32'sd9, 32'sd24, 32'sd14, 32'sd9, 32'sd6, 32'sd13, 32'sd6, 32'sd7, 32'sd3, 32'sd3, 32'sd5, 32'sd8, 32'sd9, 32'sd6, 32'sd9, 32'sd6, 32'sd7, 32'sd7, 32'sd3, 32'sd3, 32'sd5, 32'sd2, 32'sd2, 32'sd3, 32'sd9, 32'sd9, 32'sd3, 32'sd4, 32'sd4, 32'sd3, 32'sd5, 32'sd5, 32'sd12, 32'sd9, 32'sd12, 32'sd11, 32'sd11, 32'sd6, 32'sd20, 32'sd14, 32'sd16, 32'sd19, 32'sd10, 32'sd4, 32'sd21, 32'sd3, 32'sd14, 32'sd2, 32'sd9, 32'sd4, 32'sd19, 32'sd20, 32'sd2, 32'sd8, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd8, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd2, 32'sd7, 32'sd7, 32'sd3, 32'sd2, 32'sd2, 32'sd3, 32'sd10, 32'sd7, 32'sd6, 32'sd6, 32'sd2, 32'sd10, 32'sd9, 32'sd6, 32'sd5, 32'sd16, 32'sd8, 32'sd2, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd18, 32'sd18, 32'sd18, 32'sd19, 32'sd2, 32'sd5, 32'sd2, 32'sd2, 32'sd6, 32'sd11, 32'sd7, 32'sd18, 32'sd2, 32'sd18, 32'sd8, 32'sd18, 32'sd2, 32'sd2, 32'sd1, 32'sd1, 32'sd7, 32'sd9, 32'sd21, 32'sd7, 32'sd22, 32'sd12, 32'sd9, 32'sd6, 32'sd7, 32'sd7, 32'sd6, 32'sd6, 32'sd10, 32'sd3, 32'sd7, 32'sd7, 32'sd6, 32'sd3, 32'sd3, 32'sd3, 32'sd18, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd8, 32'sd9, 32'sd5, 32'sd6, 32'sd19, 32'sd4, 32'sd9, 32'sd5, 32'sd4, 32'sd6, 32'sd6, 32'sd8, 32'sd7, 32'sd10, 32'sd10, 32'sd2, 32'sd4, 32'sd4, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd9, 32'sd15, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd4, 32'sd2, 32'sd10, 32'sd4, 32'sd10, 32'sd9, 32'sd11, 32'sd6, 32'sd6, 32'sd9, 32'sd5, 32'sd6, 32'sd6, 32'sd12, 32'sd8, 32'sd8, 32'sd12, 32'sd4, 32'sd4, 32'sd4, 32'sd15, 32'sd8, 32'sd5, 32'sd6, 32'sd3, 32'sd2, 32'sd3, 32'sd20, 32'sd6, 32'sd10, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd18, 32'sd10, 32'sd4, 32'sd3, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd20, 32'sd20, 32'sd18, 32'sd6, 32'sd22, 32'sd6, 32'sd6, 32'sd24, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd18, 32'sd9, 32'sd23, 32'sd18, 32'sd9, 32'sd4, 32'sd5, 32'sd4, 32'sd3, 32'sd4, 32'sd2, 32'sd2, 32'sd6, 32'sd4, 32'sd4, 32'sd3, 32'sd3, 32'sd6, 32'sd9, 32'sd4, 32'sd11, 32'sd6, 32'sd10, 32'sd10, 32'sd5, 32'sd18, 32'sd19, 32'sd6, 32'sd11, 32'sd7, 32'sd11, 32'sd5, 32'sd3, 32'sd6, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd9, 32'sd18, 32'sd13, 32'sd4, 32'sd4, 32'sd4, 32'sd2, 32'sd3, 32'sd3, 32'sd5, 32'sd5, 32'sd6, 32'sd6, 32'sd6, 32'sd12, 32'sd1, 32'sd1, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd18, 32'sd7, 32'sd12, 32'sd9, 32'sd20, 32'sd3, 32'sd18, 32'sd18, 32'sd6, 32'sd9, 32'sd9, 32'sd3, 32'sd6, 32'sd4, 32'sd3, 32'sd4, 32'sd3, 32'sd12, 32'sd6, 32'sd6, 32'sd9, 32'sd12, 32'sd20, 32'sd4, 32'sd1, 32'sd5, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd9, 32'sd12, 32'sd2, 32'sd3, 32'sd4, 32'sd6, 32'sd8, 32'sd3, 
                                                    32'sd5, 32'sd5, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd18, 32'sd9, 32'sd5, 32'sd5, 32'sd3, 32'sd3, 32'sd5, 32'sd3, 32'sd18, 32'sd2, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd4, 32'sd5, 32'sd22, 32'sd1, 32'sd8, 32'sd10, 32'sd4, 32'sd3, 32'sd5, 32'sd20, 32'sd6, 32'sd6, 32'sd10, 32'sd4, 32'sd3, 32'sd2, 32'sd3, 32'sd2, 32'sd2, 32'sd19, 32'sd2, 32'sd2, 32'sd2, 32'sd5, 32'sd2, 32'sd2, 32'sd8, 32'sd6, 32'sd2, 32'sd6, 32'sd12, 32'sd9, 32'sd9, 32'sd18, 32'sd22, 32'sd6, 32'sd6, 32'sd16, 32'sd9, 32'sd6, 32'sd6, 32'sd2, 32'sd8, 32'sd8, 32'sd2, 32'sd18, 32'sd18, 32'sd11, 32'sd9, 32'sd7, 32'sd6, 32'sd24, 32'sd4, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd20, 32'sd6, 32'sd2, 32'sd6, 32'sd2, 32'sd1, 32'sd5, 32'sd4, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd9, 32'sd11, 32'sd5, 32'sd5, 32'sd4, 32'sd4, 32'sd5, 32'sd21, 32'sd9, 32'sd6, 32'sd6, 32'sd4, 32'sd5, 32'sd5, 32'sd4, 32'sd5, 32'sd6, 32'sd2, 32'sd3, 32'sd3, 32'sd11, 32'sd3, 32'sd4, 32'sd4, 32'sd4, 32'sd8, 32'sd18, 32'sd16, 32'sd4, 32'sd3, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd5, 32'sd7, 32'sd24, 32'sd4, 32'sd4, 32'sd12, 32'sd12, 32'sd6, 32'sd6, 32'sd4, 32'sd18, 32'sd18, 32'sd22, 32'sd12, 32'sd6, 32'sd6, 32'sd2, 32'sd9, 32'sd7, 32'sd3, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd6, 32'sd14, 32'sd17, 32'sd12, 32'sd9, 32'sd12, 32'sd9, 32'sd18, 32'sd9, 32'sd9, 32'sd24, 32'sd20, 32'sd8, 32'sd4, 32'sd10, 32'sd6, 32'sd7, 32'sd7, 32'sd3, 32'sd19, 32'sd9, 32'sd9, 32'sd10, 32'sd9, 32'sd2, 32'sd2, 32'sd4, 32'sd4, 32'sd3, 32'sd6, 32'sd10, 32'sd7, 32'sd9, 32'sd2, 32'sd3, 32'sd6, 32'sd10, 32'sd10, 32'sd5, 32'sd2, 32'sd8, 32'sd12, 32'sd2, 32'sd18, 32'sd16, 32'sd6, 32'sd7, 32'sd4, 32'sd20, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd4, 32'sd1, 32'sd3, 32'sd19, 32'sd9, 32'sd6, 32'sd2, 32'sd2, 32'sd4, 32'sd18, 32'sd14, 32'sd18, 32'sd9, 32'sd6, 32'sd7, 32'sd20, 32'sd9, 32'sd15, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd4, 32'sd8, 32'sd3, 32'sd4, 32'sd24, 32'sd6, 32'sd3, 32'sd16, 32'sd4, 32'sd5, 32'sd9, 32'sd9, 32'sd6, 32'sd20, 32'sd17, 32'sd7, 32'sd23, 32'sd2, 32'sd2, 32'sd2, 32'sd18, 32'sd3, 32'sd1, 32'sd1, 32'sd6, 32'sd5, 32'sd6, 32'sd2, 32'sd5, 32'sd5, 32'sd2, 32'sd2, 32'sd6, 32'sd18, 32'sd6, 32'sd6, 32'sd11, 32'sd5, 32'sd5, 32'sd5, 32'sd3, 32'sd5, 32'sd8, 32'sd8, 32'sd11, 32'sd4, 32'sd3, 32'sd2, 32'sd2, 32'sd7, 32'sd4, 32'sd3, 32'sd3, 32'sd4, 32'sd19, 32'sd2, 32'sd18, 32'sd5, 32'sd4, 32'sd16, 32'sd18, 32'sd5, 32'sd6, 32'sd6, 32'sd11, 32'sd3, 32'sd4, 32'sd5, 32'sd4, 32'sd4, 32'sd9, 32'sd10, 32'sd21, 32'sd11, 32'sd6, 32'sd3, 32'sd6, 32'sd6, 32'sd11, 32'sd18, 32'sd22, 32'sd6, 32'sd2, 32'sd2, 32'sd18, 32'sd3, 32'sd6, 32'sd4, 32'sd18, 32'sd6, 32'sd2, 32'sd2, 32'sd18, 32'sd2, 32'sd2, 32'sd5, 32'sd5, 32'sd5, 32'sd9, 32'sd23, 32'sd8, 32'sd6, 32'sd9, 32'sd18, 32'sd11, 32'sd11, 32'sd12, 32'sd8, 32'sd14, 32'sd21, 32'sd12, 32'sd4, 32'sd7, 32'sd6, 32'sd4, 32'sd4, 32'sd6, 32'sd3, 32'sd19, 32'sd5, 32'sd9, 32'sd2, 32'sd17, 32'sd4, 32'sd3, 32'sd16, 32'sd5, 32'sd6, 32'sd3, 32'sd20, 32'sd5, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd3, 32'sd3, 32'sd3, 32'sd7, 32'sd12, 32'sd2, 32'sd6, 32'sd2, 32'sd6, 32'sd14, 32'sd16, 32'sd2, 32'sd21, 32'sd6, 32'sd5, 32'sd8, 32'sd7, 32'sd4, 32'sd6, 32'sd6, 32'sd7, 32'sd9, 32'sd6, 32'sd8, 32'sd18, 32'sd9, 32'sd19, 32'sd24, 32'sd9, 32'sd9, 32'sd18, 32'sd18, 32'sd1, 32'sd8, 32'sd18, 32'sd1, 32'sd4, 32'sd10, 32'sd3, 32'sd10, 32'sd5, 32'sd6, 32'sd9, 32'sd4, 32'sd5, 32'sd7, 32'sd10, 32'sd4, 32'sd2, 32'sd18, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd14, 32'sd15, 32'sd4, 32'sd3, 32'sd3, 32'sd6, 32'sd4, 32'sd8, 32'sd6, 32'sd6, 32'sd12, 32'sd9, 32'sd24, 32'sd11, 32'sd9, 32'sd5, 32'sd2, 32'sd6, 32'sd6, 32'sd16, 32'sd10, 32'sd18, 32'sd9, 32'sd10, 32'sd18, 32'sd15, 32'sd15, 32'sd12, 32'sd2, 32'sd2, 32'sd3, 32'sd10, 32'sd18, 32'sd10, 32'sd5, 32'sd7, 32'sd3, 32'sd3, 32'sd3, 32'sd4, 32'sd2, 32'sd1, 32'sd8, 32'sd2, 32'sd2, 32'sd4, 32'sd4, 32'sd2, 32'sd2, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd4, 32'sd12, 32'sd12, 32'sd14, 32'sd20, 32'sd4, 32'sd13, 32'sd6, 32'sd2, 32'sd12, 32'sd15, 32'sd4, 32'sd6, 32'sd8, 32'sd1, 32'sd2, 32'sd2, 32'sd6, 32'sd17, 32'sd5, 32'sd5, 32'sd18, 32'sd4, 32'sd3, 32'sd2, 32'sd21, 32'sd3, 32'sd6, 32'sd8, 32'sd9, 32'sd5, 32'sd3, 32'sd5, 32'sd3, 32'sd3, 32'sd5, 32'sd8, 32'sd6, 32'sd3, 32'sd2, 32'sd2, 32'sd10, 32'sd18, 32'sd7, 32'sd7, 32'sd1, 32'sd5, 32'sd12, 32'sd20, 32'sd19, 32'sd9, 32'sd14, 32'sd14, 32'sd3, 32'sd18, 32'sd6, 32'sd9, 32'sd10, 32'sd10, 32'sd12, 32'sd10, 32'sd3, 32'sd3, 32'sd4, 32'sd4, 32'sd2, 32'sd10, 32'sd3, 32'sd7, 32'sd13, 32'sd4, 32'sd10, 32'sd5, 32'sd2, 32'sd6, 32'sd9, 32'sd7, 32'sd22, 32'sd18, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd2, 32'sd9, 32'sd9, 32'sd15, 32'sd3, 32'sd6, 32'sd10, 32'sd6, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd8, 32'sd2, 32'sd3, 32'sd18, 32'sd10, 32'sd10, 32'sd9, 32'sd3, 32'sd5, 32'sd4, 32'sd19, 32'sd6, 32'sd7, 32'sd16, 32'sd18, 32'sd10, 32'sd4, 32'sd6, 32'sd4, 32'sd3, 32'sd6, 32'sd6, 32'sd9, 32'sd12, 32'sd10, 32'sd10, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd10, 32'sd10, 32'sd18, 32'sd4, 32'sd24, 32'sd6, 32'sd10, 32'sd19, 32'sd10, 32'sd7, 32'sd4, 32'sd5, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd8, 32'sd8, 32'sd12, 32'sd3, 32'sd7, 32'sd7, 32'sd4, 32'sd4, 32'sd2, 32'sd1, 32'sd3, 32'sd10, 32'sd12, 32'sd4, 32'sd4, 32'sd6, 32'sd5, 32'sd7, 32'sd5, 32'sd3, 32'sd12, 32'sd4, 32'sd11, 32'sd12, 32'sd9, 32'sd23, 32'sd19, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd8, 32'sd7, 32'sd9, 32'sd2, 32'sd2, 32'sd10, 32'sd3, 32'sd5, 32'sd4, 32'sd4, 32'sd4, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd24, 32'sd10, 32'sd23, 32'sd19, 32'sd18, 32'sd9, 32'sd6, 32'sd6, 32'sd20, 32'sd3, 32'sd18, 32'sd3, 32'sd6, 32'sd6, 32'sd6, 32'sd5, 32'sd2, 32'sd2, 32'sd2, 
                                                    32'sd6, 32'sd2, 32'sd5, 32'sd2, 32'sd1, 32'sd2, 32'sd2, 32'sd19, 32'sd9, 32'sd7, 32'sd14, 32'sd8, 32'sd8, 32'sd9, 32'sd9, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd2, 32'sd4, 32'sd9, 32'sd7, 32'sd5, 32'sd10, 32'sd4, 32'sd22, 32'sd2, 32'sd3, 32'sd2, 32'sd5, 32'sd4, 32'sd6, 32'sd12, 32'sd6, 32'sd6, 32'sd2, 32'sd19, 32'sd6, 32'sd8, 32'sd6, 32'sd6, 32'sd6, 32'sd24, 32'sd10, 32'sd10, 32'sd19, 32'sd19, 32'sd16, 32'sd8, 32'sd6, 32'sd2, 32'sd18, 32'sd18, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd6, 32'sd10, 32'sd2, 32'sd3, 32'sd2, 32'sd3, 32'sd3, 32'sd15, 32'sd20, 32'sd2, 32'sd6, 32'sd2, 32'sd3, 32'sd2, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd2, 32'sd4, 32'sd18, 32'sd2, 32'sd19, 32'sd15, 32'sd7, 32'sd11, 32'sd2, 32'sd18, 32'sd3, 32'sd20, 32'sd5, 32'sd4, 32'sd3, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd1, 32'sd7, 32'sd4, 32'sd4, 32'sd5, 32'sd3, 32'sd10, 32'sd18, 32'sd15, 32'sd8, 32'sd24, 32'sd2, 32'sd4, 32'sd10, 32'sd18, 32'sd24, 32'sd2, 32'sd4, 32'sd18, 32'sd18, 32'sd9, 32'sd10, 32'sd7, 32'sd6, 32'sd7, 32'sd7, 32'sd6, 32'sd6, 32'sd2, 32'sd18, 32'sd2, 32'sd10, 32'sd11, 32'sd4, 32'sd9, 32'sd2, 32'sd4, 32'sd4, 32'sd4, 32'sd3, 32'sd4, 32'sd3, 32'sd4, 32'sd4, 32'sd14, 32'sd11, 32'sd2, 32'sd11, 32'sd9, 32'sd18, 32'sd4, 32'sd18, 32'sd18, 32'sd9, 32'sd9, 32'sd9, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd6, 32'sd2, 32'sd5, 32'sd5, 32'sd2, 32'sd3, 32'sd4, 32'sd4, 32'sd24, 32'sd7, 32'sd4, 32'sd5, 32'sd4, 32'sd2, 32'sd3, 32'sd3, 32'sd18, 32'sd16, 32'sd16, 32'sd4, 32'sd8, 32'sd4, 32'sd9, 32'sd9, 32'sd16, 32'sd19, 32'sd9, 32'sd1, 32'sd24, 32'sd5, 32'sd19, 32'sd3, 32'sd12, 32'sd9, 32'sd10, 32'sd20, 32'sd7, 32'sd7, 32'sd2, 32'sd5, 32'sd6, 32'sd3, 32'sd6, 32'sd2, 32'sd9, 32'sd11, 32'sd11, 32'sd3, 32'sd2, 32'sd6, 32'sd24, 32'sd8, 32'sd6, 32'sd2, 32'sd5, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd5, 32'sd5, 32'sd9, 32'sd14, 32'sd10, 32'sd5, 32'sd1, 32'sd3, 32'sd5, 32'sd8, 32'sd12, 32'sd2, 32'sd3, 32'sd2, 32'sd2, 32'sd19, 32'sd4, 32'sd2, 32'sd18, 32'sd10, 32'sd18, 32'sd3, 32'sd24, 32'sd4, 32'sd2, 32'sd4, 32'sd5, 32'sd9, 32'sd19, 32'sd8, 32'sd8, 32'sd10, 32'sd6, 32'sd7, 32'sd6, 32'sd6, 32'sd15, 32'sd6, 32'sd7, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd18, 32'sd18, 32'sd2, 32'sd2, 32'sd1, 32'sd8, 32'sd2, 32'sd5, 32'sd6, 32'sd7, 32'sd2, 32'sd6, 32'sd5, 32'sd9, 32'sd1, 32'sd1, 32'sd3, 32'sd3, 32'sd6, 32'sd3, 32'sd3, 32'sd5, 32'sd5, 32'sd5, 32'sd2, 32'sd2, 32'sd5, 32'sd7, 32'sd6, 32'sd24, 32'sd7, 32'sd2, 32'sd2, 32'sd7, 32'sd8, 32'sd7, 32'sd5, 32'sd3, 32'sd8, 32'sd8, 32'sd3, 32'sd3, 32'sd5, 32'sd6, 32'sd12, 32'sd5, 32'sd9, 32'sd11, 32'sd4, 32'sd9, 32'sd13, 32'sd2, 32'sd2, 32'sd10, 32'sd20, 32'sd9, 32'sd2, 32'sd2, 32'sd22, 32'sd9, 32'sd24, 32'sd16, 32'sd18, 32'sd2, 32'sd3, 32'sd3, 32'sd4, 32'sd7, 32'sd10, 32'sd19, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd6, 32'sd2, 32'sd8, 32'sd18, 32'sd5, 32'sd12, 32'sd6, 32'sd10, 32'sd24, 32'sd9, 32'sd2, 32'sd2, 32'sd8, 32'sd2, 32'sd3, 32'sd6, 32'sd5, 32'sd5, 32'sd3, 32'sd3, 32'sd7, 32'sd3, 32'sd6, 32'sd2, 32'sd16, 32'sd7, 32'sd8, 32'sd3, 32'sd3, 32'sd1, 32'sd11, 32'sd18, 32'sd6, 32'sd3, 32'sd4, 32'sd4, 32'sd10, 32'sd1, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd10, 32'sd9, 32'sd18, 32'sd3, 32'sd2, 32'sd18, 32'sd3, 32'sd10, 32'sd3, 32'sd1, 32'sd3, 32'sd11, 32'sd3, 32'sd11, 32'sd4, 32'sd10, 32'sd7, 32'sd6, 32'sd2, 32'sd4, 32'sd4, 32'sd4, 32'sd3, 32'sd4, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd5, 32'sd3, 32'sd3, 32'sd5, 32'sd8, 32'sd19, 32'sd9, 32'sd9, 32'sd6, 32'sd3, 32'sd14, 32'sd4, 32'sd7, 32'sd4, 32'sd4, 32'sd22, 32'sd6, 32'sd3, 32'sd3, 32'sd17, 32'sd6, 32'sd9, 32'sd10, 32'sd5, 32'sd8, 32'sd3, 32'sd3, 32'sd19, 32'sd6, 32'sd10, 32'sd10, 32'sd9, 32'sd18, 32'sd18, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd8, 32'sd6, 32'sd2, 32'sd6, 32'sd2, 32'sd6, 32'sd6, 32'sd3, 32'sd3, 32'sd2, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd6, 32'sd4, 32'sd4, 32'sd9, 32'sd9, 32'sd6, 32'sd9, 32'sd18, 32'sd3, 32'sd3, 32'sd3, 32'sd7, 32'sd2, 32'sd6, 32'sd6, 32'sd3, 32'sd16, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd5, 32'sd9, 32'sd18, 32'sd5, 32'sd17, 32'sd9, 32'sd24, 32'sd18, 32'sd2, 32'sd14, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd7, 32'sd4, 32'sd3, 32'sd3, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd6, 32'sd9, 32'sd10, 32'sd3, 32'sd4, 32'sd8, 32'sd5, 32'sd5, 32'sd5, 32'sd6, 32'sd5, 32'sd6, 32'sd5, 32'sd5, 32'sd6, 32'sd18, 32'sd18, 32'sd2, 32'sd4, 32'sd4, 32'sd4, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd6, 32'sd3, 32'sd2, 32'sd10, 32'sd10, 32'sd4, 32'sd1, 32'sd1, 32'sd1, 32'sd6, 32'sd5, 32'sd7, 32'sd7, 32'sd3, 32'sd4, 32'sd4, 32'sd5, 32'sd9, 32'sd9, 32'sd12, 32'sd5, 32'sd3, 32'sd2, 32'sd7, 32'sd2, 32'sd7, 32'sd19, 32'sd3, 32'sd5, 32'sd5, 32'sd4, 32'sd6, 32'sd3, 32'sd7, 32'sd7, 32'sd13, 32'sd3, 32'sd17, 32'sd17, 32'sd8, 32'sd8, 32'sd12, 32'sd5, 32'sd6, 32'sd9, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd11, 32'sd4, 32'sd4, 32'sd3, 32'sd6, 32'sd3, 32'sd3, 32'sd6, 32'sd3, 32'sd8, 32'sd5, 32'sd7, 32'sd11, 32'sd6, 32'sd4, 32'sd2, 32'sd1, 32'sd1, 32'sd9, 32'sd4, 32'sd3, 32'sd9, 32'sd1, 32'sd1, 32'sd5, 32'sd18, 32'sd20, 32'sd9, 32'sd19, 32'sd19, 32'sd9, 32'sd6, 32'sd7, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd4, 32'sd4, 32'sd2, 32'sd3, 32'sd3, 32'sd9, 32'sd8, 32'sd10, 32'sd9, 32'sd3, 32'sd5, 32'sd3, 32'sd12, 32'sd4, 32'sd4, 32'sd6, 32'sd12, 32'sd6, 32'sd6, 32'sd7, 32'sd6, 32'sd19, 32'sd6, 32'sd2, 32'sd2, 32'sd5, 32'sd5, 32'sd7, 32'sd3, 32'sd8, 32'sd10, 32'sd18, 32'sd2, 32'sd20, 32'sd2, 32'sd6, 32'sd6, 32'sd18, 32'sd15, 32'sd18, 32'sd1, 32'sd2, 32'sd2, 32'sd4, 32'sd4, 32'sd20, 32'sd13, 32'sd7, 32'sd7, 32'sd5, 32'sd5, 32'sd3, 32'sd18, 32'sd18, 32'sd9, 32'sd15, 32'sd6, 32'sd12, 32'sd3, 32'sd13, 32'sd11, 32'sd6, 32'sd6, 32'sd24, 
                                                    32'sd10, 32'sd18, 32'sd10, 32'sd1, 32'sd6, 32'sd2, 32'sd2, 32'sd18, 32'sd9, 32'sd6, 32'sd9, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd9, 32'sd9, 32'sd10, 32'sd10, 32'sd18, 32'sd18, 32'sd9, 32'sd7, 32'sd19, 32'sd16, 32'sd8, 32'sd6, 32'sd1, 32'sd1, 32'sd4, 32'sd4, 32'sd3, 32'sd6, 32'sd4, 32'sd6, 32'sd9, 32'sd9, 32'sd3, 32'sd18, 32'sd3, 32'sd3, 32'sd18, 32'sd18, 32'sd22, 32'sd7, 32'sd6, 32'sd6, 32'sd8, 32'sd16, 32'sd6, 32'sd4, 32'sd3, 32'sd3, 32'sd18, 32'sd10, 32'sd9, 32'sd9, 32'sd1, 32'sd1, 32'sd2, 32'sd6, 32'sd8, 32'sd9, 32'sd16, 32'sd18, 32'sd2, 32'sd3, 32'sd2, 32'sd2, 32'sd6, 32'sd18, 32'sd24, 32'sd9, 32'sd4, 32'sd13, 32'sd16, 32'sd14, 32'sd9, 32'sd16, 32'sd13, 32'sd13, 32'sd12, 32'sd10, 32'sd18, 32'sd18, 32'sd9, 32'sd11, 32'sd8, 32'sd8, 32'sd18, 32'sd5, 32'sd6, 32'sd9, 32'sd2, 32'sd3, 32'sd2, 32'sd2, 32'sd5, 32'sd9, 32'sd17, 32'sd12, 32'sd8, 32'sd5, 32'sd2, 32'sd2, 32'sd2, 32'sd13, 32'sd19, 32'sd6, 32'sd4, 32'sd3, 32'sd3, 32'sd3, 32'sd9, 32'sd2, 32'sd4, 32'sd4, 32'sd5, 32'sd5, 32'sd4, 32'sd4, 32'sd16, 32'sd16, 32'sd7, 32'sd3, 32'sd9, 32'sd17, 32'sd8, 32'sd8, 32'sd5, 32'sd11, 32'sd12, 32'sd6, 32'sd3, 32'sd3, 32'sd9, 32'sd11, 32'sd9, 32'sd18, 32'sd19, 32'sd18, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd1, 32'sd24, 32'sd3}

localparam logic [2912:0][31:0] rectangle2_heights = {32'sd3, 32'sd7, 32'sd3, 32'sd2, 32'sd19, 32'sd8, 32'sd3, 32'sd5, 32'sd3, 32'sd2, 32'sd7, 32'sd4, 32'sd3, 32'sd5, 32'sd5, 32'sd3, 32'sd6, 32'sd10, 32'sd10, 32'sd9, 32'sd11, 32'sd13, 32'sd9, 32'sd2, 32'sd6, 32'sd3, 32'sd3, 32'sd7, 32'sd10, 32'sd6, 32'sd3, 32'sd2, 32'sd15, 32'sd15, 32'sd15, 32'sd6, 32'sd4, 32'sd10, 32'sd10, 32'sd13, 32'sd13, 32'sd19, 32'sd9, 32'sd11, 32'sd9, 32'sd1, 32'sd9, 32'sd9, 32'sd7, 32'sd1, 32'sd11, 32'sd3, 32'sd3, 32'sd6, 32'sd5, 32'sd2, 32'sd3, 32'sd13, 32'sd13, 32'sd23, 32'sd4, 32'sd7, 32'sd3, 32'sd2, 32'sd6, 32'sd2, 32'sd1, 32'sd6, 32'sd20, 32'sd1, 32'sd7, 32'sd4, 32'sd3, 32'sd2, 32'sd2, 32'sd5, 32'sd7, 32'sd5, 32'sd3, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd4, 32'sd3, 32'sd6, 32'sd4, 32'sd6, 32'sd3, 32'sd9, 32'sd4, 32'sd9, 32'sd9, 32'sd6, 32'sd1, 32'sd5, 32'sd5, 32'sd2, 32'sd2, 32'sd1, 32'sd1, 32'sd1, 32'sd15, 32'sd10, 32'sd10, 32'sd3, 32'sd9, 32'sd9, 32'sd6, 32'sd3, 32'sd3, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd10, 32'sd3, 32'sd1, 32'sd6, 32'sd24, 32'sd5, 32'sd6, 32'sd6, 32'sd1, 32'sd4, 32'sd3, 32'sd6, 32'sd18, 32'sd14, 32'sd1, 32'sd13, 32'sd2, 32'sd10, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd2, 32'sd6, 32'sd3, 32'sd5, 32'sd3, 32'sd10, 32'sd8, 32'sd7, 32'sd22, 32'sd22, 32'sd16, 32'sd2, 32'sd4, 32'sd2, 32'sd7, 32'sd5, 32'sd11, 32'sd11, 32'sd9, 32'sd7, 32'sd8, 32'sd14, 32'sd3, 32'sd8, 32'sd6, 32'sd4, 32'sd6, 32'sd2, 32'sd6, 32'sd6, 32'sd2, 32'sd9, 32'sd2, 32'sd1, 32'sd1, 32'sd8, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd6, 32'sd17, 32'sd24, 32'sd24, 32'sd22, 32'sd22, 32'sd18, 32'sd2, 32'sd2, 32'sd1, 32'sd9, 32'sd1, 32'sd4, 32'sd3, 32'sd6, 32'sd8, 32'sd16, 32'sd3, 32'sd4, 32'sd9, 32'sd1, 32'sd1, 32'sd9, 32'sd6, 32'sd9, 32'sd6, 32'sd1, 32'sd1, 32'sd3, 32'sd2, 32'sd2, 32'sd11, 32'sd6, 32'sd5, 32'sd6, 32'sd5, 32'sd1, 32'sd3, 32'sd3, 32'sd9, 32'sd7, 32'sd13, 32'sd13, 32'sd9, 32'sd9, 32'sd2, 32'sd3, 32'sd2, 32'sd4, 32'sd9, 32'sd2, 32'sd2, 32'sd10, 32'sd7, 32'sd9, 32'sd1, 32'sd1, 32'sd2, 32'sd3, 32'sd18, 32'sd18, 32'sd10, 32'sd4, 32'sd9, 32'sd3, 32'sd4, 32'sd3, 32'sd19, 32'sd3, 32'sd4, 32'sd4, 32'sd8, 32'sd2, 32'sd2, 32'sd3, 32'sd5, 32'sd13, 32'sd14, 32'sd5, 32'sd2, 32'sd14, 32'sd4, 32'sd5, 32'sd4, 32'sd6, 32'sd3, 32'sd3, 32'sd8, 32'sd2, 32'sd9, 32'sd6, 32'sd9, 32'sd9, 32'sd2, 32'sd9, 32'sd3, 32'sd7, 32'sd4, 32'sd3, 32'sd20, 32'sd3, 32'sd21, 32'sd23, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd4, 32'sd19, 32'sd6, 32'sd10, 32'sd6, 32'sd19, 32'sd10, 32'sd6, 32'sd1, 32'sd2, 32'sd3, 32'sd2, 32'sd3, 32'sd3, 32'sd4, 32'sd9, 32'sd9, 32'sd9, 32'sd15, 32'sd15, 32'sd2, 32'sd7, 32'sd5, 32'sd4, 32'sd8, 32'sd1, 32'sd1, 32'sd9, 32'sd18, 32'sd18, 32'sd9, 32'sd14, 32'sd3, 32'sd8, 32'sd6, 32'sd8, 32'sd5, 32'sd1, 32'sd10, 32'sd4, 32'sd3, 32'sd5, 32'sd4, 32'sd5, 32'sd7, 32'sd8, 32'sd8, 32'sd1, 32'sd2, 32'sd9, 32'sd14, 32'sd12, 32'sd9, 32'sd9, 32'sd3, 32'sd2, 32'sd3, 32'sd3, 32'sd1, 32'sd2, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd15, 32'sd6, 32'sd7, 32'sd2, 32'sd4, 32'sd19, 32'sd19, 32'sd3, 32'sd1, 32'sd3, 32'sd2, 32'sd3, 32'sd11, 32'sd7, 32'sd10, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd1, 32'sd1, 32'sd2, 32'sd6, 32'sd6, 32'sd6, 32'sd3, 32'sd6, 32'sd6, 32'sd4, 32'sd9, 32'sd3, 32'sd2, 32'sd23, 32'sd2, 32'sd6, 32'sd2, 32'sd2, 32'sd4, 32'sd3, 32'sd3, 32'sd4, 32'sd6, 32'sd1, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd6, 32'sd4, 32'sd9, 32'sd10, 32'sd9, 32'sd21, 32'sd7, 32'sd9, 32'sd4, 32'sd4, 32'sd4, 32'sd9, 32'sd17, 32'sd3, 32'sd3, 32'sd19, 32'sd7, 32'sd6, 32'sd6, 32'sd6, 32'sd4, 32'sd2, 32'sd6, 32'sd14, 32'sd14, 32'sd2, 32'sd5, 32'sd11, 32'sd7, 32'sd3, 32'sd2, 32'sd3, 32'sd3, 32'sd2, 32'sd1, 32'sd3, 32'sd3, 32'sd9, 32'sd9, 32'sd7, 32'sd5, 32'sd9, 32'sd9, 32'sd1, 32'sd1, 32'sd6, 32'sd3, 32'sd2, 32'sd1, 32'sd24, 32'sd4, 32'sd3, 32'sd4, 32'sd3, 32'sd3, 32'sd8, 32'sd2, 32'sd1, 32'sd4, 32'sd3, 32'sd2, 32'sd5, 32'sd5, 32'sd2, 32'sd1, 32'sd3, 32'sd3, 32'sd1, 32'sd5, 32'sd24, 32'sd11, 32'sd6, 32'sd10, 32'sd24, 32'sd24, 32'sd7, 32'sd12, 32'sd14, 32'sd2, 32'sd9, 32'sd7, 32'sd15, 32'sd9, 32'sd7, 32'sd18, 32'sd6, 32'sd10, 32'sd9, 32'sd7, 32'sd3, 32'sd6, 32'sd6, 32'sd9, 32'sd3, 32'sd13, 32'sd3, 32'sd4, 32'sd5, 32'sd4, 32'sd3, 32'sd5, 32'sd5, 32'sd2, 32'sd3, 32'sd2, 32'sd12, 32'sd5, 32'sd5, 32'sd12, 32'sd2, 32'sd2, 32'sd8, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd1, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd5, 32'sd8, 32'sd5, 32'sd5, 32'sd10, 32'sd3, 32'sd18, 32'sd9, 32'sd7, 32'sd5, 32'sd18, 32'sd9, 32'sd2, 32'sd1, 32'sd9, 32'sd10, 32'sd12, 32'sd6, 32'sd21, 32'sd4, 32'sd4, 32'sd1, 32'sd2, 32'sd9, 32'sd9, 32'sd22, 32'sd7, 32'sd5, 32'sd7, 32'sd7, 32'sd3, 32'sd9, 32'sd16, 32'sd16, 32'sd4, 32'sd3, 32'sd1, 32'sd3, 32'sd2, 32'sd5, 32'sd6, 32'sd1, 32'sd11, 32'sd11, 32'sd9, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd17, 32'sd17, 32'sd2, 32'sd6, 32'sd6, 32'sd6, 32'sd5, 32'sd5, 32'sd2, 32'sd2, 32'sd14, 32'sd9, 32'sd15, 32'sd15, 32'sd9, 32'sd21, 32'sd4, 32'sd6, 32'sd9, 32'sd3, 32'sd1, 32'sd5, 32'sd2, 32'sd20, 32'sd4, 32'sd4, 32'sd3, 32'sd3, 32'sd2, 32'sd6, 32'sd3, 32'sd5, 32'sd7, 32'sd6, 32'sd1, 32'sd6, 32'sd6, 32'sd6, 32'sd3, 32'sd7, 32'sd2, 32'sd6, 32'sd7, 32'sd4, 32'sd2, 32'sd9, 32'sd9, 32'sd5, 32'sd1, 32'sd2, 32'sd11, 32'sd3, 32'sd9, 32'sd4, 32'sd3, 32'sd5, 32'sd8, 32'sd2, 32'sd3, 32'sd4, 32'sd8, 32'sd18, 32'sd11, 32'sd5, 32'sd1, 32'sd1, 32'sd2, 32'sd5, 32'sd1, 32'sd3, 32'sd22, 32'sd2, 32'sd2, 32'sd12, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd9, 32'sd19, 32'sd2, 32'sd19, 32'sd3, 32'sd1, 32'sd4, 32'sd5, 32'sd6, 32'sd8, 32'sd4, 32'sd3, 32'sd19, 32'sd20, 32'sd20, 32'sd6, 32'sd6, 32'sd7, 32'sd7, 32'sd7, 32'sd9, 32'sd10, 32'sd10, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd3, 32'sd3, 32'sd2, 32'sd3, 32'sd5, 32'sd5, 32'sd13, 32'sd5, 32'sd3, 32'sd2, 32'sd5, 32'sd6, 32'sd6, 32'sd1, 32'sd3, 32'sd1, 32'sd9, 32'sd1, 32'sd1, 32'sd9, 32'sd23, 
                                                    32'sd19, 32'sd9, 32'sd2, 32'sd6, 32'sd3, 32'sd5, 32'sd5, 32'sd3, 32'sd4, 32'sd3, 32'sd3, 32'sd18, 32'sd18, 32'sd2, 32'sd2, 32'sd3, 32'sd8, 32'sd5, 32'sd4, 32'sd2, 32'sd5, 32'sd4, 32'sd2, 32'sd2, 32'sd17, 32'sd9, 32'sd6, 32'sd9, 32'sd6, 32'sd1, 32'sd3, 32'sd11, 32'sd10, 32'sd17, 32'sd2, 32'sd3, 32'sd4, 32'sd4, 32'sd5, 32'sd1, 32'sd7, 32'sd3, 32'sd1, 32'sd6, 32'sd14, 32'sd9, 32'sd18, 32'sd18, 32'sd10, 32'sd11, 32'sd1, 32'sd1, 32'sd4, 32'sd4, 32'sd6, 32'sd7, 32'sd5, 32'sd1, 32'sd4, 32'sd4, 32'sd9, 32'sd9, 32'sd6, 32'sd9, 32'sd11, 32'sd6, 32'sd1, 32'sd1, 32'sd2, 32'sd5, 32'sd4, 32'sd3, 32'sd2, 32'sd2, 32'sd4, 32'sd18, 32'sd10, 32'sd5, 32'sd6, 32'sd7, 32'sd2, 32'sd2, 32'sd5, 32'sd1, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd3, 32'sd1, 32'sd2, 32'sd1, 32'sd2, 32'sd2, 32'sd1, 32'sd10, 32'sd9, 32'sd4, 32'sd4, 32'sd11, 32'sd3, 32'sd2, 32'sd6, 32'sd4, 32'sd4, 32'sd3, 32'sd4, 32'sd11, 32'sd4, 32'sd9, 32'sd9, 32'sd7, 32'sd8, 32'sd7, 32'sd10, 32'sd10, 32'sd2, 32'sd4, 32'sd9, 32'sd5, 32'sd4, 32'sd4, 32'sd5, 32'sd5, 32'sd8, 32'sd3, 32'sd4, 32'sd2, 32'sd2, 32'sd6, 32'sd6, 32'sd3, 32'sd2, 32'sd1, 32'sd3, 32'sd2, 32'sd6, 32'sd6, 32'sd8, 32'sd5, 32'sd6, 32'sd9, 32'sd4, 32'sd6, 32'sd2, 32'sd15, 32'sd1, 32'sd3, 32'sd1, 32'sd6, 32'sd1, 32'sd5, 32'sd9, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd1, 32'sd6, 32'sd6, 32'sd1, 32'sd10, 32'sd3, 32'sd3, 32'sd7, 32'sd3, 32'sd4, 32'sd6, 32'sd5, 32'sd3, 32'sd9, 32'sd6, 32'sd3, 32'sd6, 32'sd3, 32'sd3, 32'sd3, 32'sd7, 32'sd9, 32'sd7, 32'sd8, 32'sd10, 32'sd5, 32'sd1, 32'sd12, 32'sd5, 32'sd2, 32'sd12, 32'sd6, 32'sd6, 32'sd13, 32'sd13, 32'sd6, 32'sd1, 32'sd6, 32'sd7, 32'sd1, 32'sd2, 32'sd4, 32'sd9, 32'sd2, 32'sd6, 32'sd23, 32'sd23, 32'sd1, 32'sd2, 32'sd1, 32'sd2, 32'sd15, 32'sd3, 32'sd4, 32'sd4, 32'sd9, 32'sd6, 32'sd5, 32'sd3, 32'sd3, 32'sd2, 32'sd1, 32'sd6, 32'sd1, 32'sd2, 32'sd1, 32'sd8, 32'sd2, 32'sd11, 32'sd5, 32'sd6, 32'sd3, 32'sd10, 32'sd9, 32'sd10, 32'sd10, 32'sd10, 32'sd3, 32'sd1, 32'sd13, 32'sd13, 32'sd7, 32'sd3, 32'sd2, 32'sd2, 32'sd1, 32'sd8, 32'sd2, 32'sd4, 32'sd1, 32'sd6, 32'sd2, 32'sd7, 32'sd3, 32'sd9, 32'sd5, 32'sd5, 32'sd3, 32'sd3, 32'sd7, 32'sd6, 32'sd6, 32'sd9, 32'sd8, 32'sd2, 32'sd7, 32'sd1, 32'sd8, 32'sd5, 32'sd2, 32'sd7, 32'sd8, 32'sd8, 32'sd6, 32'sd6, 32'sd8, 32'sd18, 32'sd7, 32'sd7, 32'sd3, 32'sd6, 32'sd3, 32'sd9, 32'sd3, 32'sd8, 32'sd4, 32'sd8, 32'sd8, 32'sd5, 32'sd4, 32'sd1, 32'sd9, 32'sd4, 32'sd1, 32'sd11, 32'sd9, 32'sd4, 32'sd3, 32'sd1, 32'sd2, 32'sd9, 32'sd9, 32'sd19, 32'sd19, 32'sd8, 32'sd8, 32'sd1, 32'sd4, 32'sd2, 32'sd6, 32'sd7, 32'sd6, 32'sd5, 32'sd9, 32'sd9, 32'sd4, 32'sd2, 32'sd1, 32'sd6, 32'sd6, 32'sd1, 32'sd1, 32'sd7, 32'sd7, 32'sd7, 32'sd2, 32'sd3, 32'sd2, 32'sd2, 32'sd1, 32'sd3, 32'sd4, 32'sd5, 32'sd9, 32'sd10, 32'sd10, 32'sd3, 32'sd3, 32'sd19, 32'sd9, 32'sd19, 32'sd4, 32'sd9, 32'sd19, 32'sd6, 32'sd5, 32'sd18, 32'sd12, 32'sd1, 32'sd1, 32'sd2, 32'sd9, 32'sd2, 32'sd2, 32'sd6, 32'sd8, 32'sd1, 32'sd6, 32'sd5, 32'sd5, 32'sd2, 32'sd5, 32'sd4, 32'sd7, 32'sd3, 32'sd3, 32'sd2, 32'sd1, 32'sd2, 32'sd1, 32'sd2, 32'sd1, 32'sd2, 32'sd2, 32'sd3, 32'sd2, 32'sd4, 32'sd3, 32'sd6, 32'sd7, 32'sd4, 32'sd3, 32'sd2, 32'sd3, 32'sd2, 32'sd3, 32'sd5, 32'sd5, 32'sd17, 32'sd10, 32'sd4, 32'sd9, 32'sd9, 32'sd8, 32'sd2, 32'sd2, 32'sd6, 32'sd5, 32'sd6, 32'sd8, 32'sd4, 32'sd4, 32'sd2, 32'sd2, 32'sd3, 32'sd2, 32'sd2, 32'sd9, 32'sd2, 32'sd7, 32'sd3, 32'sd1, 32'sd2, 32'sd5, 32'sd1, 32'sd6, 32'sd3, 32'sd9, 32'sd3, 32'sd7, 32'sd1, 32'sd1, 32'sd13, 32'sd4, 32'sd3, 32'sd3, 32'sd10, 32'sd10, 32'sd3, 32'sd3, 32'sd21, 32'sd13, 32'sd21, 32'sd20, 32'sd2, 32'sd9, 32'sd3, 32'sd3, 32'sd9, 32'sd10, 32'sd9, 32'sd9, 32'sd2, 32'sd7, 32'sd3, 32'sd6, 32'sd10, 32'sd4, 32'sd2, 32'sd3, 32'sd7, 32'sd2, 32'sd3, 32'sd10, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd1, 32'sd1, 32'sd1, 32'sd1, 32'sd11, 32'sd6, 32'sd11, 32'sd11, 32'sd3, 32'sd2, 32'sd12, 32'sd1, 32'sd9, 32'sd1, 32'sd3, 32'sd1, 32'sd9, 32'sd9, 32'sd18, 32'sd18, 32'sd3, 32'sd2, 32'sd1, 32'sd3, 32'sd1, 32'sd8, 32'sd2, 32'sd4, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd5, 32'sd8, 32'sd15, 32'sd8, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd1, 32'sd11, 32'sd15, 32'sd13, 32'sd9, 32'sd9, 32'sd4, 32'sd4, 32'sd4, 32'sd3, 32'sd1, 32'sd10, 32'sd2, 32'sd4, 32'sd7, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd3, 32'sd9, 32'sd8, 32'sd8, 32'sd9, 32'sd16, 32'sd4, 32'sd4, 32'sd2, 32'sd11, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd5, 32'sd16, 32'sd2, 32'sd5, 32'sd2, 32'sd2, 32'sd2, 32'sd5, 32'sd3, 32'sd2, 32'sd16, 32'sd13, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd11, 32'sd5, 32'sd5, 32'sd7, 32'sd3, 32'sd6, 32'sd8, 32'sd3, 32'sd6, 32'sd9, 32'sd8, 32'sd1, 32'sd3, 32'sd2, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd1, 32'sd2, 32'sd6, 32'sd6, 32'sd11, 32'sd11, 32'sd11, 32'sd11, 32'sd9, 32'sd1, 32'sd1, 32'sd1, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd10, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd2, 32'sd1, 32'sd2, 32'sd2, 32'sd1, 32'sd2, 32'sd5, 32'sd6, 32'sd5, 32'sd12, 32'sd5, 32'sd9, 32'sd9, 32'sd4, 32'sd5, 32'sd5, 32'sd7, 32'sd19, 32'sd3, 32'sd3, 32'sd5, 32'sd4, 32'sd3, 32'sd9, 32'sd6, 32'sd4, 32'sd1, 32'sd1, 32'sd3, 32'sd2, 32'sd4, 32'sd3, 32'sd4, 32'sd7, 32'sd3, 32'sd4, 32'sd3, 32'sd9, 32'sd23, 32'sd2, 32'sd1, 32'sd7, 32'sd6, 32'sd6, 32'sd7, 32'sd9, 32'sd6, 32'sd6, 32'sd5, 32'sd5, 32'sd3, 32'sd5, 32'sd4, 32'sd2, 32'sd19, 32'sd19, 32'sd20, 32'sd20, 32'sd12, 32'sd12, 32'sd7, 32'sd4, 32'sd4, 32'sd5, 32'sd1, 32'sd6, 32'sd1, 32'sd1, 32'sd3, 32'sd2, 32'sd2, 32'sd7, 32'sd3, 32'sd9, 32'sd6, 32'sd5, 32'sd6, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd3, 32'sd1, 32'sd6, 32'sd24, 32'sd4, 32'sd6, 32'sd4, 32'sd7, 32'sd7, 32'sd5, 32'sd2, 32'sd9, 32'sd7, 32'sd5, 32'sd3, 32'sd12, 32'sd14, 32'sd4, 32'sd4, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd4, 32'sd4, 32'sd12, 32'sd11, 32'sd4, 32'sd7, 32'sd1, 
                                                    32'sd9, 32'sd7, 32'sd6, 32'sd11, 32'sd11, 32'sd18, 32'sd5, 32'sd1, 32'sd20, 32'sd4, 32'sd2, 32'sd5, 32'sd7, 32'sd4, 32'sd3, 32'sd4, 32'sd3, 32'sd2, 32'sd9, 32'sd8, 32'sd17, 32'sd6, 32'sd17, 32'sd17, 32'sd1, 32'sd9, 32'sd9, 32'sd9, 32'sd4, 32'sd9, 32'sd9, 32'sd4, 32'sd3, 32'sd9, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd1, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd3, 32'sd3, 32'sd23, 32'sd3, 32'sd4, 32'sd23, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd2, 32'sd5, 32'sd6, 32'sd9, 32'sd9, 32'sd9, 32'sd1, 32'sd3, 32'sd13, 32'sd4, 32'sd13, 32'sd18, 32'sd5, 32'sd8, 32'sd9, 32'sd9, 32'sd7, 32'sd7, 32'sd8, 32'sd10, 32'sd3, 32'sd4, 32'sd5, 32'sd5, 32'sd16, 32'sd16, 32'sd5, 32'sd1, 32'sd2, 32'sd4, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd5, 32'sd4, 32'sd3, 32'sd9, 32'sd7, 32'sd7, 32'sd6, 32'sd8, 32'sd7, 32'sd7, 32'sd9, 32'sd4, 32'sd4, 32'sd4, 32'sd10, 32'sd6, 32'sd10, 32'sd10, 32'sd7, 32'sd7, 32'sd4, 32'sd3, 32'sd5, 32'sd11, 32'sd8, 32'sd3, 32'sd3, 32'sd6, 32'sd3, 32'sd5, 32'sd1, 32'sd1, 32'sd1, 32'sd3, 32'sd3, 32'sd3, 32'sd9, 32'sd2, 32'sd6, 32'sd6, 32'sd4, 32'sd16, 32'sd9, 32'sd9, 32'sd5, 32'sd2, 32'sd4, 32'sd7, 32'sd3, 32'sd3, 32'sd5, 32'sd1, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd6, 32'sd5, 32'sd2, 32'sd4, 32'sd5, 32'sd5, 32'sd6, 32'sd4, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd9, 32'sd5, 32'sd13, 32'sd6, 32'sd3, 32'sd2, 32'sd5, 32'sd3, 32'sd9, 32'sd7, 32'sd3, 32'sd3, 32'sd2, 32'sd6, 32'sd9, 32'sd7, 32'sd3, 32'sd9, 32'sd1, 32'sd2, 32'sd3, 32'sd3, 32'sd5, 32'sd1, 32'sd6, 32'sd9, 32'sd11, 32'sd11, 32'sd5, 32'sd18, 32'sd6, 32'sd1, 32'sd2, 32'sd5, 32'sd9, 32'sd9, 32'sd5, 32'sd1, 32'sd2, 32'sd1, 32'sd2, 32'sd3, 32'sd4, 32'sd1, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd5, 32'sd4, 32'sd6, 32'sd5, 32'sd3, 32'sd4, 32'sd6, 32'sd2, 32'sd5, 32'sd4, 32'sd4, 32'sd4, 32'sd3, 32'sd4, 32'sd8, 32'sd3, 32'sd1, 32'sd9, 32'sd9, 32'sd13, 32'sd1, 32'sd6, 32'sd24, 32'sd24, 32'sd10, 32'sd6, 32'sd3, 32'sd11, 32'sd4, 32'sd18, 32'sd16, 32'sd16, 32'sd3, 32'sd1, 32'sd3, 32'sd3, 32'sd2, 32'sd4, 32'sd7, 32'sd7, 32'sd6, 32'sd4, 32'sd3, 32'sd3, 32'sd7, 32'sd5, 32'sd6, 32'sd18, 32'sd9, 32'sd3, 32'sd5, 32'sd6, 32'sd6, 32'sd5, 32'sd1, 32'sd13, 32'sd1, 32'sd4, 32'sd5, 32'sd2, 32'sd1, 32'sd4, 32'sd3, 32'sd3, 32'sd4, 32'sd6, 32'sd5, 32'sd7, 32'sd10, 32'sd10, 32'sd3, 32'sd3, 32'sd2, 32'sd8, 32'sd11, 32'sd6, 32'sd9, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd9, 32'sd9, 32'sd1, 32'sd13, 32'sd4, 32'sd6, 32'sd1, 32'sd4, 32'sd9, 32'sd13, 32'sd1, 32'sd9, 32'sd9, 32'sd4, 32'sd4, 32'sd4, 32'sd2, 32'sd5, 32'sd6, 32'sd3, 32'sd2, 32'sd1, 32'sd2, 32'sd2, 32'sd3, 32'sd4, 32'sd2, 32'sd1, 32'sd3, 32'sd5, 32'sd3, 32'sd3, 32'sd5, 32'sd5, 32'sd4, 32'sd6, 32'sd1, 32'sd5, 32'sd12, 32'sd12, 32'sd3, 32'sd11, 32'sd13, 32'sd3, 32'sd6, 32'sd3, 32'sd6, 32'sd1, 32'sd10, 32'sd9, 32'sd9, 32'sd9, 32'sd2, 32'sd9, 32'sd9, 32'sd16, 32'sd16, 32'sd3, 32'sd3, 32'sd6, 32'sd6, 32'sd8, 32'sd6, 32'sd2, 32'sd20, 32'sd3, 32'sd9, 32'sd3, 32'sd2, 32'sd6, 32'sd9, 32'sd2, 32'sd3, 32'sd4, 32'sd8, 32'sd3, 32'sd5, 32'sd4, 32'sd4, 32'sd3, 32'sd5, 32'sd21, 32'sd21, 32'sd1, 32'sd2, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd1, 32'sd1, 32'sd23, 32'sd3, 32'sd1, 32'sd23, 32'sd5, 32'sd4, 32'sd7, 32'sd3, 32'sd6, 32'sd5, 32'sd2, 32'sd5, 32'sd4, 32'sd24, 32'sd2, 32'sd5, 32'sd9, 32'sd1, 32'sd9, 32'sd9, 32'sd9, 32'sd11, 32'sd2, 32'sd4, 32'sd3, 32'sd5, 32'sd12, 32'sd12, 32'sd4, 32'sd10, 32'sd3, 32'sd9, 32'sd5, 32'sd11, 32'sd2, 32'sd4, 32'sd2, 32'sd2, 32'sd4, 32'sd9, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd1, 32'sd3, 32'sd3, 32'sd1, 32'sd2, 32'sd2, 32'sd2, 32'sd12, 32'sd9, 32'sd6, 32'sd2, 32'sd3, 32'sd3, 32'sd4, 32'sd3, 32'sd7, 32'sd6, 32'sd6, 32'sd6, 32'sd14, 32'sd18, 32'sd12, 32'sd14, 32'sd14, 32'sd20, 32'sd20, 32'sd17, 32'sd17, 32'sd2, 32'sd2, 32'sd13, 32'sd13, 32'sd9, 32'sd7, 32'sd2, 32'sd2, 32'sd3, 32'sd1, 32'sd5, 32'sd3, 32'sd6, 32'sd9, 32'sd2, 32'sd4, 32'sd5, 32'sd3, 32'sd5, 32'sd18, 32'sd14, 32'sd9, 32'sd3, 32'sd2, 32'sd4, 32'sd4, 32'sd1, 32'sd5, 32'sd6, 32'sd12, 32'sd1, 32'sd6, 32'sd3, 32'sd9, 32'sd5, 32'sd6, 32'sd6, 32'sd11, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd3, 32'sd13, 32'sd9, 32'sd9, 32'sd3, 32'sd1, 32'sd3, 32'sd3, 32'sd21, 32'sd4, 32'sd2, 32'sd1, 32'sd1, 32'sd2, 32'sd4, 32'sd6, 32'sd7, 32'sd2, 32'sd3, 32'sd2, 32'sd3, 32'sd3, 32'sd2, 32'sd4, 32'sd7, 32'sd7, 32'sd5, 32'sd5, 32'sd10, 32'sd2, 32'sd6, 32'sd3, 32'sd3, 32'sd5, 32'sd2, 32'sd4, 32'sd9, 32'sd6, 32'sd2, 32'sd3, 32'sd1, 32'sd1, 32'sd9, 32'sd9, 32'sd20, 32'sd20, 32'sd7, 32'sd9, 32'sd2, 32'sd2, 32'sd2, 32'sd6, 32'sd3, 32'sd2, 32'sd3, 32'sd7, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd6, 32'sd3, 32'sd11, 32'sd6, 32'sd1, 32'sd4, 32'sd2, 32'sd2, 32'sd6, 32'sd4, 32'sd8, 32'sd1, 32'sd3, 32'sd8, 32'sd4, 32'sd1, 32'sd7, 32'sd5, 32'sd3, 32'sd6, 32'sd9, 32'sd4, 32'sd4, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd8, 32'sd3, 32'sd2, 32'sd2, 32'sd1, 32'sd5, 32'sd2, 32'sd3, 32'sd3, 32'sd4, 32'sd2, 32'sd14, 32'sd8, 32'sd4, 32'sd9, 32'sd10, 32'sd13, 32'sd13, 32'sd6, 32'sd3, 32'sd7, 32'sd2, 32'sd6, 32'sd4, 32'sd3, 32'sd5, 32'sd5, 32'sd13, 32'sd19, 32'sd6, 32'sd2, 32'sd2, 32'sd5, 32'sd7, 32'sd3, 32'sd12, 32'sd7, 32'sd4, 32'sd6, 32'sd3, 32'sd5, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd4, 32'sd7, 32'sd3, 32'sd9, 32'sd12, 32'sd9, 32'sd9, 32'sd11, 32'sd6, 32'sd3, 32'sd2, 32'sd11, 32'sd11, 32'sd2, 32'sd7, 32'sd4, 32'sd5, 32'sd6, 32'sd6, 32'sd16, 32'sd16, 32'sd16, 32'sd16, 32'sd1, 32'sd2, 32'sd4, 32'sd1, 32'sd1, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd7, 32'sd1, 32'sd7, 32'sd5, 32'sd5, 32'sd9, 32'sd5, 32'sd9, 32'sd9, 32'sd10, 32'sd3, 32'sd10, 32'sd4, 32'sd10, 32'sd19, 32'sd10, 32'sd9, 32'sd2, 32'sd2, 32'sd3, 32'sd4, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd8, 32'sd9, 32'sd9, 32'sd9, 32'sd10, 32'sd10, 32'sd3, 32'sd9, 32'sd6, 32'sd4, 
                                                    32'sd6, 32'sd7, 32'sd2, 32'sd5, 32'sd1, 32'sd10, 32'sd6, 32'sd9, 32'sd8, 32'sd6, 32'sd7, 32'sd2, 32'sd3, 32'sd3, 32'sd10, 32'sd1, 32'sd4, 32'sd11, 32'sd4, 32'sd4, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd1, 32'sd1, 32'sd3, 32'sd5, 32'sd5, 32'sd9, 32'sd1, 32'sd1, 32'sd3, 32'sd3, 32'sd3, 32'sd5, 32'sd8, 32'sd5, 32'sd13, 32'sd13, 32'sd9, 32'sd11, 32'sd11, 32'sd2, 32'sd1, 32'sd9, 32'sd7, 32'sd9, 32'sd6, 32'sd9, 32'sd10, 32'sd3, 32'sd3, 32'sd3, 32'sd9, 32'sd15, 32'sd1, 32'sd9, 32'sd1, 32'sd2, 32'sd5, 32'sd14, 32'sd9, 32'sd1, 32'sd6, 32'sd1, 32'sd4, 32'sd5, 32'sd6, 32'sd5, 32'sd5, 32'sd3, 32'sd3, 32'sd20, 32'sd3, 32'sd13, 32'sd5, 32'sd4, 32'sd7, 32'sd2, 32'sd1, 32'sd4, 32'sd9, 32'sd1, 32'sd13, 32'sd5, 32'sd3, 32'sd1, 32'sd1, 32'sd11, 32'sd5, 32'sd1, 32'sd1, 32'sd5, 32'sd21, 32'sd3, 32'sd3, 32'sd4, 32'sd4, 32'sd3, 32'sd3, 32'sd9, 32'sd1, 32'sd9, 32'sd2, 32'sd3, 32'sd5, 32'sd2, 32'sd9, 32'sd5, 32'sd5, 32'sd5, 32'sd7, 32'sd5, 32'sd7, 32'sd5, 32'sd6, 32'sd6, 32'sd2, 32'sd10, 32'sd2, 32'sd2, 32'sd1, 32'sd13, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd2, 32'sd16, 32'sd16, 32'sd10, 32'sd10, 32'sd24, 32'sd10, 32'sd9, 32'sd9, 32'sd5, 32'sd9, 32'sd8, 32'sd8, 32'sd9, 32'sd6, 32'sd18, 32'sd18, 32'sd2, 32'sd3, 32'sd15, 32'sd14, 32'sd5, 32'sd9, 32'sd8, 32'sd8, 32'sd4, 32'sd2, 32'sd5, 32'sd5, 32'sd3, 32'sd5, 32'sd2, 32'sd2, 32'sd4, 32'sd2, 32'sd2, 32'sd23, 32'sd2, 32'sd4, 32'sd9, 32'sd6, 32'sd4, 32'sd2, 32'sd2, 32'sd1, 32'sd10, 32'sd10, 32'sd9, 32'sd12, 32'sd4, 32'sd7, 32'sd8, 32'sd9, 32'sd2, 32'sd2, 32'sd3, 32'sd6, 32'sd9, 32'sd7, 32'sd2, 32'sd10, 32'sd21, 32'sd10, 32'sd4, 32'sd9, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd9, 32'sd9, 32'sd4, 32'sd4, 32'sd2, 32'sd2, 32'sd2, 32'sd4, 32'sd19, 32'sd8, 32'sd4, 32'sd3, 32'sd2, 32'sd10, 32'sd6, 32'sd22, 32'sd22, 32'sd1, 32'sd5, 32'sd9, 32'sd1, 32'sd5, 32'sd1, 32'sd6, 32'sd7, 32'sd5, 32'sd9, 32'sd5, 32'sd5, 32'sd2, 32'sd1, 32'sd6, 32'sd8, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd4, 32'sd8, 32'sd4, 32'sd3, 32'sd3, 32'sd9, 32'sd9, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd1, 32'sd1, 32'sd11, 32'sd11, 32'sd24, 32'sd4, 32'sd9, 32'sd7, 32'sd3, 32'sd3, 32'sd10, 32'sd3, 32'sd7, 32'sd6, 32'sd24, 32'sd24, 32'sd7, 32'sd7, 32'sd19, 32'sd6, 32'sd6, 32'sd4, 32'sd5, 32'sd5, 32'sd10, 32'sd10, 32'sd4, 32'sd4, 32'sd3, 32'sd1, 32'sd10, 32'sd9, 32'sd19, 32'sd3, 32'sd10, 32'sd9, 32'sd5, 32'sd6, 32'sd10, 32'sd10, 32'sd6, 32'sd6, 32'sd4, 32'sd3, 32'sd2, 32'sd5, 32'sd2, 32'sd5, 32'sd6, 32'sd2, 32'sd2, 32'sd9, 32'sd9, 32'sd2, 32'sd1, 32'sd2, 32'sd19, 32'sd19, 32'sd1, 32'sd2, 32'sd9, 32'sd4, 32'sd2, 32'sd10, 32'sd6, 32'sd6, 32'sd5, 32'sd5, 32'sd2, 32'sd1, 32'sd9, 32'sd9, 32'sd9, 32'sd9, 32'sd5, 32'sd10, 32'sd3, 32'sd1, 32'sd6, 32'sd2, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd11, 32'sd11, 32'sd3, 32'sd9, 32'sd6, 32'sd3, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd4, 32'sd7, 32'sd4, 32'sd9, 32'sd6, 32'sd10, 32'sd6, 32'sd7, 32'sd6, 32'sd18, 32'sd7, 32'sd1, 32'sd4, 32'sd7, 32'sd6, 32'sd6, 32'sd11, 32'sd20, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd12, 32'sd4, 32'sd2, 32'sd3, 32'sd1, 32'sd8, 32'sd12, 32'sd1, 32'sd7, 32'sd2, 32'sd7, 32'sd19, 32'sd7, 32'sd3, 32'sd7, 32'sd3, 32'sd5, 32'sd19, 32'sd6, 32'sd7, 32'sd9, 32'sd5, 32'sd5, 32'sd5, 32'sd7, 32'sd5, 32'sd9, 32'sd9, 32'sd7, 32'sd7, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd8, 32'sd1, 32'sd2, 32'sd2, 32'sd5, 32'sd6, 32'sd3, 32'sd10, 32'sd3, 32'sd5, 32'sd14, 32'sd2, 32'sd3, 32'sd7, 32'sd6, 32'sd6, 32'sd3, 32'sd2, 32'sd2, 32'sd6, 32'sd3, 32'sd6, 32'sd6, 32'sd1, 32'sd3, 32'sd2, 32'sd2, 32'sd2, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd9, 32'sd12, 32'sd4, 32'sd3, 32'sd12, 32'sd3, 32'sd9, 32'sd3, 32'sd3, 32'sd10, 32'sd10, 32'sd9, 32'sd4, 32'sd3, 32'sd9, 32'sd9, 32'sd3, 32'sd10, 32'sd10, 32'sd2, 32'sd2, 32'sd3, 32'sd2, 32'sd1, 32'sd7, 32'sd6, 32'sd6, 32'sd3, 32'sd13, 32'sd3, 32'sd15, 32'sd7, 32'sd3, 32'sd6, 32'sd9, 32'sd24, 32'sd24, 32'sd4, 32'sd2, 32'sd2, 32'sd4, 32'sd2, 32'sd7, 32'sd1, 32'sd1, 32'sd9, 32'sd6, 32'sd6, 32'sd9, 32'sd10, 32'sd9, 32'sd7, 32'sd5, 32'sd8, 32'sd9, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd2, 32'sd3, 32'sd7, 32'sd8, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd9, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd7, 32'sd1, 32'sd1, 32'sd10, 32'sd24, 32'sd15, 32'sd24, 32'sd9, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd10, 32'sd23, 32'sd9, 32'sd2, 32'sd3, 32'sd5, 32'sd19, 32'sd18, 32'sd18, 32'sd3, 32'sd9, 32'sd7, 32'sd7, 32'sd6, 32'sd5, 32'sd5, 32'sd8, 32'sd2, 32'sd2, 32'sd3, 32'sd4, 32'sd6, 32'sd9, 32'sd3, 32'sd22, 32'sd3, 32'sd1, 32'sd24, 32'sd6, 32'sd7, 32'sd5, 32'sd5, 32'sd6, 32'sd7, 32'sd7, 32'sd2, 32'sd6, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd5, 32'sd8, 32'sd8, 32'sd2, 32'sd18, 32'sd19, 32'sd16, 32'sd16, 32'sd2, 32'sd5, 32'sd5, 32'sd6, 32'sd5, 32'sd7, 32'sd6, 32'sd3, 32'sd6, 32'sd10, 32'sd6, 32'sd4, 32'sd2, 32'sd4, 32'sd5, 32'sd9, 32'sd22, 32'sd22, 32'sd2, 32'sd5, 32'sd6, 32'sd13, 32'sd24, 32'sd24, 32'sd4, 32'sd1, 32'sd1, 32'sd2, 32'sd5, 32'sd1, 32'sd2, 32'sd8, 32'sd4, 32'sd16, 32'sd16, 32'sd16, 32'sd14, 32'sd14, 32'sd22, 32'sd22, 32'sd20, 32'sd20, 32'sd9, 32'sd16, 32'sd6, 32'sd3, 32'sd4, 32'sd2, 32'sd2, 32'sd6, 32'sd4, 32'sd6, 32'sd3, 32'sd6, 32'sd5, 32'sd4, 32'sd2, 32'sd3, 32'sd3, 32'sd9, 32'sd3, 32'sd1, 32'sd3, 32'sd9, 32'sd9, 32'sd5, 32'sd5, 32'sd3, 32'sd7, 32'sd5, 32'sd3, 32'sd1, 32'sd10, 32'sd1, 32'sd11, 32'sd4, 32'sd3, 32'sd1, 32'sd2, 32'sd1, 32'sd18, 32'sd10, 32'sd10, 32'sd9, 32'sd9, 32'sd1, 32'sd2, 32'sd7, 32'sd7, 32'sd6, 32'sd6, 32'sd6, 32'sd1, 32'sd1, 32'sd5, 32'sd2, 32'sd3, 32'sd3, 32'sd6, 32'sd2, 32'sd13, 32'sd3, 32'sd3, 32'sd1, 32'sd2, 32'sd1, 32'sd2, 32'sd19, 32'sd8, 32'sd9, 32'sd9, 32'sd1, 32'sd2, 32'sd3, 32'sd2, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd1, 32'sd1, 32'sd6, 32'sd3, 32'sd5, 32'sd2, 32'sd12, 32'sd15, 32'sd19, 32'sd19, 
                                                    32'sd5, 32'sd5, 32'sd6, 32'sd3, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd6, 32'sd1, 32'sd6, 32'sd6, 32'sd1, 32'sd1, 32'sd1, 32'sd10, 32'sd17, 32'sd17, 32'sd11, 32'sd3, 32'sd4, 32'sd7, 32'sd7, 32'sd7, 32'sd1, 32'sd2, 32'sd2, 32'sd2, 32'sd18, 32'sd18, 32'sd10, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd1, 32'sd9, 32'sd6, 32'sd9, 32'sd9, 32'sd3, 32'sd3, 32'sd1, 32'sd2, 32'sd5, 32'sd3, 32'sd3, 32'sd3, 32'sd2, 32'sd2, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd3, 32'sd5, 32'sd1, 32'sd5, 32'sd3, 32'sd3, 32'sd9, 32'sd6, 32'sd9, 32'sd9, 32'sd6, 32'sd12, 32'sd11, 32'sd2, 32'sd3, 32'sd9, 32'sd9, 32'sd9, 32'sd12, 32'sd2, 32'sd1, 32'sd4, 32'sd5, 32'sd7, 32'sd7, 32'sd7, 32'sd2, 32'sd10, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd5, 32'sd5, 32'sd4, 32'sd4, 32'sd3, 32'sd7, 32'sd2, 32'sd3, 32'sd5, 32'sd5, 32'sd4, 32'sd3, 32'sd4, 32'sd3, 32'sd6, 32'sd6, 32'sd2, 32'sd5, 32'sd2, 32'sd1, 32'sd1, 32'sd1, 32'sd2, 32'sd2, 32'sd2, 32'sd2, 32'sd20, 32'sd4, 32'sd11}

localparam logic [2912:0][31:0] rectangle2_weights = {32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 
                                                    32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 
                                                    32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 
                                                    32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 
                                                    32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 
                                                    32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd256, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd384, 32'sd256, 32'sd256}

localparam logic [2912:0][31:0] rectangle3_xs = {32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd12, 32'sd9, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd1, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd12, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd4, 32'sd10, 32'sd10, 32'sd3, 32'sd0, 32'sd0, 32'sd15, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd17, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd8, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd5, 32'sd0, 32'sd0, 32'sd5, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd16, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd10, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd12, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd6, 32'sd14, 32'sd6, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd20, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd7, 
                                                    32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd4, 32'sd12, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd11, 32'sd10, 32'sd0, 32'sd0, 32'sd8, 32'sd12, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd1, 32'sd0, 32'sd9, 32'sd10, 32'sd4, 32'sd0, 32'sd16, 32'sd0, 32'sd8, 32'sd0, 32'sd10, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd10, 32'sd10, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd16, 32'sd0, 32'sd16, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd8, 32'sd4, 32'sd0, 32'sd0, 32'sd17, 32'sd4, 32'sd7, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd4, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd1, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd8, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd12, 32'sd12, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd11, 32'sd5, 32'sd12, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd9, 32'sd11, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd9, 32'sd6, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd9, 32'sd0, 32'sd9, 32'sd0, 32'sd10, 32'sd0, 32'sd9, 32'sd11, 32'sd11, 32'sd0, 32'sd6, 32'sd10, 32'sd16, 32'sd11, 32'sd8, 32'sd10, 32'sd3, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd4, 32'sd0, 32'sd0, 32'sd14, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd10, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd15, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd14, 32'sd0, 
                                                    32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd4, 32'sd14, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd12, 32'sd14, 32'sd5, 32'sd0, 32'sd11, 32'sd7, 32'sd11, 32'sd10, 32'sd11, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd10, 32'sd10, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd15, 32'sd5, 32'sd11, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd12, 32'sd0, 32'sd7, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd2, 32'sd7, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd4, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd12, 32'sd6, 32'sd1, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd6, 32'sd0, 32'sd9, 32'sd0, 32'sd5, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd6, 32'sd0, 32'sd14, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd7, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd3, 32'sd11, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd12, 32'sd0, 32'sd12, 32'sd15, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd5, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd5, 32'sd0, 32'sd11, 32'sd7, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd12, 32'sd13, 32'sd9, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd11, 32'sd6, 32'sd11, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd11, 32'sd11, 32'sd5, 32'sd0, 32'sd0, 32'sd9, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd12, 32'sd7, 32'sd12, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd14, 32'sd6, 32'sd10, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd0, 32'sd19, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd9, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd11, 32'sd1, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd12, 32'sd9, 32'sd16, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd13, 32'sd12, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd14, 32'sd7, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd3, 32'sd0, 32'sd0, 32'sd11, 32'sd12, 32'sd0, 32'sd0, 32'sd20, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd20, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd9, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd15, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd12, 32'sd9, 32'sd5, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd1, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd11, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd3, 32'sd10, 32'sd12, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd4, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd3, 32'sd13, 32'sd0, 32'sd12, 32'sd9, 32'sd0, 32'sd6, 32'sd14, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd15, 32'sd5, 32'sd11, 32'sd9, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd10, 32'sd11, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd8, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd4, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd5, 32'sd0, 32'sd0, 32'sd7, 32'sd10, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd7, 32'sd0, 32'sd0, 32'sd10, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd19, 32'sd3, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd12, 32'sd7, 32'sd14, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd7, 32'sd0, 32'sd11, 32'sd10, 32'sd12, 32'sd6, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 
                                                    32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd15, 32'sd6, 32'sd3, 32'sd7, 32'sd16, 32'sd4, 32'sd13, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd18, 32'sd3, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9}

localparam logic [2912:0][31:0] rectangle3_ys = {32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd20, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd11, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd20, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd9, 32'sd11, 32'sd14, 32'sd14, 32'sd0, 32'sd0, 32'sd18, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd0, 32'sd13, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd8, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd3, 32'sd0, 32'sd18, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd0, 32'sd17, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd15, 32'sd0, 32'sd0, 32'sd19, 32'sd14, 32'sd0, 32'sd20, 32'sd20, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd8, 32'sd19, 32'sd19, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd9, 32'sd9, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd15, 32'sd11, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd15, 32'sd15, 32'sd0, 32'sd0, 32'sd7, 32'sd9, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd19, 32'sd0, 32'sd10, 32'sd10, 32'sd9, 32'sd0, 32'sd17, 32'sd0, 32'sd16, 32'sd0, 32'sd12, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd12, 32'sd12, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd16, 32'sd0, 32'sd16, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd7, 32'sd6, 32'sd0, 32'sd0, 32'sd17, 32'sd17, 32'sd13, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd14, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd20, 32'sd20, 32'sd2, 32'sd0, 32'sd7, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd11, 32'sd12, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd9, 32'sd9, 32'sd19, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd21, 32'sd22, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd11, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd13, 32'sd0, 32'sd13, 32'sd0, 32'sd15, 32'sd0, 32'sd13, 32'sd13, 32'sd17, 32'sd0, 32'sd15, 32'sd12, 32'sd19, 32'sd13, 32'sd21, 32'sd15, 32'sd12, 32'sd20, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd14, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd14, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd17, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd12, 32'sd7, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd8, 32'sd0, 32'sd20, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd16, 32'sd20, 32'sd20, 32'sd0, 32'sd20, 32'sd9, 32'sd15, 32'sd16, 32'sd16, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd10, 32'sd9, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd14, 32'sd14, 32'sd15, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd5, 32'sd0, 32'sd8, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd18, 32'sd0, 32'sd0, 32'sd18, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd12, 32'sd15, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd6, 32'sd0, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd9, 32'sd9, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd9, 32'sd0, 32'sd19, 32'sd0, 32'sd9, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd9, 32'sd0, 32'sd16, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd9, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd16, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd13, 32'sd13, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd21, 32'sd0, 32'sd12, 32'sd15, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd11, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd0, 32'sd17, 32'sd0, 32'sd12, 32'sd12, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd14, 32'sd12, 32'sd12, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd11, 32'sd20, 32'sd11, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd11, 32'sd11, 32'sd12, 32'sd0, 32'sd0, 32'sd4, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd15, 32'sd16, 
                                                    32'sd7, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd19, 32'sd19, 32'sd21, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd13, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd14, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd20, 32'sd0, 32'sd16, 32'sd16, 32'sd18, 32'sd18, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd14, 32'sd16, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd15, 32'sd15, 32'sd0, 32'sd22, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd13, 32'sd0, 32'sd0, 32'sd15, 32'sd16, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd20, 32'sd0, 32'sd0, 32'sd14, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd12, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd12, 32'sd12, 32'sd13, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd15, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd7, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd9, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd12, 32'sd0, 32'sd12, 32'sd12, 32'sd0, 32'sd12, 32'sd14, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd19, 32'sd19, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd13, 32'sd13, 32'sd0, 32'sd16, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd13, 32'sd13, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd9, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd11, 32'sd0, 32'sd0, 32'sd15, 32'sd15, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13, 32'sd12, 32'sd0, 32'sd0, 32'sd11, 32'sd16, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd15, 32'sd15, 32'sd0, 32'sd0, 32'sd21, 32'sd0, 32'sd20, 32'sd20, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19, 32'sd19, 32'sd0, 32'sd14, 32'sd10, 32'sd9, 32'sd13, 32'sd13, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd17, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd22, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd15, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd8, 32'sd8, 32'sd22, 32'sd10, 32'sd14, 32'sd14, 32'sd17, 32'sd17, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd18, 32'sd21, 32'sd0, 32'sd0, 32'sd18, 32'sd18, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12}

localparam logic [2912:0][31:0] rectangle3_widths = {32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd7, 32'sd5, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd3, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd8, 32'sd9, 32'sd4, 32'sd3, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd12, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd12, 32'sd0, 32'sd8, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd2, 32'sd0, 32'sd0, 32'sd4, 32'sd12, 32'sd0, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd6, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd4, 32'sd6, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd3, 32'sd8, 32'sd0, 32'sd0, 32'sd4, 32'sd6, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd11, 32'sd0, 32'sd5, 32'sd5, 32'sd8, 32'sd0, 32'sd4, 32'sd0, 32'sd4, 32'sd0, 32'sd4, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd4, 32'sd4, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd4, 32'sd0, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd4, 32'sd3, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd7, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd10, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd12, 32'sd0, 32'sd12, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd6, 32'sd6, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd6, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd7, 32'sd10, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd3, 32'sd9, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd4, 32'sd0, 32'sd4, 32'sd0, 32'sd2, 32'sd0, 32'sd4, 32'sd4, 32'sd3, 32'sd0, 32'sd6, 32'sd9, 32'sd4, 32'sd11, 32'sd6, 32'sd10, 32'sd10, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd3, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd3, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd3, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd4, 32'sd5, 32'sd5, 32'sd0, 32'sd5, 32'sd6, 32'sd2, 32'sd3, 32'sd3, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd4, 32'sd8, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd12, 32'sd0, 32'sd6, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd11, 32'sd4, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd3, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd7, 32'sd0, 32'sd6, 32'sd0, 32'sd7, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd7, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd3, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd10, 32'sd10, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd10, 32'sd0, 32'sd9, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd8, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd4, 32'sd0, 32'sd5, 32'sd7, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd9, 32'sd2, 32'sd2, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd2, 32'sd5, 32'sd2, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd2, 32'sd9, 32'sd0, 32'sd0, 32'sd9, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd2, 32'sd5, 32'sd4, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd4, 32'sd4, 32'sd6, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd3, 32'sd3, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd4, 32'sd5, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd3, 32'sd3, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd2, 32'sd5, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd8, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd7, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd9, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd3, 32'sd3, 32'sd5, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd9, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd2, 32'sd0, 32'sd6, 32'sd2, 32'sd0, 32'sd6, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd4, 32'sd4, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd4, 32'sd8, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd9, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd4, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd5, 32'sd0, 32'sd0, 32'sd6, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd4, 32'sd0, 32'sd6, 32'sd4, 32'sd6, 32'sd9, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd3, 32'sd9, 32'sd2, 32'sd4, 32'sd4, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd11, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3}

localparam logic [2912:0][31:0] rectangle3_heights = {32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd5, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd6, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd3, 32'sd11, 32'sd7, 32'sd10, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd8, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd2, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd9, 32'sd0, 32'sd0, 32'sd5, 32'sd2, 32'sd0, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd3, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd9, 32'sd6, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd7, 32'sd3, 32'sd0, 32'sd0, 32'sd5, 32'sd3, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd3, 32'sd0, 32'sd5, 32'sd5, 32'sd3, 32'sd0, 32'sd7, 32'sd0, 32'sd6, 32'sd0, 32'sd8, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd8, 32'sd8, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd8, 32'sd0, 32'sd8, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd4, 32'sd2, 32'sd0, 32'sd3, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd3, 32'sd6, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd4, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd2, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd6, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd5, 32'sd0, 32'sd5, 32'sd0, 32'sd9, 32'sd0, 32'sd5, 32'sd5, 32'sd7, 32'sd0, 32'sd3, 32'sd3, 32'sd5, 32'sd4, 32'sd3, 32'sd9, 32'sd6, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd7, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd7, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd4, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd8, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd0, 32'sd4, 32'sd3, 32'sd9, 32'sd7, 32'sd7, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd9, 32'sd4, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd10, 32'sd10, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd3, 32'sd0, 32'sd6, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd7, 32'sd5, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd6, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd9, 32'sd9, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd3, 32'sd0, 32'sd4, 32'sd0, 32'sd3, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd3, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd6, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd3, 32'sd3, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd2, 32'sd0, 32'sd7, 32'sd9, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd7, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd7, 32'sd0, 32'sd12, 32'sd7, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd0, 32'sd0, 32'sd2, 32'sd11, 32'sd11, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd10, 32'sd4, 32'sd10, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd10, 32'sd10, 32'sd3, 32'sd0, 32'sd0, 32'sd4, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd9, 32'sd8, 32'sd6, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd5, 32'sd5, 32'sd3, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd8, 32'sd0, 32'sd0, 32'sd2, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd6, 32'sd6, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd5, 32'sd5, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd6, 32'sd6, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd9, 32'sd7, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd10, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd10, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd11, 32'sd11, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd4, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd2, 32'sd0, 32'sd0, 32'sd12, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd6, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd2, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd10, 32'sd9, 32'sd0, 32'sd3, 32'sd9, 32'sd0, 32'sd3, 32'sd10, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd8, 32'sd4, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd2, 32'sd10, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd5, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd10, 32'sd6, 32'sd0, 32'sd0, 32'sd4, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd8, 32'sd9, 32'sd9, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd4, 32'sd4, 32'sd6, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd5, 32'sd0, 32'sd3, 32'sd5, 32'sd5, 32'sd5, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd9, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd3, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd7, 32'sd7, 32'sd7, 32'sd2, 32'sd10, 32'sd6, 32'sd6, 32'sd4, 32'sd4, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd4, 32'sd3, 32'sd0, 32'sd0, 32'sd6, 32'sd6, 32'sd0, 32'sd5, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd11}

localparam logic [2912:0][31:0] rectangle3_weights = {32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 
                                                    32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd0, 32'sd256, 32'sd256, 32'sd0, 32'sd256, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd256}

localparam logic [2912:0][31:0] feature_threshold = {-32'sd4, 32'sd2, 32'sd3, 32'sd1, 32'sd2, 32'sd13, 32'sd0, -32'sd2, 32'sd1, -32'sd3, 32'sd3, 32'sd3, 32'sd12, 32'sd5, -32'sd2, 32'sd1, 32'sd2, -32'sd1, -32'sd1, 32'sd2, -32'sd3, -32'sd18, 32'sd2, 32'sd1, 32'sd12, 32'sd9, 32'sd4, 32'sd2, 32'sd2, 32'sd0, 32'sd4, -32'sd1, 32'sd6, 32'sd6, -32'sd9, -32'sd6, 32'sd11, 32'sd0, 32'sd15, -32'sd7, -32'sd5, 32'sd48, 32'sd2, 32'sd2, 32'sd5, -32'sd1, 32'sd0, 32'sd4, -32'sd10, 32'sd0, 32'sd3, -32'sd6, -32'sd8, 32'sd2, 32'sd19, 32'sd1, 32'sd1, 32'sd2, 32'sd3, -32'sd36, 32'sd1, -32'sd5, 32'sd2, -32'sd1, 32'sd4, -32'sd5, -32'sd1, -32'sd8, -32'sd5, 32'sd0, -32'sd17, 32'sd3, -32'sd4, 32'sd3, 32'sd3, -32'sd1, 32'sd6, 32'sd7, 32'sd0, 32'sd2, -32'sd3, -32'sd1, -32'sd2, -32'sd9, 32'sd5, 32'sd24, 32'sd10, 32'sd0, 32'sd11, 32'sd1, 32'sd1, -32'sd3, 32'sd1, 32'sd4, 32'sd0, 32'sd4, -32'sd1, -32'sd1, -32'sd3, 32'sd0, -32'sd2, -32'sd1, 32'sd10, 32'sd4, 32'sd3, -32'sd4, -32'sd4, 32'sd3, 32'sd1, -32'sd5, -32'sd2, -32'sd3, -32'sd3, 32'sd2, -32'sd2, -32'sd4, 32'sd2, 32'sd0, 32'sd11, 32'sd33, -32'sd5, -32'sd2, 32'sd0, -32'sd1, 32'sd0, -32'sd6, -32'sd3, -32'sd10, 32'sd3, 32'sd0, 32'sd15, 32'sd0, 32'sd9, -32'sd6, -32'sd6, 32'sd4, 32'sd12, 32'sd2, 32'sd2, 32'sd0, 32'sd4, 32'sd0, -32'sd2, 32'sd3, 32'sd4, -32'sd6, -32'sd9, 32'sd8, 32'sd1, 32'sd5, 32'sd0, -32'sd4, -32'sd2, 32'sd5, 32'sd3, 32'sd7, -32'sd2, -32'sd23, 32'sd23, -32'sd1, 32'sd8, -32'sd4, -32'sd6, 32'sd5, -32'sd3, -32'sd8, -32'sd4, 32'sd1, 32'sd0, 32'sd3, -32'sd1, 32'sd2, -32'sd6, 32'sd3, 32'sd0, 32'sd2, -32'sd4, 32'sd9, 32'sd30, -32'sd2, 32'sd1, 32'sd2, -32'sd1, 32'sd1, 32'sd1, 32'sd2, 32'sd0, -32'sd14, 32'sd1, 32'sd4, 32'sd4, 32'sd1, 32'sd3, 32'sd2, 32'sd3, -32'sd2, -32'sd5, -32'sd1, 32'sd0, -32'sd4, 32'sd8, 32'sd1, 32'sd1, 32'sd0, 32'sd1, 32'sd1, 32'sd4, 32'sd3, 32'sd1, 32'sd4, 32'sd0, -32'sd5, -32'sd5, 32'sd0, -32'sd7, -32'sd1, 32'sd4, -32'sd14, -32'sd1, -32'sd1, -32'sd1, -32'sd2, -32'sd3, 32'sd2, -32'sd3, -32'sd5, -32'sd8, 32'sd3, 32'sd0, 32'sd6, 32'sd7, -32'sd1, -32'sd2, 32'sd3, -32'sd3, 32'sd2, -32'sd1, -32'sd1, 32'sd16, 32'sd6, 32'sd7, -32'sd5, -32'sd9, 32'sd17, -32'sd27, -32'sd8, 32'sd8, -32'sd3, -32'sd4, -32'sd2, 32'sd2, 32'sd6, 32'sd2, 32'sd2, 32'sd6, 32'sd2, -32'sd2, 32'sd5, -32'sd7, -32'sd9, 32'sd2, -32'sd1, -32'sd5, 32'sd0, -32'sd3, 32'sd0, 32'sd0, 32'sd5, 32'sd8, 32'sd0, 32'sd0, -32'sd1, -32'sd3, -32'sd13, -32'sd1, 32'sd5, -32'sd2, -32'sd6, 32'sd3, -32'sd1, 32'sd5, 32'sd0, 32'sd1, 32'sd1, -32'sd7, -32'sd29, -32'sd2, -32'sd2, -32'sd5, -32'sd1, -32'sd2, 32'sd4, 32'sd3, 32'sd1, -32'sd3, -32'sd1, -32'sd5, -32'sd3, 32'sd0, -32'sd3, -32'sd4, -32'sd2, -32'sd8, -32'sd2, -32'sd3, -32'sd4, -32'sd3, 32'sd0, -32'sd4, 32'sd2, 32'sd1, -32'sd1, 32'sd0, -32'sd1, -32'sd6, -32'sd8, -32'sd4, -32'sd19, -32'sd2, 32'sd19, 32'sd7, 32'sd0, -32'sd6, 32'sd17, -32'sd12, 32'sd2, 32'sd4, 32'sd2, 32'sd2, -32'sd4, 32'sd18, -32'sd1, 32'sd2, 32'sd3, 32'sd6, -32'sd1, 32'sd5, -32'sd4, -32'sd5, 32'sd0, 32'sd4, 32'sd4, 32'sd1, 32'sd0, 32'sd5, 32'sd3, -32'sd2, -32'sd1, 32'sd3, 32'sd8, 32'sd5, 32'sd3, -32'sd4, 32'sd1, 32'sd3, -32'sd2, 32'sd6, 32'sd0, -32'sd11, 32'sd2, 32'sd5, -32'sd26, -32'sd2, 32'sd5, 32'sd0, -32'sd2, -32'sd6, -32'sd4, -32'sd6, -32'sd4, -32'sd1, -32'sd1, 32'sd1, 32'sd7, 32'sd4, -32'sd2, -32'sd4, -32'sd10, 32'sd0, 32'sd12, 32'sd5, 32'sd7, -32'sd3, 32'sd42, 32'sd1, 32'sd21, -32'sd1, -32'sd2, 32'sd10, 32'sd2, -32'sd10, -32'sd9, -32'sd1, 32'sd4, -32'sd4, -32'sd10, 32'sd0, 32'sd4, 32'sd1, 32'sd13, -32'sd1, 32'sd1, 32'sd3, 32'sd36, -32'sd6, -32'sd2, 32'sd18, 32'sd4, 32'sd2, 32'sd3, 32'sd7, 32'sd2, 32'sd1, 32'sd4, -32'sd6, 32'sd2, 32'sd1, -32'sd6, 32'sd11, -32'sd1, 32'sd5, -32'sd1, -32'sd1, 32'sd1, 32'sd12, -32'sd4, -32'sd8, -32'sd5, -32'sd1, 32'sd6, -32'sd5, -32'sd3, 32'sd0, -32'sd4, 32'sd2, 32'sd0, 32'sd0, -32'sd12, -32'sd10, 32'sd2, -32'sd3, -32'sd2, 32'sd1, 32'sd13, -32'sd5, 32'sd3, 32'sd0, -32'sd37, 32'sd12, 32'sd15, -32'sd9, -32'sd4, -32'sd6, 32'sd23, -32'sd2, 32'sd1, 32'sd1, -32'sd3, -32'sd9, -32'sd8, 32'sd3, -32'sd2, -32'sd1, -32'sd5, -32'sd5, -32'sd2, -32'sd3, -32'sd11, -32'sd1, -32'sd5, 32'sd6, -32'sd18, -32'sd8, 32'sd1, 32'sd0, 32'sd35, -32'sd3, 32'sd5, 32'sd1, 32'sd4, -32'sd5, -32'sd12, -32'sd1, 32'sd2, -32'sd4, -32'sd3, 32'sd6, -32'sd3, -32'sd3, 32'sd8, 32'sd2, -32'sd2, -32'sd3, -32'sd3, 32'sd5, -32'sd1, -32'sd4, 32'sd5, 32'sd3, 32'sd26, 32'sd2, 32'sd5, -32'sd4, -32'sd5, -32'sd8, -32'sd2, 32'sd9, -32'sd3, -32'sd3, 32'sd0, 32'sd5, 32'sd4, 32'sd1, -32'sd1, -32'sd4, -32'sd1, -32'sd7, 32'sd1, 32'sd4, -32'sd4, 32'sd6, -32'sd1, 32'sd8, -32'sd6, 32'sd2, 32'sd4, -32'sd3, 32'sd4, 32'sd7, -32'sd4, 32'sd3, -32'sd3, 32'sd4, -32'sd1, -32'sd1, 32'sd0, -32'sd5, -32'sd4, 32'sd1, -32'sd12, 32'sd3, 32'sd0, 32'sd4, 32'sd2, 32'sd0, -32'sd6, -32'sd6, -32'sd14, -32'sd16, -32'sd6, -32'sd6, -32'sd16, -32'sd3, -32'sd2, -32'sd6, 32'sd7, -32'sd1, 32'sd2, 32'sd1, 32'sd1, 32'sd1, 32'sd1, -32'sd4, -32'sd5, -32'sd4, 32'sd0, 32'sd24, 32'sd1, 32'sd3, -32'sd3, 32'sd1, 32'sd7, 32'sd0, 32'sd2, 32'sd2, 32'sd4, 32'sd1, 32'sd18, 32'sd2, -32'sd2, -32'sd1, -32'sd2, -32'sd13, -32'sd1, 32'sd6, -32'sd15, 32'sd1, 32'sd3, -32'sd2, 32'sd7, -32'sd1, 32'sd1, -32'sd2, -32'sd3, 32'sd2, -32'sd2, 32'sd4, 32'sd12, 32'sd3, 32'sd2, 32'sd0, -32'sd1, 32'sd3, -32'sd5, -32'sd1, -32'sd3, -32'sd3, 32'sd2, 32'sd12, -32'sd4, -32'sd2, 32'sd0, 32'sd2, -32'sd2, -32'sd1, -32'sd3, -32'sd2, -32'sd5, -32'sd1, -32'sd2, -32'sd6, -32'sd8, 32'sd0, 32'sd3, 32'sd3, 32'sd3, -32'sd4, 32'sd0, 32'sd7, -32'sd12, 32'sd2, 32'sd29, -32'sd23, -32'sd9, 32'sd2, 32'sd1, -32'sd2, 32'sd2, 32'sd2, -32'sd5, 32'sd2, -32'sd3, -32'sd3, -32'sd1, 32'sd2, -32'sd4, -32'sd4, -32'sd2, 32'sd5, -32'sd2, 32'sd0, 32'sd2, 32'sd4, 32'sd0, 32'sd11, -32'sd8, 32'sd6, 32'sd5, 32'sd5, 32'sd8, -32'sd3, -32'sd21, 32'sd9, 32'sd1, 32'sd0, 
                                                    32'sd10, -32'sd7, 32'sd1, -32'sd2, 32'sd12, 32'sd1, 32'sd1, 32'sd4, -32'sd7, -32'sd9, -32'sd1, 32'sd9, -32'sd9, -32'sd3, 32'sd3, -32'sd6, 32'sd24, -32'sd6, 32'sd3, 32'sd1, 32'sd3, -32'sd12, -32'sd2, 32'sd2, 32'sd4, 32'sd1, -32'sd7, -32'sd2, 32'sd3, 32'sd6, 32'sd2, 32'sd21, 32'sd2, -32'sd2, 32'sd10, 32'sd5, 32'sd4, 32'sd2, 32'sd6, 32'sd4, 32'sd5, -32'sd2, 32'sd2, 32'sd1, 32'sd4, 32'sd0, 32'sd6, 32'sd4, 32'sd4, 32'sd1, -32'sd1, 32'sd2, 32'sd1, 32'sd0, -32'sd2, 32'sd4, 32'sd1, 32'sd1, 32'sd3, -32'sd3, 32'sd0, 32'sd1, 32'sd3, -32'sd7, -32'sd8, -32'sd4, -32'sd5, 32'sd16, -32'sd1, -32'sd8, 32'sd1, -32'sd2, 32'sd2, 32'sd1, -32'sd1, 32'sd27, -32'sd3, 32'sd8, -32'sd1, 32'sd6, -32'sd3, -32'sd1, 32'sd0, 32'sd6, 32'sd0, -32'sd4, 32'sd11, -32'sd17, -32'sd1, -32'sd2, -32'sd3, -32'sd7, -32'sd11, -32'sd7, -32'sd1, 32'sd7, -32'sd9, -32'sd3, 32'sd1, 32'sd3, -32'sd3, -32'sd3, -32'sd7, 32'sd1, -32'sd3, -32'sd11, 32'sd17, 32'sd2, 32'sd1, -32'sd6, 32'sd7, -32'sd1, -32'sd7, 32'sd6, 32'sd1, 32'sd3, -32'sd2, -32'sd5, 32'sd0, 32'sd3, 32'sd1, 32'sd4, -32'sd1, 32'sd7, -32'sd3, -32'sd2, 32'sd2, 32'sd4, 32'sd4, 32'sd0, -32'sd6, 32'sd10, 32'sd3, 32'sd0, -32'sd11, -32'sd2, -32'sd1, 32'sd12, 32'sd70, 32'sd5, 32'sd3, 32'sd7, -32'sd2, -32'sd16, 32'sd0, 32'sd15, 32'sd5, 32'sd1, -32'sd3, -32'sd4, -32'sd1, -32'sd7, -32'sd2, -32'sd1, -32'sd6, 32'sd8, -32'sd2, 32'sd6, 32'sd0, 32'sd6, 32'sd4, 32'sd4, -32'sd1, 32'sd2, 32'sd0, -32'sd7, -32'sd2, -32'sd7, 32'sd7, -32'sd3, 32'sd0, -32'sd5, -32'sd3, 32'sd4, 32'sd15, -32'sd3, 32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd5, -32'sd2, 32'sd0, -32'sd5, -32'sd4, 32'sd3, 32'sd4, -32'sd2, 32'sd2, 32'sd0, 32'sd13, 32'sd0, 32'sd1, -32'sd5, -32'sd3, 32'sd2, -32'sd1, 32'sd3, -32'sd3, 32'sd0, -32'sd5, 32'sd4, 32'sd6, 32'sd5, 32'sd6, -32'sd2, 32'sd10, 32'sd13, -32'sd2, -32'sd2, -32'sd2, -32'sd3, 32'sd1, -32'sd3, 32'sd1, -32'sd2, 32'sd3, 32'sd11, 32'sd3, -32'sd5, -32'sd10, -32'sd2, 32'sd15, 32'sd20, -32'sd6, -32'sd1, 32'sd12, 32'sd2, 32'sd0, 32'sd4, -32'sd4, 32'sd0, -32'sd8, 32'sd0, 32'sd3, -32'sd7, 32'sd1, 32'sd2, -32'sd1, 32'sd5, -32'sd51, -32'sd3, -32'sd2, -32'sd2, 32'sd3, 32'sd2, -32'sd3, 32'sd8, 32'sd14, -32'sd4, 32'sd0, -32'sd1, -32'sd1, 32'sd3, 32'sd1, -32'sd6, 32'sd0, 32'sd15, 32'sd2, 32'sd7, -32'sd1, 32'sd16, -32'sd1, 32'sd2, -32'sd6, -32'sd4, -32'sd3, -32'sd2, -32'sd2, 32'sd0, -32'sd6, 32'sd5, 32'sd1, -32'sd2, 32'sd1, 32'sd6, 32'sd1, 32'sd0, 32'sd1, -32'sd6, -32'sd3, 32'sd4, 32'sd6, 32'sd0, -32'sd3, 32'sd2, 32'sd2, 32'sd8, -32'sd5, -32'sd11, 32'sd6, 32'sd3, -32'sd1, 32'sd3, -32'sd11, 32'sd3, -32'sd2, 32'sd4, 32'sd0, 32'sd7, -32'sd14, -32'sd1, 32'sd10, -32'sd12, 32'sd6, -32'sd2, 32'sd11, 32'sd10, -32'sd4, 32'sd2, 32'sd7, 32'sd3, 32'sd1, -32'sd5, 32'sd20, -32'sd9, -32'sd4, -32'sd8, 32'sd1, -32'sd1, -32'sd17, 32'sd7, -32'sd1, 32'sd4, 32'sd5, -32'sd4, -32'sd2, -32'sd1, 32'sd1, -32'sd6, 32'sd3, 32'sd4, -32'sd9, 32'sd4, 32'sd0, 32'sd0, 32'sd4, -32'sd2, 32'sd5, 32'sd0, -32'sd5, -32'sd3, 32'sd1, -32'sd3, 32'sd3, -32'sd5, -32'sd1, 32'sd7, 32'sd3, 32'sd0, 32'sd2, 32'sd14, 32'sd5, -32'sd1, 32'sd3, -32'sd4, 32'sd3, 32'sd1, 32'sd1, 32'sd3, 32'sd10, 32'sd1, 32'sd0, 32'sd0, 32'sd4, -32'sd4, 32'sd3, -32'sd3, 32'sd1, 32'sd2, 32'sd4, 32'sd1, -32'sd1, -32'sd1, -32'sd3, -32'sd5, -32'sd2, 32'sd1, -32'sd1, 32'sd3, -32'sd3, -32'sd9, -32'sd3, -32'sd6, -32'sd14, 32'sd2, -32'sd1, -32'sd1, -32'sd5, 32'sd1, -32'sd4, 32'sd7, -32'sd5, -32'sd3, -32'sd1, 32'sd2, 32'sd1, -32'sd3, 32'sd1, 32'sd5, 32'sd2, -32'sd3, 32'sd1, 32'sd1, -32'sd1, -32'sd1, 32'sd13, 32'sd7, 32'sd2, -32'sd4, -32'sd7, -32'sd1, 32'sd4, 32'sd0, 32'sd1, 32'sd10, 32'sd7, -32'sd3, 32'sd1, -32'sd4, 32'sd5, 32'sd2, -32'sd6, -32'sd3, 32'sd2, 32'sd13, -32'sd2, 32'sd5, 32'sd3, -32'sd4, 32'sd1, -32'sd6, -32'sd5, 32'sd6, 32'sd7, 32'sd2, -32'sd12, 32'sd1, 32'sd5, 32'sd6, -32'sd2, -32'sd5, -32'sd5, 32'sd3, 32'sd1, -32'sd17, 32'sd1, 32'sd1, -32'sd8, 32'sd0, 32'sd0, 32'sd3, 32'sd1, 32'sd3, -32'sd5, 32'sd3, 32'sd2, -32'sd3, -32'sd2, 32'sd58, 32'sd2, -32'sd3, -32'sd6, -32'sd2, -32'sd3, 32'sd3, -32'sd3, 32'sd0, 32'sd2, -32'sd3, 32'sd0, 32'sd0, -32'sd4, -32'sd1, 32'sd4, -32'sd4, 32'sd2, -32'sd4, 32'sd1, 32'sd8, -32'sd8, -32'sd12, -32'sd5, 32'sd3, -32'sd3, -32'sd5, -32'sd2, 32'sd1, -32'sd1, -32'sd1, 32'sd0, -32'sd4, -32'sd2, -32'sd1, -32'sd4, 32'sd2, -32'sd2, -32'sd11, 32'sd1, -32'sd4, 32'sd0, -32'sd14, 32'sd2, 32'sd1, -32'sd3, -32'sd2, -32'sd1, 32'sd9, -32'sd2, 32'sd0, -32'sd7, -32'sd1, 32'sd27, 32'sd2, 32'sd5, 32'sd3, -32'sd4, 32'sd8, 32'sd3, -32'sd10, 32'sd2, -32'sd9, 32'sd17, -32'sd6, -32'sd4, 32'sd0, -32'sd3, 32'sd0, 32'sd2, 32'sd3, -32'sd6, -32'sd3, 32'sd3, 32'sd24, -32'sd10, -32'sd6, -32'sd2, 32'sd0, -32'sd13, -32'sd3, 32'sd8, -32'sd3, 32'sd4, 32'sd5, -32'sd3, 32'sd3, -32'sd3, -32'sd3, 32'sd0, 32'sd14, 32'sd6, 32'sd6, 32'sd0, 32'sd9, 32'sd5, -32'sd3, 32'sd54, 32'sd1, -32'sd2, -32'sd2, -32'sd2, 32'sd0, 32'sd12, -32'sd2, -32'sd3, -32'sd3, -32'sd2, 32'sd4, 32'sd7, 32'sd1, -32'sd2, 32'sd29, 32'sd14, 32'sd0, 32'sd11, 32'sd3, -32'sd2, 32'sd42, 32'sd1, 32'sd6, -32'sd5, -32'sd10, 32'sd28, 32'sd2, 32'sd7, 32'sd1, 32'sd1, -32'sd3, 32'sd0, 32'sd7, -32'sd1, -32'sd5, -32'sd3, -32'sd2, -32'sd3, 32'sd7, 32'sd0, 32'sd1, -32'sd7, -32'sd2, -32'sd4, -32'sd38, -32'sd5, -32'sd7, 32'sd4, -32'sd1, -32'sd1, 32'sd0, 32'sd7, -32'sd16, 32'sd12, 32'sd5, 32'sd0, 32'sd1, 32'sd3, -32'sd2, -32'sd1, -32'sd1, 32'sd3, -32'sd2, 32'sd2, -32'sd6, 32'sd1, 32'sd1, 32'sd2, 32'sd12, 32'sd6, 32'sd1, -32'sd5, 32'sd3, 32'sd1, 32'sd8, 32'sd1, 32'sd2, -32'sd6, 32'sd7, 32'sd3, 32'sd5, -32'sd3, -32'sd11, 32'sd1, 32'sd10, -32'sd12, -32'sd4, 32'sd1, -32'sd1, 32'sd3, -32'sd2, 32'sd3, -32'sd2, 32'sd4, -32'sd1, 32'sd3, -32'sd4, 32'sd0, 32'sd4, 32'sd1, 32'sd4, 32'sd1, 32'sd6, -32'sd4, 32'sd3, 32'sd3, 32'sd1, -32'sd7, 32'sd4, -32'sd4, 
                                                    32'sd2, -32'sd6, 32'sd11, 32'sd3, 32'sd2, -32'sd2, 32'sd0, 32'sd2, -32'sd1, -32'sd2, -32'sd13, -32'sd12, -32'sd5, 32'sd0, 32'sd14, 32'sd0, 32'sd4, 32'sd1, -32'sd2, -32'sd2, 32'sd3, 32'sd6, -32'sd3, 32'sd5, 32'sd3, -32'sd3, 32'sd10, -32'sd2, -32'sd3, -32'sd9, -32'sd1, 32'sd3, -32'sd5, 32'sd3, 32'sd6, 32'sd5, 32'sd10, 32'sd4, 32'sd1, -32'sd8, -32'sd9, -32'sd15, 32'sd0, -32'sd6, 32'sd7, -32'sd4, 32'sd3, -32'sd18, 32'sd7, 32'sd3, -32'sd2, -32'sd3, -32'sd3, 32'sd2, 32'sd7, 32'sd2, -32'sd3, 32'sd0, -32'sd1, 32'sd12, -32'sd8, 32'sd2, -32'sd3, -32'sd1, -32'sd1, -32'sd4, -32'sd3, -32'sd5, 32'sd1, 32'sd21, 32'sd12, 32'sd5, 32'sd2, 32'sd18, 32'sd2, -32'sd1, -32'sd1, 32'sd0, 32'sd4, -32'sd2, 32'sd0, 32'sd0, 32'sd0, 32'sd1, 32'sd2, -32'sd7, 32'sd12, 32'sd3, 32'sd0, -32'sd4, -32'sd3, 32'sd3, -32'sd4, -32'sd3, -32'sd2, -32'sd8, -32'sd6, -32'sd3, -32'sd1, 32'sd1, -32'sd3, -32'sd2, -32'sd2, 32'sd4, 32'sd5, -32'sd3, -32'sd8, -32'sd1, 32'sd0, -32'sd3, -32'sd2, -32'sd3, 32'sd20, 32'sd9, -32'sd1, -32'sd2, -32'sd4, 32'sd3, 32'sd12, 32'sd4, 32'sd0, -32'sd5, -32'sd3, -32'sd2, 32'sd4, -32'sd4, -32'sd1, -32'sd3, -32'sd2, -32'sd5, 32'sd4, 32'sd1, 32'sd2, 32'sd6, 32'sd0, 32'sd3, -32'sd2, 32'sd5, -32'sd10, -32'sd2, 32'sd4, -32'sd15, 32'sd15, 32'sd1, -32'sd9, 32'sd23, 32'sd1, -32'sd2, 32'sd2, 32'sd3, 32'sd8, -32'sd4, -32'sd3, 32'sd2, 32'sd4, -32'sd1, -32'sd2, -32'sd2, 32'sd9, 32'sd1, -32'sd5, 32'sd1, 32'sd22, 32'sd15, -32'sd3, -32'sd7, 32'sd29, 32'sd1, -32'sd15, 32'sd5, 32'sd3, -32'sd5, -32'sd17, -32'sd5, -32'sd4, 32'sd2, -32'sd5, -32'sd9, -32'sd3, 32'sd5, 32'sd13, -32'sd10, -32'sd3, -32'sd1, 32'sd0, 32'sd0, 32'sd2, -32'sd3, -32'sd1, 32'sd0, -32'sd6, 32'sd1, 32'sd4, -32'sd1, -32'sd3, -32'sd4, 32'sd6, 32'sd6, 32'sd3, 32'sd1, 32'sd12, 32'sd22, -32'sd6, 32'sd14, -32'sd2, 32'sd4, 32'sd3, 32'sd3, 32'sd11, 32'sd11, -32'sd7, -32'sd8, -32'sd3, 32'sd7, 32'sd0, 32'sd13, -32'sd1, 32'sd6, -32'sd1, 32'sd2, 32'sd3, -32'sd4, 32'sd0, 32'sd0, 32'sd1, 32'sd8, -32'sd4, 32'sd6, -32'sd4, 32'sd16, 32'sd1, 32'sd4, 32'sd3, 32'sd1, -32'sd2, 32'sd0, 32'sd5, -32'sd6, 32'sd4, -32'sd5, -32'sd5, 32'sd2, -32'sd3, -32'sd3, 32'sd2, -32'sd6, -32'sd1, 32'sd6, -32'sd2, 32'sd0, 32'sd0, -32'sd4, -32'sd1, -32'sd4, 32'sd1, 32'sd1, 32'sd12, -32'sd4, -32'sd2, 32'sd2, 32'sd2, -32'sd10, -32'sd2, 32'sd3, 32'sd0, -32'sd6, -32'sd1, -32'sd1, 32'sd1, 32'sd3, 32'sd3, -32'sd7, 32'sd3, 32'sd3, -32'sd2, -32'sd6, -32'sd9, 32'sd1, -32'sd4, -32'sd2, -32'sd6, 32'sd7, 32'sd5, 32'sd0, -32'sd4, 32'sd13, -32'sd5, -32'sd6, -32'sd15, -32'sd15, 32'sd9, 32'sd1, 32'sd3, 32'sd0, 32'sd4, -32'sd1, 32'sd3, 32'sd2, -32'sd1, -32'sd5, -32'sd12, -32'sd3, -32'sd3, -32'sd1, 32'sd9, 32'sd4, -32'sd6, -32'sd3, -32'sd2, -32'sd6, -32'sd3, -32'sd4, -32'sd1, -32'sd6, 32'sd2, 32'sd0, 32'sd3, -32'sd10, 32'sd6, -32'sd16, 32'sd2, 32'sd2, 32'sd5, 32'sd2, 32'sd2, 32'sd1, 32'sd5, -32'sd1, 32'sd4, -32'sd3, 32'sd3, 32'sd0, -32'sd5, 32'sd1, 32'sd6, 32'sd0, -32'sd1, -32'sd1, 32'sd0, -32'sd11, 32'sd6, 32'sd0, -32'sd2, 32'sd6, -32'sd4, -32'sd4, 32'sd1, 32'sd0, 32'sd14, 32'sd9, 32'sd0, 32'sd25, 32'sd20, -32'sd6, 32'sd7, 32'sd6, -32'sd5, -32'sd5, -32'sd5, 32'sd2, 32'sd0, 32'sd4, -32'sd1, 32'sd1, 32'sd12, 32'sd2, 32'sd1, -32'sd2, -32'sd1, 32'sd4, -32'sd2, -32'sd2, -32'sd5, 32'sd4, 32'sd8, 32'sd1, -32'sd5, 32'sd0, 32'sd1, 32'sd11, -32'sd4, -32'sd3, 32'sd5, 32'sd0, -32'sd1, 32'sd17, -32'sd2, -32'sd10, -32'sd2, -32'sd7, 32'sd0, 32'sd3, -32'sd3, -32'sd1, -32'sd5, 32'sd28, -32'sd2, 32'sd9, 32'sd7, 32'sd5, 32'sd8, 32'sd1, 32'sd8, -32'sd5, -32'sd1, 32'sd14, 32'sd2, 32'sd4, -32'sd3, -32'sd1, -32'sd1, -32'sd2, 32'sd2, 32'sd1, 32'sd2, 32'sd4, 32'sd3, 32'sd1, -32'sd7, 32'sd9, -32'sd3, -32'sd2, -32'sd5, 32'sd3, -32'sd1, 32'sd3, -32'sd9, 32'sd6, 32'sd1, 32'sd2, -32'sd1, -32'sd14, 32'sd6, -32'sd3, 32'sd2, 32'sd6, -32'sd4, 32'sd5, 32'sd24, -32'sd1, 32'sd1, -32'sd1, -32'sd1, 32'sd1, -32'sd3, 32'sd0, 32'sd0, 32'sd1, -32'sd3, 32'sd10, 32'sd2, -32'sd3, 32'sd4, 32'sd2, 32'sd11, -32'sd5, 32'sd0, -32'sd7, 32'sd3, -32'sd3, 32'sd1, 32'sd44, 32'sd1, 32'sd4, 32'sd0, 32'sd0, 32'sd7, -32'sd1, -32'sd2, -32'sd1, -32'sd1, -32'sd6, 32'sd2, 32'sd0, 32'sd0, 32'sd1, -32'sd1, 32'sd7, 32'sd2, 32'sd22, 32'sd7, -32'sd41, -32'sd3, 32'sd10, 32'sd3, 32'sd1, 32'sd4, -32'sd6, -32'sd7, 32'sd2, -32'sd6, -32'sd8, 32'sd1, 32'sd4, 32'sd8, 32'sd1, 32'sd0, 32'sd4, 32'sd4, 32'sd6, -32'sd3, -32'sd7, -32'sd3, 32'sd14, -32'sd5, 32'sd2, 32'sd3, 32'sd6, 32'sd5, 32'sd5, 32'sd2, -32'sd2, 32'sd0, -32'sd18, -32'sd1, -32'sd3, -32'sd18, -32'sd11, 32'sd0, -32'sd1, -32'sd2, -32'sd7, 32'sd2, 32'sd2, 32'sd0, -32'sd11, 32'sd4, -32'sd1, -32'sd3, 32'sd1, -32'sd4, -32'sd25, -32'sd14, -32'sd2, 32'sd0, 32'sd8, -32'sd7, -32'sd5, 32'sd11, -32'sd1, 32'sd1, 32'sd1, -32'sd2, 32'sd0, -32'sd9, -32'sd1, 32'sd0, -32'sd5, -32'sd4, -32'sd10, 32'sd5, -32'sd4, 32'sd6, 32'sd33, 32'sd0, -32'sd11, -32'sd1, -32'sd17, 32'sd5, 32'sd13, -32'sd2, -32'sd8, 32'sd3, 32'sd3, 32'sd2, 32'sd3, -32'sd5, -32'sd1, 32'sd2, -32'sd4, -32'sd2, 32'sd3, -32'sd13, -32'sd2, -32'sd2, -32'sd2, -32'sd16, 32'sd2, 32'sd4, 32'sd1, 32'sd1, 32'sd5, -32'sd10, -32'sd9, 32'sd8, 32'sd3, -32'sd10, -32'sd2, 32'sd1, -32'sd3, 32'sd0, -32'sd2, 32'sd1, 32'sd7, -32'sd14, 32'sd3, 32'sd0, 32'sd0, -32'sd3, 32'sd11, -32'sd1, 32'sd10, 32'sd1, -32'sd1, 32'sd4, -32'sd3, -32'sd7, -32'sd5, -32'sd1, 32'sd2, -32'sd5, -32'sd3, -32'sd3, -32'sd6, -32'sd3, 32'sd2, -32'sd4, 32'sd9, 32'sd0, -32'sd1, -32'sd2, -32'sd2, -32'sd1, 32'sd2, -32'sd6, -32'sd3, -32'sd3, 32'sd1, 32'sd3, 32'sd2, -32'sd1, -32'sd3, -32'sd8, -32'sd6, 32'sd1, -32'sd7, 32'sd41, 32'sd10, -32'sd2, 32'sd6, 32'sd1, -32'sd4, -32'sd4, 32'sd0, -32'sd2, -32'sd1, -32'sd7, 32'sd0, 32'sd2, 32'sd2, 32'sd2, -32'sd2, 32'sd0, -32'sd2, -32'sd2, 32'sd2, -32'sd1, -32'sd1, 32'sd1, 32'sd3, 32'sd4, -32'sd2, 32'sd3, 
                                                    32'sd53, -32'sd5, -32'sd1, 32'sd2, -32'sd1, 32'sd2, -32'sd1, -32'sd2, -32'sd6, 32'sd6, -32'sd5, 32'sd0, -32'sd6, -32'sd1, -32'sd6, 32'sd13, -32'sd2, 32'sd1, -32'sd2, 32'sd9, -32'sd2, -32'sd1, -32'sd7, 32'sd0, -32'sd6, -32'sd15, -32'sd2, -32'sd1, 32'sd7, 32'sd9, -32'sd2, -32'sd2, -32'sd5, -32'sd2, -32'sd1, -32'sd16, 32'sd6, 32'sd4, 32'sd1, -32'sd8, 32'sd0, -32'sd9, 32'sd13, 32'sd2, -32'sd1, -32'sd1, -32'sd8, 32'sd5, -32'sd5, 32'sd6, 32'sd6, 32'sd8, -32'sd8, 32'sd4, 32'sd0, -32'sd1, 32'sd6, 32'sd2, 32'sd6, 32'sd25, 32'sd2, 32'sd0, 32'sd3, -32'sd2, -32'sd1, -32'sd2, 32'sd6, 32'sd3, -32'sd2, -32'sd22, -32'sd15, -32'sd10, -32'sd2, -32'sd8, 32'sd1, 32'sd5, -32'sd5, -32'sd1, -32'sd3, 32'sd0, 32'sd2, 32'sd2, -32'sd8, 32'sd7, 32'sd3, -32'sd2, -32'sd13, 32'sd15, -32'sd2, -32'sd4, 32'sd2, -32'sd15, 32'sd0, 32'sd4, 32'sd3, -32'sd4, 32'sd5, -32'sd9, -32'sd5, 32'sd6, 32'sd8, 32'sd2, -32'sd4, -32'sd2, 32'sd9, 32'sd0, 32'sd2, 32'sd0, -32'sd1, 32'sd6, -32'sd4, 32'sd13, 32'sd0, 32'sd5, 32'sd0, 32'sd3, -32'sd1, 32'sd0, -32'sd2, -32'sd4, 32'sd0, -32'sd7, -32'sd8, 32'sd4, 32'sd4, -32'sd3, 32'sd2, 32'sd6, 32'sd24, 32'sd4, 32'sd2, -32'sd1, -32'sd1, 32'sd2, 32'sd3, -32'sd3, -32'sd2, 32'sd1, 32'sd0, -32'sd6, 32'sd7, 32'sd1, -32'sd7, 32'sd7, -32'sd2, 32'sd1, -32'sd3, -32'sd8, 32'sd0, 32'sd5, -32'sd2, -32'sd5, 32'sd13, 32'sd11, 32'sd5, 32'sd8, 32'sd19, 32'sd0, -32'sd4, 32'sd1, 32'sd6, -32'sd9, -32'sd40, 32'sd4, 32'sd1, -32'sd4, -32'sd1, 32'sd4, -32'sd4, 32'sd3, 32'sd2, -32'sd5, 32'sd1, -32'sd9, -32'sd1, -32'sd2, -32'sd2, -32'sd1, -32'sd7, 32'sd4, -32'sd1, -32'sd1, 32'sd10, -32'sd1, 32'sd4, 32'sd5, 32'sd2, -32'sd6, -32'sd2, -32'sd2, -32'sd5, 32'sd4, -32'sd1, 32'sd2, 32'sd9, 32'sd68, -32'sd2, 32'sd0, 32'sd6, -32'sd6, -32'sd12, 32'sd5, -32'sd2, -32'sd2, -32'sd7, -32'sd1, -32'sd9, -32'sd3, 32'sd2, -32'sd6, 32'sd6, 32'sd2, -32'sd12, 32'sd9, 32'sd7, -32'sd2, 32'sd3, 32'sd2, -32'sd7, -32'sd2, 32'sd1, 32'sd4, -32'sd3, 32'sd1, 32'sd11, -32'sd1, 32'sd1, -32'sd1, 32'sd1, 32'sd0, 32'sd5, -32'sd1, 32'sd4, -32'sd1, 32'sd11, 32'sd1, -32'sd2, -32'sd3, 32'sd14, -32'sd1, -32'sd7, 32'sd13, 32'sd3, -32'sd2, -32'sd41, 32'sd26, -32'sd9, 32'sd5, -32'sd9, 32'sd8, 32'sd5, 32'sd1, -32'sd6, -32'sd9, -32'sd5, 32'sd0, 32'sd2, 32'sd1, -32'sd4, 32'sd12, 32'sd0, 32'sd2, -32'sd18, -32'sd12, -32'sd1, 32'sd2, 32'sd9, -32'sd5, 32'sd66, -32'sd4, -32'sd5, 32'sd1, -32'sd2, 32'sd1, -32'sd18, 32'sd23, 32'sd1, 32'sd14, -32'sd4, -32'sd3, 32'sd0, -32'sd4, 32'sd2, 32'sd2, -32'sd2, -32'sd2, -32'sd4, -32'sd13, 32'sd5, -32'sd37, 32'sd20, 32'sd0, -32'sd3, 32'sd5, 32'sd7, 32'sd1, -32'sd7, 32'sd3, 32'sd3, 32'sd5, -32'sd13, 32'sd11, 32'sd2, 32'sd4, -32'sd8, 32'sd9, -32'sd4, -32'sd2, 32'sd3, 32'sd13, 32'sd3, 32'sd4, 32'sd5, -32'sd6, -32'sd5, 32'sd0, 32'sd5, 32'sd3, 32'sd0, -32'sd1, 32'sd2, 32'sd5, -32'sd9, -32'sd8, 32'sd4, 32'sd5, -32'sd4, -32'sd4, 32'sd0, -32'sd9, -32'sd10, 32'sd1, -32'sd5, -32'sd8, 32'sd2, -32'sd7, -32'sd6, 32'sd2, -32'sd3, -32'sd5, -32'sd5, -32'sd2, 32'sd0, -32'sd1, 32'sd5, 32'sd0, -32'sd3, 32'sd3, -32'sd2, 32'sd1, -32'sd1, 32'sd7, 32'sd7, -32'sd2, 32'sd12, -32'sd2, 32'sd4, 32'sd4, 32'sd2, -32'sd6, -32'sd1, -32'sd8, -32'sd9, 32'sd2, -32'sd1, 32'sd1, 32'sd0, 32'sd26, -32'sd2, -32'sd2, -32'sd3, -32'sd3, -32'sd3, 32'sd6, -32'sd6, 32'sd3, -32'sd6, -32'sd2, 32'sd2, 32'sd0, -32'sd6, -32'sd2, -32'sd2, -32'sd29, -32'sd16, 32'sd1, 32'sd1, 32'sd37, -32'sd30, 32'sd8, 32'sd1, -32'sd4, -32'sd2, -32'sd6, -32'sd10, 32'sd4, -32'sd12, -32'sd2, -32'sd1, 32'sd0, -32'sd1, -32'sd5, 32'sd4, -32'sd1, 32'sd0, 32'sd5, -32'sd3, 32'sd0, -32'sd2, 32'sd85, 32'sd14, 32'sd2, -32'sd3, -32'sd10, -32'sd7, -32'sd3, -32'sd6, -32'sd2, 32'sd3, 32'sd4, 32'sd3, -32'sd3, 32'sd8, 32'sd19, 32'sd7, 32'sd1, 32'sd0, -32'sd4, 32'sd3, 32'sd0, -32'sd2, -32'sd11, -32'sd2, -32'sd2, 32'sd2, -32'sd2, 32'sd2, -32'sd1, -32'sd3, -32'sd4, 32'sd1, -32'sd1, 32'sd2, 32'sd5, -32'sd7, -32'sd7, 32'sd0, 32'sd38, -32'sd11, -32'sd7, 32'sd5, -32'sd1, 32'sd0, -32'sd9, 32'sd1, -32'sd1, 32'sd2, 32'sd3, -32'sd2, -32'sd9, -32'sd2, 32'sd3, 32'sd2, -32'sd3, 32'sd1, 32'sd29, -32'sd5, -32'sd2, 32'sd5, 32'sd1, 32'sd12, -32'sd5, 32'sd1, 32'sd10, 32'sd4, -32'sd4, -32'sd1, 32'sd1, 32'sd14, -32'sd15, -32'sd5, -32'sd4, -32'sd16, 32'sd30, -32'sd4, 32'sd5, 32'sd9, 32'sd1, 32'sd7, -32'sd6, -32'sd5, -32'sd13, -32'sd16, -32'sd15, 32'sd4, 32'sd1, 32'sd7, 32'sd0, -32'sd4, -32'sd20, 32'sd1, 32'sd6, 32'sd3, 32'sd9, 32'sd1, -32'sd7, 32'sd14, 32'sd3, 32'sd4, 32'sd5, -32'sd1, 32'sd0, 32'sd3, -32'sd4, 32'sd10, -32'sd2, -32'sd2, -32'sd3, 32'sd3, 32'sd19, 32'sd0, 32'sd1, -32'sd1, -32'sd5, 32'sd3, -32'sd4, -32'sd2, -32'sd2, 32'sd1, -32'sd2, 32'sd2, -32'sd4, 32'sd0, 32'sd0, 32'sd6, -32'sd1, -32'sd6, 32'sd3, -32'sd3, 32'sd6, 32'sd8, -32'sd5, 32'sd0, 32'sd3, -32'sd2, -32'sd1, -32'sd2, -32'sd1, -32'sd16, -32'sd11, 32'sd8, -32'sd4, -32'sd10, -32'sd2, -32'sd1, -32'sd2, 32'sd0, 32'sd4, 32'sd4, 32'sd4, -32'sd2, -32'sd11, 32'sd1, 32'sd7, -32'sd1, -32'sd2, 32'sd7, -32'sd3, -32'sd9, -32'sd2, 32'sd4, 32'sd7, 32'sd5, -32'sd16, 32'sd0, 32'sd1, 32'sd6, -32'sd10, 32'sd1, -32'sd2, 32'sd4, -32'sd4, -32'sd9, -32'sd2, 32'sd6, 32'sd4, -32'sd4, 32'sd5, -32'sd3, 32'sd8, 32'sd4, 32'sd5, -32'sd3, -32'sd3, -32'sd1, -32'sd7, -32'sd3, 32'sd1, 32'sd4, -32'sd3, -32'sd1, 32'sd3, 32'sd4, 32'sd2, 32'sd14, -32'sd2, 32'sd1, -32'sd1, -32'sd11, 32'sd0, 32'sd47, 32'sd28, -32'sd2, -32'sd6, 32'sd2, -32'sd4, -32'sd1, 32'sd17, 32'sd4, 32'sd6, 32'sd0, -32'sd3, -32'sd4, 32'sd2, 32'sd0, 32'sd0, -32'sd4, -32'sd4, 32'sd20, 32'sd11, 32'sd0, 32'sd1, 32'sd5, 32'sd10, 32'sd0, -32'sd1, 32'sd15, -32'sd1, -32'sd4, 32'sd3, 32'sd6, -32'sd3, 32'sd3, 32'sd1, -32'sd30, -32'sd3, -32'sd1, 32'sd1, -32'sd5, -32'sd2, -32'sd16, 32'sd9, 32'sd11, 32'sd2, 32'sd10, 32'sd2, -32'sd11, 32'sd9, -32'sd10, 32'sd12, -32'sd5, 
                                                    -32'sd1, 32'sd0, 32'sd2, -32'sd3, 32'sd7, 32'sd0, -32'sd2, 32'sd4, 32'sd0, 32'sd11, -32'sd5, 32'sd10, 32'sd5, 32'sd3, -32'sd9, 32'sd6, 32'sd10, 32'sd8, 32'sd4, 32'sd2, 32'sd3, 32'sd4, -32'sd2, -32'sd1, -32'sd4, -32'sd1, 32'sd41, -32'sd2, -32'sd1, -32'sd4, -32'sd1, 32'sd1, 32'sd1, 32'sd25, 32'sd1, -32'sd9, -32'sd4, 32'sd1, 32'sd12, -32'sd8, -32'sd22, 32'sd1, -32'sd5, 32'sd16, 32'sd11, 32'sd11, 32'sd7, 32'sd1, 32'sd2, 32'sd7, -32'sd3, 32'sd6, 32'sd3, 32'sd1, -32'sd4, 32'sd4, 32'sd0, -32'sd12, 32'sd2, 32'sd3, 32'sd0, -32'sd1, 32'sd2, 32'sd0, -32'sd10, 32'sd6, 32'sd0, 32'sd2, 32'sd5, -32'sd2, 32'sd7, 32'sd1, 32'sd6, 32'sd3, 32'sd20, -32'sd1, 32'sd0, -32'sd3, -32'sd1, -32'sd4, -32'sd3, 32'sd0, -32'sd1, -32'sd2, -32'sd1, -32'sd1, -32'sd5, 32'sd1, -32'sd1, 32'sd1, -32'sd1, 32'sd6, 32'sd2, 32'sd21, 32'sd0, 32'sd0, -32'sd3, -32'sd2, 32'sd2, 32'sd7, -32'sd5, -32'sd4, -32'sd5, -32'sd4, -32'sd11, 32'sd54, 32'sd8, -32'sd2, -32'sd1, -32'sd7, -32'sd2, 32'sd6, 32'sd0, -32'sd11, -32'sd3, 32'sd6, 32'sd0, 32'sd1, -32'sd2, 32'sd1, 32'sd3, -32'sd3, 32'sd8, -32'sd10, 32'sd1, -32'sd3, -32'sd5, 32'sd1, -32'sd2, 32'sd1, -32'sd9, 32'sd1, 32'sd14, 32'sd5, -32'sd14, -32'sd15, 32'sd2, -32'sd1, -32'sd4, 32'sd2, -32'sd5, 32'sd3, -32'sd3, -32'sd2, -32'sd15, -32'sd11, -32'sd3, -32'sd1, 32'sd1, -32'sd4, 32'sd1, 32'sd2, -32'sd2, 32'sd36, -32'sd30, -32'sd14, 32'sd16, -32'sd8, 32'sd2, 32'sd0, 32'sd4, -32'sd6, 32'sd1, 32'sd3, -32'sd3, 32'sd4, 32'sd2, 32'sd1, 32'sd5, -32'sd2, 32'sd7, 32'sd1, -32'sd3, -32'sd1, 32'sd4, 32'sd3, -32'sd1, 32'sd4, 32'sd1, -32'sd11, -32'sd2, 32'sd0, -32'sd2, -32'sd10, -32'sd30, -32'sd13, 32'sd0, 32'sd3, -32'sd14, 32'sd2, 32'sd9, 32'sd2, 32'sd1, 32'sd1, 32'sd1, 32'sd0, 32'sd0, -32'sd4, 32'sd2, -32'sd8, -32'sd3, 32'sd4, 32'sd2, 32'sd0, -32'sd5, 32'sd2, 32'sd10, -32'sd30, 32'sd18, 32'sd1, -32'sd7, -32'sd7, -32'sd3, 32'sd3, -32'sd2, 32'sd0, 32'sd1, -32'sd1, 32'sd1, 32'sd3, -32'sd1, 32'sd1, -32'sd4, 32'sd6, -32'sd5, 32'sd5, -32'sd9, 32'sd5, -32'sd5, -32'sd3, -32'sd20, 32'sd1, 32'sd3, 32'sd10, 32'sd0, -32'sd2, -32'sd4, 32'sd6, 32'sd0, 32'sd6, 32'sd14, -32'sd5, 32'sd4, -32'sd7, 32'sd2, 32'sd9, -32'sd2, -32'sd1, 32'sd0, 32'sd2, -32'sd5, 32'sd3, 32'sd7, -32'sd2, 32'sd0, 32'sd10, -32'sd3};

localparam logic [2912:0][31:0] feature_above = {-32'sd284, 32'sd170, 32'sd136, 32'sd151, 32'sd161, -32'sd240, 32'sd56, 32'sd57, 32'sd109, -32'sd201, 32'sd151, 32'sd90, 32'sd221, -32'sd279, 32'sd58, 32'sd69, 32'sd119, -32'sd85, -32'sd38, 32'sd174, -32'sd25, -32'sd68, 32'sd146, 32'sd99, -32'sd194, 32'sd188, 32'sd128, -32'sd204, 32'sd106, 32'sd54, 32'sd135, -32'sd172, 32'sd186, 32'sd155, -32'sd59, 32'sd20, -32'sd200, 32'sd30, 32'sd164, -32'sd39, -32'sd7, 32'sd197, 32'sd120, 32'sd123, -32'sd379, -32'sd56, 32'sd51, -32'sd339, 32'sd36, 32'sd30, 32'sd138, 32'sd13, -32'sd137, 32'sd98, 32'sd177, 32'sd66, 32'sd75, 32'sd150, 32'sd122, -32'sd18, 32'sd35, 32'sd30, -32'sd172, -32'sd115, -32'sd209, 32'sd23, -32'sd49, 32'sd32, -32'sd38, 32'sd81, 32'sd7, 32'sd50, 32'sd13, -32'sd161, -32'sd305, -32'sd35, -32'sd146, -32'sd162, 32'sd35, 32'sd91, 32'sd5, -32'sd6, -32'sd45, 32'sd27, 32'sd139, 32'sd180, 32'sd95, 32'sd48, 32'sd162, 32'sd59, -32'sd123, 32'sd6, 32'sd69, -32'sd191, -32'sd67, -32'sd205, 32'sd20, -32'sd92, 32'sd9, 32'sd87, 32'sd10, -32'sd28, 32'sd168, 32'sd156, 32'sd109, 32'sd38, -32'sd42, -32'sd107, -32'sd86, 32'sd18, 32'sd10, 32'sd25, 32'sd9, 32'sd100, 32'sd16, 32'sd2, 32'sd68, 32'sd50, -32'sd271, 32'sd126, 32'sd12, -32'sd19, -32'sd74, -32'sd22, -32'sd82, 32'sd32, -32'sd35, 32'sd30, -32'sd162, 32'sd39, 32'sd68, 32'sd31, 32'sd66, -32'sd2, -32'sd33, -32'sd76, 32'sd134, 32'sd71, 32'sd82, 32'sd68, 32'sd46, 32'sd46, -32'sd64, 32'sd109, 32'sd146, -32'sd23, -32'sd40, 32'sd134, 32'sd25, -32'sd170, -32'sd90, 32'sd29, -32'sd66, 32'sd79, 32'sd61, -32'sd88, 32'sd15, -32'sd7, 32'sd106, -32'sd23, -32'sd198, 32'sd31, -32'sd41, -32'sd106, 32'sd7, 32'sd17, 32'sd5, 32'sd63, -32'sd73, 32'sd82, 32'sd8, -32'sd128, 32'sd5, -32'sd133, -32'sd69, 32'sd57, 32'sd0, -32'sd83, 32'sd103, 32'sd27, -32'sd135, -32'sd110, 32'sd8, 32'sd81, 32'sd72, -32'sd193, 32'sd48, 32'sd16, 32'sd87, 32'sd122, 32'sd63, 32'sd64, -32'sd160, 32'sd76, 32'sd39, 32'sd29, -32'sd13, 32'sd24, -32'sd60, -32'sd34, 32'sd53, 32'sd76, -32'sd59, 32'sd18, -32'sd125, 32'sd23, -32'sd170, -32'sd268, 32'sd66, -32'sd164, -32'sd59, 32'sd6, 32'sd44, 32'sd55, 32'sd21, -32'sd60, -32'sd214, 32'sd5, 32'sd30, 32'sd13, -32'sd24, -32'sd49, 32'sd25, 32'sd65, 32'sd30, -32'sd41, -32'sd2, 32'sd133, -32'sd107, 32'sd58, -32'sd192, -32'sd49, -32'sd14, -32'sd215, 32'sd31, 32'sd60, 32'sd23, 32'sd9, -32'sd198, 32'sd48, -32'sd159, 32'sd7, 32'sd29, 32'sd157, -32'sd6, -32'sd28, -32'sd243, 32'sd1, -32'sd11, 32'sd8, -32'sd98, 32'sd105, 32'sd38, 32'sd74, 32'sd115, 32'sd65, -32'sd90, 32'sd91, 32'sd34, -32'sd49, 32'sd33, -32'sd75, 32'sd22, -32'sd112, 32'sd30, -32'sd72, 32'sd49, -32'sd178, -32'sd137, 32'sd25, 32'sd56, -32'sd57, 32'sd29, -32'sd1, -32'sd67, -32'sd193, 32'sd24, 32'sd0, -32'sd284, 32'sd8, -32'sd152, 32'sd16, 32'sd91, -32'sd135, 32'sd25, -32'sd32, -32'sd27, -32'sd36, 32'sd31, 32'sd7, 32'sd25, 32'sd135, -32'sd220, 32'sd8, 32'sd4, -32'sd62, 32'sd21, 32'sd5, 32'sd41, -32'sd34, 32'sd19, 32'sd5, 32'sd20, -32'sd54, 32'sd24, 32'sd0, 32'sd40, -32'sd83, 32'sd20, 32'sd196, 32'sd83, 32'sd5, -32'sd13, -32'sd44, -32'sd2, -32'sd4, 32'sd21, 32'sd0, -32'sd23, -32'sd164, -32'sd194, 32'sd42, 32'sd19, 32'sd142, -32'sd79, 32'sd51, 32'sd37, 32'sd58, -32'sd87, 32'sd8, -32'sd221, 32'sd16, -32'sd104, 32'sd86, 32'sd108, -32'sd61, 32'sd121, -32'sd40, 32'sd23, 32'sd32, -32'sd55, -32'sd205, 32'sd48, 32'sd32, -32'sd185, -32'sd174, 32'sd35, -32'sd104, -32'sd96, 32'sd104, 32'sd110, -32'sd127, 32'sd20, -32'sd90, -32'sd52, 32'sd9, -32'sd92, 32'sd34, 32'sd19, -32'sd138, 32'sd156, 32'sd2, -32'sd20, 32'sd90, 32'sd43, 32'sd10, 32'sd6, -32'sd31, 32'sd16, -32'sd3, -32'sd15, -32'sd34, -32'sd83, -32'sd159, 32'sd130, -32'sd46, 32'sd26, -32'sd3, -32'sd38, 32'sd139, 32'sd156, -32'sd136, 32'sd22, 32'sd66, 32'sd32, -32'sd296, -32'sd42, 32'sd9, -32'sd221, 32'sd130, 32'sd19, -32'sd37, -32'sd43, -32'sd300, 32'sd20, -32'sd4, 32'sd30, 32'sd118, 32'sd40, -32'sd347, -32'sd4, 32'sd29, -32'sd134, 32'sd98, 32'sd36, -32'sd33, 32'sd140, 32'sd68, 32'sd52, 32'sd95, 32'sd94, 32'sd49, 32'sd47, 32'sd102, -32'sd42, -32'sd124, -32'sd136, 32'sd17, 32'sd77, -32'sd27, -32'sd188, 32'sd26, 32'sd13, -32'sd51, -32'sd206, -32'sd17, 32'sd1, 32'sd33, -32'sd92, -32'sd211, 32'sd3, -32'sd13, -32'sd69, 32'sd26, -32'sd129, -32'sd35, -32'sd68, 32'sd27, -32'sd5, -32'sd91, 32'sd2, -32'sd8, 32'sd102, -32'sd88, -32'sd28, 32'sd160, 32'sd19, -32'sd2, 32'sd138, 32'sd146, -32'sd1, 32'sd31, -32'sd26, -32'sd156, 32'sd7, 32'sd37, -32'sd86, 32'sd2, 32'sd3, 32'sd4, 32'sd76, 32'sd34, -32'sd43, 32'sd20, -32'sd3, -32'sd6, -32'sd57, 32'sd18, -32'sd49, 32'sd8, 32'sd102, 32'sd15, -32'sd1, 32'sd52, -32'sd49, 32'sd98, -32'sd29, -32'sd186, 32'sd33, 32'sd62, -32'sd28, 32'sd19, -32'sd26, 32'sd35, -32'sd24, 32'sd20, -32'sd210, 32'sd31, -32'sd1, -32'sd58, 32'sd56, 32'sd32, 32'sd3, 32'sd0, 32'sd195, -32'sd28, 32'sd3, 32'sd82, 32'sd74, 32'sd168, 32'sd37, 32'sd68, -32'sd57, -32'sd35, 32'sd26, 32'sd9, -32'sd67, 32'sd6, 32'sd24, -32'sd88, -32'sd108, -32'sd175, 32'sd33, 32'sd8, -32'sd2, -32'sd42, 32'sd26, 32'sd29, -32'sd137, 32'sd5, -32'sd92, -32'sd68, 32'sd125, -32'sd30, 32'sd59, -32'sd341, 32'sd3, -32'sd278, 32'sd96, 32'sd1, 32'sd127, -32'sd32, -32'sd78, 32'sd4, -32'sd17, -32'sd67, 32'sd19, 32'sd0, -32'sd79, -32'sd27, 32'sd61, 32'sd14, -32'sd192, 32'sd104, -32'sd9, 32'sd6, -32'sd1, -32'sd24, 32'sd12, -32'sd35, 32'sd20, -32'sd30, 32'sd25, 32'sd3, -32'sd2, -32'sd222, -32'sd7, -32'sd99, 32'sd86, 32'sd40, 32'sd33, 32'sd53, 32'sd2, -32'sd27, 32'sd5, 32'sd22, 32'sd105, 32'sd3, -32'sd44, 32'sd0, 32'sd32, -32'sd183, 32'sd43, 32'sd17, -32'sd40, 32'sd91, 32'sd25, -32'sd114, -32'sd35, 32'sd3, -32'sd22, -32'sd26, 32'sd15, -32'sd58, 32'sd50, -32'sd26, 32'sd26, -32'sd131, -32'sd12, -32'sd247, -32'sd9, 32'sd24, 32'sd28, -32'sd24, 32'sd48, -32'sd34, 32'sd74, 
                                                    32'sd129, 32'sd72, 32'sd40, -32'sd143, 32'sd42, 32'sd67, -32'sd4, 32'sd15, 32'sd27, -32'sd36, -32'sd90, 32'sd94, 32'sd20, -32'sd44, -32'sd17, -32'sd123, -32'sd60, -32'sd67, 32'sd28, 32'sd8, 32'sd28, 32'sd6, 32'sd22, -32'sd28, 32'sd23, 32'sd7, 32'sd67, 32'sd72, -32'sd90, 32'sd6, 32'sd33, 32'sd74, 32'sd25, 32'sd27, 32'sd99, -32'sd32, -32'sd5, 32'sd141, 32'sd92, 32'sd6, -32'sd48, 32'sd143, 32'sd25, -32'sd149, 32'sd21, -32'sd2, -32'sd11, 32'sd76, 32'sd17, -32'sd4, 32'sd2, 32'sd68, 32'sd21, -32'sd96, -32'sd84, -32'sd157, 32'sd55, -32'sd153, 32'sd18, 32'sd69, 32'sd72, -32'sd102, 32'sd190, -32'sd4, 32'sd4, 32'sd38, -32'sd49, -32'sd68, 32'sd269, -32'sd5, 32'sd46, -32'sd23, -32'sd166, 32'sd18, 32'sd50, -32'sd92, 32'sd8, -32'sd21, -32'sd21, 32'sd94, 32'sd26, -32'sd38, 32'sd52, -32'sd22, 32'sd89, 32'sd0, 32'sd69, -32'sd96, 32'sd43, -32'sd5, 32'sd2, 32'sd93, -32'sd63, 32'sd99, 32'sd9, -32'sd24, -32'sd205, 32'sd152, 32'sd50, -32'sd206, 32'sd69, -32'sd41, -32'sd132, -32'sd101, -32'sd107, -32'sd80, 32'sd201, 32'sd49, 32'sd67, -32'sd36, -32'sd39, -32'sd112, -32'sd26, 32'sd10, 32'sd73, 32'sd57, 32'sd87, 32'sd25, -32'sd91, 32'sd15, 32'sd26, 32'sd47, 32'sd16, 32'sd74, -32'sd67, 32'sd61, -32'sd199, 32'sd24, -32'sd57, -32'sd27, 32'sd67, 32'sd4, -32'sd29, 32'sd19, 32'sd2, -32'sd126, 32'sd3, 32'sd25, 32'sd49, -32'sd19, -32'sd36, 32'sd77, -32'sd48, 32'sd132, -32'sd29, -32'sd152, 32'sd6, 32'sd137, -32'sd22, -32'sd9, 32'sd51, -32'sd156, -32'sd91, 32'sd23, -32'sd198, 32'sd21, -32'sd2, 32'sd30, 32'sd7, -32'sd2, -32'sd27, 32'sd24, -32'sd51, -32'sd329, -32'sd2, 32'sd21, 32'sd42, -32'sd62, -32'sd29, 32'sd24, -32'sd27, -32'sd77, -32'sd3, 32'sd8, -32'sd197, 32'sd48, 32'sd18, -32'sd2, -32'sd157, 32'sd0, -32'sd2, -32'sd159, 32'sd66, -32'sd91, 32'sd0, 32'sd19, -32'sd60, -32'sd53, 32'sd56, -32'sd122, -32'sd39, -32'sd253, -32'sd1, -32'sd4, 32'sd50, 32'sd75, -32'sd121, 32'sd27, -32'sd4, 32'sd149, -32'sd143, 32'sd27, -32'sd20, 32'sd23, 32'sd6, -32'sd96, -32'sd214, 32'sd98, -32'sd113, -32'sd315, -32'sd38, 32'sd21, -32'sd48, 32'sd76, 32'sd71, 32'sd52, -32'sd30, 32'sd20, -32'sd44, 32'sd12, 32'sd4, -32'sd7, -32'sd3, 32'sd117, -32'sd37, 32'sd68, -32'sd57, -32'sd328, -32'sd142, 32'sd73, 32'sd16, 32'sd112, 32'sd27, 32'sd7, -32'sd1, 32'sd22, -32'sd178, 32'sd0, -32'sd53, 32'sd2, -32'sd25, 32'sd66, 32'sd90, -32'sd86, 32'sd46, 32'sd24, 32'sd34, 32'sd34, -32'sd138, -32'sd36, 32'sd31, -32'sd32, 32'sd1, 32'sd91, -32'sd184, 32'sd6, -32'sd57, 32'sd44, -32'sd172, -32'sd66, -32'sd93, -32'sd3, 32'sd25, -32'sd112, -32'sd31, -32'sd160, -32'sd11, -32'sd62, 32'sd23, 32'sd80, 32'sd118, 32'sd99, -32'sd139, -32'sd30, 32'sd79, 32'sd129, 32'sd6, 32'sd1, 32'sd2, -32'sd37, -32'sd21, -32'sd1, -32'sd38, -32'sd4, -32'sd91, -32'sd194, -32'sd50, -32'sd3, 32'sd19, -32'sd53, 32'sd53, 32'sd71, 32'sd2, -32'sd38, -32'sd59, -32'sd66, 32'sd27, 32'sd184, -32'sd5, 32'sd17, 32'sd14, 32'sd29, 32'sd48, -32'sd25, 32'sd75, -32'sd86, -32'sd10, 32'sd149, 32'sd6, -32'sd28, 32'sd26, 32'sd5, 32'sd46, 32'sd25, 32'sd31, 32'sd163, -32'sd276, -32'sd21, 32'sd27, -32'sd25, 32'sd28, -32'sd128, 32'sd63, -32'sd22, -32'sd96, 32'sd70, -32'sd65, -32'sd123, 32'sd22, -32'sd168, 32'sd2, 32'sd31, 32'sd20, -32'sd2, 32'sd8, -32'sd6, 32'sd20, 32'sd7, 32'sd1, -32'sd171, 32'sd48, -32'sd19, 32'sd33, -32'sd134, 32'sd51, 32'sd4, 32'sd48, -32'sd27, 32'sd23, -32'sd83, -32'sd127, 32'sd4, 32'sd0, 32'sd60, 32'sd73, -32'sd244, -32'sd1, -32'sd7, -32'sd157, -32'sd139, -32'sd47, 32'sd30, 32'sd20, -32'sd243, 32'sd3, 32'sd78, 32'sd24, 32'sd275, 32'sd17, -32'sd66, 32'sd158, -32'sd4, 32'sd206, -32'sd1, 32'sd122, 32'sd248, -32'sd89, 32'sd39, 32'sd73, 32'sd74, 32'sd55, -32'sd26, 32'sd141, 32'sd7, -32'sd43, 32'sd29, 32'sd8, 32'sd24, -32'sd33, 32'sd91, 32'sd10, 32'sd116, 32'sd93, 32'sd27, -32'sd2, -32'sd15, -32'sd98, 32'sd5, 32'sd76, 32'sd42, -32'sd33, -32'sd72, -32'sd67, 32'sd38, 32'sd32, -32'sd60, -32'sd145, -32'sd34, -32'sd2, 32'sd20, -32'sd90, 32'sd30, 32'sd58, 32'sd18, -32'sd33, -32'sd227, 32'sd69, 32'sd43, -32'sd149, -32'sd319, 32'sd123, -32'sd33, -32'sd129, 32'sd25, -32'sd128, 32'sd53, 32'sd50, -32'sd46, 32'sd119, 32'sd43, 32'sd12, 32'sd31, -32'sd161, 32'sd22, -32'sd112, 32'sd17, 32'sd28, -32'sd65, 32'sd59, 32'sd71, 32'sd2, -32'sd22, 32'sd1, 32'sd14, -32'sd24, 32'sd105, -32'sd44, -32'sd178, 32'sd0, 32'sd15, -32'sd3, 32'sd15, -32'sd27, 32'sd68, -32'sd40, -32'sd7, -32'sd2, 32'sd54, 32'sd5, 32'sd81, 32'sd1, -32'sd8, 32'sd11, -32'sd51, 32'sd66, 32'sd18, 32'sd80, -32'sd349, -32'sd138, 32'sd4, 32'sd56, -32'sd31, -32'sd39, 32'sd33, -32'sd251, 32'sd95, 32'sd34, 32'sd22, -32'sd33, -32'sd37, -32'sd226, -32'sd3, 32'sd132, -32'sd160, -32'sd220, 32'sd26, 32'sd26, 32'sd26, 32'sd214, -32'sd45, -32'sd23, 32'sd16, -32'sd148, -32'sd599, -32'sd19, 32'sd44, 32'sd39, 32'sd3, 32'sd28, 32'sd20, -32'sd1, -32'sd88, 32'sd156, -32'sd53, -32'sd2, 32'sd25, -32'sd54, 32'sd100, -32'sd4, 32'sd8, -32'sd24, -32'sd101, 32'sd75, -32'sd38, 32'sd53, 32'sd22, 32'sd3, -32'sd53, 32'sd46, 32'sd110, 32'sd13, -32'sd89, 32'sd5, -32'sd89, -32'sd124, 32'sd0, -32'sd42, 32'sd93, 32'sd39, -32'sd13, -32'sd28, -32'sd20, -32'sd3, -32'sd49, -32'sd35, 32'sd34, 32'sd71, 32'sd4, 32'sd8, -32'sd27, 32'sd8, 32'sd36, -32'sd113, 32'sd20, 32'sd54, 32'sd20, 32'sd16, 32'sd105, -32'sd22, 32'sd19, -32'sd4, -32'sd89, -32'sd3, 32'sd19, 32'sd5, 32'sd103, -32'sd32, 32'sd25, 32'sd17, 32'sd24, -32'sd45, 32'sd27, -32'sd2, -32'sd58, 32'sd2, 32'sd4, 32'sd35, 32'sd22, 32'sd9, 32'sd15, 32'sd142, 32'sd59, -32'sd24, 32'sd18, 32'sd1, -32'sd141, 32'sd0, 32'sd45, -32'sd4, -32'sd19, -32'sd317, -32'sd56, 32'sd90, 32'sd79, -32'sd3, -32'sd138, -32'sd91, 32'sd4, 32'sd22, 32'sd2, 32'sd144, 32'sd22, -32'sd23, -32'sd31, 32'sd0, 32'sd33, 32'sd33, 32'sd75, -32'sd28, 32'sd20, -32'sd145, 32'sd159, -32'sd24, 
                                                    32'sd16, 32'sd1, -32'sd15, -32'sd7, -32'sd5, -32'sd138, 32'sd0, -32'sd108, -32'sd102, -32'sd27, 32'sd55, 32'sd0, 32'sd29, -32'sd49, -32'sd102, 32'sd52, 32'sd102, 32'sd15, 32'sd160, 32'sd99, 32'sd20, -32'sd236, -32'sd20, 32'sd0, 32'sd22, 32'sd1, 32'sd32, -32'sd235, -32'sd49, 32'sd3, -32'sd2, -32'sd36, -32'sd180, 32'sd102, -32'sd11, -32'sd28, -32'sd165, 32'sd70, -32'sd21, 32'sd68, -32'sd22, 32'sd5, -32'sd132, 32'sd41, -32'sd209, -32'sd26, -32'sd86, 32'sd116, -32'sd164, 32'sd97, 32'sd29, 32'sd40, -32'sd49, 32'sd35, -32'sd155, -32'sd40, -32'sd26, 32'sd26, 32'sd5, 32'sd20, 32'sd151, 32'sd42, 32'sd53, 32'sd23, -32'sd57, -32'sd14, -32'sd5, -32'sd6, -32'sd26, -32'sd145, 32'sd2, 32'sd29, 32'sd5, -32'sd143, -32'sd19, -32'sd507, -32'sd126, -32'sd96, 32'sd39, 32'sd67, -32'sd1, 32'sd30, 32'sd10, -32'sd86, -32'sd27, -32'sd134, 32'sd0, 32'sd79, -32'sd109, -32'sd65, -32'sd163, 32'sd348, 32'sd20, 32'sd18, 32'sd44, 32'sd62, -32'sd257, -32'sd14, -32'sd149, 32'sd18, 32'sd79, -32'sd96, 32'sd128, -32'sd4, -32'sd24, 32'sd37, 32'sd76, 32'sd23, -32'sd27, 32'sd77, -32'sd3, 32'sd73, -32'sd35, 32'sd32, -32'sd26, -32'sd97, -32'sd33, -32'sd37, 32'sd4, -32'sd34, -32'sd147, 32'sd38, -32'sd170, 32'sd90, -32'sd58, -32'sd8, 32'sd56, 32'sd90, 32'sd31, 32'sd15, -32'sd140, 32'sd10, 32'sd15, 32'sd21, -32'sd109, 32'sd54, -32'sd83, 32'sd20, -32'sd44, 32'sd101, -32'sd29, -32'sd1, -32'sd8, 32'sd26, -32'sd29, 32'sd32, 32'sd93, 32'sd37, -32'sd143, 32'sd85, -32'sd34, 32'sd24, -32'sd141, -32'sd375, -32'sd35, -32'sd80, -32'sd47, 32'sd25, -32'sd249, 32'sd24, -32'sd20, 32'sd14, 32'sd3, 32'sd126, -32'sd6, -32'sd151, -32'sd120, -32'sd192, 32'sd200, -32'sd87, 32'sd14, 32'sd4, -32'sd22, 32'sd17, -32'sd67, 32'sd17, 32'sd62, 32'sd1, 32'sd69, -32'sd3, 32'sd64, -32'sd28, 32'sd2, 32'sd9, -32'sd1, -32'sd37, -32'sd286, 32'sd52, -32'sd26, 32'sd35, 32'sd11, -32'sd140, -32'sd19, -32'sd54, -32'sd26, 32'sd4, -32'sd28, 32'sd18, -32'sd2, 32'sd16, -32'sd81, -32'sd60, 32'sd250, -32'sd271, 32'sd63, 32'sd98, 32'sd51, -32'sd81, -32'sd74, -32'sd88, 32'sd35, 32'sd31, 32'sd35, 32'sd15, 32'sd31, -32'sd85, 32'sd54, -32'sd24, -32'sd117, 32'sd50, 32'sd57, 32'sd0, 32'sd22, -32'sd103, 32'sd23, -32'sd27, 32'sd28, -32'sd24, 32'sd19, -32'sd30, 32'sd28, -32'sd77, 32'sd20, 32'sd2, -32'sd12, -32'sd179, -32'sd63, -32'sd2, 32'sd0, -32'sd38, 32'sd26, 32'sd6, 32'sd19, -32'sd34, 32'sd133, -32'sd151, -32'sd7, -32'sd31, 32'sd22, -32'sd137, -32'sd171, 32'sd58, -32'sd48, 32'sd2, 32'sd30, -32'sd41, -32'sd131, -32'sd22, 32'sd31, -32'sd27, 32'sd22, -32'sd4, 32'sd129, -32'sd77, 32'sd48, -32'sd92, 32'sd41, -32'sd99, -32'sd8, 32'sd74, 32'sd16, -32'sd7, -32'sd81, -32'sd23, -32'sd272, 32'sd11, 32'sd2, -32'sd141, -32'sd49, -32'sd22, -32'sd49, 32'sd45, -32'sd117, -32'sd3, 32'sd0, 32'sd44, 32'sd45, 32'sd5, -32'sd7, -32'sd41, 32'sd1280, 32'sd43, 32'sd23, 32'sd21, -32'sd197, -32'sd128, 32'sd2, -32'sd26, 32'sd139, 32'sd25, 32'sd9, -32'sd108, 32'sd47, -32'sd35, 32'sd14, -32'sd30, 32'sd22, -32'sd107, -32'sd22, -32'sd19, 32'sd2, -32'sd97, 32'sd98, -32'sd1, 32'sd28, -32'sd46, 32'sd33, 32'sd4, -32'sd86, -32'sd19, 32'sd27, 32'sd6, 32'sd17, 32'sd51, -32'sd91, -32'sd37, 32'sd0, -32'sd1, -32'sd151, -32'sd238, 32'sd50, -32'sd142, 32'sd126, -32'sd89, 32'sd9, -32'sd320, 32'sd19, -32'sd274, 32'sd100, -32'sd92, -32'sd175, 32'sd93, 32'sd25, -32'sd5, 32'sd0, -32'sd233, 32'sd27, -32'sd181, -32'sd15, 32'sd33, 32'sd22, -32'sd78, 32'sd39, -32'sd29, 32'sd27, 32'sd9, 32'sd67, -32'sd63, 32'sd10, 32'sd64, -32'sd75, 32'sd77, 32'sd28, 32'sd78, 32'sd65, 32'sd53, 32'sd12, 32'sd30, 32'sd23, 32'sd5, -32'sd105, 32'sd29, -32'sd25, 32'sd103, 32'sd3, -32'sd10, 32'sd54, 32'sd20, 32'sd1, -32'sd116, -32'sd33, 32'sd34, 32'sd13, 32'sd29, -32'sd34, 32'sd18, -32'sd93, 32'sd66, -32'sd139, 32'sd19, 32'sd4, 32'sd32, 32'sd60, 32'sd17, -32'sd31, -32'sd79, 32'sd4, 32'sd22, -32'sd35, 32'sd31, 32'sd18, -32'sd31, -32'sd121, 32'sd12, -32'sd110, 32'sd49, 32'sd4, 32'sd6, -32'sd31, 32'sd32, -32'sd30, -32'sd26, -32'sd5, 32'sd77, 32'sd115, -32'sd35, 32'sd3, 32'sd82, -32'sd30, 32'sd4, 32'sd4, 32'sd21, -32'sd254, 32'sd49, -32'sd118, 32'sd29, 32'sd69, -32'sd16, 32'sd41, -32'sd78, -32'sd4, 32'sd4, -32'sd6, 32'sd1, -32'sd19, 32'sd22, 32'sd61, -32'sd45, -32'sd5, 32'sd20, -32'sd26, 32'sd11, -32'sd1, 32'sd18, 32'sd1, 32'sd19, -32'sd58, 32'sd36, 32'sd86, 32'sd12, 32'sd43, 32'sd18, -32'sd87, 32'sd69, 32'sd101, -32'sd61, -32'sd78, 32'sd53, 32'sd95, -32'sd17, 32'sd79, 32'sd19, -32'sd140, 32'sd29, 32'sd7, -32'sd27, 32'sd79, 32'sd32, 32'sd5, 32'sd0, -32'sd43, 32'sd1, 32'sd62, -32'sd22, 32'sd1, 32'sd41, -32'sd22, -32'sd1, 32'sd61, -32'sd34, -32'sd131, 32'sd73, -32'sd54, 32'sd369, 32'sd267, 32'sd18, 32'sd69, -32'sd200, -32'sd19, 32'sd17, -32'sd7, 32'sd74, 32'sd3, 32'sd48, -32'sd29, -32'sd52, -32'sd217, -32'sd59, 32'sd20, 32'sd4, -32'sd24, -32'sd61, -32'sd34, 32'sd7, -32'sd17, -32'sd87, -32'sd94, 32'sd39, -32'sd4, 32'sd42, 32'sd56, -32'sd609, -32'sd8, -32'sd4, -32'sd98, -32'sd11, -32'sd3, -32'sd285, -32'sd31, 32'sd16, -32'sd25, 32'sd18, 32'sd4, -32'sd18, -32'sd6, -32'sd9, -32'sd5, 32'sd105, -32'sd24, 32'sd78, 32'sd56, 32'sd70, 32'sd59, -32'sd126, 32'sd91, -32'sd28, 32'sd32, -32'sd138, 32'sd66, -32'sd159, 32'sd26, -32'sd45, 32'sd26, 32'sd3, 32'sd70, 32'sd34, -32'sd131, -32'sd112, 32'sd103, 32'sd29, 32'sd18, -32'sd245, -32'sd42, 32'sd0, 32'sd21, 32'sd107, -32'sd9, -32'sd148, 32'sd19, 32'sd65, 32'sd37, -32'sd114, -32'sd6, -32'sd3, 32'sd124, -32'sd22, 32'sd35, -32'sd228, -32'sd3, -32'sd90, 32'sd42, -32'sd39, 32'sd74, 32'sd6, 32'sd24, -32'sd88, 32'sd20, -32'sd77, 32'sd48, 32'sd66, 32'sd18, 32'sd151, 32'sd117, -32'sd7, -32'sd128, -32'sd1, -32'sd216, -32'sd20, -32'sd24, -32'sd2, -32'sd33, -32'sd40, 32'sd54, 32'sd119, 32'sd52, -32'sd127, 32'sd33, 32'sd15, -32'sd132, 32'sd4, 32'sd0, 
                                                    -32'sd44, 32'sd19, 32'sd4, 32'sd24, 32'sd10, 32'sd29, 32'sd8, 32'sd28, -32'sd56, 32'sd49, 32'sd51, -32'sd34, -32'sd9, 32'sd20, 32'sd99, -32'sd77, -32'sd79, -32'sd91, -32'sd9, 32'sd11, 32'sd35, -32'sd8, -32'sd8, 32'sd65, 32'sd39, -32'sd64, 32'sd50, 32'sd26, -32'sd68, -32'sd80, 32'sd182, 32'sd20, -32'sd21, 32'sd19, 32'sd54, 32'sd19, 32'sd34, 32'sd55, 32'sd89, -32'sd43, -32'sd173, -32'sd8, -32'sd5, 32'sd30, -32'sd27, 32'sd27, -32'sd1, 32'sd6, -32'sd30, 32'sd35, 32'sd10, -32'sd3, -32'sd5, 32'sd64, 32'sd34, 32'sd41, -32'sd18, -32'sd4, -32'sd2, 32'sd6, 32'sd41, 32'sd22, -32'sd19, 32'sd16, -32'sd3, 32'sd21, 32'sd144, 32'sd5, -32'sd26, 32'sd69, 32'sd0, 32'sd54, 32'sd16, 32'sd28, -32'sd53, 32'sd14, -32'sd38, 32'sd32, -32'sd30, 32'sd20, -32'sd7, -32'sd298, -32'sd1, -32'sd86, -32'sd162, 32'sd2, -32'sd3, -32'sd4, -32'sd18, 32'sd48, -32'sd434, 32'sd2, -32'sd23, -32'sd40, 32'sd42, -32'sd23, -32'sd145, 32'sd9, -32'sd2, -32'sd24, -32'sd2, 32'sd2, -32'sd53, 32'sd15, -32'sd25, -32'sd3, -32'sd3, 32'sd8, 32'sd0, 32'sd63, 32'sd65, -32'sd21, -32'sd145, 32'sd11, -32'sd19, 32'sd110, 32'sd43, 32'sd15, -32'sd31, -32'sd38, 32'sd0, -32'sd18, -32'sd36, -32'sd36, 32'sd78, -32'sd53, 32'sd38, 32'sd18, -32'sd88, 32'sd16, -32'sd131, 32'sd27, 32'sd62, 32'sd40, -32'sd38, -32'sd128, 32'sd3, -32'sd4, -32'sd34, -32'sd48, 32'sd53, 32'sd17, 32'sd0, -32'sd27, -32'sd1, -32'sd7, -32'sd94, 32'sd21, -32'sd119, 32'sd32, 32'sd9, 32'sd21, -32'sd3, -32'sd20, 32'sd94, 32'sd23, -32'sd2, -32'sd5, 32'sd54, -32'sd126, 32'sd27, 32'sd38, -32'sd31, 32'sd18, -32'sd26, 32'sd51, -32'sd7, 32'sd159, 32'sd77, 32'sd20, -32'sd58, 32'sd29, -32'sd31, 32'sd5, 32'sd18, 32'sd11, -32'sd4, 32'sd7, -32'sd43, -32'sd52, -32'sd105, -32'sd42, 32'sd6, 32'sd28, -32'sd28, 32'sd23, -32'sd112, 32'sd3, 32'sd7, 32'sd44, -32'sd84, 32'sd75, -32'sd41, -32'sd30, -32'sd206, 32'sd19, 32'sd2, 32'sd71, -32'sd48, -32'sd55, 32'sd6, 32'sd6, -32'sd23, -32'sd38, -32'sd6, 32'sd24, -32'sd23, -32'sd8, -32'sd8, -32'sd181, -32'sd7, 32'sd57, -32'sd24, 32'sd104, 32'sd0, 32'sd7, -32'sd26, 32'sd29, -32'sd33, 32'sd17, 32'sd2, 32'sd18, -32'sd72, -32'sd38, 32'sd2, 32'sd0, -32'sd5, -32'sd32, -32'sd23, 32'sd19, 32'sd44, -32'sd129, 32'sd11, 32'sd8, 32'sd11, 32'sd15, 32'sd243, 32'sd33, 32'sd6, -32'sd5, -32'sd9, 32'sd110, -32'sd20, -32'sd327, -32'sd91, 32'sd211, -32'sd22, -32'sd10, 32'sd13, 32'sd34, -32'sd109, -32'sd72, 32'sd124, -32'sd141, 32'sd105, 32'sd37, -32'sd100, 32'sd26, 32'sd8, -32'sd23, 32'sd142, 32'sd89, -32'sd32, 32'sd15, -32'sd7, 32'sd6, -32'sd44, 32'sd15, -32'sd56, -32'sd93, -32'sd23, 32'sd5, -32'sd27, 32'sd36, 32'sd70, -32'sd14, -32'sd21, -32'sd101, 32'sd85, 32'sd21, -32'sd20, -32'sd575, 32'sd2, 32'sd17, -32'sd94, 32'sd18, 32'sd10, 32'sd54, 32'sd83, 32'sd18, -32'sd300, 32'sd11, -32'sd7, 32'sd94, 32'sd89, -32'sd26, -32'sd23, 32'sd24, 32'sd420, 32'sd30, 32'sd38, -32'sd17, -32'sd37, -32'sd87, -32'sd2, 32'sd139, 32'sd25, -32'sd73, 32'sd18, -32'sd71, -32'sd29, 32'sd25, -32'sd44, 32'sd12, 32'sd0, 32'sd3, -32'sd6, -32'sd66, -32'sd153, 32'sd5, 32'sd63, 32'sd51, 32'sd88, 32'sd33, 32'sd40, -32'sd35, -32'sd35, -32'sd113, -32'sd70, 32'sd3, 32'sd27, -32'sd87, 32'sd30, -32'sd27, 32'sd86, -32'sd103, 32'sd2, 32'sd60, -32'sd8, -32'sd130, 32'sd1, 32'sd0, 32'sd32, -32'sd120, 32'sd1, -32'sd46, -32'sd209, -32'sd217, 32'sd66, 32'sd122, -32'sd148, -32'sd42, 32'sd0, -32'sd99, 32'sd95, -32'sd24, 32'sd4, -32'sd164, 32'sd85, -32'sd3, 32'sd30, 32'sd110, 32'sd4, -32'sd124, 32'sd66, -32'sd23, 32'sd41, -32'sd8, 32'sd3, -32'sd37, 32'sd30, -32'sd33, 32'sd8, 32'sd210, -32'sd57, -32'sd30, 32'sd103, -32'sd42, -32'sd182, 32'sd75, 32'sd50, -32'sd20, 32'sd1, -32'sd4, 32'sd21, 32'sd70, -32'sd2, 32'sd97, -32'sd95, 32'sd197, 32'sd26, 32'sd7, 32'sd38, -32'sd36, 32'sd11, 32'sd32, 32'sd2, -32'sd32, 32'sd11, -32'sd52, 32'sd22, -32'sd5, -32'sd103, -32'sd22, -32'sd252, -32'sd132, 32'sd16, 32'sd95, -32'sd57, -32'sd22, -32'sd16, -32'sd43, 32'sd19, -32'sd4, 32'sd42, -32'sd107, 32'sd23, 32'sd9, -32'sd48, -32'sd27, 32'sd58, 32'sd10, -32'sd36, -32'sd71, -32'sd27, 32'sd9, 32'sd97, -32'sd41, -32'sd146, 32'sd24, 32'sd21, -32'sd3, 32'sd68, -32'sd36, 32'sd8, 32'sd65, -32'sd186, 32'sd3, 32'sd15, -32'sd131, 32'sd24, -32'sd106, 32'sd18, 32'sd61, -32'sd78, 32'sd15, 32'sd8, -32'sd18, 32'sd8, -32'sd69, 32'sd50, -32'sd69, 32'sd5, 32'sd293, -32'sd77, 32'sd48, 32'sd6, -32'sd9, -32'sd6, -32'sd102, -32'sd81, -32'sd5, -32'sd202, -32'sd6, -32'sd4, 32'sd22, 32'sd21, 32'sd72, 32'sd15, 32'sd119, -32'sd21, 32'sd130, 32'sd4, -32'sd1, -32'sd15, -32'sd9, -32'sd86, -32'sd95, -32'sd3, -32'sd27, 32'sd18, -32'sd9, -32'sd290, -32'sd19, 32'sd53, -32'sd53, 32'sd8, 32'sd59, -32'sd169, 32'sd25, 32'sd10, 32'sd59, -32'sd64, -32'sd197, 32'sd15, -32'sd188, -32'sd14, 32'sd73, 32'sd12, 32'sd111, 32'sd7, -32'sd36, 32'sd38, 32'sd78, 32'sd50, 32'sd75, 32'sd82, -32'sd19, -32'sd37, 32'sd67, -32'sd114, 32'sd57, 32'sd23, -32'sd38, 32'sd205, -32'sd68, -32'sd54, 32'sd17, 32'sd126, -32'sd72, -32'sd1, 32'sd17, 32'sd12, -32'sd5, -32'sd4, 32'sd29, -32'sd4, 32'sd16, 32'sd33, 32'sd20, 32'sd0, -32'sd71, -32'sd22, 32'sd5, -32'sd2, -32'sd2, 32'sd18, 32'sd30, -32'sd166, -32'sd24, -32'sd25, -32'sd42, -32'sd1, 32'sd76, -32'sd30, 32'sd94, 32'sd140, 32'sd22, 32'sd129, -32'sd7, -32'sd120, 32'sd70, 32'sd52, 32'sd4, -32'sd45, 32'sd22, -32'sd26, -32'sd63, -32'sd2, -32'sd21, -32'sd53, 32'sd91, -32'sd39, 32'sd3, -32'sd21, 32'sd26, 32'sd1, 32'sd112, -32'sd22, -32'sd78, -32'sd25, 32'sd21, -32'sd98, -32'sd15, -32'sd5, 32'sd24, 32'sd1, 32'sd16, -32'sd25, 32'sd31, -32'sd50, -32'sd3840, -32'sd8, -32'sd90, 32'sd8, 32'sd0, -32'sd18, 32'sd0, -32'sd2, -32'sd54, -32'sd26, 32'sd23, 32'sd4, 32'sd39, -32'sd34, 32'sd9, -32'sd110, -32'sd6, -32'sd58, -32'sd60, -32'sd6, 32'sd37, -32'sd1, -32'sd451, 32'sd188, -32'sd167, -32'sd1, 32'sd11, 
                                                    -32'sd22, 32'sd32, -32'sd31, 32'sd26, -32'sd136, 32'sd64, 32'sd53, 32'sd17, 32'sd75, -32'sd403, 32'sd89, 32'sd39, -32'sd41, 32'sd7, 32'sd118, 32'sd26, 32'sd3, 32'sd17, -32'sd25, 32'sd20, -32'sd71, -32'sd6, -32'sd121, -32'sd1, -32'sd3, 32'sd14, 32'sd1, -32'sd11, 32'sd145, 32'sd98, -32'sd8, 32'sd12, 32'sd11, -32'sd141, -32'sd26, 32'sd18, -32'sd158, 32'sd2, -32'sd41, 32'sd29, 32'sd65, 32'sd9, 32'sd20, -32'sd23, 32'sd7, -32'sd9, -32'sd25, -32'sd110, -32'sd145, 32'sd20, -32'sd79, 32'sd89, -32'sd19, 32'sd22, 32'sd79, 32'sd54, 32'sd160, 32'sd18, 32'sd76, -32'sd101, -32'sd182, 32'sd4, -32'sd29, 32'sd41, 32'sd83, 32'sd14, 32'sd3, 32'sd4, -32'sd33, 32'sd116, 32'sd1, -32'sd123, 32'sd175, 32'sd28, -32'sd113, 32'sd8, -32'sd19, 32'sd16, -32'sd8, 32'sd14, 32'sd47, 32'sd35, 32'sd138, 32'sd26, 32'sd3, 32'sd7, 32'sd27, -32'sd200, 32'sd67, -32'sd168, -32'sd65, 32'sd8, 32'sd394, 32'sd50, 32'sd58, 32'sd55, -32'sd85, 32'sd36, 32'sd57, -32'sd32, 32'sd44, 32'sd4, -32'sd8, -32'sd31, -32'sd62, 32'sd92, -32'sd44, -32'sd105, 32'sd24, -32'sd4, -32'sd69, -32'sd5, 32'sd20, -32'sd28, 32'sd78, -32'sd2, -32'sd35, -32'sd5, -32'sd7, -32'sd70, 32'sd62, -32'sd42, 32'sd16, 32'sd69, 32'sd6, 32'sd53, 32'sd88, -32'sd29, -32'sd28, -32'sd93, 32'sd24, -32'sd59, 32'sd31, 32'sd4, 32'sd10, -32'sd24, -32'sd3840, -32'sd6, 32'sd20, -32'sd32, 32'sd24, -32'sd25, 32'sd29, -32'sd85, 32'sd83, 32'sd45, 32'sd27, -32'sd23, 32'sd39, 32'sd128, -32'sd8, -32'sd39, -32'sd120, -32'sd3, 32'sd11, -32'sd40, -32'sd108, -32'sd171, -32'sd78, -32'sd5, 32'sd42, 32'sd38, -32'sd192, -32'sd6, -32'sd19, -32'sd5, 32'sd77, -32'sd5, 32'sd7, -32'sd34, 32'sd46, 32'sd66, 32'sd0, 32'sd79, 32'sd23, -32'sd247, 32'sd79, 32'sd57, 32'sd31, -32'sd19, -32'sd23, -32'sd24, 32'sd29, -32'sd66, 32'sd45, -32'sd28, -32'sd37, 32'sd34, -32'sd64, -32'sd99, -32'sd41, -32'sd29, 32'sd66, 32'sd6, 32'sd1, 32'sd9, -32'sd243, -32'sd183, 32'sd23, -32'sd21, -32'sd36, -32'sd2, -32'sd1, 32'sd325, 32'sd37, 32'sd84, 32'sd35, -32'sd32, 32'sd7, 32'sd60, 32'sd33, 32'sd9, 32'sd22, -32'sd23, 32'sd306, 32'sd80, -32'sd8, 32'sd14, -32'sd117, 32'sd191, 32'sd25, 32'sd0, 32'sd134, 32'sd35, 32'sd7, -32'sd124, -32'sd45, -32'sd7, 32'sd36, 32'sd27, 32'sd15, -32'sd29, -32'sd13, 32'sd10, 32'sd21, -32'sd22, 32'sd16, -32'sd142, -32'sd617, -32'sd82, 32'sd314, -32'sd65, 32'sd14, -32'sd181, 32'sd5, 32'sd43, 32'sd6, 32'sd0, 32'sd46, 32'sd56, -32'sd6, -32'sd118, 32'sd26, -32'sd30, 32'sd34, 32'sd6, -32'sd362, -32'sd20, -32'sd255, 32'sd167, -32'sd6, -32'sd26, -32'sd122, -32'sd271, -32'sd206, 32'sd90, -32'sd51, 32'sd57, -32'sd202, -32'sd5, -32'sd2, 32'sd3, -32'sd8, -32'sd108, 32'sd21, 32'sd1, 32'sd17, -32'sd21, 32'sd71, -32'sd138, 32'sd150, 32'sd49, 32'sd14, -32'sd24, 32'sd24, 32'sd122, 32'sd5, -32'sd8, 32'sd54, -32'sd27, -32'sd272, -32'sd190, 32'sd41, 32'sd24, 32'sd36, 32'sd34, -32'sd78, 32'sd3, 32'sd62, -32'sd119, 32'sd44, -32'sd8, 32'sd82, -32'sd51, -32'sd59, 32'sd28, 32'sd54, -32'sd81, -32'sd39, 32'sd52, -32'sd100, 32'sd21, -32'sd102, 32'sd33, -32'sd91, 32'sd95, -32'sd31, -32'sd17, 32'sd18, 32'sd115, -32'sd110, 32'sd109, -32'sd38, 32'sd25, -32'sd33, 32'sd28, -32'sd6, 32'sd24, 32'sd40, 32'sd21, -32'sd80, 32'sd25, -32'sd2, -32'sd4, 32'sd27, 32'sd24, 32'sd7, 32'sd25, 32'sd122, 32'sd32, -32'sd210, -32'sd12, -32'sd46, 32'sd26, -32'sd24, 32'sd105, -32'sd59, 32'sd18, -32'sd26, 32'sd7, -32'sd28, 32'sd18, 32'sd229, -32'sd242, -32'sd7, -32'sd13, -32'sd6, -32'sd12, -32'sd183, 32'sd41, -32'sd4, -32'sd2, 32'sd140, 32'sd40, -32'sd88, -32'sd1, 32'sd16, 32'sd50, -32'sd26, 32'sd116, -32'sd25, -32'sd66, -32'sd4, 32'sd16, -32'sd81, 32'sd8, 32'sd40, 32'sd22, 32'sd45, -32'sd95, 32'sd53, 32'sd0, -32'sd21, -32'sd67, 32'sd0, 32'sd8, 32'sd19, 32'sd17, -32'sd175, -32'sd1, -32'sd40, 32'sd11, -32'sd23, 32'sd18, -32'sd30, -32'sd3, -32'sd3, 32'sd59, 32'sd51, 32'sd4, 32'sd56, 32'sd9, -32'sd27, 32'sd46, -32'sd20, 32'sd36, -32'sd47, 32'sd53, -32'sd22, -32'sd84, -32'sd59, 32'sd9, -32'sd129, 32'sd54, 32'sd34, -32'sd133, -32'sd3, 32'sd200, 32'sd19, 32'sd0, -32'sd5, -32'sd112, 32'sd76, -32'sd7, -32'sd174, 32'sd33, -32'sd18, 32'sd22, 32'sd37, 32'sd26, -32'sd20, 32'sd10, 32'sd10, -32'sd47, -32'sd118, 32'sd10, 32'sd92, -32'sd112, -32'sd76, 32'sd62, 32'sd43, 32'sd40, 32'sd23, -32'sd38, -32'sd18, 32'sd71, -32'sd8, 32'sd25, 32'sd38, 32'sd86, 32'sd0, 32'sd15, -32'sd65, -32'sd28, -32'sd19, 32'sd51, 32'sd15, 32'sd11, -32'sd24, 32'sd20, -32'sd137, 32'sd7, -32'sd8, 32'sd85, 32'sd8, -32'sd32, 32'sd51, -32'sd12, -32'sd59, 32'sd19, 32'sd202, 32'sd10, 32'sd60, 32'sd15, -32'sd107, 32'sd10, -32'sd23, 32'sd16, 32'sd35, -32'sd55, 32'sd75, -32'sd5, -32'sd3, 32'sd18, -32'sd53, 32'sd27, 32'sd81, -32'sd66, -32'sd23, 32'sd88, -32'sd20, -32'sd31, -32'sd113, 32'sd23, -32'sd21, 32'sd44, 32'sd111, 32'sd15, -32'sd115, -32'sd139, -32'sd4, 32'sd28, 32'sd215, 32'sd0}

localparam logic [2912:0][31:0] feature_below = {32'sd267, -32'sd239, -32'sd193, -32'sd112, -32'sd100, 32'sd71, -32'sd216, -32'sd189, -32'sd110, 32'sd159, -32'sd207, -32'sd249, -32'sd71, 32'sd34, -32'sd342, -32'sd139, -32'sd45, 32'sd119, 32'sd148, -32'sd54, 32'sd187, 32'sd143, -32'sd45, -32'sd78, 32'sd50, -32'sd130, -32'sd211, 32'sd59, -32'sd84, -32'sd179, -32'sd65, 32'sd47, -32'sd39, -32'sd52, 32'sd135, -32'sd208, 32'sd36, -32'sd130, -32'sd21, 32'sd194, 32'sd226, -32'sd40, -32'sd13, -32'sd52, 32'sd22, 32'sd114, -32'sd48, 32'sd8, -32'sd224, -32'sd120, -32'sd7, -32'sd234, 32'sd148, -32'sd200, -32'sd74, -32'sd187, -32'sd107, -32'sd40, -32'sd56, 32'sd191, -32'sd123, -32'sd313, 32'sd22, 32'sd62, 32'sd23, -32'sd251, 32'sd127, -32'sd330, 32'sd184, -32'sd63, -32'sd298, -32'sd108, -32'sd185, 32'sd23, 32'sd9, 32'sd50, 32'sd19, 32'sd32, -32'sd97, -32'sd47, -32'sd297, 32'sd54, 32'sd142, -32'sd426, -32'sd156, -32'sd62, -32'sd138, -32'sd154, -32'sd56, -32'sd24, 32'sd39, 32'sd160, -32'sd76, 32'sd36, 32'sd62, 32'sd34, -32'sd168, 32'sd58, -32'sd222, -32'sd25, -32'sd206, 32'sd95, -32'sd34, -32'sd8, -32'sd45, -32'sd134, 32'sd106, 32'sd26, 32'sd26, -32'sd166, -32'sd168, -32'sd135, -32'sd176, -32'sd5, -32'sd128, 32'sd185, -32'sd48, -32'sd74, 32'sd2, -32'sd10, -32'sd147, 32'sd48, 32'sd34, 32'sd97, 32'sd29, -32'sd162, 32'sd111, -32'sd178, 32'sd8, -32'sd69, -32'sd45, -32'sd75, -32'sd43, 32'sd89, 32'sd110, 32'sd25, -32'sd114, -32'sd161, -32'sd110, -32'sd96, -32'sd162, -32'sd126, 32'sd82, -32'sd31, -32'sd44, 32'sd141, 32'sd201, -32'sd35, -32'sd140, 32'sd39, 32'sd33, -32'sd158, 32'sd52, -32'sd12, -32'sd53, 32'sd32, -32'sd120, 32'sd159, -32'sd42, 32'sd45, 32'sd7, -32'sd131, 32'sd132, 32'sd28, -32'sd204, -32'sd132, -32'sd189, -32'sd31, 32'sd37, -32'sd30, -32'sd155, 32'sd31, -32'sd175, 32'sd27, 32'sd42, -32'sd36, -32'sd296, 32'sd37, -32'sd35, -32'sd196, 32'sd10, 32'sd18, -32'sd141, 32'sd2, -32'sd44, 32'sd26, -32'sd52, -32'sd285, -32'sd37, -32'sd114, -32'sd143, -32'sd129, 32'sd33, -32'sd73, -32'sd71, -32'sd165, 32'sd223, -32'sd135, 32'sd73, 32'sd167, -32'sd59, -32'sd53, 32'sd46, -32'sd114, 32'sd38, -32'sd102, 32'sd20, 32'sd4, -32'sd50, 32'sd11, 32'sd71, -32'sd237, -32'sd62, -32'sd58, -32'sd108, 32'sd45, 32'sd24, -32'sd160, -32'sd104, -32'sd119, 32'sd72, 32'sd103, -32'sd109, -32'sd52, -32'sd196, 32'sd81, 32'sd75, -32'sd33, 32'sd37, -32'sd51, 32'sd27, 32'sd56, 32'sd120, 32'sd1, -32'sd130, -32'sd48, -32'sd103, -32'sd135, 32'sd26, -32'sd49, 32'sd27, -32'sd131, -32'sd132, -32'sd27, 32'sd113, 32'sd134, 32'sd18, -32'sd213, 32'sd102, -32'sd123, 32'sd25, -32'sd133, -32'sd158, -32'sd97, -32'sd50, -32'sd92, 32'sd71, -32'sd57, -32'sd140, 32'sd107, -32'sd33, 32'sd40, -32'sd134, 32'sd21, -32'sd88, 32'sd32, -32'sd65, 32'sd5, 32'sd18, -32'sd115, -32'sd58, 32'sd43, -32'sd101, -32'sd292, 32'sd50, 32'sd4, -32'sd139, -32'sd241, 32'sd19, -32'sd130, 32'sd20, -32'sd99, -32'sd15, 32'sd9, -32'sd225, 32'sd123, 32'sd60, 32'sd91, -32'sd141, -32'sd140, -32'sd34, -32'sd28, 32'sd24, -32'sd119, 32'sd251, 32'sd27, -32'sd150, -32'sd144, -32'sd22, 32'sd106, -32'sd148, -32'sd134, -32'sd140, 32'sd54, -32'sd118, -32'sd204, -32'sd85, 32'sd25, -32'sd81, -32'sd24, -32'sd14, -32'sd138, 32'sd44, 32'sd61, 32'sd125, -32'sd278, -32'sd82, -32'sd189, 32'sd54, 32'sd3, 32'sd20, -32'sd52, -32'sd255, -32'sd80, 32'sd130, -32'sd131, -32'sd146, -32'sd73, 32'sd39, -32'sd220, 32'sd30, -32'sd156, 32'sd42, -32'sd41, -32'sd14, 32'sd51, 32'sd0, 32'sd96, -32'sd106, -32'sd76, 32'sd20, 32'sd4, -32'sd67, -32'sd68, 32'sd26, 32'sd6, -32'sd117, 32'sd12, 32'sd27, -32'sd35, -32'sd13, 32'sd8, -32'sd119, 32'sd17, 32'sd25, -32'sd146, 32'sd22, -32'sd61, -32'sd277, 32'sd6, -32'sd4, -32'sd169, 32'sd47, -32'sd33, -32'sd10, -32'sd101, 32'sd218, 32'sd99, -32'sd191, -32'sd273, 32'sd73, 32'sd87, 32'sd32, 32'sd2, -32'sd1, 32'sd58, -32'sd122, -32'sd258, 32'sd51, -32'sd32, -32'sd7, 32'sd6, -32'sd63, -32'sd38, -32'sd77, -32'sd4, 32'sd48, -32'sd128, 32'sd18, -32'sd27, -32'sd169, 32'sd63, 32'sd54, -32'sd4, -32'sd101, -32'sd288, -32'sd33, -32'sd29, -32'sd37, -32'sd4, 32'sd76, -32'sd61, 32'sd29, -32'sd33, -32'sd77, 32'sd91, -32'sd72, -32'sd91, -32'sd143, -32'sd52, -32'sd49, -32'sd90, -32'sd70, -32'sd13, 32'sd108, 32'sd34, 32'sd20, -32'sd255, -32'sd41, 32'sd76, 32'sd3, -32'sd56, -32'sd114, 32'sd27, 32'sd2, 32'sd129, -32'sd188, -32'sd104, 32'sd15, 32'sd17, -32'sd151, 32'sd81, 32'sd24, -32'sd119, 32'sd5, 32'sd47, 32'sd25, -32'sd215, -32'sd394, 32'sd27, -32'sd147, 32'sd107, -32'sd36, 32'sd23, 32'sd123, 32'sd1, -32'sd68, 32'sd105, -32'sd25, -32'sd3, -32'sd174, -32'sd83, 32'sd108, 32'sd25, -32'sd93, -32'sd46, 32'sd7, 32'sd60, -32'sd145, 32'sd126, -32'sd36, -32'sd82, 32'sd48, -32'sd167, -32'sd262, 32'sd99, 32'sd22, -32'sd192, 32'sd37, 32'sd177, -32'sd29, -32'sd203, -32'sd153, -32'sd20, 32'sd33, -32'sd11, 32'sd96, 32'sd16, -32'sd47, -32'sd10, 32'sd100, -32'sd115, 32'sd106, 32'sd2, 32'sd145, -32'sd74, -32'sd3, -32'sd70, -32'sd157, 32'sd19, -32'sd36, -32'sd31, -32'sd110, 32'sd89, -32'sd21, 32'sd56, -32'sd125, -32'sd116, -32'sd101, -32'sd39, -32'sd115, -32'sd54, 32'sd59, 32'sd117, -32'sd188, -32'sd134, 32'sd37, -32'sd165, -32'sd110, 32'sd21, 32'sd20, 32'sd3, -32'sd21, -32'sd125, 32'sd126, 32'sd61, -32'sd123, -32'sd67, 32'sd22, -32'sd145, 32'sd33, 32'sd25, -32'sd7, 32'sd136, -32'sd24, -32'sd4, 32'sd128, -32'sd4, 32'sd0, -32'sd196, 32'sd4, 32'sd98, 32'sd21, -32'sd125, 32'sd59, 32'sd33, -32'sd103, -32'sd168, 32'sd26, 32'sd125, -32'sd24, -32'sd87, 32'sd24, -32'sd30, 32'sd32, -32'sd133, 32'sd66, 32'sd207, 32'sd382, 32'sd77, -32'sd79, 32'sd85, -32'sd144, -32'sd138, 32'sd104, -32'sd3, 32'sd87, 32'sd7, -32'sd17, -32'sd48, -32'sd75, -32'sd39, 32'sd76, 32'sd124, 32'sd117, -32'sd77, 32'sd6, -32'sd120, 32'sd23, -32'sd165, -32'sd6, -32'sd2, -32'sd34, -32'sd66, 32'sd53, -32'sd32, 
                                                    -32'sd29, 32'sd8, 32'sd24, -32'sd121, 32'sd47, 32'sd123, -32'sd393, 32'sd29, 32'sd0, 32'sd122, -32'sd13, 32'sd1, 32'sd83, -32'sd5, 32'sd89, -32'sd52, -32'sd83, 32'sd125, -32'sd13, 32'sd78, -32'sd130, -32'sd53, -32'sd75, -32'sd119, 32'sd15, -32'sd74, -32'sd49, 32'sd151, -32'sd110, -32'sd96, 32'sd118, 32'sd34, -32'sd36, -32'sd79, 32'sd74, 32'sd42, 32'sd11, 32'sd44, 32'sd30, -32'sd95, -32'sd116, -32'sd44, -32'sd120, -32'sd68, 32'sd118, -32'sd91, -32'sd111, -32'sd29, -32'sd39, 32'sd34, -32'sd151, -32'sd70, -32'sd35, -32'sd117, -32'sd56, 32'sd3, 32'sd101, 32'sd103, -32'sd26, -32'sd6, -32'sd116, 32'sd45, -32'sd25, -32'sd179, 32'sd0, -32'sd63, -32'sd156, 32'sd48, -32'sd38, -32'sd184, -32'sd289, 32'sd48, -32'sd38, -32'sd128, 32'sd6, 32'sd19, -32'sd2, -32'sd18, -32'sd2, -32'sd222, -32'sd31, 32'sd1, 32'sd5, 32'sd10, -32'sd217, 32'sd81, -32'sd43, 32'sd29, 32'sd25, 32'sd12, -32'sd223, -32'sd31, 32'sd151, 32'sd18, -32'sd70, -32'sd28, 32'sd8, 32'sd88, 32'sd223, 32'sd39, -32'sd27, -32'sd102, 32'sd48, -32'sd2, 32'sd155, -32'sd3, -32'sd136, -32'sd4, 32'sd5, -32'sd10, -32'sd246, 32'sd62, -32'sd25, 32'sd25, -32'sd25, 32'sd232, 32'sd100, 32'sd20, -32'sd21, -32'sd13, -32'sd5, -32'sd7, 32'sd36, 32'sd16, 32'sd3, 32'sd24, 32'sd9, 32'sd6, -32'sd35, 32'sd7, 32'sd49, 32'sd20, 32'sd3, 32'sd21, -32'sd79, -32'sd109, -32'sd104, -32'sd47, -32'sd152, 32'sd42, -32'sd65, -32'sd134, -32'sd65, -32'sd127, -32'sd12, 32'sd30, -32'sd13, 32'sd0, -32'sd84, 32'sd36, 32'sd20, -32'sd37, 32'sd175, 32'sd156, -32'sd105, -32'sd156, 32'sd15, -32'sd150, -32'sd137, -32'sd46, 32'sd63, 32'sd75, -32'sd10, 32'sd35, -32'sd1, 32'sd105, 32'sd17, -32'sd116, 32'sd1, 32'sd228, 32'sd73, -32'sd41, 32'sd25, 32'sd9, -32'sd50, -32'sd3, -32'sd246, -32'sd164, -32'sd52, -32'sd93, 32'sd74, 32'sd117, -32'sd66, 32'sd31, 32'sd21, -32'sd175, -32'sd219, -32'sd40, 32'sd19, 32'sd95, -32'sd52, 32'sd104, 32'sd42, -32'sd161, 32'sd177, -32'sd5, -32'sd24, -32'sd57, 32'sd87, -32'sd2, 32'sd43, -32'sd136, 32'sd19, -32'sd31, 32'sd17, -32'sd134, -32'sd194, 32'sd18, 32'sd37, -32'sd35, 32'sd24, 32'sd42, 32'sd15, -32'sd142, 32'sd103, -32'sd34, 32'sd2, 32'sd2, -32'sd39, -32'sd206, 32'sd10, -32'sd1, -32'sd31, 32'sd245, -32'sd32, -32'sd89, 32'sd23, -32'sd4, 32'sd8, 32'sd1, 32'sd19, 32'sd50, -32'sd199, 32'sd28, -32'sd6, -32'sd33, -32'sd23, 32'sd70, -32'sd89, 32'sd38, 32'sd118, -32'sd102, 32'sd42, -32'sd176, 32'sd8, 32'sd46, -32'sd20, 32'sd17, 32'sd14, -32'sd1, 32'sd0, -32'sd60, -32'sd1, -32'sd44, 32'sd192, -32'sd127, -32'sd74, -32'sd4, 32'sd51, 32'sd23, 32'sd70, 32'sd87, -32'sd115, -32'sd72, 32'sd46, -32'sd71, -32'sd137, -32'sd92, -32'sd60, 32'sd27, 32'sd86, -32'sd122, 32'sd104, 32'sd158, -32'sd39, 32'sd27, -32'sd116, 32'sd29, -32'sd51, 32'sd24, 32'sd20, 32'sd28, -32'sd189, -32'sd22, 32'sd5, 32'sd43, 32'sd1, 32'sd58, 32'sd20, -32'sd167, -32'sd31, 32'sd4, -32'sd29, 32'sd26, 32'sd88, -32'sd1, -32'sd26, 32'sd61, -32'sd142, 32'sd130, 32'sd53, 32'sd27, -32'sd148, 32'sd45, -32'sd197, 32'sd26, -32'sd3, 32'sd22, -32'sd153, -32'sd140, 32'sd36, -32'sd6, -32'sd34, 32'sd77, 32'sd49, 32'sd17, 32'sd15, -32'sd44, -32'sd22, 32'sd78, -32'sd62, -32'sd515, -32'sd50, -32'sd11, 32'sd147, -32'sd3, 32'sd5, 32'sd72, -32'sd22, 32'sd162, 32'sd86, -32'sd53, -32'sd117, 32'sd0, -32'sd48, -32'sd54, -32'sd21, 32'sd19, 32'sd176, -32'sd43, 32'sd98, -32'sd89, -32'sd2, -32'sd13, 32'sd137, 32'sd24, -32'sd28, 32'sd33, -32'sd1, -32'sd37, -32'sd5, 32'sd42, -32'sd45, -32'sd184, -32'sd151, 32'sd283, -32'sd239, -32'sd98, -32'sd81, 32'sd109, -32'sd4, -32'sd25, 32'sd264, -32'sd15, -32'sd2, -32'sd5, -32'sd85, -32'sd7, 32'sd78, -32'sd73, 32'sd7, 32'sd22, -32'sd86, 32'sd38, -32'sd36, -32'sd14, -32'sd7, 32'sd58, -32'sd260, 32'sd22, -32'sd3, 32'sd39, -32'sd40, -32'sd230, -32'sd7, 32'sd27, -32'sd26, -32'sd122, -32'sd18, -32'sd140, 32'sd13, 32'sd8, -32'sd172, 32'sd6, -32'sd131, 32'sd11, -32'sd19, 32'sd84, -32'sd116, -32'sd64, -32'sd54, -32'sd61, 32'sd65, -32'sd30, 32'sd52, 32'sd58, -32'sd109, -32'sd119, -32'sd164, 32'sd75, -32'sd7, -32'sd111, -32'sd10, -32'sd32, -32'sd144, -32'sd186, 32'sd69, 32'sd9, 32'sd146, -32'sd32, -32'sd5, 32'sd75, 32'sd20, 32'sd22, -32'sd19, -32'sd51, 32'sd36, 32'sd0, 32'sd53, -32'sd183, -32'sd32, 32'sd6, -32'sd120, -32'sd35, -32'sd132, 32'sd81, 32'sd21, -32'sd32, -32'sd37, -32'sd1, 32'sd14, -32'sd25, 32'sd40, -32'sd1, -32'sd59, -32'sd2, -32'sd10, -32'sd34, 32'sd23, -32'sd24, -32'sd19, -32'sd67, -32'sd49, -32'sd1, -32'sd74, 32'sd3, -32'sd83, -32'sd43, 32'sd19, -32'sd32, -32'sd14, -32'sd125, 32'sd49, -32'sd133, -32'sd705, 32'sd122, 32'sd1, 32'sd29, 32'sd21, -32'sd111, -32'sd361, -32'sd166, -32'sd104, 32'sd84, 32'sd1, 32'sd39, 32'sd33, -32'sd184, -32'sd22, -32'sd83, -32'sd7, -32'sd118, 32'sd69, -32'sd70, 32'sd20, -32'sd31, -32'sd65, -32'sd28, 32'sd15, -32'sd2, 32'sd156, -32'sd32, 32'sd29, 32'sd32, -32'sd42, -32'sd7, 32'sd0, -32'sd39, -32'sd31, 32'sd60, 32'sd49, -32'sd6, 32'sd27, -32'sd22, 32'sd15, -32'sd6, -32'sd52, -32'sd42, -32'sd93, -32'sd20, 32'sd25, 32'sd105, -32'sd55, -32'sd4, 32'sd14, 32'sd279, -32'sd6, -32'sd42, 32'sd147, -32'sd50, -32'sd215, -32'sd125, 32'sd27, -32'sd21, 32'sd30, -32'sd119, -32'sd94, 32'sd18, 32'sd1, -32'sd152, 32'sd311, 32'sd92, 32'sd20, -32'sd104, 32'sd119, -32'sd72, -32'sd101, -32'sd181, 32'sd49, -32'sd52, -32'sd31, -32'sd112, 32'sd20, -32'sd147, 32'sd20, 32'sd5, 32'sd56, 32'sd56, -32'sd12, -32'sd49, 32'sd114, 32'sd110, 32'sd77, -32'sd203, 32'sd22, 32'sd65, -32'sd55, -32'sd40, 32'sd135, -32'sd92, 32'sd32, -32'sd88, -32'sd76, 32'sd6, -32'sd79, -32'sd39, -32'sd176, -32'sd72, 32'sd1, 32'sd200, -32'sd202, -32'sd199, 32'sd22, -32'sd167, -32'sd177, -32'sd91, -32'sd5, 32'sd74, -32'sd63, -32'sd63, -32'sd77, 32'sd30, -32'sd10, -32'sd154, 32'sd30, -32'sd104, 32'sd79, -32'sd38, -32'sd78, 
                                                    -32'sd68, -32'sd165, -32'sd22, -32'sd14, 32'sd131, -32'sd100, -32'sd113, 32'sd15, -32'sd104, -32'sd9, -32'sd165, 32'sd61, -32'sd8, 32'sd22, -32'sd26, -32'sd9, -32'sd163, 32'sd16, 32'sd2, 32'sd79, -32'sd46, 32'sd67, -32'sd22, -32'sd152, 32'sd107, 32'sd45, -32'sd113, -32'sd18, -32'sd37, -32'sd4, 32'sd89, -32'sd83, -32'sd4, -32'sd1, 32'sd109, -32'sd266, -32'sd110, 32'sd49, -32'sd221, 32'sd70, -32'sd5, 32'sd75, -32'sd2, 32'sd19, 32'sd66, -32'sd3, -32'sd110, -32'sd58, 32'sd17, 32'sd17, -32'sd32, 32'sd3, -32'sd50, 32'sd11, -32'sd23, -32'sd79, -32'sd6, 32'sd23, -32'sd108, -32'sd24, -32'sd102, -32'sd30, -32'sd7, 32'sd34, -32'sd86, 32'sd86, 32'sd39, 32'sd19, -32'sd24, 32'sd24, 32'sd58, 32'sd17, -32'sd27, 32'sd41, -32'sd26, 32'sd20, -32'sd80, 32'sd21, -32'sd32, 32'sd20, 32'sd73, 32'sd73, -32'sd49, 32'sd28, -32'sd37, -32'sd83, -32'sd37, 32'sd58, -32'sd66, 32'sd2, 32'sd50, 32'sd152, -32'sd87, -32'sd109, -32'sd141, -32'sd25, -32'sd52, -32'sd38, -32'sd167, 32'sd30, 32'sd37, -32'sd310, 32'sd113, 32'sd103, 32'sd19, -32'sd104, -32'sd91, -32'sd93, 32'sd22, 32'sd354, 32'sd15, -32'sd1, 32'sd30, -32'sd40, -32'sd6, -32'sd149, -32'sd35, -32'sd69, 32'sd23, 32'sd80, 32'sd31, -32'sd120, -32'sd10, 32'sd5, 32'sd22, -32'sd4, 32'sd12, -32'sd51, -32'sd29, -32'sd35, -32'sd14, -32'sd6, 32'sd19, -32'sd3, -32'sd103, -32'sd27, 32'sd26, -32'sd23, 32'sd64, 32'sd150, -32'sd8, -32'sd30, -32'sd105, 32'sd78, -32'sd5, -32'sd147, -32'sd1, 32'sd48, -32'sd13, 32'sd86, 32'sd20, 32'sd49, 32'sd19, -32'sd87, 32'sd33, -32'sd4, -32'sd45, -32'sd5, -32'sd3, 32'sd14, 32'sd60, -32'sd36, -32'sd3, -32'sd42, -32'sd157, -32'sd2, 32'sd84, -32'sd67, -32'sd100, 32'sd0, -32'sd7, 32'sd2, -32'sd80, 32'sd23, 32'sd6, 32'sd58, 32'sd43, -32'sd299, -32'sd85, 32'sd59, -32'sd34, -32'sd24, -32'sd3, -32'sd4, 32'sd1, 32'sd54, -32'sd3, -32'sd4, 32'sd14, 32'sd37, 32'sd15, 32'sd19, -32'sd69, -32'sd8, -32'sd58, 32'sd155, -32'sd295, -32'sd92, 32'sd9, -32'sd157, 32'sd17, -32'sd4, 32'sd17, -32'sd19, 32'sd25, -32'sd48, 32'sd104, 32'sd107, -32'sd121, 32'sd6, -32'sd249, -32'sd27, 32'sd77, -32'sd28, 32'sd81, -32'sd30, 32'sd23, -32'sd89, 32'sd44, -32'sd112, 32'sd30, -32'sd8, -32'sd25, 32'sd124, -32'sd8, -32'sd58, 32'sd15, 32'sd232, 32'sd30, 32'sd63, 32'sd78, 32'sd51, -32'sd109, -32'sd101, -32'sd86, 32'sd5, 32'sd18, -32'sd18, 32'sd18, -32'sd26, -32'sd60, -32'sd121, 32'sd42, 32'sd35, 32'sd30, -32'sd74, -32'sd78, -32'sd72, -32'sd103, -32'sd104, 32'sd18, -32'sd21, 32'sd185, 32'sd17, -32'sd43, -32'sd15, -32'sd127, -32'sd62, 32'sd5, -32'sd139, 32'sd122, -32'sd133, 32'sd115, -32'sd130, 32'sd79, -32'sd11, 32'sd8, -32'sd120, -32'sd108, 32'sd78, -32'sd4, 32'sd17, -32'sd145, 32'sd97, 32'sd38, 32'sd3, -32'sd109, -32'sd8, 32'sd46, 32'sd0, -32'sd4, 32'sd76, 32'sd76, -32'sd150, -32'sd2, 32'sd21, -32'sd29, 32'sd35, -32'sd97, -32'sd29, 32'sd25, 32'sd21, 32'sd164, -32'sd69, 32'sd81, -32'sd64, -32'sd152, 32'sd3, 32'sd4, -32'sd27, 32'sd0, -32'sd28, -32'sd1, 32'sd57, -32'sd26, -32'sd98, -32'sd181, 32'sd25, 32'sd108, 32'sd16, -32'sd60, 32'sd66, -32'sd4, 32'sd31, 32'sd125, 32'sd26, -32'sd33, 32'sd22, -32'sd110, 32'sd72, -32'sd33, 32'sd1, -32'sd77, 32'sd54, 32'sd29, 32'sd12, -32'sd34, -32'sd93, -32'sd45, 32'sd15, -32'sd1, 32'sd26, 32'sd74, 32'sd2, -32'sd42, 32'sd176, 32'sd0, -32'sd2, 32'sd48, -32'sd352, 32'sd61, -32'sd74, -32'sd1, 32'sd45, 32'sd182, 32'sd31, -32'sd1, -32'sd2, -32'sd116, -32'sd27, 32'sd25, -32'sd12, -32'sd71, 32'sd24, 32'sd248, -32'sd34, -32'sd70, -32'sd328, -32'sd32, 32'sd21, 32'sd28, 32'sd40, -32'sd122, 32'sd16, -32'sd8, 32'sd5, -32'sd6, 32'sd5, 32'sd4, 32'sd132, -32'sd9, -32'sd76, -32'sd8, 32'sd7, -32'sd1, 32'sd19, -32'sd23, -32'sd76, -32'sd138, 32'sd100, -32'sd8, -32'sd2, -32'sd7, 32'sd44, -32'sd34, -32'sd17, 32'sd4, 32'sd3, 32'sd58, -32'sd25, -32'sd69, -32'sd2, 32'sd9, 32'sd87, -32'sd26, 32'sd91, -32'sd47, -32'sd110, -32'sd35, -32'sd44, -32'sd41, -32'sd88, -32'sd27, -32'sd63, 32'sd172, 32'sd6, -32'sd91, 32'sd129, -32'sd2, -32'sd105, 32'sd69, -32'sd43, -32'sd153, -32'sd114, 32'sd21, 32'sd80, -32'sd36, -32'sd82, -32'sd98, 32'sd58, -32'sd98, 32'sd6, -32'sd6, -32'sd3, -32'sd123, -32'sd90, -32'sd36, -32'sd32, -32'sd89, 32'sd59, 32'sd23, -32'sd81, -32'sd132, 32'sd44, -32'sd37, -32'sd57, 32'sd23, -32'sd1, 32'sd212, -32'sd1, 32'sd0, -32'sd79, 32'sd90, 32'sd50, -32'sd3, 32'sd60, 32'sd41, -32'sd157, 32'sd6, -32'sd21, 32'sd43, -32'sd109, 32'sd7, 32'sd67, 32'sd80, -32'sd79, -32'sd108, -32'sd8, -32'sd23, -32'sd4, -32'sd31, -32'sd30, 32'sd50, -32'sd34, 32'sd22, -32'sd139, 32'sd92, -32'sd152, 32'sd81, 32'sd169, -32'sd43, -32'sd33, 32'sd18, -32'sd149, -32'sd51, 32'sd63, 32'sd240, -32'sd114, -32'sd149, -32'sd86, -32'sd61, 32'sd15, -32'sd10, -32'sd26, 32'sd118, -32'sd34, -32'sd69, 32'sd2, -32'sd2, -32'sd23, 32'sd27, 32'sd3, -32'sd2, -32'sd24, 32'sd52, -32'sd26, -32'sd217, -32'sd4, -32'sd26, -32'sd58, 32'sd30, -32'sd23, -32'sd35, -32'sd59, 32'sd53, 32'sd19, 32'sd96, -32'sd24, 32'sd45, -32'sd82, 32'sd2, 32'sd135, 32'sd38, -32'sd28, 32'sd31, -32'sd4, -32'sd1, 32'sd10, 32'sd10, -32'sd18, -32'sd238, -32'sd24, 32'sd18, 32'sd206, -32'sd104, -32'sd178, 32'sd4, -32'sd71, 32'sd3, 32'sd57, 32'sd23, -32'sd8, 32'sd26, -32'sd41, 32'sd111, 32'sd82, 32'sd22, 32'sd31, 32'sd69, 32'sd306, 32'sd20, 32'sd0, -32'sd15, -32'sd135, -32'sd26, -32'sd27, 32'sd14, -32'sd220, 32'sd83, -32'sd1, 32'sd25, -32'sd111, 32'sd18, 32'sd43, -32'sd320, 32'sd65, -32'sd375, -32'sd77, 32'sd43, -32'sd142, 32'sd57, -32'sd133, 32'sd4, 32'sd68, -32'sd69, -32'sd64, -32'sd42, -32'sd41, 32'sd14, -32'sd18, 32'sd121, -32'sd70, 32'sd2, -32'sd40, -32'sd1, -32'sd98, 32'sd31, -32'sd12, -32'sd101, -32'sd13, -32'sd52, 32'sd26, 32'sd0, -32'sd1, -32'sd47, -32'sd183, -32'sd5, 32'sd34, -32'sd107, -32'sd63, -32'sd24, 32'sd30, -32'sd5, -32'sd228, -32'sd28, 
                                                    -32'sd23, -32'sd1, 32'sd39, -32'sd122, 32'sd4, 32'sd125, -32'sd3, -32'sd7, 32'sd84, 32'sd3, -32'sd1, 32'sd44, -32'sd1, -32'sd67, -32'sd75, 32'sd3, -32'sd47, 32'sd5, -32'sd19, -32'sd28, -32'sd139, -32'sd20, 32'sd6, -32'sd198, 32'sd21, -32'sd99, 32'sd14, 32'sd142, 32'sd35, -32'sd103, 32'sd18, 32'sd25, -32'sd6, -32'sd21, -32'sd16, -32'sd4, -32'sd8, -32'sd47, 32'sd15, -32'sd67, 32'sd83, 32'sd22, -32'sd25, -32'sd65, -32'sd9, -32'sd52, -32'sd27, -32'sd64, -32'sd26, 32'sd23, 32'sd2, -32'sd27, 32'sd32, -32'sd244, -32'sd91, -32'sd22, 32'sd24, 32'sd1, 32'sd22, -32'sd289, 32'sd308, -32'sd35, 32'sd40, -32'sd186, -32'sd2, -32'sd30, 32'sd18, -32'sd28, -32'sd15, 32'sd3, 32'sd23, -32'sd19, -32'sd67, 32'sd113, -32'sd62, -32'sd27, -32'sd9, -32'sd32, 32'sd1, -32'sd23, 32'sd17, -32'sd6, 32'sd22, -32'sd145, -32'sd29, 32'sd58, -32'sd19, -32'sd87, 32'sd83, 32'sd57, -32'sd11, -32'sd60, 32'sd37, -32'sd155, -32'sd6, -32'sd34, -32'sd17, 32'sd249, 32'sd20, -32'sd91, 32'sd118, -32'sd29, -32'sd93, 32'sd160, -32'sd185, -32'sd100, -32'sd109, -32'sd19, 32'sd70, 32'sd47, -32'sd4, -32'sd79, -32'sd8, -32'sd44, -32'sd39, 32'sd10, -32'sd125, 32'sd24, -32'sd8, 32'sd42, -32'sd38, -32'sd155, 32'sd17, -32'sd85, 32'sd21, -32'sd7, 32'sd26, -32'sd101, 32'sd37, 32'sd221, 32'sd2, -32'sd10, 32'sd41, 32'sd98, 32'sd24, -32'sd30, 32'sd22, -32'sd6, 32'sd103, -32'sd105, 32'sd19, -32'sd93, 32'sd73, 32'sd5, -32'sd254, 32'sd64, 32'sd51, -32'sd98, 32'sd111, -32'sd72, 32'sd5, -32'sd25, 32'sd24, -32'sd6, 32'sd181, 32'sd169, 32'sd6, -32'sd27, -32'sd160, 32'sd33, 32'sd29, -32'sd110, 32'sd40, 32'sd32, 32'sd34, -32'sd69, 32'sd92, -32'sd75, -32'sd95, 32'sd23, -32'sd138, 32'sd3, -32'sd58, -32'sd35, -32'sd63, 32'sd53, 32'sd21, -32'sd141, 32'sd83, 32'sd54, 32'sd45, -32'sd37, -32'sd169, -32'sd112, 32'sd33, -32'sd127, 32'sd81, 32'sd3, -32'sd72, 32'sd0, -32'sd12, -32'sd84, -32'sd60, -32'sd136, 32'sd65, -32'sd39, -32'sd143, -32'sd111, 32'sd84, -32'sd29, 32'sd23, -32'sd42, -32'sd15, 32'sd49, -32'sd114, 32'sd69, -32'sd7, -32'sd195, 32'sd10, -32'sd25, -32'sd82, 32'sd11, -32'sd55, 32'sd51, 32'sd68, -32'sd50, 32'sd112, -32'sd149, 32'sd140, 32'sd18, 32'sd17, -32'sd2, 32'sd23, -32'sd68, -32'sd14, 32'sd50, -32'sd33, -32'sd3, 32'sd101, -32'sd61, -32'sd22, 32'sd0, 32'sd2, 32'sd26, 32'sd24, -32'sd8, -32'sd42, -32'sd80, -32'sd4, 32'sd25, 32'sd26, -32'sd73, 32'sd96, 32'sd109, 32'sd21, -32'sd170, -32'sd8, 32'sd98, 32'sd29, -32'sd204, 32'sd15, -32'sd168, 32'sd0, 32'sd84, 32'sd9, -32'sd86, 32'sd43, 32'sd58, -32'sd6, 32'sd34, -32'sd106, -32'sd86, -32'sd9, 32'sd4, 32'sd17, -32'sd76, 32'sd52, -32'sd139, 32'sd37, 32'sd84, -32'sd251, -32'sd29, 32'sd20, -32'sd50, 32'sd220, -32'sd49, -32'sd396, -32'sd18, -32'sd8, -32'sd72, 32'sd32, -32'sd335, 32'sd8, 32'sd120, 32'sd18, -32'sd2, 32'sd8, 32'sd91, 32'sd19, -32'sd48, -32'sd30, -32'sd4, 32'sd24, -32'sd20, 32'sd19, -32'sd21, -32'sd9, -32'sd3, -32'sd23, -32'sd58, 32'sd34, -32'sd20, 32'sd9, 32'sd35, -32'sd394, -32'sd187, 32'sd113, 32'sd18, -32'sd132, 32'sd10, 32'sd15, 32'sd86, 32'sd27, 32'sd57, 32'sd5, -32'sd25, 32'sd17, 32'sd108, 32'sd22, -32'sd23, -32'sd18, 32'sd134, 32'sd14, -32'sd101, -32'sd78, -32'sd2, -32'sd262, -32'sd54, 32'sd3, -32'sd22, -32'sd28, -32'sd9, 32'sd165, -32'sd149, 32'sd9, -32'sd23, 32'sd28, 32'sd79, -32'sd59, -32'sd16, -32'sd39, -32'sd29, 32'sd32, 32'sd37, 32'sd25, -32'sd97, 32'sd11, -32'sd34, 32'sd17, -32'sd52, 32'sd21, 32'sd40, -32'sd34, 32'sd20, 32'sd147, -32'sd91, 32'sd53, -32'sd171, 32'sd18, -32'sd6, 32'sd82, -32'sd28, -32'sd103, -32'sd41, -32'sd82, -32'sd59, 32'sd59, 32'sd47, 32'sd3, 32'sd22, -32'sd123, -32'sd91, 32'sd9, -32'sd96, 32'sd87, -32'sd16, 32'sd9, 32'sd122, -32'sd36, 32'sd49, 32'sd0, 32'sd109, -32'sd118, -32'sd70, -32'sd1, 32'sd92, 32'sd25, 32'sd15, -32'sd7, -32'sd14, -32'sd23, 32'sd21, 32'sd26, 32'sd120, 32'sd0, 32'sd0, 32'sd93, 32'sd128, -32'sd6, 32'sd2, -32'sd121, -32'sd56, -32'sd23, 32'sd74, -32'sd3, -32'sd18, 32'sd125, -32'sd11, -32'sd265, 32'sd56, 32'sd37, -32'sd73, 32'sd44, 32'sd72, -32'sd19, 32'sd31, 32'sd55, 32'sd3, 32'sd23, 32'sd19, -32'sd25, 32'sd0, 32'sd162, 32'sd83, -32'sd132, -32'sd61, -32'sd27, 32'sd66, -32'sd27, 32'sd23, -32'sd19, -32'sd36, -32'sd57, 32'sd5, 32'sd51, 32'sd282, -32'sd36, 32'sd44, 32'sd37, 32'sd82, 32'sd10, -32'sd57, -32'sd126, 32'sd29, 32'sd107, 32'sd15, -32'sd5, -32'sd173, -32'sd23, 32'sd16, 32'sd103, 32'sd21, 32'sd20, -32'sd236, -32'sd103, -32'sd18, -32'sd3, -32'sd94, -32'sd58, 32'sd27, 32'sd51, -32'sd3, -32'sd64, 32'sd23, 32'sd6, 32'sd22, -32'sd59, 32'sd7, 32'sd19, 32'sd18, -32'sd37, -32'sd39, -32'sd126, 32'sd6, 32'sd30, 32'sd60, -32'sd27, 32'sd21, -32'sd72, -32'sd456, -32'sd5, -32'sd72, -32'sd4, -32'sd68, -32'sd28, 32'sd18, -32'sd44, 32'sd123, 32'sd223, 32'sd178, 32'sd7, -32'sd12, 32'sd5, 32'sd122, -32'sd17, 32'sd29, -32'sd28, 32'sd165, -32'sd506, 32'sd48, -32'sd3, 32'sd22, -32'sd120, 32'sd17, -32'sd146, 32'sd63, -32'sd40, -32'sd49, -32'sd24, -32'sd76, -32'sd20, 32'sd41, -32'sd20, 32'sd97, -32'sd113, 32'sd31, -32'sd240, 32'sd17, -32'sd3, 32'sd60, 32'sd51, -32'sd200, -32'sd246, 32'sd17, 32'sd131, -32'sd12, 32'sd14, 32'sd77, -32'sd24, 32'sd15, -32'sd36, 32'sd93, -32'sd25, 32'sd20, -32'sd7, -32'sd206, -32'sd8, 32'sd21, -32'sd23, 32'sd595, -32'sd22, 32'sd117, 32'sd28, -32'sd115, -32'sd48, -32'sd49, -32'sd23, -32'sd29, 32'sd91, 32'sd61, -32'sd24, 32'sd5, -32'sd30, -32'sd59, 32'sd43, -32'sd21, 32'sd29, 32'sd19, -32'sd190, -32'sd25, 32'sd17, -32'sd139, -32'sd76, -32'sd63, 32'sd76, -32'sd151, -32'sd78, -32'sd146, -32'sd211, -32'sd40, -32'sd89, -32'sd92, 32'sd29, 32'sd132, 32'sd58, -32'sd109, 32'sd74, -32'sd48, -32'sd34, -32'sd4, 32'sd26, 32'sd86, 32'sd22, -32'sd107, -32'sd4, 32'sd54, 32'sd9, -32'sd20, -32'sd91, -32'sd21, 32'sd50, 32'sd2, 32'sd6, -32'sd35, 32'sd108, 32'sd20, -32'sd119, 
                                                    32'sd66, 32'sd18, -32'sd115, 32'sd25, 32'sd12, -32'sd8, 32'sd31, 32'sd78, 32'sd116, -32'sd40, -32'sd85, 32'sd8, 32'sd102, 32'sd24, 32'sd75, -32'sd33, -32'sd2, 32'sd26, -32'sd137, -32'sd74, -32'sd85, -32'sd62, 32'sd74, -32'sd7, 32'sd16, 32'sd14, -32'sd222, 32'sd17, -32'sd60, 32'sd89, 32'sd216, 32'sd102, -32'sd130, 32'sd18, 32'sd65, -32'sd20, -32'sd70, -32'sd22, 32'sd32, 32'sd119, -32'sd4, 32'sd45, 32'sd9, 32'sd18, -32'sd132, -32'sd25, -32'sd99, 32'sd17, -32'sd20, 32'sd19, -32'sd91, 32'sd142, 32'sd119, -32'sd25, 32'sd54, -32'sd66, -32'sd6, 32'sd7, -32'sd30, -32'sd113, -32'sd26, 32'sd17, -32'sd22, 32'sd7, 32'sd20, 32'sd91, -32'sd20, -32'sd44, -32'sd71, -32'sd462, 32'sd66, -32'sd11, 32'sd4, 32'sd30, -32'sd5, 32'sd59, -32'sd98, -32'sd479, -32'sd82, 32'sd25, -32'sd21, 32'sd3, -32'sd217, 32'sd152, -32'sd52, 32'sd20, 32'sd63, -32'sd31, -32'sd6, 32'sd56, 32'sd24, -32'sd56, -32'sd26, 32'sd40, -32'sd40, 32'sd18, -32'sd65, 32'sd61, 32'sd58, 32'sd17, -32'sd5, -32'sd44, 32'sd1, 32'sd10, 32'sd149, -32'sd41, -32'sd23, 32'sd0, -32'sd19, -32'sd51, -32'sd23, 32'sd19, -32'sd8, 32'sd44, 32'sd40, -32'sd5, -32'sd23, -32'sd129, -32'sd69, 32'sd62, 32'sd34, 32'sd5, -32'sd77, 32'sd20, -32'sd19, 32'sd2, -32'sd2, 32'sd46, 32'sd153, -32'sd79, -32'sd234, -32'sd3840, -32'sd31, -32'sd4, -32'sd20, -32'sd8, -32'sd83, 32'sd139, -32'sd33, 32'sd18, -32'sd27, 32'sd19, 32'sd4, 32'sd162, -32'sd16, -32'sd88, -32'sd61, -32'sd60, 32'sd33, -32'sd62, -32'sd31, 32'sd97, -32'sd45, -32'sd101, 32'sd60, 32'sd86, 32'sd32, -32'sd28, 32'sd36, 32'sd7, -32'sd128, -32'sd153, 32'sd19, -32'sd182, -32'sd36, 32'sd61, -32'sd8, -32'sd110, 32'sd21, -32'sd150, 32'sd34, 32'sd5, -32'sd5, 32'sd37, -32'sd180, -32'sd27, 32'sd43, -32'sd32, 32'sd5, 32'sd68, 32'sd32, 32'sd1, -32'sd64, 32'sd11, -32'sd67, -32'sd81, 32'sd165, 32'sd107, 32'sd14, -32'sd173, -32'sd173, 32'sd52, -32'sd34, 32'sd75, -32'sd21, 32'sd2, -32'sd2, -32'sd31, -32'sd69, 32'sd96, -32'sd21, -32'sd22, 32'sd30, 32'sd32, 32'sd17, -32'sd107, 32'sd302, 32'sd24, 32'sd19, -32'sd6, 32'sd23, -32'sd126, -32'sd21, -32'sd31, 32'sd18, -32'sd133, 32'sd25, -32'sd116, -32'sd4, -32'sd128, 32'sd94, 32'sd36, 32'sd1, -32'sd26, 32'sd83, -32'sd24, -32'sd37, -32'sd9, -32'sd2, -32'sd27, -32'sd46, 32'sd139, 32'sd27, 32'sd66, -32'sd56, 32'sd4, 32'sd2, 32'sd44, 32'sd42, -32'sd32, 32'sd18, -32'sd2, 32'sd24, 32'sd45, -32'sd5, -32'sd55, 32'sd85, -32'sd63, 32'sd17, -32'sd7, -32'sd74, 32'sd125, 32'sd23, -32'sd104, 32'sd36, -32'sd17, -32'sd9, -32'sd23, -32'sd20, 32'sd37, 32'sd57, -32'sd25, -32'sd1, -32'sd54, -32'sd109, 32'sd107, 32'sd13, -32'sd24, 32'sd32, -32'sd45, 32'sd21, -32'sd19, -32'sd27, -32'sd91, 32'sd4, -32'sd35, 32'sd46, -32'sd6, 32'sd17, -32'sd138, 32'sd3, -32'sd33, -32'sd227, 32'sd38, 32'sd25, -32'sd55, -32'sd65, 32'sd100, -32'sd81, -32'sd6, 32'sd15, -32'sd2, 32'sd11, 32'sd5, -32'sd243, -32'sd8, 32'sd114, -32'sd28, 32'sd74, -32'sd69, -32'sd10, -32'sd26, 32'sd53, -32'sd4, -32'sd15, 32'sd42, -32'sd3, -32'sd56, 32'sd15, 32'sd117, 32'sd14, -32'sd18, 32'sd26, 32'sd42, 32'sd20, -32'sd10, 32'sd15, -32'sd21, 32'sd29, -32'sd25, 32'sd15, -32'sd115, 32'sd46, -32'sd59, 32'sd30, -32'sd4, -32'sd65, -32'sd69, -32'sd114, 32'sd103, 32'sd2, -32'sd6, 32'sd9, -32'sd25, -32'sd696, 32'sd57, -32'sd2, -32'sd19, 32'sd59, -32'sd211, -32'sd5, 32'sd44, 32'sd16, -32'sd8, 32'sd2, -32'sd35, -32'sd23, -32'sd41, 32'sd16, -32'sd64, 32'sd6, -32'sd5, 32'sd0, -32'sd196, 32'sd5, 32'sd13, 32'sd80, -32'sd119, -32'sd52, 32'sd12, 32'sd48, -32'sd30, 32'sd5, -32'sd64, 32'sd4, -32'sd64, 32'sd5, -32'sd8, 32'sd62, 32'sd17, -32'sd57, 32'sd4, 32'sd2, 32'sd2, 32'sd37, -32'sd52, 32'sd42, -32'sd68, -32'sd185, -32'sd101, -32'sd34, -32'sd70, 32'sd3, -32'sd64, -32'sd101, 32'sd102, -32'sd42, -32'sd35, -32'sd68, -32'sd72, -32'sd22, -32'sd12, -32'sd7, 32'sd30, 32'sd23, -32'sd55, 32'sd74, 32'sd4, 32'sd9, -32'sd161, 32'sd68, 32'sd149, 32'sd50, -32'sd94, -32'sd18, 32'sd15, -32'sd181, 32'sd57, -32'sd178, 32'sd66, -32'sd7, -32'sd10, -32'sd111, 32'sd67, -32'sd21, -32'sd22, -32'sd1, 32'sd81, -32'sd43, -32'sd4, 32'sd83, 32'sd7, 32'sd84, 32'sd25, -32'sd119, -32'sd87, 32'sd2, 32'sd129, -32'sd30, -32'sd93, -32'sd28, 32'sd21, -32'sd31, 32'sd65, 32'sd116, 32'sd18, -32'sd85, 32'sd103, -32'sd43, -32'sd71, -32'sd8, 32'sd44, 32'sd36, 32'sd150, 32'sd105, -32'sd24, 32'sd42, 32'sd25, -32'sd120, 32'sd3, -32'sd27, 32'sd95, -32'sd25, 32'sd89, 32'sd50, -32'sd9, 32'sd122, -32'sd7, 32'sd10, 32'sd7, 32'sd92, 32'sd18, 32'sd5, 32'sd69, -32'sd6, 32'sd4, -32'sd33, 32'sd20, -32'sd94, 32'sd11, -32'sd45, 32'sd36, -32'sd108, 32'sd19, -32'sd24, 32'sd57, -32'sd7, -32'sd40, 32'sd210, -32'sd100, -32'sd30, -32'sd46, 32'sd100, 32'sd151, -32'sd60, 32'sd28, -32'sd5, 32'sd54, -32'sd21, 32'sd20, -32'sd1, -32'sd4, -32'sd29, -32'sd8, -32'sd38, 32'sd28, 32'sd156, 32'sd2, -32'sd191, -32'sd49, -32'sd27, 32'sd0, -32'sd80, -32'sd54, 32'sd3, 32'sd17, 32'sd151, 32'sd4, -32'sd41, 32'sd108, 32'sd47, -32'sd67, -32'sd8, 32'sd101, -32'sd150, 32'sd5, -32'sd46, 32'sd27, -32'sd24, 32'sd33, 32'sd4, -32'sd127, -32'sd17, 32'sd43, -32'sd23, -32'sd126, -32'sd4, 32'sd149, 32'sd82, -32'sd30, -32'sd28, 32'sd21, -32'sd22, 32'sd33, -32'sd98, -32'sd35, 32'sd10, -32'sd5, -32'sd23, 32'sd24, 32'sd90, 32'sd9, 32'sd96, 32'sd25, -32'sd6, -32'sd57, 32'sd83, -32'sd7, -32'sd20, -32'sd78, -32'sd6, 32'sd14, -32'sd102, -32'sd24, -32'sd17, 32'sd62}

