320 x 240 - 63936 windows
266 x 199 - 42350 windows
222 x 166
185 x 138
154 x 115
128 x 96
107 x 80
89 x 66
74 x 55
62 x 46
51 x 38
43 x 32
35 x 26