`include "vj_weights.vh"

module vj_pipeline(
  input  logic clock, reset,
  input  logic [`WINDOW_SIZE:0][`WINDOW_SIZE:0][31:0] scan_win,
  input  logic [31:0] input_std_dev,
  input  logic [1:0][31:0] scan_win_index,
  output logic [1:0][31:0] top_left,
  output logic top_left_ready);

  logic [`WINDOW_SIZE:0][`WINDOW_SIZE:0][31:0] scan_win0, scan_win1,scan_win2,scan_win3,scan_win4,scan_win5,scan_win6,scan_win7,scan_win8,scan_win9,scan_win10,scan_win11,scan_win12,scan_win13,scan_win14,scan_win15,scan_win16,scan_win17,scan_win18,scan_win19,scan_win20,scan_win21,scan_win22,scan_win23,scan_win24,scan_win25,scan_win26,scan_win27,scan_win28,scan_win29,scan_win30,scan_win31,scan_win32,scan_win33,scan_win34,scan_win35,scan_win36,scan_win37,scan_win38,scan_win39,scan_win40,scan_win41,scan_win42,scan_win43,scan_win44,scan_win45,scan_win46,scan_win47,scan_win48,scan_win49,scan_win50,scan_win51,scan_win52,scan_win53,scan_win54,scan_win55,scan_win56,scan_win57,scan_win58,scan_win59,scan_win60,scan_win61,scan_win62,scan_win63,scan_win64,scan_win65,scan_win66,scan_win67,scan_win68,scan_win69,scan_win70,scan_win71,scan_win72,scan_win73,scan_win74,scan_win75,scan_win76,scan_win77,scan_win78,scan_win79,scan_win80,scan_win81,scan_win82,scan_win83,scan_win84,scan_win85,scan_win86,scan_win87,scan_win88,scan_win89,scan_win90,scan_win91,scan_win92,scan_win93,scan_win94,scan_win95,scan_win96,scan_win97,scan_win98,scan_win99,scan_win100,scan_win101,scan_win102,scan_win103,scan_win104,scan_win105,scan_win106,scan_win107,scan_win108,scan_win109,scan_win110,scan_win111,scan_win112,scan_win113,scan_win114,scan_win115,scan_win116,scan_win117,scan_win118,scan_win119,scan_win120,scan_win121,scan_win122,scan_win123,scan_win124,scan_win125,scan_win126,scan_win127,scan_win128,scan_win129,scan_win130,scan_win131,scan_win132,scan_win133,scan_win134,scan_win135,scan_win136,scan_win137,scan_win138,scan_win139,scan_win140,scan_win141,scan_win142,scan_win143,scan_win144,scan_win145,scan_win146,scan_win147,scan_win148,scan_win149,scan_win150,scan_win151,scan_win152,scan_win153,scan_win154,scan_win155,scan_win156,scan_win157,scan_win158,scan_win159,scan_win160,scan_win161,scan_win162,scan_win163,scan_win164,scan_win165,scan_win166,scan_win167,scan_win168,scan_win169,scan_win170,scan_win171,scan_win172,scan_win173,scan_win174,scan_win175,scan_win176,scan_win177,scan_win178,scan_win179,scan_win180,scan_win181,scan_win182,scan_win183,scan_win184,scan_win185,scan_win186,scan_win187,scan_win188,scan_win189,scan_win190,scan_win191,scan_win192,scan_win193,scan_win194,scan_win195,scan_win196,scan_win197,scan_win198,scan_win199,scan_win200,
  scan_win201,scan_win202,scan_win203,scan_win204,scan_win205,scan_win206,scan_win207,scan_win208,scan_win209,scan_win210,scan_win211,scan_win212,scan_win213,scan_win214,scan_win215,scan_win216,scan_win217,scan_win218,scan_win219,scan_win220,scan_win221,scan_win222,scan_win223,scan_win224,scan_win225,scan_win226,scan_win227,scan_win228,scan_win229,scan_win230,scan_win231,scan_win232,scan_win233,scan_win234,scan_win235,scan_win236,scan_win237,scan_win238,scan_win239,scan_win240,scan_win241,scan_win242,scan_win243,scan_win244,scan_win245,scan_win246,scan_win247,scan_win248,scan_win249,scan_win250,scan_win251,scan_win252,scan_win253,scan_win254,scan_win255,scan_win256,scan_win257,scan_win258,scan_win259,scan_win260,scan_win261,scan_win262,scan_win263,scan_win264,scan_win265,scan_win266,scan_win267,scan_win268,scan_win269,scan_win270,scan_win271,scan_win272,scan_win273,scan_win274,scan_win275,scan_win276,scan_win277,scan_win278,scan_win279,scan_win280,scan_win281,scan_win282,scan_win283,scan_win284,scan_win285,scan_win286,scan_win287,scan_win288,scan_win289,scan_win290,scan_win291,scan_win292,scan_win293,scan_win294,scan_win295,scan_win296,scan_win297,scan_win298,scan_win299,scan_win300,scan_win301,scan_win302,scan_win303,scan_win304,scan_win305,scan_win306,scan_win307,scan_win308,scan_win309,scan_win310,scan_win311,scan_win312,scan_win313,scan_win314,scan_win315,scan_win316,scan_win317,scan_win318,scan_win319,scan_win320,scan_win321,scan_win322,scan_win323,scan_win324,scan_win325,scan_win326,scan_win327,scan_win328,scan_win329,scan_win330,scan_win331,scan_win332,scan_win333,scan_win334,scan_win335,scan_win336,scan_win337,scan_win338,scan_win339,scan_win340,scan_win341,scan_win342,scan_win343,scan_win344,scan_win345,scan_win346,scan_win347,scan_win348,scan_win349,scan_win350,scan_win351,scan_win352,scan_win353,scan_win354,scan_win355,scan_win356,scan_win357,scan_win358,scan_win359,scan_win360,scan_win361,scan_win362,scan_win363,scan_win364,scan_win365,scan_win366,scan_win367,scan_win368,scan_win369,scan_win370,scan_win371,scan_win372,scan_win373,scan_win374,scan_win375,scan_win376,scan_win377,scan_win378,scan_win379,scan_win380,scan_win381,scan_win382,scan_win383,scan_win384,scan_win385,scan_win386,scan_win387,scan_win388,scan_win389,scan_win390,scan_win391,scan_win392,scan_win393,scan_win394,scan_win395,scan_win396,scan_win397,scan_win398,scan_win399,scan_win400,
  scan_win401,scan_win402,scan_win403,scan_win404,scan_win405,scan_win406,scan_win407,scan_win408,scan_win409,scan_win410,scan_win411,scan_win412,scan_win413,scan_win414,scan_win415,scan_win416,scan_win417,scan_win418,scan_win419,scan_win420,scan_win421,scan_win422,scan_win423,scan_win424,scan_win425,scan_win426,scan_win427,scan_win428,scan_win429,scan_win430,scan_win431,scan_win432,scan_win433,scan_win434,scan_win435,scan_win436,scan_win437,scan_win438,scan_win439,scan_win440,scan_win441,scan_win442,scan_win443,scan_win444,scan_win445,scan_win446,scan_win447,scan_win448,scan_win449,scan_win450,scan_win451,scan_win452,scan_win453,scan_win454,scan_win455,scan_win456,scan_win457,scan_win458,scan_win459,scan_win460,scan_win461,scan_win462,scan_win463,scan_win464,scan_win465,scan_win466,scan_win467,scan_win468,scan_win469,scan_win470,scan_win471,scan_win472,scan_win473,scan_win474,scan_win475,scan_win476,scan_win477,scan_win478,scan_win479,scan_win480,scan_win481,scan_win482,scan_win483,scan_win484,scan_win485,scan_win486,scan_win487,scan_win488,scan_win489,scan_win490,scan_win491,scan_win492,scan_win493,scan_win494,scan_win495,scan_win496,scan_win497,scan_win498,scan_win499,scan_win500,scan_win501,scan_win502,scan_win503,scan_win504,scan_win505,scan_win506,scan_win507,scan_win508,scan_win509,scan_win510,scan_win511,scan_win512,scan_win513,scan_win514,scan_win515,scan_win516,scan_win517,scan_win518,scan_win519,scan_win520,scan_win521,scan_win522,scan_win523,scan_win524,scan_win525,scan_win526,scan_win527,scan_win528,scan_win529,scan_win530,scan_win531,scan_win532,scan_win533,scan_win534,scan_win535,scan_win536,scan_win537,scan_win538,scan_win539,scan_win540,scan_win541,scan_win542,scan_win543,scan_win544,scan_win545,scan_win546,scan_win547,scan_win548,scan_win549,scan_win550,scan_win551,scan_win552,scan_win553,scan_win554,scan_win555,scan_win556,scan_win557,scan_win558,scan_win559,scan_win560,scan_win561,scan_win562,scan_win563,scan_win564,scan_win565,scan_win566,scan_win567,scan_win568,scan_win569,scan_win570,scan_win571,scan_win572,scan_win573,scan_win574,scan_win575,scan_win576,scan_win577,scan_win578,scan_win579,scan_win580,scan_win581,scan_win582,scan_win583,scan_win584,scan_win585,scan_win586,scan_win587,scan_win588,scan_win589,scan_win590,scan_win591,scan_win592,scan_win593,scan_win594,scan_win595,scan_win596,scan_win597,scan_win598,scan_win599,scan_win600,
  scan_win601,scan_win602,scan_win603,scan_win604,scan_win605,scan_win606,scan_win607,scan_win608,scan_win609,scan_win610,scan_win611,scan_win612,scan_win613,scan_win614,scan_win615,scan_win616,scan_win617,scan_win618,scan_win619,scan_win620,scan_win621,scan_win622,scan_win623,scan_win624,scan_win625,scan_win626,scan_win627,scan_win628,scan_win629,scan_win630,scan_win631,scan_win632,scan_win633,scan_win634,scan_win635,scan_win636,scan_win637,scan_win638,scan_win639,scan_win640,scan_win641,scan_win642,scan_win643,scan_win644,scan_win645,scan_win646,scan_win647,scan_win648,scan_win649,scan_win650,scan_win651,scan_win652,scan_win653,scan_win654,scan_win655,scan_win656,scan_win657,scan_win658,scan_win659,scan_win660,scan_win661,scan_win662,scan_win663,scan_win664,scan_win665,scan_win666,scan_win667,scan_win668,scan_win669,scan_win670,scan_win671,scan_win672,scan_win673,scan_win674,scan_win675,scan_win676,scan_win677,scan_win678,scan_win679,scan_win680,scan_win681,scan_win682,scan_win683,scan_win684,scan_win685,scan_win686,scan_win687,scan_win688,scan_win689,scan_win690,scan_win691,scan_win692,scan_win693,scan_win694,scan_win695,scan_win696,scan_win697,scan_win698,scan_win699,scan_win700,scan_win701,scan_win702,scan_win703,scan_win704,scan_win705,scan_win706,scan_win707,scan_win708,scan_win709,scan_win710,scan_win711,scan_win712,scan_win713,scan_win714,scan_win715,scan_win716,scan_win717,scan_win718,scan_win719,scan_win720,scan_win721,scan_win722,scan_win723,scan_win724,scan_win725,scan_win726,scan_win727,scan_win728,scan_win729,scan_win730,scan_win731,scan_win732,scan_win733,scan_win734,scan_win735,scan_win736,scan_win737,scan_win738,scan_win739,scan_win740,scan_win741,scan_win742,scan_win743,scan_win744,scan_win745,scan_win746,scan_win747,scan_win748,scan_win749,scan_win750,scan_win751,scan_win752,scan_win753,scan_win754,scan_win755,scan_win756,scan_win757,scan_win758,scan_win759,scan_win760,scan_win761,scan_win762,scan_win763,scan_win764,scan_win765,scan_win766,scan_win767,scan_win768,scan_win769,scan_win770,scan_win771,scan_win772,scan_win773,scan_win774,scan_win775,scan_win776,scan_win777,scan_win778,scan_win779,scan_win780,scan_win781,scan_win782,scan_win783,scan_win784,scan_win785,scan_win786,scan_win787,scan_win788,scan_win789,scan_win790,scan_win791,scan_win792,scan_win793,scan_win794,scan_win795,scan_win796,scan_win797,scan_win798,scan_win799,scan_win800,
  scan_win801,scan_win802,scan_win803,scan_win804,scan_win805,scan_win806,scan_win807,scan_win808,scan_win809,scan_win810,scan_win811,scan_win812,scan_win813,scan_win814,scan_win815,scan_win816,scan_win817,scan_win818,scan_win819,scan_win820,scan_win821,scan_win822,scan_win823,scan_win824,scan_win825,scan_win826,scan_win827,scan_win828,scan_win829,scan_win830,scan_win831,scan_win832,scan_win833,scan_win834,scan_win835,scan_win836,scan_win837,scan_win838,scan_win839,scan_win840,scan_win841,scan_win842,scan_win843,scan_win844,scan_win845,scan_win846,scan_win847,scan_win848,scan_win849,scan_win850,scan_win851,scan_win852,scan_win853,scan_win854,scan_win855,scan_win856,scan_win857,scan_win858,scan_win859,scan_win860,scan_win861,scan_win862,scan_win863,scan_win864,scan_win865,scan_win866,scan_win867,scan_win868,scan_win869,scan_win870,scan_win871,scan_win872,scan_win873,scan_win874,scan_win875,scan_win876,scan_win877,scan_win878,scan_win879,scan_win880,scan_win881,scan_win882,scan_win883,scan_win884,scan_win885,scan_win886,scan_win887,scan_win888,scan_win889,scan_win890,scan_win891,scan_win892,scan_win893,scan_win894,scan_win895,scan_win896,scan_win897,scan_win898,scan_win899,scan_win900,scan_win901,scan_win902,scan_win903,scan_win904,scan_win905,scan_win906,scan_win907,scan_win908,scan_win909,scan_win910,scan_win911,scan_win912,scan_win913,scan_win914,scan_win915,scan_win916,scan_win917,scan_win918,scan_win919,scan_win920,scan_win921,scan_win922,scan_win923,scan_win924,scan_win925,scan_win926,scan_win927,scan_win928,scan_win929,scan_win930,scan_win931,scan_win932,scan_win933,scan_win934,scan_win935,scan_win936,scan_win937,scan_win938,scan_win939,scan_win940,scan_win941,scan_win942,scan_win943,scan_win944,scan_win945,scan_win946,scan_win947,scan_win948,scan_win949,scan_win950,scan_win951,scan_win952,scan_win953,scan_win954,scan_win955,scan_win956,scan_win957,scan_win958,scan_win959,scan_win960,scan_win961,scan_win962,scan_win963,scan_win964,scan_win965,scan_win966,scan_win967,scan_win968,scan_win969,scan_win970,scan_win971,scan_win972,scan_win973,scan_win974,scan_win975,scan_win976,scan_win977,scan_win978,scan_win979,scan_win980,scan_win981,scan_win982,scan_win983,scan_win984,scan_win985,scan_win986,scan_win987,scan_win988,scan_win989,scan_win990,scan_win991,scan_win992,scan_win993,scan_win994,scan_win995,scan_win996,scan_win997,scan_win998,scan_win999,scan_win1000,
  scan_win1001,scan_win1002,scan_win1003,scan_win1004,scan_win1005,scan_win1006,scan_win1007,scan_win1008,scan_win1009,scan_win1010,scan_win1011,scan_win1012,scan_win1013,scan_win1014,scan_win1015,scan_win1016,scan_win1017,scan_win1018,scan_win1019,scan_win1020,scan_win1021,scan_win1022,scan_win1023,scan_win1024,scan_win1025,scan_win1026,scan_win1027,scan_win1028,scan_win1029,scan_win1030,scan_win1031,scan_win1032,scan_win1033,scan_win1034,scan_win1035,scan_win1036,scan_win1037,scan_win1038,scan_win1039,scan_win1040,scan_win1041,scan_win1042,scan_win1043,scan_win1044,scan_win1045,scan_win1046,scan_win1047,scan_win1048,scan_win1049,scan_win1050,scan_win1051,scan_win1052,scan_win1053,scan_win1054,scan_win1055,scan_win1056,scan_win1057,scan_win1058,scan_win1059,scan_win1060,scan_win1061,scan_win1062,scan_win1063,scan_win1064,scan_win1065,scan_win1066,scan_win1067,scan_win1068,scan_win1069,scan_win1070,scan_win1071,scan_win1072,scan_win1073,scan_win1074,scan_win1075,scan_win1076,scan_win1077,scan_win1078,scan_win1079,scan_win1080,scan_win1081,scan_win1082,scan_win1083,scan_win1084,scan_win1085,scan_win1086,scan_win1087,scan_win1088,scan_win1089,scan_win1090,scan_win1091,scan_win1092,scan_win1093,scan_win1094,scan_win1095,scan_win1096,scan_win1097,scan_win1098,scan_win1099,scan_win1100,scan_win1101,scan_win1102,scan_win1103,scan_win1104,scan_win1105,scan_win1106,scan_win1107,scan_win1108,scan_win1109,scan_win1110,scan_win1111,scan_win1112,scan_win1113,scan_win1114,scan_win1115,scan_win1116,scan_win1117,scan_win1118,scan_win1119,scan_win1120,scan_win1121,scan_win1122,scan_win1123,scan_win1124,scan_win1125,scan_win1126,scan_win1127,scan_win1128,scan_win1129,scan_win1130,scan_win1131,scan_win1132,scan_win1133,scan_win1134,scan_win1135,scan_win1136,scan_win1137,scan_win1138,scan_win1139,scan_win1140,scan_win1141,scan_win1142,scan_win1143,scan_win1144,scan_win1145,scan_win1146,scan_win1147,scan_win1148,scan_win1149,scan_win1150,scan_win1151,scan_win1152,scan_win1153,scan_win1154,scan_win1155,scan_win1156,scan_win1157,scan_win1158,scan_win1159,scan_win1160,scan_win1161,scan_win1162,scan_win1163,scan_win1164,scan_win1165,scan_win1166,scan_win1167,scan_win1168,scan_win1169,scan_win1170,scan_win1171,scan_win1172,scan_win1173,scan_win1174,scan_win1175,scan_win1176,scan_win1177,scan_win1178,scan_win1179,scan_win1180,scan_win1181,scan_win1182,scan_win1183,scan_win1184,scan_win1185,scan_win1186,scan_win1187,scan_win1188,scan_win1189,scan_win1190,scan_win1191,scan_win1192,scan_win1193,scan_win1194,scan_win1195,scan_win1196,scan_win1197,scan_win1198,scan_win1199,scan_win1200,
  scan_win1201,scan_win1202,scan_win1203,scan_win1204,scan_win1205,scan_win1206,scan_win1207,scan_win1208,scan_win1209,scan_win1210,scan_win1211,scan_win1212,scan_win1213,scan_win1214,scan_win1215,scan_win1216,scan_win1217,scan_win1218,scan_win1219,scan_win1220,scan_win1221,scan_win1222,scan_win1223,scan_win1224,scan_win1225,scan_win1226,scan_win1227,scan_win1228,scan_win1229,scan_win1230,scan_win1231,scan_win1232,scan_win1233,scan_win1234,scan_win1235,scan_win1236,scan_win1237,scan_win1238,scan_win1239,scan_win1240,scan_win1241,scan_win1242,scan_win1243,scan_win1244,scan_win1245,scan_win1246,scan_win1247,scan_win1248,scan_win1249,scan_win1250,scan_win1251,scan_win1252,scan_win1253,scan_win1254,scan_win1255,scan_win1256,scan_win1257,scan_win1258,scan_win1259,scan_win1260,scan_win1261,scan_win1262,scan_win1263,scan_win1264,scan_win1265,scan_win1266,scan_win1267,scan_win1268,scan_win1269,scan_win1270,scan_win1271,scan_win1272,scan_win1273,scan_win1274,scan_win1275,scan_win1276,scan_win1277,scan_win1278,scan_win1279,scan_win1280,scan_win1281,scan_win1282,scan_win1283,scan_win1284,scan_win1285,scan_win1286,scan_win1287,scan_win1288,scan_win1289,scan_win1290,scan_win1291,scan_win1292,scan_win1293,scan_win1294,scan_win1295,scan_win1296,scan_win1297,scan_win1298,scan_win1299,scan_win1300,scan_win1301,scan_win1302,scan_win1303,scan_win1304,scan_win1305,scan_win1306,scan_win1307,scan_win1308,scan_win1309,scan_win1310,scan_win1311,scan_win1312,scan_win1313,scan_win1314,scan_win1315,scan_win1316,scan_win1317,scan_win1318,scan_win1319,scan_win1320,scan_win1321,scan_win1322,scan_win1323,scan_win1324,scan_win1325,scan_win1326,scan_win1327,scan_win1328,scan_win1329,scan_win1330,scan_win1331,scan_win1332,scan_win1333,scan_win1334,scan_win1335,scan_win1336,scan_win1337,scan_win1338,scan_win1339,scan_win1340,scan_win1341,scan_win1342,scan_win1343,scan_win1344,scan_win1345,scan_win1346,scan_win1347,scan_win1348,scan_win1349,scan_win1350,scan_win1351,scan_win1352,scan_win1353,scan_win1354,scan_win1355,scan_win1356,scan_win1357,scan_win1358,scan_win1359,scan_win1360,scan_win1361,scan_win1362,scan_win1363,scan_win1364,scan_win1365,scan_win1366,scan_win1367,scan_win1368,scan_win1369,scan_win1370,scan_win1371,scan_win1372,scan_win1373,scan_win1374,scan_win1375,scan_win1376,scan_win1377,scan_win1378,scan_win1379,scan_win1380,scan_win1381,scan_win1382,scan_win1383,scan_win1384,scan_win1385,scan_win1386,scan_win1387,scan_win1388,scan_win1389,scan_win1390,scan_win1391,scan_win1392,scan_win1393,scan_win1394,scan_win1395,scan_win1396,scan_win1397,scan_win1398,scan_win1399,scan_win1400,
  scan_win1401,scan_win1402,scan_win1403,scan_win1404,scan_win1405,scan_win1406,scan_win1407,scan_win1408,scan_win1409,scan_win1410,scan_win1411,scan_win1412,scan_win1413,scan_win1414,scan_win1415,scan_win1416,scan_win1417,scan_win1418,scan_win1419,scan_win1420,scan_win1421,scan_win1422,scan_win1423,scan_win1424,scan_win1425,scan_win1426,scan_win1427,scan_win1428,scan_win1429,scan_win1430,scan_win1431,scan_win1432,scan_win1433,scan_win1434,scan_win1435,scan_win1436,scan_win1437,scan_win1438,scan_win1439,scan_win1440,scan_win1441,scan_win1442,scan_win1443,scan_win1444,scan_win1445,scan_win1446,scan_win1447,scan_win1448,scan_win1449,scan_win1450,scan_win1451,scan_win1452,scan_win1453,scan_win1454,scan_win1455,scan_win1456,scan_win1457,scan_win1458,scan_win1459,scan_win1460,scan_win1461,scan_win1462,scan_win1463,scan_win1464,scan_win1465,scan_win1466,scan_win1467,scan_win1468,scan_win1469,scan_win1470,scan_win1471,scan_win1472,scan_win1473,scan_win1474,scan_win1475,scan_win1476,scan_win1477,scan_win1478,scan_win1479,scan_win1480,scan_win1481,scan_win1482,scan_win1483,scan_win1484,scan_win1485,scan_win1486,scan_win1487,scan_win1488,scan_win1489,scan_win1490,scan_win1491,scan_win1492,scan_win1493,scan_win1494,scan_win1495,scan_win1496,scan_win1497,scan_win1498,scan_win1499,scan_win1500,scan_win1501,scan_win1502,scan_win1503,scan_win1504,scan_win1505,scan_win1506,scan_win1507,scan_win1508,scan_win1509,scan_win1510,scan_win1511,scan_win1512,scan_win1513,scan_win1514,scan_win1515,scan_win1516,scan_win1517,scan_win1518,scan_win1519,scan_win1520,scan_win1521,scan_win1522,scan_win1523,scan_win1524,scan_win1525,scan_win1526,scan_win1527,scan_win1528,scan_win1529,scan_win1530,scan_win1531,scan_win1532,scan_win1533,scan_win1534,scan_win1535,scan_win1536,scan_win1537,scan_win1538,scan_win1539,scan_win1540,scan_win1541,scan_win1542,scan_win1543,scan_win1544,scan_win1545,scan_win1546,scan_win1547,scan_win1548,scan_win1549,scan_win1550,scan_win1551,scan_win1552,scan_win1553,scan_win1554,scan_win1555,scan_win1556,scan_win1557,scan_win1558,scan_win1559,scan_win1560,scan_win1561,scan_win1562,scan_win1563,scan_win1564,scan_win1565,scan_win1566,scan_win1567,scan_win1568,scan_win1569,scan_win1570,scan_win1571,scan_win1572,scan_win1573,scan_win1574,scan_win1575,scan_win1576,scan_win1577,scan_win1578,scan_win1579,scan_win1580,scan_win1581,scan_win1582,scan_win1583,scan_win1584,scan_win1585,scan_win1586,scan_win1587,scan_win1588,scan_win1589,scan_win1590,scan_win1591,scan_win1592,scan_win1593,scan_win1594,scan_win1595,scan_win1596,scan_win1597,scan_win1598,scan_win1599,scan_win1600,
  scan_win1601,scan_win1602,scan_win1603,scan_win1604,scan_win1605,scan_win1606,scan_win1607,scan_win1608,scan_win1609,scan_win1610,scan_win1611,scan_win1612,scan_win1613,scan_win1614,scan_win1615,scan_win1616,scan_win1617,scan_win1618,scan_win1619,scan_win1620,scan_win1621,scan_win1622,scan_win1623,scan_win1624,scan_win1625,scan_win1626,scan_win1627,scan_win1628,scan_win1629,scan_win1630,scan_win1631,scan_win1632,scan_win1633,scan_win1634,scan_win1635,scan_win1636,scan_win1637,scan_win1638,scan_win1639,scan_win1640,scan_win1641,scan_win1642,scan_win1643,scan_win1644,scan_win1645,scan_win1646,scan_win1647,scan_win1648,scan_win1649,scan_win1650,scan_win1651,scan_win1652,scan_win1653,scan_win1654,scan_win1655,scan_win1656,scan_win1657,scan_win1658,scan_win1659,scan_win1660,scan_win1661,scan_win1662,scan_win1663,scan_win1664,scan_win1665,scan_win1666,scan_win1667,scan_win1668,scan_win1669,scan_win1670,scan_win1671,scan_win1672,scan_win1673,scan_win1674,scan_win1675,scan_win1676,scan_win1677,scan_win1678,scan_win1679,scan_win1680,scan_win1681,scan_win1682,scan_win1683,scan_win1684,scan_win1685,scan_win1686,scan_win1687,scan_win1688,scan_win1689,scan_win1690,scan_win1691,scan_win1692,scan_win1693,scan_win1694,scan_win1695,scan_win1696,scan_win1697,scan_win1698,scan_win1699,scan_win1700,scan_win1701,scan_win1702,scan_win1703,scan_win1704,scan_win1705,scan_win1706,scan_win1707,scan_win1708,scan_win1709,scan_win1710,scan_win1711,scan_win1712,scan_win1713,scan_win1714,scan_win1715,scan_win1716,scan_win1717,scan_win1718,scan_win1719,scan_win1720,scan_win1721,scan_win1722,scan_win1723,scan_win1724,scan_win1725,scan_win1726,scan_win1727,scan_win1728,scan_win1729,scan_win1730,scan_win1731,scan_win1732,scan_win1733,scan_win1734,scan_win1735,scan_win1736,scan_win1737,scan_win1738,scan_win1739,scan_win1740,scan_win1741,scan_win1742,scan_win1743,scan_win1744,scan_win1745,scan_win1746,scan_win1747,scan_win1748,scan_win1749,scan_win1750,scan_win1751,scan_win1752,scan_win1753,scan_win1754,scan_win1755,scan_win1756,scan_win1757,scan_win1758,scan_win1759,scan_win1760,scan_win1761,scan_win1762,scan_win1763,scan_win1764,scan_win1765,scan_win1766,scan_win1767,scan_win1768,scan_win1769,scan_win1770,scan_win1771,scan_win1772,scan_win1773,scan_win1774,scan_win1775,scan_win1776,scan_win1777,scan_win1778,scan_win1779,scan_win1780,scan_win1781,scan_win1782,scan_win1783,scan_win1784,scan_win1785,scan_win1786,scan_win1787,scan_win1788,scan_win1789,scan_win1790,scan_win1791,scan_win1792,scan_win1793,scan_win1794,scan_win1795,scan_win1796,scan_win1797,scan_win1798,scan_win1799,scan_win1800,
  scan_win1801,scan_win1802,scan_win1803,scan_win1804,scan_win1805,scan_win1806,scan_win1807,scan_win1808,scan_win1809,scan_win1810,scan_win1811,scan_win1812,scan_win1813,scan_win1814,scan_win1815,scan_win1816,scan_win1817,scan_win1818,scan_win1819,scan_win1820,scan_win1821,scan_win1822,scan_win1823,scan_win1824,scan_win1825,scan_win1826,scan_win1827,scan_win1828,scan_win1829,scan_win1830,scan_win1831,scan_win1832,scan_win1833,scan_win1834,scan_win1835,scan_win1836,scan_win1837,scan_win1838,scan_win1839,scan_win1840,scan_win1841,scan_win1842,scan_win1843,scan_win1844,scan_win1845,scan_win1846,scan_win1847,scan_win1848,scan_win1849,scan_win1850,scan_win1851,scan_win1852,scan_win1853,scan_win1854,scan_win1855,scan_win1856,scan_win1857,scan_win1858,scan_win1859,scan_win1860,scan_win1861,scan_win1862,scan_win1863,scan_win1864,scan_win1865,scan_win1866,scan_win1867,scan_win1868,scan_win1869,scan_win1870,scan_win1871,scan_win1872,scan_win1873,scan_win1874,scan_win1875,scan_win1876,scan_win1877,scan_win1878,scan_win1879,scan_win1880,scan_win1881,scan_win1882,scan_win1883,scan_win1884,scan_win1885,scan_win1886,scan_win1887,scan_win1888,scan_win1889,scan_win1890,scan_win1891,scan_win1892,scan_win1893,scan_win1894,scan_win1895,scan_win1896,scan_win1897,scan_win1898,scan_win1899,scan_win1900,scan_win1901,scan_win1902,scan_win1903,scan_win1904,scan_win1905,scan_win1906,scan_win1907,scan_win1908,scan_win1909,scan_win1910,scan_win1911,scan_win1912,scan_win1913,scan_win1914,scan_win1915,scan_win1916,scan_win1917,scan_win1918,scan_win1919,scan_win1920,scan_win1921,scan_win1922,scan_win1923,scan_win1924,scan_win1925,scan_win1926,scan_win1927,scan_win1928,scan_win1929,scan_win1930,scan_win1931,scan_win1932,scan_win1933,scan_win1934,scan_win1935,scan_win1936,scan_win1937,scan_win1938,scan_win1939,scan_win1940,scan_win1941,scan_win1942,scan_win1943,scan_win1944,scan_win1945,scan_win1946,scan_win1947,scan_win1948,scan_win1949,scan_win1950,scan_win1951,scan_win1952,scan_win1953,scan_win1954,scan_win1955,scan_win1956,scan_win1957,scan_win1958,scan_win1959,scan_win1960,scan_win1961,scan_win1962,scan_win1963,scan_win1964,scan_win1965,scan_win1966,scan_win1967,scan_win1968,scan_win1969,scan_win1970,scan_win1971,scan_win1972,scan_win1973,scan_win1974,scan_win1975,scan_win1976,scan_win1977,scan_win1978,scan_win1979,scan_win1980,scan_win1981,scan_win1982,scan_win1983,scan_win1984,scan_win1985,scan_win1986,scan_win1987,scan_win1988,scan_win1989,scan_win1990,scan_win1991,scan_win1992,scan_win1993,scan_win1994,scan_win1995,scan_win1996,scan_win1997,scan_win1998,scan_win1999,scan_win2000,
  scan_win2001,scan_win2002,scan_win2003,scan_win2004,scan_win2005,scan_win2006,scan_win2007,scan_win2008,scan_win2009,scan_win2010,scan_win2011,scan_win2012,scan_win2013,scan_win2014,scan_win2015,scan_win2016,scan_win2017,scan_win2018,scan_win2019,scan_win2020,scan_win2021,scan_win2022,scan_win2023,scan_win2024,scan_win2025,scan_win2026,scan_win2027,scan_win2028,scan_win2029,scan_win2030,scan_win2031,scan_win2032,scan_win2033,scan_win2034,scan_win2035,scan_win2036,scan_win2037,scan_win2038,scan_win2039,scan_win2040,scan_win2041,scan_win2042,scan_win2043,scan_win2044,scan_win2045,scan_win2046,scan_win2047,scan_win2048,scan_win2049,scan_win2050,scan_win2051,scan_win2052,scan_win2053,scan_win2054,scan_win2055,scan_win2056,scan_win2057,scan_win2058,scan_win2059,scan_win2060,scan_win2061,scan_win2062,scan_win2063,scan_win2064,scan_win2065,scan_win2066,scan_win2067,scan_win2068,scan_win2069,scan_win2070,scan_win2071,scan_win2072,scan_win2073,scan_win2074,scan_win2075,scan_win2076,scan_win2077,scan_win2078,scan_win2079,scan_win2080,scan_win2081,scan_win2082,scan_win2083,scan_win2084,scan_win2085,scan_win2086,scan_win2087,scan_win2088,scan_win2089,scan_win2090,scan_win2091,scan_win2092,scan_win2093,scan_win2094,scan_win2095,scan_win2096,scan_win2097,scan_win2098,scan_win2099,scan_win2100,scan_win2101,scan_win2102,scan_win2103,scan_win2104,scan_win2105,scan_win2106,scan_win2107,scan_win2108,scan_win2109,scan_win2110,scan_win2111,scan_win2112,scan_win2113,scan_win2114,scan_win2115,scan_win2116,scan_win2117,scan_win2118,scan_win2119,scan_win2120,scan_win2121,scan_win2122,scan_win2123,scan_win2124,scan_win2125,scan_win2126,scan_win2127,scan_win2128,scan_win2129,scan_win2130,scan_win2131,scan_win2132,scan_win2133,scan_win2134,scan_win2135,scan_win2136,scan_win2137,scan_win2138,scan_win2139,scan_win2140,scan_win2141,scan_win2142,scan_win2143,scan_win2144,scan_win2145,scan_win2146,scan_win2147,scan_win2148,scan_win2149,scan_win2150,scan_win2151,scan_win2152,scan_win2153,scan_win2154,scan_win2155,scan_win2156,scan_win2157,scan_win2158,scan_win2159,scan_win2160,scan_win2161,scan_win2162,scan_win2163,scan_win2164,scan_win2165,scan_win2166,scan_win2167,scan_win2168,scan_win2169,scan_win2170,scan_win2171,scan_win2172,scan_win2173,scan_win2174,scan_win2175,scan_win2176,scan_win2177,scan_win2178,scan_win2179,scan_win2180,scan_win2181,scan_win2182,scan_win2183,scan_win2184,scan_win2185,scan_win2186,scan_win2187,scan_win2188,scan_win2189,scan_win2190,scan_win2191,scan_win2192,scan_win2193,scan_win2194,scan_win2195,scan_win2196,scan_win2197,scan_win2198,scan_win2199,scan_win2200,
  scan_win2201,scan_win2202,scan_win2203,scan_win2204,scan_win2205,scan_win2206,scan_win2207,scan_win2208,scan_win2209,scan_win2210,scan_win2211,scan_win2212,scan_win2213,scan_win2214,scan_win2215,scan_win2216,scan_win2217,scan_win2218,scan_win2219,scan_win2220,scan_win2221,scan_win2222,scan_win2223,scan_win2224,scan_win2225,scan_win2226,scan_win2227,scan_win2228,scan_win2229,scan_win2230,scan_win2231,scan_win2232,scan_win2233,scan_win2234,scan_win2235,scan_win2236,scan_win2237,scan_win2238,scan_win2239,scan_win2240,scan_win2241,scan_win2242,scan_win2243,scan_win2244,scan_win2245,scan_win2246,scan_win2247,scan_win2248,scan_win2249,scan_win2250,scan_win2251,scan_win2252,scan_win2253,scan_win2254,scan_win2255,scan_win2256,scan_win2257,scan_win2258,scan_win2259,scan_win2260,scan_win2261,scan_win2262,scan_win2263,scan_win2264,scan_win2265,scan_win2266,scan_win2267,scan_win2268,scan_win2269,scan_win2270,scan_win2271,scan_win2272,scan_win2273,scan_win2274,scan_win2275,scan_win2276,scan_win2277,scan_win2278,scan_win2279,scan_win2280,scan_win2281,scan_win2282,scan_win2283,scan_win2284,scan_win2285,scan_win2286,scan_win2287,scan_win2288,scan_win2289,scan_win2290,scan_win2291,scan_win2292,scan_win2293,scan_win2294,scan_win2295,scan_win2296,scan_win2297,scan_win2298,scan_win2299,scan_win2300,scan_win2301,scan_win2302,scan_win2303,scan_win2304,scan_win2305,scan_win2306,scan_win2307,scan_win2308,scan_win2309,scan_win2310,scan_win2311,scan_win2312,scan_win2313,scan_win2314,scan_win2315,scan_win2316,scan_win2317,scan_win2318,scan_win2319,scan_win2320,scan_win2321,scan_win2322,scan_win2323,scan_win2324,scan_win2325,scan_win2326,scan_win2327,scan_win2328,scan_win2329,scan_win2330,scan_win2331,scan_win2332,scan_win2333,scan_win2334,scan_win2335,scan_win2336,scan_win2337,scan_win2338,scan_win2339,scan_win2340,scan_win2341,scan_win2342,scan_win2343,scan_win2344,scan_win2345,scan_win2346,scan_win2347,scan_win2348,scan_win2349,scan_win2350,scan_win2351,scan_win2352,scan_win2353,scan_win2354,scan_win2355,scan_win2356,scan_win2357,scan_win2358,scan_win2359,scan_win2360,scan_win2361,scan_win2362,scan_win2363,scan_win2364,scan_win2365,scan_win2366,scan_win2367,scan_win2368,scan_win2369,scan_win2370,scan_win2371,scan_win2372,scan_win2373,scan_win2374,scan_win2375,scan_win2376,scan_win2377,scan_win2378,scan_win2379,scan_win2380,scan_win2381,scan_win2382,scan_win2383,scan_win2384,scan_win2385,scan_win2386,scan_win2387,scan_win2388,scan_win2389,scan_win2390,scan_win2391,scan_win2392,scan_win2393,scan_win2394,scan_win2395,scan_win2396,scan_win2397,scan_win2398,scan_win2399,scan_win2400,
  scan_win2401,scan_win2402,scan_win2403,scan_win2404,scan_win2405,scan_win2406,scan_win2407,scan_win2408,scan_win2409,scan_win2410,scan_win2411,scan_win2412,scan_win2413,scan_win2414,scan_win2415,scan_win2416,scan_win2417,scan_win2418,scan_win2419,scan_win2420,scan_win2421,scan_win2422,scan_win2423,scan_win2424,scan_win2425,scan_win2426,scan_win2427,scan_win2428,scan_win2429,scan_win2430,scan_win2431,scan_win2432,scan_win2433,scan_win2434,scan_win2435,scan_win2436,scan_win2437,scan_win2438,scan_win2439,scan_win2440,scan_win2441,scan_win2442,scan_win2443,scan_win2444,scan_win2445,scan_win2446,scan_win2447,scan_win2448,scan_win2449,scan_win2450,scan_win2451,scan_win2452,scan_win2453,scan_win2454,scan_win2455,scan_win2456,scan_win2457,scan_win2458,scan_win2459,scan_win2460,scan_win2461,scan_win2462,scan_win2463,scan_win2464,scan_win2465,scan_win2466,scan_win2467,scan_win2468,scan_win2469,scan_win2470,scan_win2471,scan_win2472,scan_win2473,scan_win2474,scan_win2475,scan_win2476,scan_win2477,scan_win2478,scan_win2479,scan_win2480,scan_win2481,scan_win2482,scan_win2483,scan_win2484,scan_win2485,scan_win2486,scan_win2487,scan_win2488,scan_win2489,scan_win2490,scan_win2491,scan_win2492,scan_win2493,scan_win2494,scan_win2495,scan_win2496,scan_win2497,scan_win2498,scan_win2499,scan_win2500,scan_win2501,scan_win2502,scan_win2503,scan_win2504,scan_win2505,scan_win2506,scan_win2507,scan_win2508,scan_win2509,scan_win2510,scan_win2511,scan_win2512,scan_win2513,scan_win2514,scan_win2515,scan_win2516,scan_win2517,scan_win2518,scan_win2519,scan_win2520,scan_win2521,scan_win2522,scan_win2523,scan_win2524,scan_win2525,scan_win2526,scan_win2527,scan_win2528,scan_win2529,scan_win2530,scan_win2531,scan_win2532,scan_win2533,scan_win2534,scan_win2535,scan_win2536,scan_win2537,scan_win2538,scan_win2539,scan_win2540,scan_win2541,scan_win2542,scan_win2543,scan_win2544,scan_win2545,scan_win2546,scan_win2547,scan_win2548,scan_win2549,scan_win2550,scan_win2551,scan_win2552,scan_win2553,scan_win2554,scan_win2555,scan_win2556,scan_win2557,scan_win2558,scan_win2559,scan_win2560,scan_win2561,scan_win2562,scan_win2563,scan_win2564,scan_win2565,scan_win2566,scan_win2567,scan_win2568,scan_win2569,scan_win2570,scan_win2571,scan_win2572,scan_win2573,scan_win2574,scan_win2575,scan_win2576,scan_win2577,scan_win2578,scan_win2579,scan_win2580,scan_win2581,scan_win2582,scan_win2583,scan_win2584,scan_win2585,scan_win2586,scan_win2587,scan_win2588,scan_win2589,scan_win2590,scan_win2591,scan_win2592,scan_win2593,scan_win2594,scan_win2595,scan_win2596,scan_win2597,scan_win2598,scan_win2599,scan_win2600,
  scan_win2601,scan_win2602,scan_win2603,scan_win2604,scan_win2605,scan_win2606,scan_win2607,scan_win2608,scan_win2609,scan_win2610,scan_win2611,scan_win2612,scan_win2613,scan_win2614,scan_win2615,scan_win2616,scan_win2617,scan_win2618,scan_win2619,scan_win2620,scan_win2621,scan_win2622,scan_win2623,scan_win2624,scan_win2625,scan_win2626,scan_win2627,scan_win2628,scan_win2629,scan_win2630,scan_win2631,scan_win2632,scan_win2633,scan_win2634,scan_win2635,scan_win2636,scan_win2637,scan_win2638,scan_win2639,scan_win2640,scan_win2641,scan_win2642,scan_win2643,scan_win2644,scan_win2645,scan_win2646,scan_win2647,scan_win2648,scan_win2649,scan_win2650,scan_win2651,scan_win2652,scan_win2653,scan_win2654,scan_win2655,scan_win2656,scan_win2657,scan_win2658,scan_win2659,scan_win2660,scan_win2661,scan_win2662,scan_win2663,scan_win2664,scan_win2665,scan_win2666,scan_win2667,scan_win2668,scan_win2669,scan_win2670,scan_win2671,scan_win2672,scan_win2673,scan_win2674,scan_win2675,scan_win2676,scan_win2677,scan_win2678,scan_win2679,scan_win2680,scan_win2681,scan_win2682,scan_win2683,scan_win2684,scan_win2685,scan_win2686,scan_win2687,scan_win2688,scan_win2689,scan_win2690,scan_win2691,scan_win2692,scan_win2693,scan_win2694,scan_win2695,scan_win2696,scan_win2697,scan_win2698,scan_win2699,scan_win2700,scan_win2701,scan_win2702,scan_win2703,scan_win2704,scan_win2705,scan_win2706,scan_win2707,scan_win2708,scan_win2709,scan_win2710,scan_win2711,scan_win2712,scan_win2713,scan_win2714,scan_win2715,scan_win2716,scan_win2717,scan_win2718,scan_win2719,scan_win2720,scan_win2721,scan_win2722,scan_win2723,scan_win2724,scan_win2725,scan_win2726,scan_win2727,scan_win2728,scan_win2729,scan_win2730,scan_win2731,scan_win2732,scan_win2733,scan_win2734,scan_win2735,scan_win2736,scan_win2737,scan_win2738,scan_win2739,scan_win2740,scan_win2741,scan_win2742,scan_win2743,scan_win2744,scan_win2745,scan_win2746,scan_win2747,scan_win2748,scan_win2749,scan_win2750,scan_win2751,scan_win2752,scan_win2753,scan_win2754,scan_win2755,scan_win2756,scan_win2757,scan_win2758,scan_win2759,scan_win2760,scan_win2761,scan_win2762,scan_win2763,scan_win2764,scan_win2765,scan_win2766,scan_win2767,scan_win2768,scan_win2769,scan_win2770,scan_win2771,scan_win2772,scan_win2773,scan_win2774,scan_win2775,scan_win2776,scan_win2777,scan_win2778,scan_win2779,scan_win2780,scan_win2781,scan_win2782,scan_win2783,scan_win2784,scan_win2785,scan_win2786,scan_win2787,scan_win2788,scan_win2789,scan_win2790,scan_win2791,scan_win2792,scan_win2793,scan_win2794,scan_win2795,scan_win2796,scan_win2797,scan_win2798,scan_win2799,scan_win2800,
  scan_win2801,scan_win2802,scan_win2803,scan_win2804,scan_win2805,scan_win2806,scan_win2807,scan_win2808,scan_win2809,scan_win2810,scan_win2811,scan_win2812,scan_win2813,scan_win2814,scan_win2815,scan_win2816,scan_win2817,scan_win2818,scan_win2819,scan_win2820,scan_win2821,scan_win2822,scan_win2823,scan_win2824,scan_win2825,scan_win2826,scan_win2827,scan_win2828,scan_win2829,scan_win2830,scan_win2831,scan_win2832,scan_win2833,scan_win2834,scan_win2835,scan_win2836,scan_win2837,scan_win2838,scan_win2839,scan_win2840,scan_win2841,scan_win2842,scan_win2843,scan_win2844,scan_win2845,scan_win2846,scan_win2847,scan_win2848,scan_win2849,scan_win2850,scan_win2851,scan_win2852,scan_win2853,scan_win2854,scan_win2855,scan_win2856,scan_win2857,scan_win2858,scan_win2859,scan_win2860,scan_win2861,scan_win2862,scan_win2863,scan_win2864,scan_win2865,scan_win2866,scan_win2867,scan_win2868,scan_win2869,scan_win2870,scan_win2871,scan_win2872,scan_win2873,scan_win2874,scan_win2875,scan_win2876,scan_win2877,scan_win2878,scan_win2879,scan_win2880,scan_win2881,scan_win2882,scan_win2883,scan_win2884,scan_win2885,scan_win2886,scan_win2887,scan_win2888,scan_win2889,scan_win2890,scan_win2891,scan_win2892,scan_win2893,scan_win2894,scan_win2895,scan_win2896,scan_win2897,scan_win2898,scan_win2899,scan_win2900,scan_win2901,scan_win2902,scan_win2903,scan_win2904,scan_win2905,scan_win2906,scan_win2907,scan_win2908,scan_win2909,scan_win2910,scan_win2911,scan_win2912;
  logic [`NUM_FEATURE-1:0][1:0][31:0] scan_coords;
  logic [`NUM_FEATURE-1:0][31:0] scan_win_std_dev;

  localparam [`NUM_STAGE:0][31:0] stage_num_feature = `STAGE_NUM_FEATURE;
  localparam [`NUM_STAGE-1:0][31:0] stage_threshold = `STAGE_THRESHOLD;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle1_xs = `RECTANGLE1_XS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle1_ys = `RECTANGLE1_YS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle1_widths = `RECTANGLE1_WIDTHS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle1_heights = `RECTANGLE1_HEIGHTS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle1_weights = `RECTANGLE1_WEIGHTS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle2_xs = `RECTANGLE2_XS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle2_ys = `RECTANGLE2_YS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle2_widths = `RECTANGLE2_WIDTHS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle2_heights = `RECTANGLE2_HEIGHTS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle2_weights = `RECTANGLE2_WEIGHTS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle3_xs = `RECTANGLE3_XS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle3_ys = `RECTANGLE3_YS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle3_widths = `RECTANGLE3_WIDTHS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle3_heights = `RECTANGLE3_HEIGHTS;
  localparam [`NUM_FEATURE-1:0][31:0] rectangle3_weights = `RECTANGLE3_WEIGHTS;
  localparam [`NUM_FEATURE-1:0][31:0] feature_thresholds = `FEATURE_THRESHOLD;
  localparam [`NUM_FEATURE-1:0][31:0] feature_aboves = `FEATURE_ABOVE;
  localparam [`NUM_FEATURE-1:0][31:0] feature_belows = `FEATURE_BELOW;

  always_ff @(posedge clock, posedge reset) begin: set_scan_coords_and_scan_win_std_devs
    if (reset) begin: reset_scanning_windows
       scan_coords <= 'd0;
       scan_win_std_dev <= 'd0;
       top_left <= 'd0;
    end else begin: move_scan_coords_and_scan_win_std_devs
      scan_coords[0] <= scan_win_index;
      scan_win_std_dev[0] <= input_std_dev;
      for (int i = 0; i < `NUM_FEATURE-1; i++) begin
        scan_coords[i+1] <= scan_coords[i];
        scan_win_std_dev[i+1] <= scan_win_std_dev[i];
      end
      top_left <= scan_coords[`NUM_FEATURE-1];
    end
  end

  logic [`NUM_FEATURE-1:0][31:0] rectangle1_vals, rectangle2_vals, rectangle3_vals,
                                rectangle1_products, rectangle2_products, rectangle3_products,
                                feature_sums, feature_products,
                                feature_accums;
  logic [`NUM_FEATURE-1:0] feature_comparisons;

  logic [`NUM_FEATURE:0][31:0] stage_accums; // stage_accums[0] is wire to zero and stage_accums[2913] is reg to zero
  logic [`NUM_FEATURE:0] is_feature; // is_feature[0] is wire to one and is_feature[2913] is reg to face_coords_ready
  logic [`NUM_STAGE:1] stage_comparisons;
  assign top_left_ready = is_feature[`NUM_FEATURE];

  always_ff @(posedge clock, posedge reset) begin: set_accums_and_is_feature
    if (reset) begin
      stage_accums <= 'd0;
      is_feature <= 'd0;
    end else begin
      stage_accums[0] <= 32'd0;
      is_feature[0] <= 1'd1;
      for (int k = 1; k < 26; k++) begin
        for (int l = stage_num_feature[k-1]; l < stage_num_feature[k] - 1; l++) begin
          stage_accums[l+1] <= stage_accums[l] + feature_accums[l];
          is_feature[l+1] <= is_feature[l];
        end
        is_feature[stage_num_feature[k]] <= stage_comparisons[k] & is_feature[stage_num_feature[k] - 1];
        stage_accums[stage_num_feature[k]] <= 32'd0;
      end
    end
  end

  genvar m;
  generate
    for (m = 1; m < `NUM_STAGE+1; m=m+1) begin: stage_threshold_check
      signed_comparator stage_c(.gt(stage_comparisons[m]), .A(stage_accums[stage_num_feature[m] - 1] + feature_accums[stage_num_feature[m] - 1]), .B(stage_threshold[m-1]));
    end
  endgenerate

  always_ff @(posedge clock, posedge reset) begin : set_scan_wins
    if (reset) begin: reset_scan_wins
      scan_win0 <= 32'd0; 
      scan_win1 <= 32'd0; scan_win2 <= 32'd0; scan_win3 <= 32'd0; scan_win4 <= 32'd0; scan_win5 <= 32'd0; scan_win6 <= 32'd0; scan_win7 <= 32'd0; scan_win8 <= 32'd0; scan_win9 <= 32'd0; scan_win10 <= 32'd0; scan_win11 <= 32'd0; scan_win12 <= 32'd0; scan_win13 <= 32'd0; scan_win14 <= 32'd0; scan_win15 <= 32'd0; scan_win16 <= 32'd0; scan_win17 <= 32'd0; scan_win18 <= 32'd0; scan_win19 <= 32'd0; scan_win20 <= 32'd0; scan_win21 <= 32'd0; scan_win22 <= 32'd0; scan_win23 <= 32'd0; scan_win24 <= 32'd0; scan_win25 <= 32'd0; scan_win26 <= 32'd0; scan_win27 <= 32'd0; scan_win28 <= 32'd0; scan_win29 <= 32'd0; scan_win30 <= 32'd0; scan_win31 <= 32'd0; scan_win32 <= 32'd0; scan_win33 <= 32'd0; scan_win34 <= 32'd0; scan_win35 <= 32'd0; scan_win36 <= 32'd0; scan_win37 <= 32'd0; scan_win38 <= 32'd0; scan_win39 <= 32'd0; scan_win40 <= 32'd0; scan_win41 <= 32'd0; scan_win42 <= 32'd0; scan_win43 <= 32'd0; scan_win44 <= 32'd0; scan_win45 <= 32'd0; scan_win46 <= 32'd0; scan_win47 <= 32'd0; scan_win48 <= 32'd0; scan_win49 <= 32'd0; scan_win50 <= 32'd0; scan_win51 <= 32'd0; scan_win52 <= 32'd0; scan_win53 <= 32'd0; scan_win54 <= 32'd0; scan_win55 <= 32'd0; scan_win56 <= 32'd0; scan_win57 <= 32'd0; scan_win58 <= 32'd0; scan_win59 <= 32'd0; scan_win60 <= 32'd0; scan_win61 <= 32'd0; scan_win62 <= 32'd0; scan_win63 <= 32'd0; scan_win64 <= 32'd0; scan_win65 <= 32'd0; scan_win66 <= 32'd0; scan_win67 <= 32'd0; scan_win68 <= 32'd0; scan_win69 <= 32'd0; scan_win70 <= 32'd0; scan_win71 <= 32'd0; scan_win72 <= 32'd0; scan_win73 <= 32'd0; scan_win74 <= 32'd0; scan_win75 <= 32'd0; scan_win76 <= 32'd0; scan_win77 <= 32'd0; scan_win78 <= 32'd0; scan_win79 <= 32'd0; scan_win80 <= 32'd0; scan_win81 <= 32'd0; scan_win82 <= 32'd0; scan_win83 <= 32'd0; scan_win84 <= 32'd0; scan_win85 <= 32'd0; scan_win86 <= 32'd0; scan_win87 <= 32'd0; scan_win88 <= 32'd0; scan_win89 <= 32'd0; scan_win90 <= 32'd0; scan_win91 <= 32'd0; scan_win92 <= 32'd0; scan_win93 <= 32'd0; scan_win94 <= 32'd0; scan_win95 <= 32'd0; scan_win96 <= 32'd0; scan_win97 <= 32'd0; scan_win98 <= 32'd0; scan_win99 <= 32'd0; scan_win100 <= 32'd0; scan_win101 <= 32'd0; scan_win102 <= 32'd0; scan_win103 <= 32'd0; scan_win104 <= 32'd0; scan_win105 <= 32'd0; scan_win106 <= 32'd0; scan_win107 <= 32'd0; scan_win108 <= 32'd0; scan_win109 <= 32'd0; scan_win110 <= 32'd0; scan_win111 <= 32'd0; scan_win112 <= 32'd0; scan_win113 <= 32'd0; scan_win114 <= 32'd0; scan_win115 <= 32'd0; scan_win116 <= 32'd0; scan_win117 <= 32'd0; scan_win118 <= 32'd0; scan_win119 <= 32'd0; scan_win120 <= 32'd0; scan_win121 <= 32'd0; scan_win122 <= 32'd0; scan_win123 <= 32'd0; scan_win124 <= 32'd0; scan_win125 <= 32'd0; scan_win126 <= 32'd0; scan_win127 <= 32'd0; scan_win128 <= 32'd0; scan_win129 <= 32'd0; scan_win130 <= 32'd0; scan_win131 <= 32'd0; scan_win132 <= 32'd0; scan_win133 <= 32'd0; scan_win134 <= 32'd0; scan_win135 <= 32'd0; scan_win136 <= 32'd0; scan_win137 <= 32'd0; scan_win138 <= 32'd0; scan_win139 <= 32'd0; scan_win140 <= 32'd0; scan_win141 <= 32'd0; scan_win142 <= 32'd0; scan_win143 <= 32'd0; scan_win144 <= 32'd0; scan_win145 <= 32'd0; scan_win146 <= 32'd0; scan_win147 <= 32'd0; scan_win148 <= 32'd0; scan_win149 <= 32'd0; scan_win150 <= 32'd0; scan_win151 <= 32'd0; scan_win152 <= 32'd0; scan_win153 <= 32'd0; scan_win154 <= 32'd0; scan_win155 <= 32'd0; scan_win156 <= 32'd0; scan_win157 <= 32'd0; scan_win158 <= 32'd0; scan_win159 <= 32'd0; scan_win160 <= 32'd0; scan_win161 <= 32'd0; scan_win162 <= 32'd0; scan_win163 <= 32'd0; scan_win164 <= 32'd0; scan_win165 <= 32'd0; scan_win166 <= 32'd0; scan_win167 <= 32'd0; scan_win168 <= 32'd0; scan_win169 <= 32'd0; scan_win170 <= 32'd0; scan_win171 <= 32'd0; scan_win172 <= 32'd0; scan_win173 <= 32'd0; scan_win174 <= 32'd0; scan_win175 <= 32'd0; scan_win176 <= 32'd0; scan_win177 <= 32'd0; scan_win178 <= 32'd0; scan_win179 <= 32'd0; scan_win180 <= 32'd0; scan_win181 <= 32'd0; scan_win182 <= 32'd0; scan_win183 <= 32'd0; scan_win184 <= 32'd0; scan_win185 <= 32'd0; scan_win186 <= 32'd0; scan_win187 <= 32'd0; scan_win188 <= 32'd0; scan_win189 <= 32'd0; scan_win190 <= 32'd0; scan_win191 <= 32'd0; scan_win192 <= 32'd0; scan_win193 <= 32'd0; scan_win194 <= 32'd0; scan_win195 <= 32'd0; scan_win196 <= 32'd0; scan_win197 <= 32'd0; scan_win198 <= 32'd0; scan_win199 <= 32'd0; scan_win200 <= 32'd0; 
      scan_win201 <= 32'd0; scan_win202 <= 32'd0; scan_win203 <= 32'd0; scan_win204 <= 32'd0; scan_win205 <= 32'd0; scan_win206 <= 32'd0; scan_win207 <= 32'd0; scan_win208 <= 32'd0; scan_win209 <= 32'd0; scan_win210 <= 32'd0; scan_win211 <= 32'd0; scan_win212 <= 32'd0; scan_win213 <= 32'd0; scan_win214 <= 32'd0; scan_win215 <= 32'd0; scan_win216 <= 32'd0; scan_win217 <= 32'd0; scan_win218 <= 32'd0; scan_win219 <= 32'd0; scan_win220 <= 32'd0; scan_win221 <= 32'd0; scan_win222 <= 32'd0; scan_win223 <= 32'd0; scan_win224 <= 32'd0; scan_win225 <= 32'd0; scan_win226 <= 32'd0; scan_win227 <= 32'd0; scan_win228 <= 32'd0; scan_win229 <= 32'd0; scan_win230 <= 32'd0; scan_win231 <= 32'd0; scan_win232 <= 32'd0; scan_win233 <= 32'd0; scan_win234 <= 32'd0; scan_win235 <= 32'd0; scan_win236 <= 32'd0; scan_win237 <= 32'd0; scan_win238 <= 32'd0; scan_win239 <= 32'd0; scan_win240 <= 32'd0; scan_win241 <= 32'd0; scan_win242 <= 32'd0; scan_win243 <= 32'd0; scan_win244 <= 32'd0; scan_win245 <= 32'd0; scan_win246 <= 32'd0; scan_win247 <= 32'd0; scan_win248 <= 32'd0; scan_win249 <= 32'd0; scan_win250 <= 32'd0; scan_win251 <= 32'd0; scan_win252 <= 32'd0; scan_win253 <= 32'd0; scan_win254 <= 32'd0; scan_win255 <= 32'd0; scan_win256 <= 32'd0; scan_win257 <= 32'd0; scan_win258 <= 32'd0; scan_win259 <= 32'd0; scan_win260 <= 32'd0; scan_win261 <= 32'd0; scan_win262 <= 32'd0; scan_win263 <= 32'd0; scan_win264 <= 32'd0; scan_win265 <= 32'd0; scan_win266 <= 32'd0; scan_win267 <= 32'd0; scan_win268 <= 32'd0; scan_win269 <= 32'd0; scan_win270 <= 32'd0; scan_win271 <= 32'd0; scan_win272 <= 32'd0; scan_win273 <= 32'd0; scan_win274 <= 32'd0; scan_win275 <= 32'd0; scan_win276 <= 32'd0; scan_win277 <= 32'd0; scan_win278 <= 32'd0; scan_win279 <= 32'd0; scan_win280 <= 32'd0; scan_win281 <= 32'd0; scan_win282 <= 32'd0; scan_win283 <= 32'd0; scan_win284 <= 32'd0; scan_win285 <= 32'd0; scan_win286 <= 32'd0; scan_win287 <= 32'd0; scan_win288 <= 32'd0; scan_win289 <= 32'd0; scan_win290 <= 32'd0; scan_win291 <= 32'd0; scan_win292 <= 32'd0; scan_win293 <= 32'd0; scan_win294 <= 32'd0; scan_win295 <= 32'd0; scan_win296 <= 32'd0; scan_win297 <= 32'd0; scan_win298 <= 32'd0; scan_win299 <= 32'd0; scan_win300 <= 32'd0; scan_win301 <= 32'd0; scan_win302 <= 32'd0; scan_win303 <= 32'd0; scan_win304 <= 32'd0; scan_win305 <= 32'd0; scan_win306 <= 32'd0; scan_win307 <= 32'd0; scan_win308 <= 32'd0; scan_win309 <= 32'd0; scan_win310 <= 32'd0; scan_win311 <= 32'd0; scan_win312 <= 32'd0; scan_win313 <= 32'd0; scan_win314 <= 32'd0; scan_win315 <= 32'd0; scan_win316 <= 32'd0; scan_win317 <= 32'd0; scan_win318 <= 32'd0; scan_win319 <= 32'd0; scan_win320 <= 32'd0; scan_win321 <= 32'd0; scan_win322 <= 32'd0; scan_win323 <= 32'd0; scan_win324 <= 32'd0; scan_win325 <= 32'd0; scan_win326 <= 32'd0; scan_win327 <= 32'd0; scan_win328 <= 32'd0; scan_win329 <= 32'd0; scan_win330 <= 32'd0; scan_win331 <= 32'd0; scan_win332 <= 32'd0; scan_win333 <= 32'd0; scan_win334 <= 32'd0; scan_win335 <= 32'd0; scan_win336 <= 32'd0; scan_win337 <= 32'd0; scan_win338 <= 32'd0; scan_win339 <= 32'd0; scan_win340 <= 32'd0; scan_win341 <= 32'd0; scan_win342 <= 32'd0; scan_win343 <= 32'd0; scan_win344 <= 32'd0; scan_win345 <= 32'd0; scan_win346 <= 32'd0; scan_win347 <= 32'd0; scan_win348 <= 32'd0; scan_win349 <= 32'd0; scan_win350 <= 32'd0; scan_win351 <= 32'd0; scan_win352 <= 32'd0; scan_win353 <= 32'd0; scan_win354 <= 32'd0; scan_win355 <= 32'd0; scan_win356 <= 32'd0; scan_win357 <= 32'd0; scan_win358 <= 32'd0; scan_win359 <= 32'd0; scan_win360 <= 32'd0; scan_win361 <= 32'd0; scan_win362 <= 32'd0; scan_win363 <= 32'd0; scan_win364 <= 32'd0; scan_win365 <= 32'd0; scan_win366 <= 32'd0; scan_win367 <= 32'd0; scan_win368 <= 32'd0; scan_win369 <= 32'd0; scan_win370 <= 32'd0; scan_win371 <= 32'd0; scan_win372 <= 32'd0; scan_win373 <= 32'd0; scan_win374 <= 32'd0; scan_win375 <= 32'd0; scan_win376 <= 32'd0; scan_win377 <= 32'd0; scan_win378 <= 32'd0; scan_win379 <= 32'd0; scan_win380 <= 32'd0; scan_win381 <= 32'd0; scan_win382 <= 32'd0; scan_win383 <= 32'd0; scan_win384 <= 32'd0; scan_win385 <= 32'd0; scan_win386 <= 32'd0; scan_win387 <= 32'd0; scan_win388 <= 32'd0; scan_win389 <= 32'd0; scan_win390 <= 32'd0; scan_win391 <= 32'd0; scan_win392 <= 32'd0; scan_win393 <= 32'd0; scan_win394 <= 32'd0; scan_win395 <= 32'd0; scan_win396 <= 32'd0; scan_win397 <= 32'd0; scan_win398 <= 32'd0; scan_win399 <= 32'd0; scan_win400 <= 32'd0; 
      scan_win401 <= 32'd0; scan_win402 <= 32'd0; scan_win403 <= 32'd0; scan_win404 <= 32'd0; scan_win405 <= 32'd0; scan_win406 <= 32'd0; scan_win407 <= 32'd0; scan_win408 <= 32'd0; scan_win409 <= 32'd0; scan_win410 <= 32'd0; scan_win411 <= 32'd0; scan_win412 <= 32'd0; scan_win413 <= 32'd0; scan_win414 <= 32'd0; scan_win415 <= 32'd0; scan_win416 <= 32'd0; scan_win417 <= 32'd0; scan_win418 <= 32'd0; scan_win419 <= 32'd0; scan_win420 <= 32'd0; scan_win421 <= 32'd0; scan_win422 <= 32'd0; scan_win423 <= 32'd0; scan_win424 <= 32'd0; scan_win425 <= 32'd0; scan_win426 <= 32'd0; scan_win427 <= 32'd0; scan_win428 <= 32'd0; scan_win429 <= 32'd0; scan_win430 <= 32'd0; scan_win431 <= 32'd0; scan_win432 <= 32'd0; scan_win433 <= 32'd0; scan_win434 <= 32'd0; scan_win435 <= 32'd0; scan_win436 <= 32'd0; scan_win437 <= 32'd0; scan_win438 <= 32'd0; scan_win439 <= 32'd0; scan_win440 <= 32'd0; scan_win441 <= 32'd0; scan_win442 <= 32'd0; scan_win443 <= 32'd0; scan_win444 <= 32'd0; scan_win445 <= 32'd0; scan_win446 <= 32'd0; scan_win447 <= 32'd0; scan_win448 <= 32'd0; scan_win449 <= 32'd0; scan_win450 <= 32'd0; scan_win451 <= 32'd0; scan_win452 <= 32'd0; scan_win453 <= 32'd0; scan_win454 <= 32'd0; scan_win455 <= 32'd0; scan_win456 <= 32'd0; scan_win457 <= 32'd0; scan_win458 <= 32'd0; scan_win459 <= 32'd0; scan_win460 <= 32'd0; scan_win461 <= 32'd0; scan_win462 <= 32'd0; scan_win463 <= 32'd0; scan_win464 <= 32'd0; scan_win465 <= 32'd0; scan_win466 <= 32'd0; scan_win467 <= 32'd0; scan_win468 <= 32'd0; scan_win469 <= 32'd0; scan_win470 <= 32'd0; scan_win471 <= 32'd0; scan_win472 <= 32'd0; scan_win473 <= 32'd0; scan_win474 <= 32'd0; scan_win475 <= 32'd0; scan_win476 <= 32'd0; scan_win477 <= 32'd0; scan_win478 <= 32'd0; scan_win479 <= 32'd0; scan_win480 <= 32'd0; scan_win481 <= 32'd0; scan_win482 <= 32'd0; scan_win483 <= 32'd0; scan_win484 <= 32'd0; scan_win485 <= 32'd0; scan_win486 <= 32'd0; scan_win487 <= 32'd0; scan_win488 <= 32'd0; scan_win489 <= 32'd0; scan_win490 <= 32'd0; scan_win491 <= 32'd0; scan_win492 <= 32'd0; scan_win493 <= 32'd0; scan_win494 <= 32'd0; scan_win495 <= 32'd0; scan_win496 <= 32'd0; scan_win497 <= 32'd0; scan_win498 <= 32'd0; scan_win499 <= 32'd0; scan_win500 <= 32'd0; scan_win501 <= 32'd0; scan_win502 <= 32'd0; scan_win503 <= 32'd0; scan_win504 <= 32'd0; scan_win505 <= 32'd0; scan_win506 <= 32'd0; scan_win507 <= 32'd0; scan_win508 <= 32'd0; scan_win509 <= 32'd0; scan_win510 <= 32'd0; scan_win511 <= 32'd0; scan_win512 <= 32'd0; scan_win513 <= 32'd0; scan_win514 <= 32'd0; scan_win515 <= 32'd0; scan_win516 <= 32'd0; scan_win517 <= 32'd0; scan_win518 <= 32'd0; scan_win519 <= 32'd0; scan_win520 <= 32'd0; scan_win521 <= 32'd0; scan_win522 <= 32'd0; scan_win523 <= 32'd0; scan_win524 <= 32'd0; scan_win525 <= 32'd0; scan_win526 <= 32'd0; scan_win527 <= 32'd0; scan_win528 <= 32'd0; scan_win529 <= 32'd0; scan_win530 <= 32'd0; scan_win531 <= 32'd0; scan_win532 <= 32'd0; scan_win533 <= 32'd0; scan_win534 <= 32'd0; scan_win535 <= 32'd0; scan_win536 <= 32'd0; scan_win537 <= 32'd0; scan_win538 <= 32'd0; scan_win539 <= 32'd0; scan_win540 <= 32'd0; scan_win541 <= 32'd0; scan_win542 <= 32'd0; scan_win543 <= 32'd0; scan_win544 <= 32'd0; scan_win545 <= 32'd0; scan_win546 <= 32'd0; scan_win547 <= 32'd0; scan_win548 <= 32'd0; scan_win549 <= 32'd0; scan_win550 <= 32'd0; scan_win551 <= 32'd0; scan_win552 <= 32'd0; scan_win553 <= 32'd0; scan_win554 <= 32'd0; scan_win555 <= 32'd0; scan_win556 <= 32'd0; scan_win557 <= 32'd0; scan_win558 <= 32'd0; scan_win559 <= 32'd0; scan_win560 <= 32'd0; scan_win561 <= 32'd0; scan_win562 <= 32'd0; scan_win563 <= 32'd0; scan_win564 <= 32'd0; scan_win565 <= 32'd0; scan_win566 <= 32'd0; scan_win567 <= 32'd0; scan_win568 <= 32'd0; scan_win569 <= 32'd0; scan_win570 <= 32'd0; scan_win571 <= 32'd0; scan_win572 <= 32'd0; scan_win573 <= 32'd0; scan_win574 <= 32'd0; scan_win575 <= 32'd0; scan_win576 <= 32'd0; scan_win577 <= 32'd0; scan_win578 <= 32'd0; scan_win579 <= 32'd0; scan_win580 <= 32'd0; scan_win581 <= 32'd0; scan_win582 <= 32'd0; scan_win583 <= 32'd0; scan_win584 <= 32'd0; scan_win585 <= 32'd0; scan_win586 <= 32'd0; scan_win587 <= 32'd0; scan_win588 <= 32'd0; scan_win589 <= 32'd0; scan_win590 <= 32'd0; scan_win591 <= 32'd0; scan_win592 <= 32'd0; scan_win593 <= 32'd0; scan_win594 <= 32'd0; scan_win595 <= 32'd0; scan_win596 <= 32'd0; scan_win597 <= 32'd0; scan_win598 <= 32'd0; scan_win599 <= 32'd0; scan_win600 <= 32'd0; 
      scan_win601 <= 32'd0; scan_win602 <= 32'd0; scan_win603 <= 32'd0; scan_win604 <= 32'd0; scan_win605 <= 32'd0; scan_win606 <= 32'd0; scan_win607 <= 32'd0; scan_win608 <= 32'd0; scan_win609 <= 32'd0; scan_win610 <= 32'd0; scan_win611 <= 32'd0; scan_win612 <= 32'd0; scan_win613 <= 32'd0; scan_win614 <= 32'd0; scan_win615 <= 32'd0; scan_win616 <= 32'd0; scan_win617 <= 32'd0; scan_win618 <= 32'd0; scan_win619 <= 32'd0; scan_win620 <= 32'd0; scan_win621 <= 32'd0; scan_win622 <= 32'd0; scan_win623 <= 32'd0; scan_win624 <= 32'd0; scan_win625 <= 32'd0; scan_win626 <= 32'd0; scan_win627 <= 32'd0; scan_win628 <= 32'd0; scan_win629 <= 32'd0; scan_win630 <= 32'd0; scan_win631 <= 32'd0; scan_win632 <= 32'd0; scan_win633 <= 32'd0; scan_win634 <= 32'd0; scan_win635 <= 32'd0; scan_win636 <= 32'd0; scan_win637 <= 32'd0; scan_win638 <= 32'd0; scan_win639 <= 32'd0; scan_win640 <= 32'd0; scan_win641 <= 32'd0; scan_win642 <= 32'd0; scan_win643 <= 32'd0; scan_win644 <= 32'd0; scan_win645 <= 32'd0; scan_win646 <= 32'd0; scan_win647 <= 32'd0; scan_win648 <= 32'd0; scan_win649 <= 32'd0; scan_win650 <= 32'd0; scan_win651 <= 32'd0; scan_win652 <= 32'd0; scan_win653 <= 32'd0; scan_win654 <= 32'd0; scan_win655 <= 32'd0; scan_win656 <= 32'd0; scan_win657 <= 32'd0; scan_win658 <= 32'd0; scan_win659 <= 32'd0; scan_win660 <= 32'd0; scan_win661 <= 32'd0; scan_win662 <= 32'd0; scan_win663 <= 32'd0; scan_win664 <= 32'd0; scan_win665 <= 32'd0; scan_win666 <= 32'd0; scan_win667 <= 32'd0; scan_win668 <= 32'd0; scan_win669 <= 32'd0; scan_win670 <= 32'd0; scan_win671 <= 32'd0; scan_win672 <= 32'd0; scan_win673 <= 32'd0; scan_win674 <= 32'd0; scan_win675 <= 32'd0; scan_win676 <= 32'd0; scan_win677 <= 32'd0; scan_win678 <= 32'd0; scan_win679 <= 32'd0; scan_win680 <= 32'd0; scan_win681 <= 32'd0; scan_win682 <= 32'd0; scan_win683 <= 32'd0; scan_win684 <= 32'd0; scan_win685 <= 32'd0; scan_win686 <= 32'd0; scan_win687 <= 32'd0; scan_win688 <= 32'd0; scan_win689 <= 32'd0; scan_win690 <= 32'd0; scan_win691 <= 32'd0; scan_win692 <= 32'd0; scan_win693 <= 32'd0; scan_win694 <= 32'd0; scan_win695 <= 32'd0; scan_win696 <= 32'd0; scan_win697 <= 32'd0; scan_win698 <= 32'd0; scan_win699 <= 32'd0; scan_win700 <= 32'd0; scan_win701 <= 32'd0; scan_win702 <= 32'd0; scan_win703 <= 32'd0; scan_win704 <= 32'd0; scan_win705 <= 32'd0; scan_win706 <= 32'd0; scan_win707 <= 32'd0; scan_win708 <= 32'd0; scan_win709 <= 32'd0; scan_win710 <= 32'd0; scan_win711 <= 32'd0; scan_win712 <= 32'd0; scan_win713 <= 32'd0; scan_win714 <= 32'd0; scan_win715 <= 32'd0; scan_win716 <= 32'd0; scan_win717 <= 32'd0; scan_win718 <= 32'd0; scan_win719 <= 32'd0; scan_win720 <= 32'd0; scan_win721 <= 32'd0; scan_win722 <= 32'd0; scan_win723 <= 32'd0; scan_win724 <= 32'd0; scan_win725 <= 32'd0; scan_win726 <= 32'd0; scan_win727 <= 32'd0; scan_win728 <= 32'd0; scan_win729 <= 32'd0; scan_win730 <= 32'd0; scan_win731 <= 32'd0; scan_win732 <= 32'd0; scan_win733 <= 32'd0; scan_win734 <= 32'd0; scan_win735 <= 32'd0; scan_win736 <= 32'd0; scan_win737 <= 32'd0; scan_win738 <= 32'd0; scan_win739 <= 32'd0; scan_win740 <= 32'd0; scan_win741 <= 32'd0; scan_win742 <= 32'd0; scan_win743 <= 32'd0; scan_win744 <= 32'd0; scan_win745 <= 32'd0; scan_win746 <= 32'd0; scan_win747 <= 32'd0; scan_win748 <= 32'd0; scan_win749 <= 32'd0; scan_win750 <= 32'd0; scan_win751 <= 32'd0; scan_win752 <= 32'd0; scan_win753 <= 32'd0; scan_win754 <= 32'd0; scan_win755 <= 32'd0; scan_win756 <= 32'd0; scan_win757 <= 32'd0; scan_win758 <= 32'd0; scan_win759 <= 32'd0; scan_win760 <= 32'd0; scan_win761 <= 32'd0; scan_win762 <= 32'd0; scan_win763 <= 32'd0; scan_win764 <= 32'd0; scan_win765 <= 32'd0; scan_win766 <= 32'd0; scan_win767 <= 32'd0; scan_win768 <= 32'd0; scan_win769 <= 32'd0; scan_win770 <= 32'd0; scan_win771 <= 32'd0; scan_win772 <= 32'd0; scan_win773 <= 32'd0; scan_win774 <= 32'd0; scan_win775 <= 32'd0; scan_win776 <= 32'd0; scan_win777 <= 32'd0; scan_win778 <= 32'd0; scan_win779 <= 32'd0; scan_win780 <= 32'd0; scan_win781 <= 32'd0; scan_win782 <= 32'd0; scan_win783 <= 32'd0; scan_win784 <= 32'd0; scan_win785 <= 32'd0; scan_win786 <= 32'd0; scan_win787 <= 32'd0; scan_win788 <= 32'd0; scan_win789 <= 32'd0; scan_win790 <= 32'd0; scan_win791 <= 32'd0; scan_win792 <= 32'd0; scan_win793 <= 32'd0; scan_win794 <= 32'd0; scan_win795 <= 32'd0; scan_win796 <= 32'd0; scan_win797 <= 32'd0; scan_win798 <= 32'd0; scan_win799 <= 32'd0; scan_win800 <= 32'd0; 
      scan_win801 <= 32'd0; scan_win802 <= 32'd0; scan_win803 <= 32'd0; scan_win804 <= 32'd0; scan_win805 <= 32'd0; scan_win806 <= 32'd0; scan_win807 <= 32'd0; scan_win808 <= 32'd0; scan_win809 <= 32'd0; scan_win810 <= 32'd0; scan_win811 <= 32'd0; scan_win812 <= 32'd0; scan_win813 <= 32'd0; scan_win814 <= 32'd0; scan_win815 <= 32'd0; scan_win816 <= 32'd0; scan_win817 <= 32'd0; scan_win818 <= 32'd0; scan_win819 <= 32'd0; scan_win820 <= 32'd0; scan_win821 <= 32'd0; scan_win822 <= 32'd0; scan_win823 <= 32'd0; scan_win824 <= 32'd0; scan_win825 <= 32'd0; scan_win826 <= 32'd0; scan_win827 <= 32'd0; scan_win828 <= 32'd0; scan_win829 <= 32'd0; scan_win830 <= 32'd0; scan_win831 <= 32'd0; scan_win832 <= 32'd0; scan_win833 <= 32'd0; scan_win834 <= 32'd0; scan_win835 <= 32'd0; scan_win836 <= 32'd0; scan_win837 <= 32'd0; scan_win838 <= 32'd0; scan_win839 <= 32'd0; scan_win840 <= 32'd0; scan_win841 <= 32'd0; scan_win842 <= 32'd0; scan_win843 <= 32'd0; scan_win844 <= 32'd0; scan_win845 <= 32'd0; scan_win846 <= 32'd0; scan_win847 <= 32'd0; scan_win848 <= 32'd0; scan_win849 <= 32'd0; scan_win850 <= 32'd0; scan_win851 <= 32'd0; scan_win852 <= 32'd0; scan_win853 <= 32'd0; scan_win854 <= 32'd0; scan_win855 <= 32'd0; scan_win856 <= 32'd0; scan_win857 <= 32'd0; scan_win858 <= 32'd0; scan_win859 <= 32'd0; scan_win860 <= 32'd0; scan_win861 <= 32'd0; scan_win862 <= 32'd0; scan_win863 <= 32'd0; scan_win864 <= 32'd0; scan_win865 <= 32'd0; scan_win866 <= 32'd0; scan_win867 <= 32'd0; scan_win868 <= 32'd0; scan_win869 <= 32'd0; scan_win870 <= 32'd0; scan_win871 <= 32'd0; scan_win872 <= 32'd0; scan_win873 <= 32'd0; scan_win874 <= 32'd0; scan_win875 <= 32'd0; scan_win876 <= 32'd0; scan_win877 <= 32'd0; scan_win878 <= 32'd0; scan_win879 <= 32'd0; scan_win880 <= 32'd0; scan_win881 <= 32'd0; scan_win882 <= 32'd0; scan_win883 <= 32'd0; scan_win884 <= 32'd0; scan_win885 <= 32'd0; scan_win886 <= 32'd0; scan_win887 <= 32'd0; scan_win888 <= 32'd0; scan_win889 <= 32'd0; scan_win890 <= 32'd0; scan_win891 <= 32'd0; scan_win892 <= 32'd0; scan_win893 <= 32'd0; scan_win894 <= 32'd0; scan_win895 <= 32'd0; scan_win896 <= 32'd0; scan_win897 <= 32'd0; scan_win898 <= 32'd0; scan_win899 <= 32'd0; scan_win900 <= 32'd0; scan_win901 <= 32'd0; scan_win902 <= 32'd0; scan_win903 <= 32'd0; scan_win904 <= 32'd0; scan_win905 <= 32'd0; scan_win906 <= 32'd0; scan_win907 <= 32'd0; scan_win908 <= 32'd0; scan_win909 <= 32'd0; scan_win910 <= 32'd0; scan_win911 <= 32'd0; scan_win912 <= 32'd0; scan_win913 <= 32'd0; scan_win914 <= 32'd0; scan_win915 <= 32'd0; scan_win916 <= 32'd0; scan_win917 <= 32'd0; scan_win918 <= 32'd0; scan_win919 <= 32'd0; scan_win920 <= 32'd0; scan_win921 <= 32'd0; scan_win922 <= 32'd0; scan_win923 <= 32'd0; scan_win924 <= 32'd0; scan_win925 <= 32'd0; scan_win926 <= 32'd0; scan_win927 <= 32'd0; scan_win928 <= 32'd0; scan_win929 <= 32'd0; scan_win930 <= 32'd0; scan_win931 <= 32'd0; scan_win932 <= 32'd0; scan_win933 <= 32'd0; scan_win934 <= 32'd0; scan_win935 <= 32'd0; scan_win936 <= 32'd0; scan_win937 <= 32'd0; scan_win938 <= 32'd0; scan_win939 <= 32'd0; scan_win940 <= 32'd0; scan_win941 <= 32'd0; scan_win942 <= 32'd0; scan_win943 <= 32'd0; scan_win944 <= 32'd0; scan_win945 <= 32'd0; scan_win946 <= 32'd0; scan_win947 <= 32'd0; scan_win948 <= 32'd0; scan_win949 <= 32'd0; scan_win950 <= 32'd0; scan_win951 <= 32'd0; scan_win952 <= 32'd0; scan_win953 <= 32'd0; scan_win954 <= 32'd0; scan_win955 <= 32'd0; scan_win956 <= 32'd0; scan_win957 <= 32'd0; scan_win958 <= 32'd0; scan_win959 <= 32'd0; scan_win960 <= 32'd0; scan_win961 <= 32'd0; scan_win962 <= 32'd0; scan_win963 <= 32'd0; scan_win964 <= 32'd0; scan_win965 <= 32'd0; scan_win966 <= 32'd0; scan_win967 <= 32'd0; scan_win968 <= 32'd0; scan_win969 <= 32'd0; scan_win970 <= 32'd0; scan_win971 <= 32'd0; scan_win972 <= 32'd0; scan_win973 <= 32'd0; scan_win974 <= 32'd0; scan_win975 <= 32'd0; scan_win976 <= 32'd0; scan_win977 <= 32'd0; scan_win978 <= 32'd0; scan_win979 <= 32'd0; scan_win980 <= 32'd0; scan_win981 <= 32'd0; scan_win982 <= 32'd0; scan_win983 <= 32'd0; scan_win984 <= 32'd0; scan_win985 <= 32'd0; scan_win986 <= 32'd0; scan_win987 <= 32'd0; scan_win988 <= 32'd0; scan_win989 <= 32'd0; scan_win990 <= 32'd0; scan_win991 <= 32'd0; scan_win992 <= 32'd0; scan_win993 <= 32'd0; scan_win994 <= 32'd0; scan_win995 <= 32'd0; scan_win996 <= 32'd0; scan_win997 <= 32'd0; scan_win998 <= 32'd0; scan_win999 <= 32'd0; scan_win1000 <= 32'd0; 
      scan_win1001 <= 32'd0; scan_win1002 <= 32'd0; scan_win1003 <= 32'd0; scan_win1004 <= 32'd0; scan_win1005 <= 32'd0; scan_win1006 <= 32'd0; scan_win1007 <= 32'd0; scan_win1008 <= 32'd0; scan_win1009 <= 32'd0; scan_win1010 <= 32'd0; scan_win1011 <= 32'd0; scan_win1012 <= 32'd0; scan_win1013 <= 32'd0; scan_win1014 <= 32'd0; scan_win1015 <= 32'd0; scan_win1016 <= 32'd0; scan_win1017 <= 32'd0; scan_win1018 <= 32'd0; scan_win1019 <= 32'd0; scan_win1020 <= 32'd0; scan_win1021 <= 32'd0; scan_win1022 <= 32'd0; scan_win1023 <= 32'd0; scan_win1024 <= 32'd0; scan_win1025 <= 32'd0; scan_win1026 <= 32'd0; scan_win1027 <= 32'd0; scan_win1028 <= 32'd0; scan_win1029 <= 32'd0; scan_win1030 <= 32'd0; scan_win1031 <= 32'd0; scan_win1032 <= 32'd0; scan_win1033 <= 32'd0; scan_win1034 <= 32'd0; scan_win1035 <= 32'd0; scan_win1036 <= 32'd0; scan_win1037 <= 32'd0; scan_win1038 <= 32'd0; scan_win1039 <= 32'd0; scan_win1040 <= 32'd0; scan_win1041 <= 32'd0; scan_win1042 <= 32'd0; scan_win1043 <= 32'd0; scan_win1044 <= 32'd0; scan_win1045 <= 32'd0; scan_win1046 <= 32'd0; scan_win1047 <= 32'd0; scan_win1048 <= 32'd0; scan_win1049 <= 32'd0; scan_win1050 <= 32'd0; scan_win1051 <= 32'd0; scan_win1052 <= 32'd0; scan_win1053 <= 32'd0; scan_win1054 <= 32'd0; scan_win1055 <= 32'd0; scan_win1056 <= 32'd0; scan_win1057 <= 32'd0; scan_win1058 <= 32'd0; scan_win1059 <= 32'd0; scan_win1060 <= 32'd0; scan_win1061 <= 32'd0; scan_win1062 <= 32'd0; scan_win1063 <= 32'd0; scan_win1064 <= 32'd0; scan_win1065 <= 32'd0; scan_win1066 <= 32'd0; scan_win1067 <= 32'd0; scan_win1068 <= 32'd0; scan_win1069 <= 32'd0; scan_win1070 <= 32'd0; scan_win1071 <= 32'd0; scan_win1072 <= 32'd0; scan_win1073 <= 32'd0; scan_win1074 <= 32'd0; scan_win1075 <= 32'd0; scan_win1076 <= 32'd0; scan_win1077 <= 32'd0; scan_win1078 <= 32'd0; scan_win1079 <= 32'd0; scan_win1080 <= 32'd0; scan_win1081 <= 32'd0; scan_win1082 <= 32'd0; scan_win1083 <= 32'd0; scan_win1084 <= 32'd0; scan_win1085 <= 32'd0; scan_win1086 <= 32'd0; scan_win1087 <= 32'd0; scan_win1088 <= 32'd0; scan_win1089 <= 32'd0; scan_win1090 <= 32'd0; scan_win1091 <= 32'd0; scan_win1092 <= 32'd0; scan_win1093 <= 32'd0; scan_win1094 <= 32'd0; scan_win1095 <= 32'd0; scan_win1096 <= 32'd0; scan_win1097 <= 32'd0; scan_win1098 <= 32'd0; scan_win1099 <= 32'd0; scan_win1100 <= 32'd0; scan_win1101 <= 32'd0; scan_win1102 <= 32'd0; scan_win1103 <= 32'd0; scan_win1104 <= 32'd0; scan_win1105 <= 32'd0; scan_win1106 <= 32'd0; scan_win1107 <= 32'd0; scan_win1108 <= 32'd0; scan_win1109 <= 32'd0; scan_win1110 <= 32'd0; scan_win1111 <= 32'd0; scan_win1112 <= 32'd0; scan_win1113 <= 32'd0; scan_win1114 <= 32'd0; scan_win1115 <= 32'd0; scan_win1116 <= 32'd0; scan_win1117 <= 32'd0; scan_win1118 <= 32'd0; scan_win1119 <= 32'd0; scan_win1120 <= 32'd0; scan_win1121 <= 32'd0; scan_win1122 <= 32'd0; scan_win1123 <= 32'd0; scan_win1124 <= 32'd0; scan_win1125 <= 32'd0; scan_win1126 <= 32'd0; scan_win1127 <= 32'd0; scan_win1128 <= 32'd0; scan_win1129 <= 32'd0; scan_win1130 <= 32'd0; scan_win1131 <= 32'd0; scan_win1132 <= 32'd0; scan_win1133 <= 32'd0; scan_win1134 <= 32'd0; scan_win1135 <= 32'd0; scan_win1136 <= 32'd0; scan_win1137 <= 32'd0; scan_win1138 <= 32'd0; scan_win1139 <= 32'd0; scan_win1140 <= 32'd0; scan_win1141 <= 32'd0; scan_win1142 <= 32'd0; scan_win1143 <= 32'd0; scan_win1144 <= 32'd0; scan_win1145 <= 32'd0; scan_win1146 <= 32'd0; scan_win1147 <= 32'd0; scan_win1148 <= 32'd0; scan_win1149 <= 32'd0; scan_win1150 <= 32'd0; scan_win1151 <= 32'd0; scan_win1152 <= 32'd0; scan_win1153 <= 32'd0; scan_win1154 <= 32'd0; scan_win1155 <= 32'd0; scan_win1156 <= 32'd0; scan_win1157 <= 32'd0; scan_win1158 <= 32'd0; scan_win1159 <= 32'd0; scan_win1160 <= 32'd0; scan_win1161 <= 32'd0; scan_win1162 <= 32'd0; scan_win1163 <= 32'd0; scan_win1164 <= 32'd0; scan_win1165 <= 32'd0; scan_win1166 <= 32'd0; scan_win1167 <= 32'd0; scan_win1168 <= 32'd0; scan_win1169 <= 32'd0; scan_win1170 <= 32'd0; scan_win1171 <= 32'd0; scan_win1172 <= 32'd0; scan_win1173 <= 32'd0; scan_win1174 <= 32'd0; scan_win1175 <= 32'd0; scan_win1176 <= 32'd0; scan_win1177 <= 32'd0; scan_win1178 <= 32'd0; scan_win1179 <= 32'd0; scan_win1180 <= 32'd0; scan_win1181 <= 32'd0; scan_win1182 <= 32'd0; scan_win1183 <= 32'd0; scan_win1184 <= 32'd0; scan_win1185 <= 32'd0; scan_win1186 <= 32'd0; scan_win1187 <= 32'd0; scan_win1188 <= 32'd0; scan_win1189 <= 32'd0; scan_win1190 <= 32'd0; scan_win1191 <= 32'd0; scan_win1192 <= 32'd0; scan_win1193 <= 32'd0; scan_win1194 <= 32'd0; scan_win1195 <= 32'd0; scan_win1196 <= 32'd0; scan_win1197 <= 32'd0; scan_win1198 <= 32'd0; scan_win1199 <= 32'd0; scan_win1200 <= 32'd0; 
      scan_win1201 <= 32'd0; scan_win1202 <= 32'd0; scan_win1203 <= 32'd0; scan_win1204 <= 32'd0; scan_win1205 <= 32'd0; scan_win1206 <= 32'd0; scan_win1207 <= 32'd0; scan_win1208 <= 32'd0; scan_win1209 <= 32'd0; scan_win1210 <= 32'd0; scan_win1211 <= 32'd0; scan_win1212 <= 32'd0; scan_win1213 <= 32'd0; scan_win1214 <= 32'd0; scan_win1215 <= 32'd0; scan_win1216 <= 32'd0; scan_win1217 <= 32'd0; scan_win1218 <= 32'd0; scan_win1219 <= 32'd0; scan_win1220 <= 32'd0; scan_win1221 <= 32'd0; scan_win1222 <= 32'd0; scan_win1223 <= 32'd0; scan_win1224 <= 32'd0; scan_win1225 <= 32'd0; scan_win1226 <= 32'd0; scan_win1227 <= 32'd0; scan_win1228 <= 32'd0; scan_win1229 <= 32'd0; scan_win1230 <= 32'd0; scan_win1231 <= 32'd0; scan_win1232 <= 32'd0; scan_win1233 <= 32'd0; scan_win1234 <= 32'd0; scan_win1235 <= 32'd0; scan_win1236 <= 32'd0; scan_win1237 <= 32'd0; scan_win1238 <= 32'd0; scan_win1239 <= 32'd0; scan_win1240 <= 32'd0; scan_win1241 <= 32'd0; scan_win1242 <= 32'd0; scan_win1243 <= 32'd0; scan_win1244 <= 32'd0; scan_win1245 <= 32'd0; scan_win1246 <= 32'd0; scan_win1247 <= 32'd0; scan_win1248 <= 32'd0; scan_win1249 <= 32'd0; scan_win1250 <= 32'd0; scan_win1251 <= 32'd0; scan_win1252 <= 32'd0; scan_win1253 <= 32'd0; scan_win1254 <= 32'd0; scan_win1255 <= 32'd0; scan_win1256 <= 32'd0; scan_win1257 <= 32'd0; scan_win1258 <= 32'd0; scan_win1259 <= 32'd0; scan_win1260 <= 32'd0; scan_win1261 <= 32'd0; scan_win1262 <= 32'd0; scan_win1263 <= 32'd0; scan_win1264 <= 32'd0; scan_win1265 <= 32'd0; scan_win1266 <= 32'd0; scan_win1267 <= 32'd0; scan_win1268 <= 32'd0; scan_win1269 <= 32'd0; scan_win1270 <= 32'd0; scan_win1271 <= 32'd0; scan_win1272 <= 32'd0; scan_win1273 <= 32'd0; scan_win1274 <= 32'd0; scan_win1275 <= 32'd0; scan_win1276 <= 32'd0; scan_win1277 <= 32'd0; scan_win1278 <= 32'd0; scan_win1279 <= 32'd0; scan_win1280 <= 32'd0; scan_win1281 <= 32'd0; scan_win1282 <= 32'd0; scan_win1283 <= 32'd0; scan_win1284 <= 32'd0; scan_win1285 <= 32'd0; scan_win1286 <= 32'd0; scan_win1287 <= 32'd0; scan_win1288 <= 32'd0; scan_win1289 <= 32'd0; scan_win1290 <= 32'd0; scan_win1291 <= 32'd0; scan_win1292 <= 32'd0; scan_win1293 <= 32'd0; scan_win1294 <= 32'd0; scan_win1295 <= 32'd0; scan_win1296 <= 32'd0; scan_win1297 <= 32'd0; scan_win1298 <= 32'd0; scan_win1299 <= 32'd0; scan_win1300 <= 32'd0; scan_win1301 <= 32'd0; scan_win1302 <= 32'd0; scan_win1303 <= 32'd0; scan_win1304 <= 32'd0; scan_win1305 <= 32'd0; scan_win1306 <= 32'd0; scan_win1307 <= 32'd0; scan_win1308 <= 32'd0; scan_win1309 <= 32'd0; scan_win1310 <= 32'd0; scan_win1311 <= 32'd0; scan_win1312 <= 32'd0; scan_win1313 <= 32'd0; scan_win1314 <= 32'd0; scan_win1315 <= 32'd0; scan_win1316 <= 32'd0; scan_win1317 <= 32'd0; scan_win1318 <= 32'd0; scan_win1319 <= 32'd0; scan_win1320 <= 32'd0; scan_win1321 <= 32'd0; scan_win1322 <= 32'd0; scan_win1323 <= 32'd0; scan_win1324 <= 32'd0; scan_win1325 <= 32'd0; scan_win1326 <= 32'd0; scan_win1327 <= 32'd0; scan_win1328 <= 32'd0; scan_win1329 <= 32'd0; scan_win1330 <= 32'd0; scan_win1331 <= 32'd0; scan_win1332 <= 32'd0; scan_win1333 <= 32'd0; scan_win1334 <= 32'd0; scan_win1335 <= 32'd0; scan_win1336 <= 32'd0; scan_win1337 <= 32'd0; scan_win1338 <= 32'd0; scan_win1339 <= 32'd0; scan_win1340 <= 32'd0; scan_win1341 <= 32'd0; scan_win1342 <= 32'd0; scan_win1343 <= 32'd0; scan_win1344 <= 32'd0; scan_win1345 <= 32'd0; scan_win1346 <= 32'd0; scan_win1347 <= 32'd0; scan_win1348 <= 32'd0; scan_win1349 <= 32'd0; scan_win1350 <= 32'd0; scan_win1351 <= 32'd0; scan_win1352 <= 32'd0; scan_win1353 <= 32'd0; scan_win1354 <= 32'd0; scan_win1355 <= 32'd0; scan_win1356 <= 32'd0; scan_win1357 <= 32'd0; scan_win1358 <= 32'd0; scan_win1359 <= 32'd0; scan_win1360 <= 32'd0; scan_win1361 <= 32'd0; scan_win1362 <= 32'd0; scan_win1363 <= 32'd0; scan_win1364 <= 32'd0; scan_win1365 <= 32'd0; scan_win1366 <= 32'd0; scan_win1367 <= 32'd0; scan_win1368 <= 32'd0; scan_win1369 <= 32'd0; scan_win1370 <= 32'd0; scan_win1371 <= 32'd0; scan_win1372 <= 32'd0; scan_win1373 <= 32'd0; scan_win1374 <= 32'd0; scan_win1375 <= 32'd0; scan_win1376 <= 32'd0; scan_win1377 <= 32'd0; scan_win1378 <= 32'd0; scan_win1379 <= 32'd0; scan_win1380 <= 32'd0; scan_win1381 <= 32'd0; scan_win1382 <= 32'd0; scan_win1383 <= 32'd0; scan_win1384 <= 32'd0; scan_win1385 <= 32'd0; scan_win1386 <= 32'd0; scan_win1387 <= 32'd0; scan_win1388 <= 32'd0; scan_win1389 <= 32'd0; scan_win1390 <= 32'd0; scan_win1391 <= 32'd0; scan_win1392 <= 32'd0; scan_win1393 <= 32'd0; scan_win1394 <= 32'd0; scan_win1395 <= 32'd0; scan_win1396 <= 32'd0; scan_win1397 <= 32'd0; scan_win1398 <= 32'd0; scan_win1399 <= 32'd0; scan_win1400 <= 32'd0; 
      scan_win1401 <= 32'd0; scan_win1402 <= 32'd0; scan_win1403 <= 32'd0; scan_win1404 <= 32'd0; scan_win1405 <= 32'd0; scan_win1406 <= 32'd0; scan_win1407 <= 32'd0; scan_win1408 <= 32'd0; scan_win1409 <= 32'd0; scan_win1410 <= 32'd0; scan_win1411 <= 32'd0; scan_win1412 <= 32'd0; scan_win1413 <= 32'd0; scan_win1414 <= 32'd0; scan_win1415 <= 32'd0; scan_win1416 <= 32'd0; scan_win1417 <= 32'd0; scan_win1418 <= 32'd0; scan_win1419 <= 32'd0; scan_win1420 <= 32'd0; scan_win1421 <= 32'd0; scan_win1422 <= 32'd0; scan_win1423 <= 32'd0; scan_win1424 <= 32'd0; scan_win1425 <= 32'd0; scan_win1426 <= 32'd0; scan_win1427 <= 32'd0; scan_win1428 <= 32'd0; scan_win1429 <= 32'd0; scan_win1430 <= 32'd0; scan_win1431 <= 32'd0; scan_win1432 <= 32'd0; scan_win1433 <= 32'd0; scan_win1434 <= 32'd0; scan_win1435 <= 32'd0; scan_win1436 <= 32'd0; scan_win1437 <= 32'd0; scan_win1438 <= 32'd0; scan_win1439 <= 32'd0; scan_win1440 <= 32'd0; scan_win1441 <= 32'd0; scan_win1442 <= 32'd0; scan_win1443 <= 32'd0; scan_win1444 <= 32'd0; scan_win1445 <= 32'd0; scan_win1446 <= 32'd0; scan_win1447 <= 32'd0; scan_win1448 <= 32'd0; scan_win1449 <= 32'd0; scan_win1450 <= 32'd0; scan_win1451 <= 32'd0; scan_win1452 <= 32'd0; scan_win1453 <= 32'd0; scan_win1454 <= 32'd0; scan_win1455 <= 32'd0; scan_win1456 <= 32'd0; scan_win1457 <= 32'd0; scan_win1458 <= 32'd0; scan_win1459 <= 32'd0; scan_win1460 <= 32'd0; scan_win1461 <= 32'd0; scan_win1462 <= 32'd0; scan_win1463 <= 32'd0; scan_win1464 <= 32'd0; scan_win1465 <= 32'd0; scan_win1466 <= 32'd0; scan_win1467 <= 32'd0; scan_win1468 <= 32'd0; scan_win1469 <= 32'd0; scan_win1470 <= 32'd0; scan_win1471 <= 32'd0; scan_win1472 <= 32'd0; scan_win1473 <= 32'd0; scan_win1474 <= 32'd0; scan_win1475 <= 32'd0; scan_win1476 <= 32'd0; scan_win1477 <= 32'd0; scan_win1478 <= 32'd0; scan_win1479 <= 32'd0; scan_win1480 <= 32'd0; scan_win1481 <= 32'd0; scan_win1482 <= 32'd0; scan_win1483 <= 32'd0; scan_win1484 <= 32'd0; scan_win1485 <= 32'd0; scan_win1486 <= 32'd0; scan_win1487 <= 32'd0; scan_win1488 <= 32'd0; scan_win1489 <= 32'd0; scan_win1490 <= 32'd0; scan_win1491 <= 32'd0; scan_win1492 <= 32'd0; scan_win1493 <= 32'd0; scan_win1494 <= 32'd0; scan_win1495 <= 32'd0; scan_win1496 <= 32'd0; scan_win1497 <= 32'd0; scan_win1498 <= 32'd0; scan_win1499 <= 32'd0; scan_win1500 <= 32'd0; scan_win1501 <= 32'd0; scan_win1502 <= 32'd0; scan_win1503 <= 32'd0; scan_win1504 <= 32'd0; scan_win1505 <= 32'd0; scan_win1506 <= 32'd0; scan_win1507 <= 32'd0; scan_win1508 <= 32'd0; scan_win1509 <= 32'd0; scan_win1510 <= 32'd0; scan_win1511 <= 32'd0; scan_win1512 <= 32'd0; scan_win1513 <= 32'd0; scan_win1514 <= 32'd0; scan_win1515 <= 32'd0; scan_win1516 <= 32'd0; scan_win1517 <= 32'd0; scan_win1518 <= 32'd0; scan_win1519 <= 32'd0; scan_win1520 <= 32'd0; scan_win1521 <= 32'd0; scan_win1522 <= 32'd0; scan_win1523 <= 32'd0; scan_win1524 <= 32'd0; scan_win1525 <= 32'd0; scan_win1526 <= 32'd0; scan_win1527 <= 32'd0; scan_win1528 <= 32'd0; scan_win1529 <= 32'd0; scan_win1530 <= 32'd0; scan_win1531 <= 32'd0; scan_win1532 <= 32'd0; scan_win1533 <= 32'd0; scan_win1534 <= 32'd0; scan_win1535 <= 32'd0; scan_win1536 <= 32'd0; scan_win1537 <= 32'd0; scan_win1538 <= 32'd0; scan_win1539 <= 32'd0; scan_win1540 <= 32'd0; scan_win1541 <= 32'd0; scan_win1542 <= 32'd0; scan_win1543 <= 32'd0; scan_win1544 <= 32'd0; scan_win1545 <= 32'd0; scan_win1546 <= 32'd0; scan_win1547 <= 32'd0; scan_win1548 <= 32'd0; scan_win1549 <= 32'd0; scan_win1550 <= 32'd0; scan_win1551 <= 32'd0; scan_win1552 <= 32'd0; scan_win1553 <= 32'd0; scan_win1554 <= 32'd0; scan_win1555 <= 32'd0; scan_win1556 <= 32'd0; scan_win1557 <= 32'd0; scan_win1558 <= 32'd0; scan_win1559 <= 32'd0; scan_win1560 <= 32'd0; scan_win1561 <= 32'd0; scan_win1562 <= 32'd0; scan_win1563 <= 32'd0; scan_win1564 <= 32'd0; scan_win1565 <= 32'd0; scan_win1566 <= 32'd0; scan_win1567 <= 32'd0; scan_win1568 <= 32'd0; scan_win1569 <= 32'd0; scan_win1570 <= 32'd0; scan_win1571 <= 32'd0; scan_win1572 <= 32'd0; scan_win1573 <= 32'd0; scan_win1574 <= 32'd0; scan_win1575 <= 32'd0; scan_win1576 <= 32'd0; scan_win1577 <= 32'd0; scan_win1578 <= 32'd0; scan_win1579 <= 32'd0; scan_win1580 <= 32'd0; scan_win1581 <= 32'd0; scan_win1582 <= 32'd0; scan_win1583 <= 32'd0; scan_win1584 <= 32'd0; scan_win1585 <= 32'd0; scan_win1586 <= 32'd0; scan_win1587 <= 32'd0; scan_win1588 <= 32'd0; scan_win1589 <= 32'd0; scan_win1590 <= 32'd0; scan_win1591 <= 32'd0; scan_win1592 <= 32'd0; scan_win1593 <= 32'd0; scan_win1594 <= 32'd0; scan_win1595 <= 32'd0; scan_win1596 <= 32'd0; scan_win1597 <= 32'd0; scan_win1598 <= 32'd0; scan_win1599 <= 32'd0; scan_win1600 <= 32'd0; 
      scan_win1601 <= 32'd0; scan_win1602 <= 32'd0; scan_win1603 <= 32'd0; scan_win1604 <= 32'd0; scan_win1605 <= 32'd0; scan_win1606 <= 32'd0; scan_win1607 <= 32'd0; scan_win1608 <= 32'd0; scan_win1609 <= 32'd0; scan_win1610 <= 32'd0; scan_win1611 <= 32'd0; scan_win1612 <= 32'd0; scan_win1613 <= 32'd0; scan_win1614 <= 32'd0; scan_win1615 <= 32'd0; scan_win1616 <= 32'd0; scan_win1617 <= 32'd0; scan_win1618 <= 32'd0; scan_win1619 <= 32'd0; scan_win1620 <= 32'd0; scan_win1621 <= 32'd0; scan_win1622 <= 32'd0; scan_win1623 <= 32'd0; scan_win1624 <= 32'd0; scan_win1625 <= 32'd0; scan_win1626 <= 32'd0; scan_win1627 <= 32'd0; scan_win1628 <= 32'd0; scan_win1629 <= 32'd0; scan_win1630 <= 32'd0; scan_win1631 <= 32'd0; scan_win1632 <= 32'd0; scan_win1633 <= 32'd0; scan_win1634 <= 32'd0; scan_win1635 <= 32'd0; scan_win1636 <= 32'd0; scan_win1637 <= 32'd0; scan_win1638 <= 32'd0; scan_win1639 <= 32'd0; scan_win1640 <= 32'd0; scan_win1641 <= 32'd0; scan_win1642 <= 32'd0; scan_win1643 <= 32'd0; scan_win1644 <= 32'd0; scan_win1645 <= 32'd0; scan_win1646 <= 32'd0; scan_win1647 <= 32'd0; scan_win1648 <= 32'd0; scan_win1649 <= 32'd0; scan_win1650 <= 32'd0; scan_win1651 <= 32'd0; scan_win1652 <= 32'd0; scan_win1653 <= 32'd0; scan_win1654 <= 32'd0; scan_win1655 <= 32'd0; scan_win1656 <= 32'd0; scan_win1657 <= 32'd0; scan_win1658 <= 32'd0; scan_win1659 <= 32'd0; scan_win1660 <= 32'd0; scan_win1661 <= 32'd0; scan_win1662 <= 32'd0; scan_win1663 <= 32'd0; scan_win1664 <= 32'd0; scan_win1665 <= 32'd0; scan_win1666 <= 32'd0; scan_win1667 <= 32'd0; scan_win1668 <= 32'd0; scan_win1669 <= 32'd0; scan_win1670 <= 32'd0; scan_win1671 <= 32'd0; scan_win1672 <= 32'd0; scan_win1673 <= 32'd0; scan_win1674 <= 32'd0; scan_win1675 <= 32'd0; scan_win1676 <= 32'd0; scan_win1677 <= 32'd0; scan_win1678 <= 32'd0; scan_win1679 <= 32'd0; scan_win1680 <= 32'd0; scan_win1681 <= 32'd0; scan_win1682 <= 32'd0; scan_win1683 <= 32'd0; scan_win1684 <= 32'd0; scan_win1685 <= 32'd0; scan_win1686 <= 32'd0; scan_win1687 <= 32'd0; scan_win1688 <= 32'd0; scan_win1689 <= 32'd0; scan_win1690 <= 32'd0; scan_win1691 <= 32'd0; scan_win1692 <= 32'd0; scan_win1693 <= 32'd0; scan_win1694 <= 32'd0; scan_win1695 <= 32'd0; scan_win1696 <= 32'd0; scan_win1697 <= 32'd0; scan_win1698 <= 32'd0; scan_win1699 <= 32'd0; scan_win1700 <= 32'd0; scan_win1701 <= 32'd0; scan_win1702 <= 32'd0; scan_win1703 <= 32'd0; scan_win1704 <= 32'd0; scan_win1705 <= 32'd0; scan_win1706 <= 32'd0; scan_win1707 <= 32'd0; scan_win1708 <= 32'd0; scan_win1709 <= 32'd0; scan_win1710 <= 32'd0; scan_win1711 <= 32'd0; scan_win1712 <= 32'd0; scan_win1713 <= 32'd0; scan_win1714 <= 32'd0; scan_win1715 <= 32'd0; scan_win1716 <= 32'd0; scan_win1717 <= 32'd0; scan_win1718 <= 32'd0; scan_win1719 <= 32'd0; scan_win1720 <= 32'd0; scan_win1721 <= 32'd0; scan_win1722 <= 32'd0; scan_win1723 <= 32'd0; scan_win1724 <= 32'd0; scan_win1725 <= 32'd0; scan_win1726 <= 32'd0; scan_win1727 <= 32'd0; scan_win1728 <= 32'd0; scan_win1729 <= 32'd0; scan_win1730 <= 32'd0; scan_win1731 <= 32'd0; scan_win1732 <= 32'd0; scan_win1733 <= 32'd0; scan_win1734 <= 32'd0; scan_win1735 <= 32'd0; scan_win1736 <= 32'd0; scan_win1737 <= 32'd0; scan_win1738 <= 32'd0; scan_win1739 <= 32'd0; scan_win1740 <= 32'd0; scan_win1741 <= 32'd0; scan_win1742 <= 32'd0; scan_win1743 <= 32'd0; scan_win1744 <= 32'd0; scan_win1745 <= 32'd0; scan_win1746 <= 32'd0; scan_win1747 <= 32'd0; scan_win1748 <= 32'd0; scan_win1749 <= 32'd0; scan_win1750 <= 32'd0; scan_win1751 <= 32'd0; scan_win1752 <= 32'd0; scan_win1753 <= 32'd0; scan_win1754 <= 32'd0; scan_win1755 <= 32'd0; scan_win1756 <= 32'd0; scan_win1757 <= 32'd0; scan_win1758 <= 32'd0; scan_win1759 <= 32'd0; scan_win1760 <= 32'd0; scan_win1761 <= 32'd0; scan_win1762 <= 32'd0; scan_win1763 <= 32'd0; scan_win1764 <= 32'd0; scan_win1765 <= 32'd0; scan_win1766 <= 32'd0; scan_win1767 <= 32'd0; scan_win1768 <= 32'd0; scan_win1769 <= 32'd0; scan_win1770 <= 32'd0; scan_win1771 <= 32'd0; scan_win1772 <= 32'd0; scan_win1773 <= 32'd0; scan_win1774 <= 32'd0; scan_win1775 <= 32'd0; scan_win1776 <= 32'd0; scan_win1777 <= 32'd0; scan_win1778 <= 32'd0; scan_win1779 <= 32'd0; scan_win1780 <= 32'd0; scan_win1781 <= 32'd0; scan_win1782 <= 32'd0; scan_win1783 <= 32'd0; scan_win1784 <= 32'd0; scan_win1785 <= 32'd0; scan_win1786 <= 32'd0; scan_win1787 <= 32'd0; scan_win1788 <= 32'd0; scan_win1789 <= 32'd0; scan_win1790 <= 32'd0; scan_win1791 <= 32'd0; scan_win1792 <= 32'd0; scan_win1793 <= 32'd0; scan_win1794 <= 32'd0; scan_win1795 <= 32'd0; scan_win1796 <= 32'd0; scan_win1797 <= 32'd0; scan_win1798 <= 32'd0; scan_win1799 <= 32'd0; scan_win1800 <= 32'd0; 
      scan_win1801 <= 32'd0; scan_win1802 <= 32'd0; scan_win1803 <= 32'd0; scan_win1804 <= 32'd0; scan_win1805 <= 32'd0; scan_win1806 <= 32'd0; scan_win1807 <= 32'd0; scan_win1808 <= 32'd0; scan_win1809 <= 32'd0; scan_win1810 <= 32'd0; scan_win1811 <= 32'd0; scan_win1812 <= 32'd0; scan_win1813 <= 32'd0; scan_win1814 <= 32'd0; scan_win1815 <= 32'd0; scan_win1816 <= 32'd0; scan_win1817 <= 32'd0; scan_win1818 <= 32'd0; scan_win1819 <= 32'd0; scan_win1820 <= 32'd0; scan_win1821 <= 32'd0; scan_win1822 <= 32'd0; scan_win1823 <= 32'd0; scan_win1824 <= 32'd0; scan_win1825 <= 32'd0; scan_win1826 <= 32'd0; scan_win1827 <= 32'd0; scan_win1828 <= 32'd0; scan_win1829 <= 32'd0; scan_win1830 <= 32'd0; scan_win1831 <= 32'd0; scan_win1832 <= 32'd0; scan_win1833 <= 32'd0; scan_win1834 <= 32'd0; scan_win1835 <= 32'd0; scan_win1836 <= 32'd0; scan_win1837 <= 32'd0; scan_win1838 <= 32'd0; scan_win1839 <= 32'd0; scan_win1840 <= 32'd0; scan_win1841 <= 32'd0; scan_win1842 <= 32'd0; scan_win1843 <= 32'd0; scan_win1844 <= 32'd0; scan_win1845 <= 32'd0; scan_win1846 <= 32'd0; scan_win1847 <= 32'd0; scan_win1848 <= 32'd0; scan_win1849 <= 32'd0; scan_win1850 <= 32'd0; scan_win1851 <= 32'd0; scan_win1852 <= 32'd0; scan_win1853 <= 32'd0; scan_win1854 <= 32'd0; scan_win1855 <= 32'd0; scan_win1856 <= 32'd0; scan_win1857 <= 32'd0; scan_win1858 <= 32'd0; scan_win1859 <= 32'd0; scan_win1860 <= 32'd0; scan_win1861 <= 32'd0; scan_win1862 <= 32'd0; scan_win1863 <= 32'd0; scan_win1864 <= 32'd0; scan_win1865 <= 32'd0; scan_win1866 <= 32'd0; scan_win1867 <= 32'd0; scan_win1868 <= 32'd0; scan_win1869 <= 32'd0; scan_win1870 <= 32'd0; scan_win1871 <= 32'd0; scan_win1872 <= 32'd0; scan_win1873 <= 32'd0; scan_win1874 <= 32'd0; scan_win1875 <= 32'd0; scan_win1876 <= 32'd0; scan_win1877 <= 32'd0; scan_win1878 <= 32'd0; scan_win1879 <= 32'd0; scan_win1880 <= 32'd0; scan_win1881 <= 32'd0; scan_win1882 <= 32'd0; scan_win1883 <= 32'd0; scan_win1884 <= 32'd0; scan_win1885 <= 32'd0; scan_win1886 <= 32'd0; scan_win1887 <= 32'd0; scan_win1888 <= 32'd0; scan_win1889 <= 32'd0; scan_win1890 <= 32'd0; scan_win1891 <= 32'd0; scan_win1892 <= 32'd0; scan_win1893 <= 32'd0; scan_win1894 <= 32'd0; scan_win1895 <= 32'd0; scan_win1896 <= 32'd0; scan_win1897 <= 32'd0; scan_win1898 <= 32'd0; scan_win1899 <= 32'd0; scan_win1900 <= 32'd0; scan_win1901 <= 32'd0; scan_win1902 <= 32'd0; scan_win1903 <= 32'd0; scan_win1904 <= 32'd0; scan_win1905 <= 32'd0; scan_win1906 <= 32'd0; scan_win1907 <= 32'd0; scan_win1908 <= 32'd0; scan_win1909 <= 32'd0; scan_win1910 <= 32'd0; scan_win1911 <= 32'd0; scan_win1912 <= 32'd0; scan_win1913 <= 32'd0; scan_win1914 <= 32'd0; scan_win1915 <= 32'd0; scan_win1916 <= 32'd0; scan_win1917 <= 32'd0; scan_win1918 <= 32'd0; scan_win1919 <= 32'd0; scan_win1920 <= 32'd0; scan_win1921 <= 32'd0; scan_win1922 <= 32'd0; scan_win1923 <= 32'd0; scan_win1924 <= 32'd0; scan_win1925 <= 32'd0; scan_win1926 <= 32'd0; scan_win1927 <= 32'd0; scan_win1928 <= 32'd0; scan_win1929 <= 32'd0; scan_win1930 <= 32'd0; scan_win1931 <= 32'd0; scan_win1932 <= 32'd0; scan_win1933 <= 32'd0; scan_win1934 <= 32'd0; scan_win1935 <= 32'd0; scan_win1936 <= 32'd0; scan_win1937 <= 32'd0; scan_win1938 <= 32'd0; scan_win1939 <= 32'd0; scan_win1940 <= 32'd0; scan_win1941 <= 32'd0; scan_win1942 <= 32'd0; scan_win1943 <= 32'd0; scan_win1944 <= 32'd0; scan_win1945 <= 32'd0; scan_win1946 <= 32'd0; scan_win1947 <= 32'd0; scan_win1948 <= 32'd0; scan_win1949 <= 32'd0; scan_win1950 <= 32'd0; scan_win1951 <= 32'd0; scan_win1952 <= 32'd0; scan_win1953 <= 32'd0; scan_win1954 <= 32'd0; scan_win1955 <= 32'd0; scan_win1956 <= 32'd0; scan_win1957 <= 32'd0; scan_win1958 <= 32'd0; scan_win1959 <= 32'd0; scan_win1960 <= 32'd0; scan_win1961 <= 32'd0; scan_win1962 <= 32'd0; scan_win1963 <= 32'd0; scan_win1964 <= 32'd0; scan_win1965 <= 32'd0; scan_win1966 <= 32'd0; scan_win1967 <= 32'd0; scan_win1968 <= 32'd0; scan_win1969 <= 32'd0; scan_win1970 <= 32'd0; scan_win1971 <= 32'd0; scan_win1972 <= 32'd0; scan_win1973 <= 32'd0; scan_win1974 <= 32'd0; scan_win1975 <= 32'd0; scan_win1976 <= 32'd0; scan_win1977 <= 32'd0; scan_win1978 <= 32'd0; scan_win1979 <= 32'd0; scan_win1980 <= 32'd0; scan_win1981 <= 32'd0; scan_win1982 <= 32'd0; scan_win1983 <= 32'd0; scan_win1984 <= 32'd0; scan_win1985 <= 32'd0; scan_win1986 <= 32'd0; scan_win1987 <= 32'd0; scan_win1988 <= 32'd0; scan_win1989 <= 32'd0; scan_win1990 <= 32'd0; scan_win1991 <= 32'd0; scan_win1992 <= 32'd0; scan_win1993 <= 32'd0; scan_win1994 <= 32'd0; scan_win1995 <= 32'd0; scan_win1996 <= 32'd0; scan_win1997 <= 32'd0; scan_win1998 <= 32'd0; scan_win1999 <= 32'd0; scan_win2000 <= 32'd0; 
      scan_win2001 <= 32'd0; scan_win2002 <= 32'd0; scan_win2003 <= 32'd0; scan_win2004 <= 32'd0; scan_win2005 <= 32'd0; scan_win2006 <= 32'd0; scan_win2007 <= 32'd0; scan_win2008 <= 32'd0; scan_win2009 <= 32'd0; scan_win2010 <= 32'd0; scan_win2011 <= 32'd0; scan_win2012 <= 32'd0; scan_win2013 <= 32'd0; scan_win2014 <= 32'd0; scan_win2015 <= 32'd0; scan_win2016 <= 32'd0; scan_win2017 <= 32'd0; scan_win2018 <= 32'd0; scan_win2019 <= 32'd0; scan_win2020 <= 32'd0; scan_win2021 <= 32'd0; scan_win2022 <= 32'd0; scan_win2023 <= 32'd0; scan_win2024 <= 32'd0; scan_win2025 <= 32'd0; scan_win2026 <= 32'd0; scan_win2027 <= 32'd0; scan_win2028 <= 32'd0; scan_win2029 <= 32'd0; scan_win2030 <= 32'd0; scan_win2031 <= 32'd0; scan_win2032 <= 32'd0; scan_win2033 <= 32'd0; scan_win2034 <= 32'd0; scan_win2035 <= 32'd0; scan_win2036 <= 32'd0; scan_win2037 <= 32'd0; scan_win2038 <= 32'd0; scan_win2039 <= 32'd0; scan_win2040 <= 32'd0; scan_win2041 <= 32'd0; scan_win2042 <= 32'd0; scan_win2043 <= 32'd0; scan_win2044 <= 32'd0; scan_win2045 <= 32'd0; scan_win2046 <= 32'd0; scan_win2047 <= 32'd0; scan_win2048 <= 32'd0; scan_win2049 <= 32'd0; scan_win2050 <= 32'd0; scan_win2051 <= 32'd0; scan_win2052 <= 32'd0; scan_win2053 <= 32'd0; scan_win2054 <= 32'd0; scan_win2055 <= 32'd0; scan_win2056 <= 32'd0; scan_win2057 <= 32'd0; scan_win2058 <= 32'd0; scan_win2059 <= 32'd0; scan_win2060 <= 32'd0; scan_win2061 <= 32'd0; scan_win2062 <= 32'd0; scan_win2063 <= 32'd0; scan_win2064 <= 32'd0; scan_win2065 <= 32'd0; scan_win2066 <= 32'd0; scan_win2067 <= 32'd0; scan_win2068 <= 32'd0; scan_win2069 <= 32'd0; scan_win2070 <= 32'd0; scan_win2071 <= 32'd0; scan_win2072 <= 32'd0; scan_win2073 <= 32'd0; scan_win2074 <= 32'd0; scan_win2075 <= 32'd0; scan_win2076 <= 32'd0; scan_win2077 <= 32'd0; scan_win2078 <= 32'd0; scan_win2079 <= 32'd0; scan_win2080 <= 32'd0; scan_win2081 <= 32'd0; scan_win2082 <= 32'd0; scan_win2083 <= 32'd0; scan_win2084 <= 32'd0; scan_win2085 <= 32'd0; scan_win2086 <= 32'd0; scan_win2087 <= 32'd0; scan_win2088 <= 32'd0; scan_win2089 <= 32'd0; scan_win2090 <= 32'd0; scan_win2091 <= 32'd0; scan_win2092 <= 32'd0; scan_win2093 <= 32'd0; scan_win2094 <= 32'd0; scan_win2095 <= 32'd0; scan_win2096 <= 32'd0; scan_win2097 <= 32'd0; scan_win2098 <= 32'd0; scan_win2099 <= 32'd0; scan_win2100 <= 32'd0; scan_win2101 <= 32'd0; scan_win2102 <= 32'd0; scan_win2103 <= 32'd0; scan_win2104 <= 32'd0; scan_win2105 <= 32'd0; scan_win2106 <= 32'd0; scan_win2107 <= 32'd0; scan_win2108 <= 32'd0; scan_win2109 <= 32'd0; scan_win2110 <= 32'd0; scan_win2111 <= 32'd0; scan_win2112 <= 32'd0; scan_win2113 <= 32'd0; scan_win2114 <= 32'd0; scan_win2115 <= 32'd0; scan_win2116 <= 32'd0; scan_win2117 <= 32'd0; scan_win2118 <= 32'd0; scan_win2119 <= 32'd0; scan_win2120 <= 32'd0; scan_win2121 <= 32'd0; scan_win2122 <= 32'd0; scan_win2123 <= 32'd0; scan_win2124 <= 32'd0; scan_win2125 <= 32'd0; scan_win2126 <= 32'd0; scan_win2127 <= 32'd0; scan_win2128 <= 32'd0; scan_win2129 <= 32'd0; scan_win2130 <= 32'd0; scan_win2131 <= 32'd0; scan_win2132 <= 32'd0; scan_win2133 <= 32'd0; scan_win2134 <= 32'd0; scan_win2135 <= 32'd0; scan_win2136 <= 32'd0; scan_win2137 <= 32'd0; scan_win2138 <= 32'd0; scan_win2139 <= 32'd0; scan_win2140 <= 32'd0; scan_win2141 <= 32'd0; scan_win2142 <= 32'd0; scan_win2143 <= 32'd0; scan_win2144 <= 32'd0; scan_win2145 <= 32'd0; scan_win2146 <= 32'd0; scan_win2147 <= 32'd0; scan_win2148 <= 32'd0; scan_win2149 <= 32'd0; scan_win2150 <= 32'd0; scan_win2151 <= 32'd0; scan_win2152 <= 32'd0; scan_win2153 <= 32'd0; scan_win2154 <= 32'd0; scan_win2155 <= 32'd0; scan_win2156 <= 32'd0; scan_win2157 <= 32'd0; scan_win2158 <= 32'd0; scan_win2159 <= 32'd0; scan_win2160 <= 32'd0; scan_win2161 <= 32'd0; scan_win2162 <= 32'd0; scan_win2163 <= 32'd0; scan_win2164 <= 32'd0; scan_win2165 <= 32'd0; scan_win2166 <= 32'd0; scan_win2167 <= 32'd0; scan_win2168 <= 32'd0; scan_win2169 <= 32'd0; scan_win2170 <= 32'd0; scan_win2171 <= 32'd0; scan_win2172 <= 32'd0; scan_win2173 <= 32'd0; scan_win2174 <= 32'd0; scan_win2175 <= 32'd0; scan_win2176 <= 32'd0; scan_win2177 <= 32'd0; scan_win2178 <= 32'd0; scan_win2179 <= 32'd0; scan_win2180 <= 32'd0; scan_win2181 <= 32'd0; scan_win2182 <= 32'd0; scan_win2183 <= 32'd0; scan_win2184 <= 32'd0; scan_win2185 <= 32'd0; scan_win2186 <= 32'd0; scan_win2187 <= 32'd0; scan_win2188 <= 32'd0; scan_win2189 <= 32'd0; scan_win2190 <= 32'd0; scan_win2191 <= 32'd0; scan_win2192 <= 32'd0; scan_win2193 <= 32'd0; scan_win2194 <= 32'd0; scan_win2195 <= 32'd0; scan_win2196 <= 32'd0; scan_win2197 <= 32'd0; scan_win2198 <= 32'd0; scan_win2199 <= 32'd0; scan_win2200 <= 32'd0; 
      scan_win2201 <= 32'd0; scan_win2202 <= 32'd0; scan_win2203 <= 32'd0; scan_win2204 <= 32'd0; scan_win2205 <= 32'd0; scan_win2206 <= 32'd0; scan_win2207 <= 32'd0; scan_win2208 <= 32'd0; scan_win2209 <= 32'd0; scan_win2210 <= 32'd0; scan_win2211 <= 32'd0; scan_win2212 <= 32'd0; scan_win2213 <= 32'd0; scan_win2214 <= 32'd0; scan_win2215 <= 32'd0; scan_win2216 <= 32'd0; scan_win2217 <= 32'd0; scan_win2218 <= 32'd0; scan_win2219 <= 32'd0; scan_win2220 <= 32'd0; scan_win2221 <= 32'd0; scan_win2222 <= 32'd0; scan_win2223 <= 32'd0; scan_win2224 <= 32'd0; scan_win2225 <= 32'd0; scan_win2226 <= 32'd0; scan_win2227 <= 32'd0; scan_win2228 <= 32'd0; scan_win2229 <= 32'd0; scan_win2230 <= 32'd0; scan_win2231 <= 32'd0; scan_win2232 <= 32'd0; scan_win2233 <= 32'd0; scan_win2234 <= 32'd0; scan_win2235 <= 32'd0; scan_win2236 <= 32'd0; scan_win2237 <= 32'd0; scan_win2238 <= 32'd0; scan_win2239 <= 32'd0; scan_win2240 <= 32'd0; scan_win2241 <= 32'd0; scan_win2242 <= 32'd0; scan_win2243 <= 32'd0; scan_win2244 <= 32'd0; scan_win2245 <= 32'd0; scan_win2246 <= 32'd0; scan_win2247 <= 32'd0; scan_win2248 <= 32'd0; scan_win2249 <= 32'd0; scan_win2250 <= 32'd0; scan_win2251 <= 32'd0; scan_win2252 <= 32'd0; scan_win2253 <= 32'd0; scan_win2254 <= 32'd0; scan_win2255 <= 32'd0; scan_win2256 <= 32'd0; scan_win2257 <= 32'd0; scan_win2258 <= 32'd0; scan_win2259 <= 32'd0; scan_win2260 <= 32'd0; scan_win2261 <= 32'd0; scan_win2262 <= 32'd0; scan_win2263 <= 32'd0; scan_win2264 <= 32'd0; scan_win2265 <= 32'd0; scan_win2266 <= 32'd0; scan_win2267 <= 32'd0; scan_win2268 <= 32'd0; scan_win2269 <= 32'd0; scan_win2270 <= 32'd0; scan_win2271 <= 32'd0; scan_win2272 <= 32'd0; scan_win2273 <= 32'd0; scan_win2274 <= 32'd0; scan_win2275 <= 32'd0; scan_win2276 <= 32'd0; scan_win2277 <= 32'd0; scan_win2278 <= 32'd0; scan_win2279 <= 32'd0; scan_win2280 <= 32'd0; scan_win2281 <= 32'd0; scan_win2282 <= 32'd0; scan_win2283 <= 32'd0; scan_win2284 <= 32'd0; scan_win2285 <= 32'd0; scan_win2286 <= 32'd0; scan_win2287 <= 32'd0; scan_win2288 <= 32'd0; scan_win2289 <= 32'd0; scan_win2290 <= 32'd0; scan_win2291 <= 32'd0; scan_win2292 <= 32'd0; scan_win2293 <= 32'd0; scan_win2294 <= 32'd0; scan_win2295 <= 32'd0; scan_win2296 <= 32'd0; scan_win2297 <= 32'd0; scan_win2298 <= 32'd0; scan_win2299 <= 32'd0; scan_win2300 <= 32'd0; scan_win2301 <= 32'd0; scan_win2302 <= 32'd0; scan_win2303 <= 32'd0; scan_win2304 <= 32'd0; scan_win2305 <= 32'd0; scan_win2306 <= 32'd0; scan_win2307 <= 32'd0; scan_win2308 <= 32'd0; scan_win2309 <= 32'd0; scan_win2310 <= 32'd0; scan_win2311 <= 32'd0; scan_win2312 <= 32'd0; scan_win2313 <= 32'd0; scan_win2314 <= 32'd0; scan_win2315 <= 32'd0; scan_win2316 <= 32'd0; scan_win2317 <= 32'd0; scan_win2318 <= 32'd0; scan_win2319 <= 32'd0; scan_win2320 <= 32'd0; scan_win2321 <= 32'd0; scan_win2322 <= 32'd0; scan_win2323 <= 32'd0; scan_win2324 <= 32'd0; scan_win2325 <= 32'd0; scan_win2326 <= 32'd0; scan_win2327 <= 32'd0; scan_win2328 <= 32'd0; scan_win2329 <= 32'd0; scan_win2330 <= 32'd0; scan_win2331 <= 32'd0; scan_win2332 <= 32'd0; scan_win2333 <= 32'd0; scan_win2334 <= 32'd0; scan_win2335 <= 32'd0; scan_win2336 <= 32'd0; scan_win2337 <= 32'd0; scan_win2338 <= 32'd0; scan_win2339 <= 32'd0; scan_win2340 <= 32'd0; scan_win2341 <= 32'd0; scan_win2342 <= 32'd0; scan_win2343 <= 32'd0; scan_win2344 <= 32'd0; scan_win2345 <= 32'd0; scan_win2346 <= 32'd0; scan_win2347 <= 32'd0; scan_win2348 <= 32'd0; scan_win2349 <= 32'd0; scan_win2350 <= 32'd0; scan_win2351 <= 32'd0; scan_win2352 <= 32'd0; scan_win2353 <= 32'd0; scan_win2354 <= 32'd0; scan_win2355 <= 32'd0; scan_win2356 <= 32'd0; scan_win2357 <= 32'd0; scan_win2358 <= 32'd0; scan_win2359 <= 32'd0; scan_win2360 <= 32'd0; scan_win2361 <= 32'd0; scan_win2362 <= 32'd0; scan_win2363 <= 32'd0; scan_win2364 <= 32'd0; scan_win2365 <= 32'd0; scan_win2366 <= 32'd0; scan_win2367 <= 32'd0; scan_win2368 <= 32'd0; scan_win2369 <= 32'd0; scan_win2370 <= 32'd0; scan_win2371 <= 32'd0; scan_win2372 <= 32'd0; scan_win2373 <= 32'd0; scan_win2374 <= 32'd0; scan_win2375 <= 32'd0; scan_win2376 <= 32'd0; scan_win2377 <= 32'd0; scan_win2378 <= 32'd0; scan_win2379 <= 32'd0; scan_win2380 <= 32'd0; scan_win2381 <= 32'd0; scan_win2382 <= 32'd0; scan_win2383 <= 32'd0; scan_win2384 <= 32'd0; scan_win2385 <= 32'd0; scan_win2386 <= 32'd0; scan_win2387 <= 32'd0; scan_win2388 <= 32'd0; scan_win2389 <= 32'd0; scan_win2390 <= 32'd0; scan_win2391 <= 32'd0; scan_win2392 <= 32'd0; scan_win2393 <= 32'd0; scan_win2394 <= 32'd0; scan_win2395 <= 32'd0; scan_win2396 <= 32'd0; scan_win2397 <= 32'd0; scan_win2398 <= 32'd0; scan_win2399 <= 32'd0; scan_win2400 <= 32'd0; 
      scan_win2401 <= 32'd0; scan_win2402 <= 32'd0; scan_win2403 <= 32'd0; scan_win2404 <= 32'd0; scan_win2405 <= 32'd0; scan_win2406 <= 32'd0; scan_win2407 <= 32'd0; scan_win2408 <= 32'd0; scan_win2409 <= 32'd0; scan_win2410 <= 32'd0; scan_win2411 <= 32'd0; scan_win2412 <= 32'd0; scan_win2413 <= 32'd0; scan_win2414 <= 32'd0; scan_win2415 <= 32'd0; scan_win2416 <= 32'd0; scan_win2417 <= 32'd0; scan_win2418 <= 32'd0; scan_win2419 <= 32'd0; scan_win2420 <= 32'd0; scan_win2421 <= 32'd0; scan_win2422 <= 32'd0; scan_win2423 <= 32'd0; scan_win2424 <= 32'd0; scan_win2425 <= 32'd0; scan_win2426 <= 32'd0; scan_win2427 <= 32'd0; scan_win2428 <= 32'd0; scan_win2429 <= 32'd0; scan_win2430 <= 32'd0; scan_win2431 <= 32'd0; scan_win2432 <= 32'd0; scan_win2433 <= 32'd0; scan_win2434 <= 32'd0; scan_win2435 <= 32'd0; scan_win2436 <= 32'd0; scan_win2437 <= 32'd0; scan_win2438 <= 32'd0; scan_win2439 <= 32'd0; scan_win2440 <= 32'd0; scan_win2441 <= 32'd0; scan_win2442 <= 32'd0; scan_win2443 <= 32'd0; scan_win2444 <= 32'd0; scan_win2445 <= 32'd0; scan_win2446 <= 32'd0; scan_win2447 <= 32'd0; scan_win2448 <= 32'd0; scan_win2449 <= 32'd0; scan_win2450 <= 32'd0; scan_win2451 <= 32'd0; scan_win2452 <= 32'd0; scan_win2453 <= 32'd0; scan_win2454 <= 32'd0; scan_win2455 <= 32'd0; scan_win2456 <= 32'd0; scan_win2457 <= 32'd0; scan_win2458 <= 32'd0; scan_win2459 <= 32'd0; scan_win2460 <= 32'd0; scan_win2461 <= 32'd0; scan_win2462 <= 32'd0; scan_win2463 <= 32'd0; scan_win2464 <= 32'd0; scan_win2465 <= 32'd0; scan_win2466 <= 32'd0; scan_win2467 <= 32'd0; scan_win2468 <= 32'd0; scan_win2469 <= 32'd0; scan_win2470 <= 32'd0; scan_win2471 <= 32'd0; scan_win2472 <= 32'd0; scan_win2473 <= 32'd0; scan_win2474 <= 32'd0; scan_win2475 <= 32'd0; scan_win2476 <= 32'd0; scan_win2477 <= 32'd0; scan_win2478 <= 32'd0; scan_win2479 <= 32'd0; scan_win2480 <= 32'd0; scan_win2481 <= 32'd0; scan_win2482 <= 32'd0; scan_win2483 <= 32'd0; scan_win2484 <= 32'd0; scan_win2485 <= 32'd0; scan_win2486 <= 32'd0; scan_win2487 <= 32'd0; scan_win2488 <= 32'd0; scan_win2489 <= 32'd0; scan_win2490 <= 32'd0; scan_win2491 <= 32'd0; scan_win2492 <= 32'd0; scan_win2493 <= 32'd0; scan_win2494 <= 32'd0; scan_win2495 <= 32'd0; scan_win2496 <= 32'd0; scan_win2497 <= 32'd0; scan_win2498 <= 32'd0; scan_win2499 <= 32'd0; scan_win2500 <= 32'd0; scan_win2501 <= 32'd0; scan_win2502 <= 32'd0; scan_win2503 <= 32'd0; scan_win2504 <= 32'd0; scan_win2505 <= 32'd0; scan_win2506 <= 32'd0; scan_win2507 <= 32'd0; scan_win2508 <= 32'd0; scan_win2509 <= 32'd0; scan_win2510 <= 32'd0; scan_win2511 <= 32'd0; scan_win2512 <= 32'd0; scan_win2513 <= 32'd0; scan_win2514 <= 32'd0; scan_win2515 <= 32'd0; scan_win2516 <= 32'd0; scan_win2517 <= 32'd0; scan_win2518 <= 32'd0; scan_win2519 <= 32'd0; scan_win2520 <= 32'd0; scan_win2521 <= 32'd0; scan_win2522 <= 32'd0; scan_win2523 <= 32'd0; scan_win2524 <= 32'd0; scan_win2525 <= 32'd0; scan_win2526 <= 32'd0; scan_win2527 <= 32'd0; scan_win2528 <= 32'd0; scan_win2529 <= 32'd0; scan_win2530 <= 32'd0; scan_win2531 <= 32'd0; scan_win2532 <= 32'd0; scan_win2533 <= 32'd0; scan_win2534 <= 32'd0; scan_win2535 <= 32'd0; scan_win2536 <= 32'd0; scan_win2537 <= 32'd0; scan_win2538 <= 32'd0; scan_win2539 <= 32'd0; scan_win2540 <= 32'd0; scan_win2541 <= 32'd0; scan_win2542 <= 32'd0; scan_win2543 <= 32'd0; scan_win2544 <= 32'd0; scan_win2545 <= 32'd0; scan_win2546 <= 32'd0; scan_win2547 <= 32'd0; scan_win2548 <= 32'd0; scan_win2549 <= 32'd0; scan_win2550 <= 32'd0; scan_win2551 <= 32'd0; scan_win2552 <= 32'd0; scan_win2553 <= 32'd0; scan_win2554 <= 32'd0; scan_win2555 <= 32'd0; scan_win2556 <= 32'd0; scan_win2557 <= 32'd0; scan_win2558 <= 32'd0; scan_win2559 <= 32'd0; scan_win2560 <= 32'd0; scan_win2561 <= 32'd0; scan_win2562 <= 32'd0; scan_win2563 <= 32'd0; scan_win2564 <= 32'd0; scan_win2565 <= 32'd0; scan_win2566 <= 32'd0; scan_win2567 <= 32'd0; scan_win2568 <= 32'd0; scan_win2569 <= 32'd0; scan_win2570 <= 32'd0; scan_win2571 <= 32'd0; scan_win2572 <= 32'd0; scan_win2573 <= 32'd0; scan_win2574 <= 32'd0; scan_win2575 <= 32'd0; scan_win2576 <= 32'd0; scan_win2577 <= 32'd0; scan_win2578 <= 32'd0; scan_win2579 <= 32'd0; scan_win2580 <= 32'd0; scan_win2581 <= 32'd0; scan_win2582 <= 32'd0; scan_win2583 <= 32'd0; scan_win2584 <= 32'd0; scan_win2585 <= 32'd0; scan_win2586 <= 32'd0; scan_win2587 <= 32'd0; scan_win2588 <= 32'd0; scan_win2589 <= 32'd0; scan_win2590 <= 32'd0; scan_win2591 <= 32'd0; scan_win2592 <= 32'd0; scan_win2593 <= 32'd0; scan_win2594 <= 32'd0; scan_win2595 <= 32'd0; scan_win2596 <= 32'd0; scan_win2597 <= 32'd0; scan_win2598 <= 32'd0; scan_win2599 <= 32'd0; scan_win2600 <= 32'd0; 
      scan_win2601 <= 32'd0; scan_win2602 <= 32'd0; scan_win2603 <= 32'd0; scan_win2604 <= 32'd0; scan_win2605 <= 32'd0; scan_win2606 <= 32'd0; scan_win2607 <= 32'd0; scan_win2608 <= 32'd0; scan_win2609 <= 32'd0; scan_win2610 <= 32'd0; scan_win2611 <= 32'd0; scan_win2612 <= 32'd0; scan_win2613 <= 32'd0; scan_win2614 <= 32'd0; scan_win2615 <= 32'd0; scan_win2616 <= 32'd0; scan_win2617 <= 32'd0; scan_win2618 <= 32'd0; scan_win2619 <= 32'd0; scan_win2620 <= 32'd0; scan_win2621 <= 32'd0; scan_win2622 <= 32'd0; scan_win2623 <= 32'd0; scan_win2624 <= 32'd0; scan_win2625 <= 32'd0; scan_win2626 <= 32'd0; scan_win2627 <= 32'd0; scan_win2628 <= 32'd0; scan_win2629 <= 32'd0; scan_win2630 <= 32'd0; scan_win2631 <= 32'd0; scan_win2632 <= 32'd0; scan_win2633 <= 32'd0; scan_win2634 <= 32'd0; scan_win2635 <= 32'd0; scan_win2636 <= 32'd0; scan_win2637 <= 32'd0; scan_win2638 <= 32'd0; scan_win2639 <= 32'd0; scan_win2640 <= 32'd0; scan_win2641 <= 32'd0; scan_win2642 <= 32'd0; scan_win2643 <= 32'd0; scan_win2644 <= 32'd0; scan_win2645 <= 32'd0; scan_win2646 <= 32'd0; scan_win2647 <= 32'd0; scan_win2648 <= 32'd0; scan_win2649 <= 32'd0; scan_win2650 <= 32'd0; scan_win2651 <= 32'd0; scan_win2652 <= 32'd0; scan_win2653 <= 32'd0; scan_win2654 <= 32'd0; scan_win2655 <= 32'd0; scan_win2656 <= 32'd0; scan_win2657 <= 32'd0; scan_win2658 <= 32'd0; scan_win2659 <= 32'd0; scan_win2660 <= 32'd0; scan_win2661 <= 32'd0; scan_win2662 <= 32'd0; scan_win2663 <= 32'd0; scan_win2664 <= 32'd0; scan_win2665 <= 32'd0; scan_win2666 <= 32'd0; scan_win2667 <= 32'd0; scan_win2668 <= 32'd0; scan_win2669 <= 32'd0; scan_win2670 <= 32'd0; scan_win2671 <= 32'd0; scan_win2672 <= 32'd0; scan_win2673 <= 32'd0; scan_win2674 <= 32'd0; scan_win2675 <= 32'd0; scan_win2676 <= 32'd0; scan_win2677 <= 32'd0; scan_win2678 <= 32'd0; scan_win2679 <= 32'd0; scan_win2680 <= 32'd0; scan_win2681 <= 32'd0; scan_win2682 <= 32'd0; scan_win2683 <= 32'd0; scan_win2684 <= 32'd0; scan_win2685 <= 32'd0; scan_win2686 <= 32'd0; scan_win2687 <= 32'd0; scan_win2688 <= 32'd0; scan_win2689 <= 32'd0; scan_win2690 <= 32'd0; scan_win2691 <= 32'd0; scan_win2692 <= 32'd0; scan_win2693 <= 32'd0; scan_win2694 <= 32'd0; scan_win2695 <= 32'd0; scan_win2696 <= 32'd0; scan_win2697 <= 32'd0; scan_win2698 <= 32'd0; scan_win2699 <= 32'd0; scan_win2700 <= 32'd0; scan_win2701 <= 32'd0; scan_win2702 <= 32'd0; scan_win2703 <= 32'd0; scan_win2704 <= 32'd0; scan_win2705 <= 32'd0; scan_win2706 <= 32'd0; scan_win2707 <= 32'd0; scan_win2708 <= 32'd0; scan_win2709 <= 32'd0; scan_win2710 <= 32'd0; scan_win2711 <= 32'd0; scan_win2712 <= 32'd0; scan_win2713 <= 32'd0; scan_win2714 <= 32'd0; scan_win2715 <= 32'd0; scan_win2716 <= 32'd0; scan_win2717 <= 32'd0; scan_win2718 <= 32'd0; scan_win2719 <= 32'd0; scan_win2720 <= 32'd0; scan_win2721 <= 32'd0; scan_win2722 <= 32'd0; scan_win2723 <= 32'd0; scan_win2724 <= 32'd0; scan_win2725 <= 32'd0; scan_win2726 <= 32'd0; scan_win2727 <= 32'd0; scan_win2728 <= 32'd0; scan_win2729 <= 32'd0; scan_win2730 <= 32'd0; scan_win2731 <= 32'd0; scan_win2732 <= 32'd0; scan_win2733 <= 32'd0; scan_win2734 <= 32'd0; scan_win2735 <= 32'd0; scan_win2736 <= 32'd0; scan_win2737 <= 32'd0; scan_win2738 <= 32'd0; scan_win2739 <= 32'd0; scan_win2740 <= 32'd0; scan_win2741 <= 32'd0; scan_win2742 <= 32'd0; scan_win2743 <= 32'd0; scan_win2744 <= 32'd0; scan_win2745 <= 32'd0; scan_win2746 <= 32'd0; scan_win2747 <= 32'd0; scan_win2748 <= 32'd0; scan_win2749 <= 32'd0; scan_win2750 <= 32'd0; scan_win2751 <= 32'd0; scan_win2752 <= 32'd0; scan_win2753 <= 32'd0; scan_win2754 <= 32'd0; scan_win2755 <= 32'd0; scan_win2756 <= 32'd0; scan_win2757 <= 32'd0; scan_win2758 <= 32'd0; scan_win2759 <= 32'd0; scan_win2760 <= 32'd0; scan_win2761 <= 32'd0; scan_win2762 <= 32'd0; scan_win2763 <= 32'd0; scan_win2764 <= 32'd0; scan_win2765 <= 32'd0; scan_win2766 <= 32'd0; scan_win2767 <= 32'd0; scan_win2768 <= 32'd0; scan_win2769 <= 32'd0; scan_win2770 <= 32'd0; scan_win2771 <= 32'd0; scan_win2772 <= 32'd0; scan_win2773 <= 32'd0; scan_win2774 <= 32'd0; scan_win2775 <= 32'd0; scan_win2776 <= 32'd0; scan_win2777 <= 32'd0; scan_win2778 <= 32'd0; scan_win2779 <= 32'd0; scan_win2780 <= 32'd0; scan_win2781 <= 32'd0; scan_win2782 <= 32'd0; scan_win2783 <= 32'd0; scan_win2784 <= 32'd0; scan_win2785 <= 32'd0; scan_win2786 <= 32'd0; scan_win2787 <= 32'd0; scan_win2788 <= 32'd0; scan_win2789 <= 32'd0; scan_win2790 <= 32'd0; scan_win2791 <= 32'd0; scan_win2792 <= 32'd0; scan_win2793 <= 32'd0; scan_win2794 <= 32'd0; scan_win2795 <= 32'd0; scan_win2796 <= 32'd0; scan_win2797 <= 32'd0; scan_win2798 <= 32'd0; scan_win2799 <= 32'd0; scan_win2800 <= 32'd0; 
      scan_win2801 <= 32'd0; scan_win2802 <= 32'd0; scan_win2803 <= 32'd0; scan_win2804 <= 32'd0; scan_win2805 <= 32'd0; scan_win2806 <= 32'd0; scan_win2807 <= 32'd0; scan_win2808 <= 32'd0; scan_win2809 <= 32'd0; scan_win2810 <= 32'd0; scan_win2811 <= 32'd0; scan_win2812 <= 32'd0; scan_win2813 <= 32'd0; scan_win2814 <= 32'd0; scan_win2815 <= 32'd0; scan_win2816 <= 32'd0; scan_win2817 <= 32'd0; scan_win2818 <= 32'd0; scan_win2819 <= 32'd0; scan_win2820 <= 32'd0; scan_win2821 <= 32'd0; scan_win2822 <= 32'd0; scan_win2823 <= 32'd0; scan_win2824 <= 32'd0; scan_win2825 <= 32'd0; scan_win2826 <= 32'd0; scan_win2827 <= 32'd0; scan_win2828 <= 32'd0; scan_win2829 <= 32'd0; scan_win2830 <= 32'd0; scan_win2831 <= 32'd0; scan_win2832 <= 32'd0; scan_win2833 <= 32'd0; scan_win2834 <= 32'd0; scan_win2835 <= 32'd0; scan_win2836 <= 32'd0; scan_win2837 <= 32'd0; scan_win2838 <= 32'd0; scan_win2839 <= 32'd0; scan_win2840 <= 32'd0; scan_win2841 <= 32'd0; scan_win2842 <= 32'd0; scan_win2843 <= 32'd0; scan_win2844 <= 32'd0; scan_win2845 <= 32'd0; scan_win2846 <= 32'd0; scan_win2847 <= 32'd0; scan_win2848 <= 32'd0; scan_win2849 <= 32'd0; scan_win2850 <= 32'd0; scan_win2851 <= 32'd0; scan_win2852 <= 32'd0; scan_win2853 <= 32'd0; scan_win2854 <= 32'd0; scan_win2855 <= 32'd0; scan_win2856 <= 32'd0; scan_win2857 <= 32'd0; scan_win2858 <= 32'd0; scan_win2859 <= 32'd0; scan_win2860 <= 32'd0; scan_win2861 <= 32'd0; scan_win2862 <= 32'd0; scan_win2863 <= 32'd0; scan_win2864 <= 32'd0; scan_win2865 <= 32'd0; scan_win2866 <= 32'd0; scan_win2867 <= 32'd0; scan_win2868 <= 32'd0; scan_win2869 <= 32'd0; scan_win2870 <= 32'd0; scan_win2871 <= 32'd0; scan_win2872 <= 32'd0; scan_win2873 <= 32'd0; scan_win2874 <= 32'd0; scan_win2875 <= 32'd0; scan_win2876 <= 32'd0; scan_win2877 <= 32'd0; scan_win2878 <= 32'd0; scan_win2879 <= 32'd0; scan_win2880 <= 32'd0; scan_win2881 <= 32'd0; scan_win2882 <= 32'd0; scan_win2883 <= 32'd0; scan_win2884 <= 32'd0; scan_win2885 <= 32'd0; scan_win2886 <= 32'd0; scan_win2887 <= 32'd0; scan_win2888 <= 32'd0; scan_win2889 <= 32'd0; scan_win2890 <= 32'd0; scan_win2891 <= 32'd0; scan_win2892 <= 32'd0; scan_win2893 <= 32'd0; scan_win2894 <= 32'd0; scan_win2895 <= 32'd0; scan_win2896 <= 32'd0; scan_win2897 <= 32'd0; scan_win2898 <= 32'd0; scan_win2899 <= 32'd0; scan_win2900 <= 32'd0; scan_win2901 <= 32'd0; scan_win2902 <= 32'd0; scan_win2903 <= 32'd0; scan_win2904 <= 32'd0; scan_win2905 <= 32'd0; scan_win2906 <= 32'd0; scan_win2907 <= 32'd0; scan_win2908 <= 32'd0; scan_win2909 <= 32'd0; scan_win2910 <= 32'd0; scan_win2911 <= 32'd0; scan_win2912 <= 32'd0;
    end else begin: move_scan_wins
      scan_win0 <= scan_win;
      scan_win1 <= scan_win0; scan_win2 <= scan_win1; scan_win3 <= scan_win2; scan_win4 <= scan_win3; scan_win5 <= scan_win4; scan_win6 <= scan_win5; scan_win7 <= scan_win6; scan_win8 <= scan_win7; scan_win9 <= scan_win8; scan_win10 <= scan_win9; scan_win11 <= scan_win10; scan_win12 <= scan_win11; scan_win13 <= scan_win12; scan_win14 <= scan_win13; scan_win15 <= scan_win14; scan_win16 <= scan_win15; scan_win17 <= scan_win16; scan_win18 <= scan_win17; scan_win19 <= scan_win18; scan_win20 <= scan_win19; scan_win21 <= scan_win20; scan_win22 <= scan_win21; scan_win23 <= scan_win22; scan_win24 <= scan_win23; scan_win25 <= scan_win24; scan_win26 <= scan_win25; scan_win27 <= scan_win26; scan_win28 <= scan_win27; scan_win29 <= scan_win28; scan_win30 <= scan_win29; scan_win31 <= scan_win30; scan_win32 <= scan_win31; scan_win33 <= scan_win32; scan_win34 <= scan_win33; scan_win35 <= scan_win34; scan_win36 <= scan_win35; scan_win37 <= scan_win36; scan_win38 <= scan_win37; scan_win39 <= scan_win38; scan_win40 <= scan_win39; scan_win41 <= scan_win40; scan_win42 <= scan_win41; scan_win43 <= scan_win42; scan_win44 <= scan_win43; scan_win45 <= scan_win44; scan_win46 <= scan_win45; scan_win47 <= scan_win46; scan_win48 <= scan_win47; scan_win49 <= scan_win48; scan_win50 <= scan_win49; scan_win51 <= scan_win50; scan_win52 <= scan_win51; scan_win53 <= scan_win52; scan_win54 <= scan_win53; scan_win55 <= scan_win54; scan_win56 <= scan_win55; scan_win57 <= scan_win56; scan_win58 <= scan_win57; scan_win59 <= scan_win58; scan_win60 <= scan_win59; scan_win61 <= scan_win60; scan_win62 <= scan_win61; scan_win63 <= scan_win62; scan_win64 <= scan_win63; scan_win65 <= scan_win64; scan_win66 <= scan_win65; scan_win67 <= scan_win66; scan_win68 <= scan_win67; scan_win69 <= scan_win68; scan_win70 <= scan_win69; scan_win71 <= scan_win70; scan_win72 <= scan_win71; scan_win73 <= scan_win72; scan_win74 <= scan_win73; scan_win75 <= scan_win74; scan_win76 <= scan_win75; scan_win77 <= scan_win76; scan_win78 <= scan_win77; scan_win79 <= scan_win78; scan_win80 <= scan_win79; scan_win81 <= scan_win80; scan_win82 <= scan_win81; scan_win83 <= scan_win82; scan_win84 <= scan_win83; scan_win85 <= scan_win84; scan_win86 <= scan_win85; scan_win87 <= scan_win86; scan_win88 <= scan_win87; scan_win89 <= scan_win88; scan_win90 <= scan_win89; scan_win91 <= scan_win90; scan_win92 <= scan_win91; scan_win93 <= scan_win92; scan_win94 <= scan_win93; scan_win95 <= scan_win94; scan_win96 <= scan_win95; scan_win97 <= scan_win96; scan_win98 <= scan_win97; scan_win99 <= scan_win98; scan_win100 <= scan_win99; scan_win101 <= scan_win100; scan_win102 <= scan_win101; scan_win103 <= scan_win102; scan_win104 <= scan_win103; scan_win105 <= scan_win104; scan_win106 <= scan_win105; scan_win107 <= scan_win106; scan_win108 <= scan_win107; scan_win109 <= scan_win108; scan_win110 <= scan_win109; scan_win111 <= scan_win110; scan_win112 <= scan_win111; scan_win113 <= scan_win112; scan_win114 <= scan_win113; scan_win115 <= scan_win114; scan_win116 <= scan_win115; scan_win117 <= scan_win116; scan_win118 <= scan_win117; scan_win119 <= scan_win118; scan_win120 <= scan_win119; scan_win121 <= scan_win120; scan_win122 <= scan_win121; scan_win123 <= scan_win122; scan_win124 <= scan_win123; scan_win125 <= scan_win124; scan_win126 <= scan_win125; scan_win127 <= scan_win126; scan_win128 <= scan_win127; scan_win129 <= scan_win128; scan_win130 <= scan_win129; scan_win131 <= scan_win130; scan_win132 <= scan_win131; scan_win133 <= scan_win132; scan_win134 <= scan_win133; scan_win135 <= scan_win134; scan_win136 <= scan_win135; scan_win137 <= scan_win136; scan_win138 <= scan_win137; scan_win139 <= scan_win138; scan_win140 <= scan_win139; scan_win141 <= scan_win140; scan_win142 <= scan_win141; scan_win143 <= scan_win142; scan_win144 <= scan_win143; scan_win145 <= scan_win144; scan_win146 <= scan_win145; scan_win147 <= scan_win146; scan_win148 <= scan_win147; scan_win149 <= scan_win148; scan_win150 <= scan_win149; scan_win151 <= scan_win150; scan_win152 <= scan_win151; scan_win153 <= scan_win152; scan_win154 <= scan_win153; scan_win155 <= scan_win154; scan_win156 <= scan_win155; scan_win157 <= scan_win156; scan_win158 <= scan_win157; scan_win159 <= scan_win158; scan_win160 <= scan_win159; scan_win161 <= scan_win160; scan_win162 <= scan_win161; scan_win163 <= scan_win162; scan_win164 <= scan_win163; scan_win165 <= scan_win164; scan_win166 <= scan_win165; scan_win167 <= scan_win166; scan_win168 <= scan_win167; scan_win169 <= scan_win168; scan_win170 <= scan_win169; scan_win171 <= scan_win170; scan_win172 <= scan_win171; scan_win173 <= scan_win172; scan_win174 <= scan_win173; scan_win175 <= scan_win174; scan_win176 <= scan_win175; scan_win177 <= scan_win176; scan_win178 <= scan_win177; scan_win179 <= scan_win178; scan_win180 <= scan_win179; scan_win181 <= scan_win180; scan_win182 <= scan_win181; scan_win183 <= scan_win182; scan_win184 <= scan_win183; scan_win185 <= scan_win184; scan_win186 <= scan_win185; scan_win187 <= scan_win186; scan_win188 <= scan_win187; scan_win189 <= scan_win188; scan_win190 <= scan_win189; scan_win191 <= scan_win190; scan_win192 <= scan_win191; scan_win193 <= scan_win192; scan_win194 <= scan_win193; scan_win195 <= scan_win194; scan_win196 <= scan_win195; scan_win197 <= scan_win196; scan_win198 <= scan_win197; scan_win199 <= scan_win198; scan_win200 <= scan_win199; 
      scan_win201 <= scan_win200; scan_win202 <= scan_win201; scan_win203 <= scan_win202; scan_win204 <= scan_win203; scan_win205 <= scan_win204; scan_win206 <= scan_win205; scan_win207 <= scan_win206; scan_win208 <= scan_win207; scan_win209 <= scan_win208; scan_win210 <= scan_win209; scan_win211 <= scan_win210; scan_win212 <= scan_win211; scan_win213 <= scan_win212; scan_win214 <= scan_win213; scan_win215 <= scan_win214; scan_win216 <= scan_win215; scan_win217 <= scan_win216; scan_win218 <= scan_win217; scan_win219 <= scan_win218; scan_win220 <= scan_win219; scan_win221 <= scan_win220; scan_win222 <= scan_win221; scan_win223 <= scan_win222; scan_win224 <= scan_win223; scan_win225 <= scan_win224; scan_win226 <= scan_win225; scan_win227 <= scan_win226; scan_win228 <= scan_win227; scan_win229 <= scan_win228; scan_win230 <= scan_win229; scan_win231 <= scan_win230; scan_win232 <= scan_win231; scan_win233 <= scan_win232; scan_win234 <= scan_win233; scan_win235 <= scan_win234; scan_win236 <= scan_win235; scan_win237 <= scan_win236; scan_win238 <= scan_win237; scan_win239 <= scan_win238; scan_win240 <= scan_win239; scan_win241 <= scan_win240; scan_win242 <= scan_win241; scan_win243 <= scan_win242; scan_win244 <= scan_win243; scan_win245 <= scan_win244; scan_win246 <= scan_win245; scan_win247 <= scan_win246; scan_win248 <= scan_win247; scan_win249 <= scan_win248; scan_win250 <= scan_win249; scan_win251 <= scan_win250; scan_win252 <= scan_win251; scan_win253 <= scan_win252; scan_win254 <= scan_win253; scan_win255 <= scan_win254; scan_win256 <= scan_win255; scan_win257 <= scan_win256; scan_win258 <= scan_win257; scan_win259 <= scan_win258; scan_win260 <= scan_win259; scan_win261 <= scan_win260; scan_win262 <= scan_win261; scan_win263 <= scan_win262; scan_win264 <= scan_win263; scan_win265 <= scan_win264; scan_win266 <= scan_win265; scan_win267 <= scan_win266; scan_win268 <= scan_win267; scan_win269 <= scan_win268; scan_win270 <= scan_win269; scan_win271 <= scan_win270; scan_win272 <= scan_win271; scan_win273 <= scan_win272; scan_win274 <= scan_win273; scan_win275 <= scan_win274; scan_win276 <= scan_win275; scan_win277 <= scan_win276; scan_win278 <= scan_win277; scan_win279 <= scan_win278; scan_win280 <= scan_win279; scan_win281 <= scan_win280; scan_win282 <= scan_win281; scan_win283 <= scan_win282; scan_win284 <= scan_win283; scan_win285 <= scan_win284; scan_win286 <= scan_win285; scan_win287 <= scan_win286; scan_win288 <= scan_win287; scan_win289 <= scan_win288; scan_win290 <= scan_win289; scan_win291 <= scan_win290; scan_win292 <= scan_win291; scan_win293 <= scan_win292; scan_win294 <= scan_win293; scan_win295 <= scan_win294; scan_win296 <= scan_win295; scan_win297 <= scan_win296; scan_win298 <= scan_win297; scan_win299 <= scan_win298; scan_win300 <= scan_win299; scan_win301 <= scan_win300; scan_win302 <= scan_win301; scan_win303 <= scan_win302; scan_win304 <= scan_win303; scan_win305 <= scan_win304; scan_win306 <= scan_win305; scan_win307 <= scan_win306; scan_win308 <= scan_win307; scan_win309 <= scan_win308; scan_win310 <= scan_win309; scan_win311 <= scan_win310; scan_win312 <= scan_win311; scan_win313 <= scan_win312; scan_win314 <= scan_win313; scan_win315 <= scan_win314; scan_win316 <= scan_win315; scan_win317 <= scan_win316; scan_win318 <= scan_win317; scan_win319 <= scan_win318; scan_win320 <= scan_win319; scan_win321 <= scan_win320; scan_win322 <= scan_win321; scan_win323 <= scan_win322; scan_win324 <= scan_win323; scan_win325 <= scan_win324; scan_win326 <= scan_win325; scan_win327 <= scan_win326; scan_win328 <= scan_win327; scan_win329 <= scan_win328; scan_win330 <= scan_win329; scan_win331 <= scan_win330; scan_win332 <= scan_win331; scan_win333 <= scan_win332; scan_win334 <= scan_win333; scan_win335 <= scan_win334; scan_win336 <= scan_win335; scan_win337 <= scan_win336; scan_win338 <= scan_win337; scan_win339 <= scan_win338; scan_win340 <= scan_win339; scan_win341 <= scan_win340; scan_win342 <= scan_win341; scan_win343 <= scan_win342; scan_win344 <= scan_win343; scan_win345 <= scan_win344; scan_win346 <= scan_win345; scan_win347 <= scan_win346; scan_win348 <= scan_win347; scan_win349 <= scan_win348; scan_win350 <= scan_win349; scan_win351 <= scan_win350; scan_win352 <= scan_win351; scan_win353 <= scan_win352; scan_win354 <= scan_win353; scan_win355 <= scan_win354; scan_win356 <= scan_win355; scan_win357 <= scan_win356; scan_win358 <= scan_win357; scan_win359 <= scan_win358; scan_win360 <= scan_win359; scan_win361 <= scan_win360; scan_win362 <= scan_win361; scan_win363 <= scan_win362; scan_win364 <= scan_win363; scan_win365 <= scan_win364; scan_win366 <= scan_win365; scan_win367 <= scan_win366; scan_win368 <= scan_win367; scan_win369 <= scan_win368; scan_win370 <= scan_win369; scan_win371 <= scan_win370; scan_win372 <= scan_win371; scan_win373 <= scan_win372; scan_win374 <= scan_win373; scan_win375 <= scan_win374; scan_win376 <= scan_win375; scan_win377 <= scan_win376; scan_win378 <= scan_win377; scan_win379 <= scan_win378; scan_win380 <= scan_win379; scan_win381 <= scan_win380; scan_win382 <= scan_win381; scan_win383 <= scan_win382; scan_win384 <= scan_win383; scan_win385 <= scan_win384; scan_win386 <= scan_win385; scan_win387 <= scan_win386; scan_win388 <= scan_win387; scan_win389 <= scan_win388; scan_win390 <= scan_win389; scan_win391 <= scan_win390; scan_win392 <= scan_win391; scan_win393 <= scan_win392; scan_win394 <= scan_win393; scan_win395 <= scan_win394; scan_win396 <= scan_win395; scan_win397 <= scan_win396; scan_win398 <= scan_win397; scan_win399 <= scan_win398; scan_win400 <= scan_win399; 
      scan_win401 <= scan_win400; scan_win402 <= scan_win401; scan_win403 <= scan_win402; scan_win404 <= scan_win403; scan_win405 <= scan_win404; scan_win406 <= scan_win405; scan_win407 <= scan_win406; scan_win408 <= scan_win407; scan_win409 <= scan_win408; scan_win410 <= scan_win409; scan_win411 <= scan_win410; scan_win412 <= scan_win411; scan_win413 <= scan_win412; scan_win414 <= scan_win413; scan_win415 <= scan_win414; scan_win416 <= scan_win415; scan_win417 <= scan_win416; scan_win418 <= scan_win417; scan_win419 <= scan_win418; scan_win420 <= scan_win419; scan_win421 <= scan_win420; scan_win422 <= scan_win421; scan_win423 <= scan_win422; scan_win424 <= scan_win423; scan_win425 <= scan_win424; scan_win426 <= scan_win425; scan_win427 <= scan_win426; scan_win428 <= scan_win427; scan_win429 <= scan_win428; scan_win430 <= scan_win429; scan_win431 <= scan_win430; scan_win432 <= scan_win431; scan_win433 <= scan_win432; scan_win434 <= scan_win433; scan_win435 <= scan_win434; scan_win436 <= scan_win435; scan_win437 <= scan_win436; scan_win438 <= scan_win437; scan_win439 <= scan_win438; scan_win440 <= scan_win439; scan_win441 <= scan_win440; scan_win442 <= scan_win441; scan_win443 <= scan_win442; scan_win444 <= scan_win443; scan_win445 <= scan_win444; scan_win446 <= scan_win445; scan_win447 <= scan_win446; scan_win448 <= scan_win447; scan_win449 <= scan_win448; scan_win450 <= scan_win449; scan_win451 <= scan_win450; scan_win452 <= scan_win451; scan_win453 <= scan_win452; scan_win454 <= scan_win453; scan_win455 <= scan_win454; scan_win456 <= scan_win455; scan_win457 <= scan_win456; scan_win458 <= scan_win457; scan_win459 <= scan_win458; scan_win460 <= scan_win459; scan_win461 <= scan_win460; scan_win462 <= scan_win461; scan_win463 <= scan_win462; scan_win464 <= scan_win463; scan_win465 <= scan_win464; scan_win466 <= scan_win465; scan_win467 <= scan_win466; scan_win468 <= scan_win467; scan_win469 <= scan_win468; scan_win470 <= scan_win469; scan_win471 <= scan_win470; scan_win472 <= scan_win471; scan_win473 <= scan_win472; scan_win474 <= scan_win473; scan_win475 <= scan_win474; scan_win476 <= scan_win475; scan_win477 <= scan_win476; scan_win478 <= scan_win477; scan_win479 <= scan_win478; scan_win480 <= scan_win479; scan_win481 <= scan_win480; scan_win482 <= scan_win481; scan_win483 <= scan_win482; scan_win484 <= scan_win483; scan_win485 <= scan_win484; scan_win486 <= scan_win485; scan_win487 <= scan_win486; scan_win488 <= scan_win487; scan_win489 <= scan_win488; scan_win490 <= scan_win489; scan_win491 <= scan_win490; scan_win492 <= scan_win491; scan_win493 <= scan_win492; scan_win494 <= scan_win493; scan_win495 <= scan_win494; scan_win496 <= scan_win495; scan_win497 <= scan_win496; scan_win498 <= scan_win497; scan_win499 <= scan_win498; scan_win500 <= scan_win499; scan_win501 <= scan_win500; scan_win502 <= scan_win501; scan_win503 <= scan_win502; scan_win504 <= scan_win503; scan_win505 <= scan_win504; scan_win506 <= scan_win505; scan_win507 <= scan_win506; scan_win508 <= scan_win507; scan_win509 <= scan_win508; scan_win510 <= scan_win509; scan_win511 <= scan_win510; scan_win512 <= scan_win511; scan_win513 <= scan_win512; scan_win514 <= scan_win513; scan_win515 <= scan_win514; scan_win516 <= scan_win515; scan_win517 <= scan_win516; scan_win518 <= scan_win517; scan_win519 <= scan_win518; scan_win520 <= scan_win519; scan_win521 <= scan_win520; scan_win522 <= scan_win521; scan_win523 <= scan_win522; scan_win524 <= scan_win523; scan_win525 <= scan_win524; scan_win526 <= scan_win525; scan_win527 <= scan_win526; scan_win528 <= scan_win527; scan_win529 <= scan_win528; scan_win530 <= scan_win529; scan_win531 <= scan_win530; scan_win532 <= scan_win531; scan_win533 <= scan_win532; scan_win534 <= scan_win533; scan_win535 <= scan_win534; scan_win536 <= scan_win535; scan_win537 <= scan_win536; scan_win538 <= scan_win537; scan_win539 <= scan_win538; scan_win540 <= scan_win539; scan_win541 <= scan_win540; scan_win542 <= scan_win541; scan_win543 <= scan_win542; scan_win544 <= scan_win543; scan_win545 <= scan_win544; scan_win546 <= scan_win545; scan_win547 <= scan_win546; scan_win548 <= scan_win547; scan_win549 <= scan_win548; scan_win550 <= scan_win549; scan_win551 <= scan_win550; scan_win552 <= scan_win551; scan_win553 <= scan_win552; scan_win554 <= scan_win553; scan_win555 <= scan_win554; scan_win556 <= scan_win555; scan_win557 <= scan_win556; scan_win558 <= scan_win557; scan_win559 <= scan_win558; scan_win560 <= scan_win559; scan_win561 <= scan_win560; scan_win562 <= scan_win561; scan_win563 <= scan_win562; scan_win564 <= scan_win563; scan_win565 <= scan_win564; scan_win566 <= scan_win565; scan_win567 <= scan_win566; scan_win568 <= scan_win567; scan_win569 <= scan_win568; scan_win570 <= scan_win569; scan_win571 <= scan_win570; scan_win572 <= scan_win571; scan_win573 <= scan_win572; scan_win574 <= scan_win573; scan_win575 <= scan_win574; scan_win576 <= scan_win575; scan_win577 <= scan_win576; scan_win578 <= scan_win577; scan_win579 <= scan_win578; scan_win580 <= scan_win579; scan_win581 <= scan_win580; scan_win582 <= scan_win581; scan_win583 <= scan_win582; scan_win584 <= scan_win583; scan_win585 <= scan_win584; scan_win586 <= scan_win585; scan_win587 <= scan_win586; scan_win588 <= scan_win587; scan_win589 <= scan_win588; scan_win590 <= scan_win589; scan_win591 <= scan_win590; scan_win592 <= scan_win591; scan_win593 <= scan_win592; scan_win594 <= scan_win593; scan_win595 <= scan_win594; scan_win596 <= scan_win595; scan_win597 <= scan_win596; scan_win598 <= scan_win597; scan_win599 <= scan_win598; scan_win600 <= scan_win599; 
      scan_win601 <= scan_win600; scan_win602 <= scan_win601; scan_win603 <= scan_win602; scan_win604 <= scan_win603; scan_win605 <= scan_win604; scan_win606 <= scan_win605; scan_win607 <= scan_win606; scan_win608 <= scan_win607; scan_win609 <= scan_win608; scan_win610 <= scan_win609; scan_win611 <= scan_win610; scan_win612 <= scan_win611; scan_win613 <= scan_win612; scan_win614 <= scan_win613; scan_win615 <= scan_win614; scan_win616 <= scan_win615; scan_win617 <= scan_win616; scan_win618 <= scan_win617; scan_win619 <= scan_win618; scan_win620 <= scan_win619; scan_win621 <= scan_win620; scan_win622 <= scan_win621; scan_win623 <= scan_win622; scan_win624 <= scan_win623; scan_win625 <= scan_win624; scan_win626 <= scan_win625; scan_win627 <= scan_win626; scan_win628 <= scan_win627; scan_win629 <= scan_win628; scan_win630 <= scan_win629; scan_win631 <= scan_win630; scan_win632 <= scan_win631; scan_win633 <= scan_win632; scan_win634 <= scan_win633; scan_win635 <= scan_win634; scan_win636 <= scan_win635; scan_win637 <= scan_win636; scan_win638 <= scan_win637; scan_win639 <= scan_win638; scan_win640 <= scan_win639; scan_win641 <= scan_win640; scan_win642 <= scan_win641; scan_win643 <= scan_win642; scan_win644 <= scan_win643; scan_win645 <= scan_win644; scan_win646 <= scan_win645; scan_win647 <= scan_win646; scan_win648 <= scan_win647; scan_win649 <= scan_win648; scan_win650 <= scan_win649; scan_win651 <= scan_win650; scan_win652 <= scan_win651; scan_win653 <= scan_win652; scan_win654 <= scan_win653; scan_win655 <= scan_win654; scan_win656 <= scan_win655; scan_win657 <= scan_win656; scan_win658 <= scan_win657; scan_win659 <= scan_win658; scan_win660 <= scan_win659; scan_win661 <= scan_win660; scan_win662 <= scan_win661; scan_win663 <= scan_win662; scan_win664 <= scan_win663; scan_win665 <= scan_win664; scan_win666 <= scan_win665; scan_win667 <= scan_win666; scan_win668 <= scan_win667; scan_win669 <= scan_win668; scan_win670 <= scan_win669; scan_win671 <= scan_win670; scan_win672 <= scan_win671; scan_win673 <= scan_win672; scan_win674 <= scan_win673; scan_win675 <= scan_win674; scan_win676 <= scan_win675; scan_win677 <= scan_win676; scan_win678 <= scan_win677; scan_win679 <= scan_win678; scan_win680 <= scan_win679; scan_win681 <= scan_win680; scan_win682 <= scan_win681; scan_win683 <= scan_win682; scan_win684 <= scan_win683; scan_win685 <= scan_win684; scan_win686 <= scan_win685; scan_win687 <= scan_win686; scan_win688 <= scan_win687; scan_win689 <= scan_win688; scan_win690 <= scan_win689; scan_win691 <= scan_win690; scan_win692 <= scan_win691; scan_win693 <= scan_win692; scan_win694 <= scan_win693; scan_win695 <= scan_win694; scan_win696 <= scan_win695; scan_win697 <= scan_win696; scan_win698 <= scan_win697; scan_win699 <= scan_win698; scan_win700 <= scan_win699; scan_win701 <= scan_win700; scan_win702 <= scan_win701; scan_win703 <= scan_win702; scan_win704 <= scan_win703; scan_win705 <= scan_win704; scan_win706 <= scan_win705; scan_win707 <= scan_win706; scan_win708 <= scan_win707; scan_win709 <= scan_win708; scan_win710 <= scan_win709; scan_win711 <= scan_win710; scan_win712 <= scan_win711; scan_win713 <= scan_win712; scan_win714 <= scan_win713; scan_win715 <= scan_win714; scan_win716 <= scan_win715; scan_win717 <= scan_win716; scan_win718 <= scan_win717; scan_win719 <= scan_win718; scan_win720 <= scan_win719; scan_win721 <= scan_win720; scan_win722 <= scan_win721; scan_win723 <= scan_win722; scan_win724 <= scan_win723; scan_win725 <= scan_win724; scan_win726 <= scan_win725; scan_win727 <= scan_win726; scan_win728 <= scan_win727; scan_win729 <= scan_win728; scan_win730 <= scan_win729; scan_win731 <= scan_win730; scan_win732 <= scan_win731; scan_win733 <= scan_win732; scan_win734 <= scan_win733; scan_win735 <= scan_win734; scan_win736 <= scan_win735; scan_win737 <= scan_win736; scan_win738 <= scan_win737; scan_win739 <= scan_win738; scan_win740 <= scan_win739; scan_win741 <= scan_win740; scan_win742 <= scan_win741; scan_win743 <= scan_win742; scan_win744 <= scan_win743; scan_win745 <= scan_win744; scan_win746 <= scan_win745; scan_win747 <= scan_win746; scan_win748 <= scan_win747; scan_win749 <= scan_win748; scan_win750 <= scan_win749; scan_win751 <= scan_win750; scan_win752 <= scan_win751; scan_win753 <= scan_win752; scan_win754 <= scan_win753; scan_win755 <= scan_win754; scan_win756 <= scan_win755; scan_win757 <= scan_win756; scan_win758 <= scan_win757; scan_win759 <= scan_win758; scan_win760 <= scan_win759; scan_win761 <= scan_win760; scan_win762 <= scan_win761; scan_win763 <= scan_win762; scan_win764 <= scan_win763; scan_win765 <= scan_win764; scan_win766 <= scan_win765; scan_win767 <= scan_win766; scan_win768 <= scan_win767; scan_win769 <= scan_win768; scan_win770 <= scan_win769; scan_win771 <= scan_win770; scan_win772 <= scan_win771; scan_win773 <= scan_win772; scan_win774 <= scan_win773; scan_win775 <= scan_win774; scan_win776 <= scan_win775; scan_win777 <= scan_win776; scan_win778 <= scan_win777; scan_win779 <= scan_win778; scan_win780 <= scan_win779; scan_win781 <= scan_win780; scan_win782 <= scan_win781; scan_win783 <= scan_win782; scan_win784 <= scan_win783; scan_win785 <= scan_win784; scan_win786 <= scan_win785; scan_win787 <= scan_win786; scan_win788 <= scan_win787; scan_win789 <= scan_win788; scan_win790 <= scan_win789; scan_win791 <= scan_win790; scan_win792 <= scan_win791; scan_win793 <= scan_win792; scan_win794 <= scan_win793; scan_win795 <= scan_win794; scan_win796 <= scan_win795; scan_win797 <= scan_win796; scan_win798 <= scan_win797; scan_win799 <= scan_win798; scan_win800 <= scan_win799; 
      scan_win801 <= scan_win800; scan_win802 <= scan_win801; scan_win803 <= scan_win802; scan_win804 <= scan_win803; scan_win805 <= scan_win804; scan_win806 <= scan_win805; scan_win807 <= scan_win806; scan_win808 <= scan_win807; scan_win809 <= scan_win808; scan_win810 <= scan_win809; scan_win811 <= scan_win810; scan_win812 <= scan_win811; scan_win813 <= scan_win812; scan_win814 <= scan_win813; scan_win815 <= scan_win814; scan_win816 <= scan_win815; scan_win817 <= scan_win816; scan_win818 <= scan_win817; scan_win819 <= scan_win818; scan_win820 <= scan_win819; scan_win821 <= scan_win820; scan_win822 <= scan_win821; scan_win823 <= scan_win822; scan_win824 <= scan_win823; scan_win825 <= scan_win824; scan_win826 <= scan_win825; scan_win827 <= scan_win826; scan_win828 <= scan_win827; scan_win829 <= scan_win828; scan_win830 <= scan_win829; scan_win831 <= scan_win830; scan_win832 <= scan_win831; scan_win833 <= scan_win832; scan_win834 <= scan_win833; scan_win835 <= scan_win834; scan_win836 <= scan_win835; scan_win837 <= scan_win836; scan_win838 <= scan_win837; scan_win839 <= scan_win838; scan_win840 <= scan_win839; scan_win841 <= scan_win840; scan_win842 <= scan_win841; scan_win843 <= scan_win842; scan_win844 <= scan_win843; scan_win845 <= scan_win844; scan_win846 <= scan_win845; scan_win847 <= scan_win846; scan_win848 <= scan_win847; scan_win849 <= scan_win848; scan_win850 <= scan_win849; scan_win851 <= scan_win850; scan_win852 <= scan_win851; scan_win853 <= scan_win852; scan_win854 <= scan_win853; scan_win855 <= scan_win854; scan_win856 <= scan_win855; scan_win857 <= scan_win856; scan_win858 <= scan_win857; scan_win859 <= scan_win858; scan_win860 <= scan_win859; scan_win861 <= scan_win860; scan_win862 <= scan_win861; scan_win863 <= scan_win862; scan_win864 <= scan_win863; scan_win865 <= scan_win864; scan_win866 <= scan_win865; scan_win867 <= scan_win866; scan_win868 <= scan_win867; scan_win869 <= scan_win868; scan_win870 <= scan_win869; scan_win871 <= scan_win870; scan_win872 <= scan_win871; scan_win873 <= scan_win872; scan_win874 <= scan_win873; scan_win875 <= scan_win874; scan_win876 <= scan_win875; scan_win877 <= scan_win876; scan_win878 <= scan_win877; scan_win879 <= scan_win878; scan_win880 <= scan_win879; scan_win881 <= scan_win880; scan_win882 <= scan_win881; scan_win883 <= scan_win882; scan_win884 <= scan_win883; scan_win885 <= scan_win884; scan_win886 <= scan_win885; scan_win887 <= scan_win886; scan_win888 <= scan_win887; scan_win889 <= scan_win888; scan_win890 <= scan_win889; scan_win891 <= scan_win890; scan_win892 <= scan_win891; scan_win893 <= scan_win892; scan_win894 <= scan_win893; scan_win895 <= scan_win894; scan_win896 <= scan_win895; scan_win897 <= scan_win896; scan_win898 <= scan_win897; scan_win899 <= scan_win898; scan_win900 <= scan_win899; scan_win901 <= scan_win900; scan_win902 <= scan_win901; scan_win903 <= scan_win902; scan_win904 <= scan_win903; scan_win905 <= scan_win904; scan_win906 <= scan_win905; scan_win907 <= scan_win906; scan_win908 <= scan_win907; scan_win909 <= scan_win908; scan_win910 <= scan_win909; scan_win911 <= scan_win910; scan_win912 <= scan_win911; scan_win913 <= scan_win912; scan_win914 <= scan_win913; scan_win915 <= scan_win914; scan_win916 <= scan_win915; scan_win917 <= scan_win916; scan_win918 <= scan_win917; scan_win919 <= scan_win918; scan_win920 <= scan_win919; scan_win921 <= scan_win920; scan_win922 <= scan_win921; scan_win923 <= scan_win922; scan_win924 <= scan_win923; scan_win925 <= scan_win924; scan_win926 <= scan_win925; scan_win927 <= scan_win926; scan_win928 <= scan_win927; scan_win929 <= scan_win928; scan_win930 <= scan_win929; scan_win931 <= scan_win930; scan_win932 <= scan_win931; scan_win933 <= scan_win932; scan_win934 <= scan_win933; scan_win935 <= scan_win934; scan_win936 <= scan_win935; scan_win937 <= scan_win936; scan_win938 <= scan_win937; scan_win939 <= scan_win938; scan_win940 <= scan_win939; scan_win941 <= scan_win940; scan_win942 <= scan_win941; scan_win943 <= scan_win942; scan_win944 <= scan_win943; scan_win945 <= scan_win944; scan_win946 <= scan_win945; scan_win947 <= scan_win946; scan_win948 <= scan_win947; scan_win949 <= scan_win948; scan_win950 <= scan_win949; scan_win951 <= scan_win950; scan_win952 <= scan_win951; scan_win953 <= scan_win952; scan_win954 <= scan_win953; scan_win955 <= scan_win954; scan_win956 <= scan_win955; scan_win957 <= scan_win956; scan_win958 <= scan_win957; scan_win959 <= scan_win958; scan_win960 <= scan_win959; scan_win961 <= scan_win960; scan_win962 <= scan_win961; scan_win963 <= scan_win962; scan_win964 <= scan_win963; scan_win965 <= scan_win964; scan_win966 <= scan_win965; scan_win967 <= scan_win966; scan_win968 <= scan_win967; scan_win969 <= scan_win968; scan_win970 <= scan_win969; scan_win971 <= scan_win970; scan_win972 <= scan_win971; scan_win973 <= scan_win972; scan_win974 <= scan_win973; scan_win975 <= scan_win974; scan_win976 <= scan_win975; scan_win977 <= scan_win976; scan_win978 <= scan_win977; scan_win979 <= scan_win978; scan_win980 <= scan_win979; scan_win981 <= scan_win980; scan_win982 <= scan_win981; scan_win983 <= scan_win982; scan_win984 <= scan_win983; scan_win985 <= scan_win984; scan_win986 <= scan_win985; scan_win987 <= scan_win986; scan_win988 <= scan_win987; scan_win989 <= scan_win988; scan_win990 <= scan_win989; scan_win991 <= scan_win990; scan_win992 <= scan_win991; scan_win993 <= scan_win992; scan_win994 <= scan_win993; scan_win995 <= scan_win994; scan_win996 <= scan_win995; scan_win997 <= scan_win996; scan_win998 <= scan_win997; scan_win999 <= scan_win998; scan_win1000 <= scan_win999; 
      scan_win1001 <= scan_win1000; scan_win1002 <= scan_win1001; scan_win1003 <= scan_win1002; scan_win1004 <= scan_win1003; scan_win1005 <= scan_win1004; scan_win1006 <= scan_win1005; scan_win1007 <= scan_win1006; scan_win1008 <= scan_win1007; scan_win1009 <= scan_win1008; scan_win1010 <= scan_win1009; scan_win1011 <= scan_win1010; scan_win1012 <= scan_win1011; scan_win1013 <= scan_win1012; scan_win1014 <= scan_win1013; scan_win1015 <= scan_win1014; scan_win1016 <= scan_win1015; scan_win1017 <= scan_win1016; scan_win1018 <= scan_win1017; scan_win1019 <= scan_win1018; scan_win1020 <= scan_win1019; scan_win1021 <= scan_win1020; scan_win1022 <= scan_win1021; scan_win1023 <= scan_win1022; scan_win1024 <= scan_win1023; scan_win1025 <= scan_win1024; scan_win1026 <= scan_win1025; scan_win1027 <= scan_win1026; scan_win1028 <= scan_win1027; scan_win1029 <= scan_win1028; scan_win1030 <= scan_win1029; scan_win1031 <= scan_win1030; scan_win1032 <= scan_win1031; scan_win1033 <= scan_win1032; scan_win1034 <= scan_win1033; scan_win1035 <= scan_win1034; scan_win1036 <= scan_win1035; scan_win1037 <= scan_win1036; scan_win1038 <= scan_win1037; scan_win1039 <= scan_win1038; scan_win1040 <= scan_win1039; scan_win1041 <= scan_win1040; scan_win1042 <= scan_win1041; scan_win1043 <= scan_win1042; scan_win1044 <= scan_win1043; scan_win1045 <= scan_win1044; scan_win1046 <= scan_win1045; scan_win1047 <= scan_win1046; scan_win1048 <= scan_win1047; scan_win1049 <= scan_win1048; scan_win1050 <= scan_win1049; scan_win1051 <= scan_win1050; scan_win1052 <= scan_win1051; scan_win1053 <= scan_win1052; scan_win1054 <= scan_win1053; scan_win1055 <= scan_win1054; scan_win1056 <= scan_win1055; scan_win1057 <= scan_win1056; scan_win1058 <= scan_win1057; scan_win1059 <= scan_win1058; scan_win1060 <= scan_win1059; scan_win1061 <= scan_win1060; scan_win1062 <= scan_win1061; scan_win1063 <= scan_win1062; scan_win1064 <= scan_win1063; scan_win1065 <= scan_win1064; scan_win1066 <= scan_win1065; scan_win1067 <= scan_win1066; scan_win1068 <= scan_win1067; scan_win1069 <= scan_win1068; scan_win1070 <= scan_win1069; scan_win1071 <= scan_win1070; scan_win1072 <= scan_win1071; scan_win1073 <= scan_win1072; scan_win1074 <= scan_win1073; scan_win1075 <= scan_win1074; scan_win1076 <= scan_win1075; scan_win1077 <= scan_win1076; scan_win1078 <= scan_win1077; scan_win1079 <= scan_win1078; scan_win1080 <= scan_win1079; scan_win1081 <= scan_win1080; scan_win1082 <= scan_win1081; scan_win1083 <= scan_win1082; scan_win1084 <= scan_win1083; scan_win1085 <= scan_win1084; scan_win1086 <= scan_win1085; scan_win1087 <= scan_win1086; scan_win1088 <= scan_win1087; scan_win1089 <= scan_win1088; scan_win1090 <= scan_win1089; scan_win1091 <= scan_win1090; scan_win1092 <= scan_win1091; scan_win1093 <= scan_win1092; scan_win1094 <= scan_win1093; scan_win1095 <= scan_win1094; scan_win1096 <= scan_win1095; scan_win1097 <= scan_win1096; scan_win1098 <= scan_win1097; scan_win1099 <= scan_win1098; scan_win1100 <= scan_win1099; scan_win1101 <= scan_win1100; scan_win1102 <= scan_win1101; scan_win1103 <= scan_win1102; scan_win1104 <= scan_win1103; scan_win1105 <= scan_win1104; scan_win1106 <= scan_win1105; scan_win1107 <= scan_win1106; scan_win1108 <= scan_win1107; scan_win1109 <= scan_win1108; scan_win1110 <= scan_win1109; scan_win1111 <= scan_win1110; scan_win1112 <= scan_win1111; scan_win1113 <= scan_win1112; scan_win1114 <= scan_win1113; scan_win1115 <= scan_win1114; scan_win1116 <= scan_win1115; scan_win1117 <= scan_win1116; scan_win1118 <= scan_win1117; scan_win1119 <= scan_win1118; scan_win1120 <= scan_win1119; scan_win1121 <= scan_win1120; scan_win1122 <= scan_win1121; scan_win1123 <= scan_win1122; scan_win1124 <= scan_win1123; scan_win1125 <= scan_win1124; scan_win1126 <= scan_win1125; scan_win1127 <= scan_win1126; scan_win1128 <= scan_win1127; scan_win1129 <= scan_win1128; scan_win1130 <= scan_win1129; scan_win1131 <= scan_win1130; scan_win1132 <= scan_win1131; scan_win1133 <= scan_win1132; scan_win1134 <= scan_win1133; scan_win1135 <= scan_win1134; scan_win1136 <= scan_win1135; scan_win1137 <= scan_win1136; scan_win1138 <= scan_win1137; scan_win1139 <= scan_win1138; scan_win1140 <= scan_win1139; scan_win1141 <= scan_win1140; scan_win1142 <= scan_win1141; scan_win1143 <= scan_win1142; scan_win1144 <= scan_win1143; scan_win1145 <= scan_win1144; scan_win1146 <= scan_win1145; scan_win1147 <= scan_win1146; scan_win1148 <= scan_win1147; scan_win1149 <= scan_win1148; scan_win1150 <= scan_win1149; scan_win1151 <= scan_win1150; scan_win1152 <= scan_win1151; scan_win1153 <= scan_win1152; scan_win1154 <= scan_win1153; scan_win1155 <= scan_win1154; scan_win1156 <= scan_win1155; scan_win1157 <= scan_win1156; scan_win1158 <= scan_win1157; scan_win1159 <= scan_win1158; scan_win1160 <= scan_win1159; scan_win1161 <= scan_win1160; scan_win1162 <= scan_win1161; scan_win1163 <= scan_win1162; scan_win1164 <= scan_win1163; scan_win1165 <= scan_win1164; scan_win1166 <= scan_win1165; scan_win1167 <= scan_win1166; scan_win1168 <= scan_win1167; scan_win1169 <= scan_win1168; scan_win1170 <= scan_win1169; scan_win1171 <= scan_win1170; scan_win1172 <= scan_win1171; scan_win1173 <= scan_win1172; scan_win1174 <= scan_win1173; scan_win1175 <= scan_win1174; scan_win1176 <= scan_win1175; scan_win1177 <= scan_win1176; scan_win1178 <= scan_win1177; scan_win1179 <= scan_win1178; scan_win1180 <= scan_win1179; scan_win1181 <= scan_win1180; scan_win1182 <= scan_win1181; scan_win1183 <= scan_win1182; scan_win1184 <= scan_win1183; scan_win1185 <= scan_win1184; scan_win1186 <= scan_win1185; scan_win1187 <= scan_win1186; scan_win1188 <= scan_win1187; scan_win1189 <= scan_win1188; scan_win1190 <= scan_win1189; scan_win1191 <= scan_win1190; scan_win1192 <= scan_win1191; scan_win1193 <= scan_win1192; scan_win1194 <= scan_win1193; scan_win1195 <= scan_win1194; scan_win1196 <= scan_win1195; scan_win1197 <= scan_win1196; scan_win1198 <= scan_win1197; scan_win1199 <= scan_win1198; scan_win1200 <= scan_win1199; 
      scan_win1201 <= scan_win1200; scan_win1202 <= scan_win1201; scan_win1203 <= scan_win1202; scan_win1204 <= scan_win1203; scan_win1205 <= scan_win1204; scan_win1206 <= scan_win1205; scan_win1207 <= scan_win1206; scan_win1208 <= scan_win1207; scan_win1209 <= scan_win1208; scan_win1210 <= scan_win1209; scan_win1211 <= scan_win1210; scan_win1212 <= scan_win1211; scan_win1213 <= scan_win1212; scan_win1214 <= scan_win1213; scan_win1215 <= scan_win1214; scan_win1216 <= scan_win1215; scan_win1217 <= scan_win1216; scan_win1218 <= scan_win1217; scan_win1219 <= scan_win1218; scan_win1220 <= scan_win1219; scan_win1221 <= scan_win1220; scan_win1222 <= scan_win1221; scan_win1223 <= scan_win1222; scan_win1224 <= scan_win1223; scan_win1225 <= scan_win1224; scan_win1226 <= scan_win1225; scan_win1227 <= scan_win1226; scan_win1228 <= scan_win1227; scan_win1229 <= scan_win1228; scan_win1230 <= scan_win1229; scan_win1231 <= scan_win1230; scan_win1232 <= scan_win1231; scan_win1233 <= scan_win1232; scan_win1234 <= scan_win1233; scan_win1235 <= scan_win1234; scan_win1236 <= scan_win1235; scan_win1237 <= scan_win1236; scan_win1238 <= scan_win1237; scan_win1239 <= scan_win1238; scan_win1240 <= scan_win1239; scan_win1241 <= scan_win1240; scan_win1242 <= scan_win1241; scan_win1243 <= scan_win1242; scan_win1244 <= scan_win1243; scan_win1245 <= scan_win1244; scan_win1246 <= scan_win1245; scan_win1247 <= scan_win1246; scan_win1248 <= scan_win1247; scan_win1249 <= scan_win1248; scan_win1250 <= scan_win1249; scan_win1251 <= scan_win1250; scan_win1252 <= scan_win1251; scan_win1253 <= scan_win1252; scan_win1254 <= scan_win1253; scan_win1255 <= scan_win1254; scan_win1256 <= scan_win1255; scan_win1257 <= scan_win1256; scan_win1258 <= scan_win1257; scan_win1259 <= scan_win1258; scan_win1260 <= scan_win1259; scan_win1261 <= scan_win1260; scan_win1262 <= scan_win1261; scan_win1263 <= scan_win1262; scan_win1264 <= scan_win1263; scan_win1265 <= scan_win1264; scan_win1266 <= scan_win1265; scan_win1267 <= scan_win1266; scan_win1268 <= scan_win1267; scan_win1269 <= scan_win1268; scan_win1270 <= scan_win1269; scan_win1271 <= scan_win1270; scan_win1272 <= scan_win1271; scan_win1273 <= scan_win1272; scan_win1274 <= scan_win1273; scan_win1275 <= scan_win1274; scan_win1276 <= scan_win1275; scan_win1277 <= scan_win1276; scan_win1278 <= scan_win1277; scan_win1279 <= scan_win1278; scan_win1280 <= scan_win1279; scan_win1281 <= scan_win1280; scan_win1282 <= scan_win1281; scan_win1283 <= scan_win1282; scan_win1284 <= scan_win1283; scan_win1285 <= scan_win1284; scan_win1286 <= scan_win1285; scan_win1287 <= scan_win1286; scan_win1288 <= scan_win1287; scan_win1289 <= scan_win1288; scan_win1290 <= scan_win1289; scan_win1291 <= scan_win1290; scan_win1292 <= scan_win1291; scan_win1293 <= scan_win1292; scan_win1294 <= scan_win1293; scan_win1295 <= scan_win1294; scan_win1296 <= scan_win1295; scan_win1297 <= scan_win1296; scan_win1298 <= scan_win1297; scan_win1299 <= scan_win1298; scan_win1300 <= scan_win1299; scan_win1301 <= scan_win1300; scan_win1302 <= scan_win1301; scan_win1303 <= scan_win1302; scan_win1304 <= scan_win1303; scan_win1305 <= scan_win1304; scan_win1306 <= scan_win1305; scan_win1307 <= scan_win1306; scan_win1308 <= scan_win1307; scan_win1309 <= scan_win1308; scan_win1310 <= scan_win1309; scan_win1311 <= scan_win1310; scan_win1312 <= scan_win1311; scan_win1313 <= scan_win1312; scan_win1314 <= scan_win1313; scan_win1315 <= scan_win1314; scan_win1316 <= scan_win1315; scan_win1317 <= scan_win1316; scan_win1318 <= scan_win1317; scan_win1319 <= scan_win1318; scan_win1320 <= scan_win1319; scan_win1321 <= scan_win1320; scan_win1322 <= scan_win1321; scan_win1323 <= scan_win1322; scan_win1324 <= scan_win1323; scan_win1325 <= scan_win1324; scan_win1326 <= scan_win1325; scan_win1327 <= scan_win1326; scan_win1328 <= scan_win1327; scan_win1329 <= scan_win1328; scan_win1330 <= scan_win1329; scan_win1331 <= scan_win1330; scan_win1332 <= scan_win1331; scan_win1333 <= scan_win1332; scan_win1334 <= scan_win1333; scan_win1335 <= scan_win1334; scan_win1336 <= scan_win1335; scan_win1337 <= scan_win1336; scan_win1338 <= scan_win1337; scan_win1339 <= scan_win1338; scan_win1340 <= scan_win1339; scan_win1341 <= scan_win1340; scan_win1342 <= scan_win1341; scan_win1343 <= scan_win1342; scan_win1344 <= scan_win1343; scan_win1345 <= scan_win1344; scan_win1346 <= scan_win1345; scan_win1347 <= scan_win1346; scan_win1348 <= scan_win1347; scan_win1349 <= scan_win1348; scan_win1350 <= scan_win1349; scan_win1351 <= scan_win1350; scan_win1352 <= scan_win1351; scan_win1353 <= scan_win1352; scan_win1354 <= scan_win1353; scan_win1355 <= scan_win1354; scan_win1356 <= scan_win1355; scan_win1357 <= scan_win1356; scan_win1358 <= scan_win1357; scan_win1359 <= scan_win1358; scan_win1360 <= scan_win1359; scan_win1361 <= scan_win1360; scan_win1362 <= scan_win1361; scan_win1363 <= scan_win1362; scan_win1364 <= scan_win1363; scan_win1365 <= scan_win1364; scan_win1366 <= scan_win1365; scan_win1367 <= scan_win1366; scan_win1368 <= scan_win1367; scan_win1369 <= scan_win1368; scan_win1370 <= scan_win1369; scan_win1371 <= scan_win1370; scan_win1372 <= scan_win1371; scan_win1373 <= scan_win1372; scan_win1374 <= scan_win1373; scan_win1375 <= scan_win1374; scan_win1376 <= scan_win1375; scan_win1377 <= scan_win1376; scan_win1378 <= scan_win1377; scan_win1379 <= scan_win1378; scan_win1380 <= scan_win1379; scan_win1381 <= scan_win1380; scan_win1382 <= scan_win1381; scan_win1383 <= scan_win1382; scan_win1384 <= scan_win1383; scan_win1385 <= scan_win1384; scan_win1386 <= scan_win1385; scan_win1387 <= scan_win1386; scan_win1388 <= scan_win1387; scan_win1389 <= scan_win1388; scan_win1390 <= scan_win1389; scan_win1391 <= scan_win1390; scan_win1392 <= scan_win1391; scan_win1393 <= scan_win1392; scan_win1394 <= scan_win1393; scan_win1395 <= scan_win1394; scan_win1396 <= scan_win1395; scan_win1397 <= scan_win1396; scan_win1398 <= scan_win1397; scan_win1399 <= scan_win1398; scan_win1400 <= scan_win1399; 
      scan_win1401 <= scan_win1400; scan_win1402 <= scan_win1401; scan_win1403 <= scan_win1402; scan_win1404 <= scan_win1403; scan_win1405 <= scan_win1404; scan_win1406 <= scan_win1405; scan_win1407 <= scan_win1406; scan_win1408 <= scan_win1407; scan_win1409 <= scan_win1408; scan_win1410 <= scan_win1409; scan_win1411 <= scan_win1410; scan_win1412 <= scan_win1411; scan_win1413 <= scan_win1412; scan_win1414 <= scan_win1413; scan_win1415 <= scan_win1414; scan_win1416 <= scan_win1415; scan_win1417 <= scan_win1416; scan_win1418 <= scan_win1417; scan_win1419 <= scan_win1418; scan_win1420 <= scan_win1419; scan_win1421 <= scan_win1420; scan_win1422 <= scan_win1421; scan_win1423 <= scan_win1422; scan_win1424 <= scan_win1423; scan_win1425 <= scan_win1424; scan_win1426 <= scan_win1425; scan_win1427 <= scan_win1426; scan_win1428 <= scan_win1427; scan_win1429 <= scan_win1428; scan_win1430 <= scan_win1429; scan_win1431 <= scan_win1430; scan_win1432 <= scan_win1431; scan_win1433 <= scan_win1432; scan_win1434 <= scan_win1433; scan_win1435 <= scan_win1434; scan_win1436 <= scan_win1435; scan_win1437 <= scan_win1436; scan_win1438 <= scan_win1437; scan_win1439 <= scan_win1438; scan_win1440 <= scan_win1439; scan_win1441 <= scan_win1440; scan_win1442 <= scan_win1441; scan_win1443 <= scan_win1442; scan_win1444 <= scan_win1443; scan_win1445 <= scan_win1444; scan_win1446 <= scan_win1445; scan_win1447 <= scan_win1446; scan_win1448 <= scan_win1447; scan_win1449 <= scan_win1448; scan_win1450 <= scan_win1449; scan_win1451 <= scan_win1450; scan_win1452 <= scan_win1451; scan_win1453 <= scan_win1452; scan_win1454 <= scan_win1453; scan_win1455 <= scan_win1454; scan_win1456 <= scan_win1455; scan_win1457 <= scan_win1456; scan_win1458 <= scan_win1457; scan_win1459 <= scan_win1458; scan_win1460 <= scan_win1459; scan_win1461 <= scan_win1460; scan_win1462 <= scan_win1461; scan_win1463 <= scan_win1462; scan_win1464 <= scan_win1463; scan_win1465 <= scan_win1464; scan_win1466 <= scan_win1465; scan_win1467 <= scan_win1466; scan_win1468 <= scan_win1467; scan_win1469 <= scan_win1468; scan_win1470 <= scan_win1469; scan_win1471 <= scan_win1470; scan_win1472 <= scan_win1471; scan_win1473 <= scan_win1472; scan_win1474 <= scan_win1473; scan_win1475 <= scan_win1474; scan_win1476 <= scan_win1475; scan_win1477 <= scan_win1476; scan_win1478 <= scan_win1477; scan_win1479 <= scan_win1478; scan_win1480 <= scan_win1479; scan_win1481 <= scan_win1480; scan_win1482 <= scan_win1481; scan_win1483 <= scan_win1482; scan_win1484 <= scan_win1483; scan_win1485 <= scan_win1484; scan_win1486 <= scan_win1485; scan_win1487 <= scan_win1486; scan_win1488 <= scan_win1487; scan_win1489 <= scan_win1488; scan_win1490 <= scan_win1489; scan_win1491 <= scan_win1490; scan_win1492 <= scan_win1491; scan_win1493 <= scan_win1492; scan_win1494 <= scan_win1493; scan_win1495 <= scan_win1494; scan_win1496 <= scan_win1495; scan_win1497 <= scan_win1496; scan_win1498 <= scan_win1497; scan_win1499 <= scan_win1498; scan_win1500 <= scan_win1499; scan_win1501 <= scan_win1500; scan_win1502 <= scan_win1501; scan_win1503 <= scan_win1502; scan_win1504 <= scan_win1503; scan_win1505 <= scan_win1504; scan_win1506 <= scan_win1505; scan_win1507 <= scan_win1506; scan_win1508 <= scan_win1507; scan_win1509 <= scan_win1508; scan_win1510 <= scan_win1509; scan_win1511 <= scan_win1510; scan_win1512 <= scan_win1511; scan_win1513 <= scan_win1512; scan_win1514 <= scan_win1513; scan_win1515 <= scan_win1514; scan_win1516 <= scan_win1515; scan_win1517 <= scan_win1516; scan_win1518 <= scan_win1517; scan_win1519 <= scan_win1518; scan_win1520 <= scan_win1519; scan_win1521 <= scan_win1520; scan_win1522 <= scan_win1521; scan_win1523 <= scan_win1522; scan_win1524 <= scan_win1523; scan_win1525 <= scan_win1524; scan_win1526 <= scan_win1525; scan_win1527 <= scan_win1526; scan_win1528 <= scan_win1527; scan_win1529 <= scan_win1528; scan_win1530 <= scan_win1529; scan_win1531 <= scan_win1530; scan_win1532 <= scan_win1531; scan_win1533 <= scan_win1532; scan_win1534 <= scan_win1533; scan_win1535 <= scan_win1534; scan_win1536 <= scan_win1535; scan_win1537 <= scan_win1536; scan_win1538 <= scan_win1537; scan_win1539 <= scan_win1538; scan_win1540 <= scan_win1539; scan_win1541 <= scan_win1540; scan_win1542 <= scan_win1541; scan_win1543 <= scan_win1542; scan_win1544 <= scan_win1543; scan_win1545 <= scan_win1544; scan_win1546 <= scan_win1545; scan_win1547 <= scan_win1546; scan_win1548 <= scan_win1547; scan_win1549 <= scan_win1548; scan_win1550 <= scan_win1549; scan_win1551 <= scan_win1550; scan_win1552 <= scan_win1551; scan_win1553 <= scan_win1552; scan_win1554 <= scan_win1553; scan_win1555 <= scan_win1554; scan_win1556 <= scan_win1555; scan_win1557 <= scan_win1556; scan_win1558 <= scan_win1557; scan_win1559 <= scan_win1558; scan_win1560 <= scan_win1559; scan_win1561 <= scan_win1560; scan_win1562 <= scan_win1561; scan_win1563 <= scan_win1562; scan_win1564 <= scan_win1563; scan_win1565 <= scan_win1564; scan_win1566 <= scan_win1565; scan_win1567 <= scan_win1566; scan_win1568 <= scan_win1567; scan_win1569 <= scan_win1568; scan_win1570 <= scan_win1569; scan_win1571 <= scan_win1570; scan_win1572 <= scan_win1571; scan_win1573 <= scan_win1572; scan_win1574 <= scan_win1573; scan_win1575 <= scan_win1574; scan_win1576 <= scan_win1575; scan_win1577 <= scan_win1576; scan_win1578 <= scan_win1577; scan_win1579 <= scan_win1578; scan_win1580 <= scan_win1579; scan_win1581 <= scan_win1580; scan_win1582 <= scan_win1581; scan_win1583 <= scan_win1582; scan_win1584 <= scan_win1583; scan_win1585 <= scan_win1584; scan_win1586 <= scan_win1585; scan_win1587 <= scan_win1586; scan_win1588 <= scan_win1587; scan_win1589 <= scan_win1588; scan_win1590 <= scan_win1589; scan_win1591 <= scan_win1590; scan_win1592 <= scan_win1591; scan_win1593 <= scan_win1592; scan_win1594 <= scan_win1593; scan_win1595 <= scan_win1594; scan_win1596 <= scan_win1595; scan_win1597 <= scan_win1596; scan_win1598 <= scan_win1597; scan_win1599 <= scan_win1598; scan_win1600 <= scan_win1599; 
      scan_win1601 <= scan_win1600; scan_win1602 <= scan_win1601; scan_win1603 <= scan_win1602; scan_win1604 <= scan_win1603; scan_win1605 <= scan_win1604; scan_win1606 <= scan_win1605; scan_win1607 <= scan_win1606; scan_win1608 <= scan_win1607; scan_win1609 <= scan_win1608; scan_win1610 <= scan_win1609; scan_win1611 <= scan_win1610; scan_win1612 <= scan_win1611; scan_win1613 <= scan_win1612; scan_win1614 <= scan_win1613; scan_win1615 <= scan_win1614; scan_win1616 <= scan_win1615; scan_win1617 <= scan_win1616; scan_win1618 <= scan_win1617; scan_win1619 <= scan_win1618; scan_win1620 <= scan_win1619; scan_win1621 <= scan_win1620; scan_win1622 <= scan_win1621; scan_win1623 <= scan_win1622; scan_win1624 <= scan_win1623; scan_win1625 <= scan_win1624; scan_win1626 <= scan_win1625; scan_win1627 <= scan_win1626; scan_win1628 <= scan_win1627; scan_win1629 <= scan_win1628; scan_win1630 <= scan_win1629; scan_win1631 <= scan_win1630; scan_win1632 <= scan_win1631; scan_win1633 <= scan_win1632; scan_win1634 <= scan_win1633; scan_win1635 <= scan_win1634; scan_win1636 <= scan_win1635; scan_win1637 <= scan_win1636; scan_win1638 <= scan_win1637; scan_win1639 <= scan_win1638; scan_win1640 <= scan_win1639; scan_win1641 <= scan_win1640; scan_win1642 <= scan_win1641; scan_win1643 <= scan_win1642; scan_win1644 <= scan_win1643; scan_win1645 <= scan_win1644; scan_win1646 <= scan_win1645; scan_win1647 <= scan_win1646; scan_win1648 <= scan_win1647; scan_win1649 <= scan_win1648; scan_win1650 <= scan_win1649; scan_win1651 <= scan_win1650; scan_win1652 <= scan_win1651; scan_win1653 <= scan_win1652; scan_win1654 <= scan_win1653; scan_win1655 <= scan_win1654; scan_win1656 <= scan_win1655; scan_win1657 <= scan_win1656; scan_win1658 <= scan_win1657; scan_win1659 <= scan_win1658; scan_win1660 <= scan_win1659; scan_win1661 <= scan_win1660; scan_win1662 <= scan_win1661; scan_win1663 <= scan_win1662; scan_win1664 <= scan_win1663; scan_win1665 <= scan_win1664; scan_win1666 <= scan_win1665; scan_win1667 <= scan_win1666; scan_win1668 <= scan_win1667; scan_win1669 <= scan_win1668; scan_win1670 <= scan_win1669; scan_win1671 <= scan_win1670; scan_win1672 <= scan_win1671; scan_win1673 <= scan_win1672; scan_win1674 <= scan_win1673; scan_win1675 <= scan_win1674; scan_win1676 <= scan_win1675; scan_win1677 <= scan_win1676; scan_win1678 <= scan_win1677; scan_win1679 <= scan_win1678; scan_win1680 <= scan_win1679; scan_win1681 <= scan_win1680; scan_win1682 <= scan_win1681; scan_win1683 <= scan_win1682; scan_win1684 <= scan_win1683; scan_win1685 <= scan_win1684; scan_win1686 <= scan_win1685; scan_win1687 <= scan_win1686; scan_win1688 <= scan_win1687; scan_win1689 <= scan_win1688; scan_win1690 <= scan_win1689; scan_win1691 <= scan_win1690; scan_win1692 <= scan_win1691; scan_win1693 <= scan_win1692; scan_win1694 <= scan_win1693; scan_win1695 <= scan_win1694; scan_win1696 <= scan_win1695; scan_win1697 <= scan_win1696; scan_win1698 <= scan_win1697; scan_win1699 <= scan_win1698; scan_win1700 <= scan_win1699; scan_win1701 <= scan_win1700; scan_win1702 <= scan_win1701; scan_win1703 <= scan_win1702; scan_win1704 <= scan_win1703; scan_win1705 <= scan_win1704; scan_win1706 <= scan_win1705; scan_win1707 <= scan_win1706; scan_win1708 <= scan_win1707; scan_win1709 <= scan_win1708; scan_win1710 <= scan_win1709; scan_win1711 <= scan_win1710; scan_win1712 <= scan_win1711; scan_win1713 <= scan_win1712; scan_win1714 <= scan_win1713; scan_win1715 <= scan_win1714; scan_win1716 <= scan_win1715; scan_win1717 <= scan_win1716; scan_win1718 <= scan_win1717; scan_win1719 <= scan_win1718; scan_win1720 <= scan_win1719; scan_win1721 <= scan_win1720; scan_win1722 <= scan_win1721; scan_win1723 <= scan_win1722; scan_win1724 <= scan_win1723; scan_win1725 <= scan_win1724; scan_win1726 <= scan_win1725; scan_win1727 <= scan_win1726; scan_win1728 <= scan_win1727; scan_win1729 <= scan_win1728; scan_win1730 <= scan_win1729; scan_win1731 <= scan_win1730; scan_win1732 <= scan_win1731; scan_win1733 <= scan_win1732; scan_win1734 <= scan_win1733; scan_win1735 <= scan_win1734; scan_win1736 <= scan_win1735; scan_win1737 <= scan_win1736; scan_win1738 <= scan_win1737; scan_win1739 <= scan_win1738; scan_win1740 <= scan_win1739; scan_win1741 <= scan_win1740; scan_win1742 <= scan_win1741; scan_win1743 <= scan_win1742; scan_win1744 <= scan_win1743; scan_win1745 <= scan_win1744; scan_win1746 <= scan_win1745; scan_win1747 <= scan_win1746; scan_win1748 <= scan_win1747; scan_win1749 <= scan_win1748; scan_win1750 <= scan_win1749; scan_win1751 <= scan_win1750; scan_win1752 <= scan_win1751; scan_win1753 <= scan_win1752; scan_win1754 <= scan_win1753; scan_win1755 <= scan_win1754; scan_win1756 <= scan_win1755; scan_win1757 <= scan_win1756; scan_win1758 <= scan_win1757; scan_win1759 <= scan_win1758; scan_win1760 <= scan_win1759; scan_win1761 <= scan_win1760; scan_win1762 <= scan_win1761; scan_win1763 <= scan_win1762; scan_win1764 <= scan_win1763; scan_win1765 <= scan_win1764; scan_win1766 <= scan_win1765; scan_win1767 <= scan_win1766; scan_win1768 <= scan_win1767; scan_win1769 <= scan_win1768; scan_win1770 <= scan_win1769; scan_win1771 <= scan_win1770; scan_win1772 <= scan_win1771; scan_win1773 <= scan_win1772; scan_win1774 <= scan_win1773; scan_win1775 <= scan_win1774; scan_win1776 <= scan_win1775; scan_win1777 <= scan_win1776; scan_win1778 <= scan_win1777; scan_win1779 <= scan_win1778; scan_win1780 <= scan_win1779; scan_win1781 <= scan_win1780; scan_win1782 <= scan_win1781; scan_win1783 <= scan_win1782; scan_win1784 <= scan_win1783; scan_win1785 <= scan_win1784; scan_win1786 <= scan_win1785; scan_win1787 <= scan_win1786; scan_win1788 <= scan_win1787; scan_win1789 <= scan_win1788; scan_win1790 <= scan_win1789; scan_win1791 <= scan_win1790; scan_win1792 <= scan_win1791; scan_win1793 <= scan_win1792; scan_win1794 <= scan_win1793; scan_win1795 <= scan_win1794; scan_win1796 <= scan_win1795; scan_win1797 <= scan_win1796; scan_win1798 <= scan_win1797; scan_win1799 <= scan_win1798; scan_win1800 <= scan_win1799; 
      scan_win1801 <= scan_win1800; scan_win1802 <= scan_win1801; scan_win1803 <= scan_win1802; scan_win1804 <= scan_win1803; scan_win1805 <= scan_win1804; scan_win1806 <= scan_win1805; scan_win1807 <= scan_win1806; scan_win1808 <= scan_win1807; scan_win1809 <= scan_win1808; scan_win1810 <= scan_win1809; scan_win1811 <= scan_win1810; scan_win1812 <= scan_win1811; scan_win1813 <= scan_win1812; scan_win1814 <= scan_win1813; scan_win1815 <= scan_win1814; scan_win1816 <= scan_win1815; scan_win1817 <= scan_win1816; scan_win1818 <= scan_win1817; scan_win1819 <= scan_win1818; scan_win1820 <= scan_win1819; scan_win1821 <= scan_win1820; scan_win1822 <= scan_win1821; scan_win1823 <= scan_win1822; scan_win1824 <= scan_win1823; scan_win1825 <= scan_win1824; scan_win1826 <= scan_win1825; scan_win1827 <= scan_win1826; scan_win1828 <= scan_win1827; scan_win1829 <= scan_win1828; scan_win1830 <= scan_win1829; scan_win1831 <= scan_win1830; scan_win1832 <= scan_win1831; scan_win1833 <= scan_win1832; scan_win1834 <= scan_win1833; scan_win1835 <= scan_win1834; scan_win1836 <= scan_win1835; scan_win1837 <= scan_win1836; scan_win1838 <= scan_win1837; scan_win1839 <= scan_win1838; scan_win1840 <= scan_win1839; scan_win1841 <= scan_win1840; scan_win1842 <= scan_win1841; scan_win1843 <= scan_win1842; scan_win1844 <= scan_win1843; scan_win1845 <= scan_win1844; scan_win1846 <= scan_win1845; scan_win1847 <= scan_win1846; scan_win1848 <= scan_win1847; scan_win1849 <= scan_win1848; scan_win1850 <= scan_win1849; scan_win1851 <= scan_win1850; scan_win1852 <= scan_win1851; scan_win1853 <= scan_win1852; scan_win1854 <= scan_win1853; scan_win1855 <= scan_win1854; scan_win1856 <= scan_win1855; scan_win1857 <= scan_win1856; scan_win1858 <= scan_win1857; scan_win1859 <= scan_win1858; scan_win1860 <= scan_win1859; scan_win1861 <= scan_win1860; scan_win1862 <= scan_win1861; scan_win1863 <= scan_win1862; scan_win1864 <= scan_win1863; scan_win1865 <= scan_win1864; scan_win1866 <= scan_win1865; scan_win1867 <= scan_win1866; scan_win1868 <= scan_win1867; scan_win1869 <= scan_win1868; scan_win1870 <= scan_win1869; scan_win1871 <= scan_win1870; scan_win1872 <= scan_win1871; scan_win1873 <= scan_win1872; scan_win1874 <= scan_win1873; scan_win1875 <= scan_win1874; scan_win1876 <= scan_win1875; scan_win1877 <= scan_win1876; scan_win1878 <= scan_win1877; scan_win1879 <= scan_win1878; scan_win1880 <= scan_win1879; scan_win1881 <= scan_win1880; scan_win1882 <= scan_win1881; scan_win1883 <= scan_win1882; scan_win1884 <= scan_win1883; scan_win1885 <= scan_win1884; scan_win1886 <= scan_win1885; scan_win1887 <= scan_win1886; scan_win1888 <= scan_win1887; scan_win1889 <= scan_win1888; scan_win1890 <= scan_win1889; scan_win1891 <= scan_win1890; scan_win1892 <= scan_win1891; scan_win1893 <= scan_win1892; scan_win1894 <= scan_win1893; scan_win1895 <= scan_win1894; scan_win1896 <= scan_win1895; scan_win1897 <= scan_win1896; scan_win1898 <= scan_win1897; scan_win1899 <= scan_win1898; scan_win1900 <= scan_win1899; scan_win1901 <= scan_win1900; scan_win1902 <= scan_win1901; scan_win1903 <= scan_win1902; scan_win1904 <= scan_win1903; scan_win1905 <= scan_win1904; scan_win1906 <= scan_win1905; scan_win1907 <= scan_win1906; scan_win1908 <= scan_win1907; scan_win1909 <= scan_win1908; scan_win1910 <= scan_win1909; scan_win1911 <= scan_win1910; scan_win1912 <= scan_win1911; scan_win1913 <= scan_win1912; scan_win1914 <= scan_win1913; scan_win1915 <= scan_win1914; scan_win1916 <= scan_win1915; scan_win1917 <= scan_win1916; scan_win1918 <= scan_win1917; scan_win1919 <= scan_win1918; scan_win1920 <= scan_win1919; scan_win1921 <= scan_win1920; scan_win1922 <= scan_win1921; scan_win1923 <= scan_win1922; scan_win1924 <= scan_win1923; scan_win1925 <= scan_win1924; scan_win1926 <= scan_win1925; scan_win1927 <= scan_win1926; scan_win1928 <= scan_win1927; scan_win1929 <= scan_win1928; scan_win1930 <= scan_win1929; scan_win1931 <= scan_win1930; scan_win1932 <= scan_win1931; scan_win1933 <= scan_win1932; scan_win1934 <= scan_win1933; scan_win1935 <= scan_win1934; scan_win1936 <= scan_win1935; scan_win1937 <= scan_win1936; scan_win1938 <= scan_win1937; scan_win1939 <= scan_win1938; scan_win1940 <= scan_win1939; scan_win1941 <= scan_win1940; scan_win1942 <= scan_win1941; scan_win1943 <= scan_win1942; scan_win1944 <= scan_win1943; scan_win1945 <= scan_win1944; scan_win1946 <= scan_win1945; scan_win1947 <= scan_win1946; scan_win1948 <= scan_win1947; scan_win1949 <= scan_win1948; scan_win1950 <= scan_win1949; scan_win1951 <= scan_win1950; scan_win1952 <= scan_win1951; scan_win1953 <= scan_win1952; scan_win1954 <= scan_win1953; scan_win1955 <= scan_win1954; scan_win1956 <= scan_win1955; scan_win1957 <= scan_win1956; scan_win1958 <= scan_win1957; scan_win1959 <= scan_win1958; scan_win1960 <= scan_win1959; scan_win1961 <= scan_win1960; scan_win1962 <= scan_win1961; scan_win1963 <= scan_win1962; scan_win1964 <= scan_win1963; scan_win1965 <= scan_win1964; scan_win1966 <= scan_win1965; scan_win1967 <= scan_win1966; scan_win1968 <= scan_win1967; scan_win1969 <= scan_win1968; scan_win1970 <= scan_win1969; scan_win1971 <= scan_win1970; scan_win1972 <= scan_win1971; scan_win1973 <= scan_win1972; scan_win1974 <= scan_win1973; scan_win1975 <= scan_win1974; scan_win1976 <= scan_win1975; scan_win1977 <= scan_win1976; scan_win1978 <= scan_win1977; scan_win1979 <= scan_win1978; scan_win1980 <= scan_win1979; scan_win1981 <= scan_win1980; scan_win1982 <= scan_win1981; scan_win1983 <= scan_win1982; scan_win1984 <= scan_win1983; scan_win1985 <= scan_win1984; scan_win1986 <= scan_win1985; scan_win1987 <= scan_win1986; scan_win1988 <= scan_win1987; scan_win1989 <= scan_win1988; scan_win1990 <= scan_win1989; scan_win1991 <= scan_win1990; scan_win1992 <= scan_win1991; scan_win1993 <= scan_win1992; scan_win1994 <= scan_win1993; scan_win1995 <= scan_win1994; scan_win1996 <= scan_win1995; scan_win1997 <= scan_win1996; scan_win1998 <= scan_win1997; scan_win1999 <= scan_win1998; scan_win2000 <= scan_win1999; 
      scan_win2001 <= scan_win2000; scan_win2002 <= scan_win2001; scan_win2003 <= scan_win2002; scan_win2004 <= scan_win2003; scan_win2005 <= scan_win2004; scan_win2006 <= scan_win2005; scan_win2007 <= scan_win2006; scan_win2008 <= scan_win2007; scan_win2009 <= scan_win2008; scan_win2010 <= scan_win2009; scan_win2011 <= scan_win2010; scan_win2012 <= scan_win2011; scan_win2013 <= scan_win2012; scan_win2014 <= scan_win2013; scan_win2015 <= scan_win2014; scan_win2016 <= scan_win2015; scan_win2017 <= scan_win2016; scan_win2018 <= scan_win2017; scan_win2019 <= scan_win2018; scan_win2020 <= scan_win2019; scan_win2021 <= scan_win2020; scan_win2022 <= scan_win2021; scan_win2023 <= scan_win2022; scan_win2024 <= scan_win2023; scan_win2025 <= scan_win2024; scan_win2026 <= scan_win2025; scan_win2027 <= scan_win2026; scan_win2028 <= scan_win2027; scan_win2029 <= scan_win2028; scan_win2030 <= scan_win2029; scan_win2031 <= scan_win2030; scan_win2032 <= scan_win2031; scan_win2033 <= scan_win2032; scan_win2034 <= scan_win2033; scan_win2035 <= scan_win2034; scan_win2036 <= scan_win2035; scan_win2037 <= scan_win2036; scan_win2038 <= scan_win2037; scan_win2039 <= scan_win2038; scan_win2040 <= scan_win2039; scan_win2041 <= scan_win2040; scan_win2042 <= scan_win2041; scan_win2043 <= scan_win2042; scan_win2044 <= scan_win2043; scan_win2045 <= scan_win2044; scan_win2046 <= scan_win2045; scan_win2047 <= scan_win2046; scan_win2048 <= scan_win2047; scan_win2049 <= scan_win2048; scan_win2050 <= scan_win2049; scan_win2051 <= scan_win2050; scan_win2052 <= scan_win2051; scan_win2053 <= scan_win2052; scan_win2054 <= scan_win2053; scan_win2055 <= scan_win2054; scan_win2056 <= scan_win2055; scan_win2057 <= scan_win2056; scan_win2058 <= scan_win2057; scan_win2059 <= scan_win2058; scan_win2060 <= scan_win2059; scan_win2061 <= scan_win2060; scan_win2062 <= scan_win2061; scan_win2063 <= scan_win2062; scan_win2064 <= scan_win2063; scan_win2065 <= scan_win2064; scan_win2066 <= scan_win2065; scan_win2067 <= scan_win2066; scan_win2068 <= scan_win2067; scan_win2069 <= scan_win2068; scan_win2070 <= scan_win2069; scan_win2071 <= scan_win2070; scan_win2072 <= scan_win2071; scan_win2073 <= scan_win2072; scan_win2074 <= scan_win2073; scan_win2075 <= scan_win2074; scan_win2076 <= scan_win2075; scan_win2077 <= scan_win2076; scan_win2078 <= scan_win2077; scan_win2079 <= scan_win2078; scan_win2080 <= scan_win2079; scan_win2081 <= scan_win2080; scan_win2082 <= scan_win2081; scan_win2083 <= scan_win2082; scan_win2084 <= scan_win2083; scan_win2085 <= scan_win2084; scan_win2086 <= scan_win2085; scan_win2087 <= scan_win2086; scan_win2088 <= scan_win2087; scan_win2089 <= scan_win2088; scan_win2090 <= scan_win2089; scan_win2091 <= scan_win2090; scan_win2092 <= scan_win2091; scan_win2093 <= scan_win2092; scan_win2094 <= scan_win2093; scan_win2095 <= scan_win2094; scan_win2096 <= scan_win2095; scan_win2097 <= scan_win2096; scan_win2098 <= scan_win2097; scan_win2099 <= scan_win2098; scan_win2100 <= scan_win2099; scan_win2101 <= scan_win2100; scan_win2102 <= scan_win2101; scan_win2103 <= scan_win2102; scan_win2104 <= scan_win2103; scan_win2105 <= scan_win2104; scan_win2106 <= scan_win2105; scan_win2107 <= scan_win2106; scan_win2108 <= scan_win2107; scan_win2109 <= scan_win2108; scan_win2110 <= scan_win2109; scan_win2111 <= scan_win2110; scan_win2112 <= scan_win2111; scan_win2113 <= scan_win2112; scan_win2114 <= scan_win2113; scan_win2115 <= scan_win2114; scan_win2116 <= scan_win2115; scan_win2117 <= scan_win2116; scan_win2118 <= scan_win2117; scan_win2119 <= scan_win2118; scan_win2120 <= scan_win2119; scan_win2121 <= scan_win2120; scan_win2122 <= scan_win2121; scan_win2123 <= scan_win2122; scan_win2124 <= scan_win2123; scan_win2125 <= scan_win2124; scan_win2126 <= scan_win2125; scan_win2127 <= scan_win2126; scan_win2128 <= scan_win2127; scan_win2129 <= scan_win2128; scan_win2130 <= scan_win2129; scan_win2131 <= scan_win2130; scan_win2132 <= scan_win2131; scan_win2133 <= scan_win2132; scan_win2134 <= scan_win2133; scan_win2135 <= scan_win2134; scan_win2136 <= scan_win2135; scan_win2137 <= scan_win2136; scan_win2138 <= scan_win2137; scan_win2139 <= scan_win2138; scan_win2140 <= scan_win2139; scan_win2141 <= scan_win2140; scan_win2142 <= scan_win2141; scan_win2143 <= scan_win2142; scan_win2144 <= scan_win2143; scan_win2145 <= scan_win2144; scan_win2146 <= scan_win2145; scan_win2147 <= scan_win2146; scan_win2148 <= scan_win2147; scan_win2149 <= scan_win2148; scan_win2150 <= scan_win2149; scan_win2151 <= scan_win2150; scan_win2152 <= scan_win2151; scan_win2153 <= scan_win2152; scan_win2154 <= scan_win2153; scan_win2155 <= scan_win2154; scan_win2156 <= scan_win2155; scan_win2157 <= scan_win2156; scan_win2158 <= scan_win2157; scan_win2159 <= scan_win2158; scan_win2160 <= scan_win2159; scan_win2161 <= scan_win2160; scan_win2162 <= scan_win2161; scan_win2163 <= scan_win2162; scan_win2164 <= scan_win2163; scan_win2165 <= scan_win2164; scan_win2166 <= scan_win2165; scan_win2167 <= scan_win2166; scan_win2168 <= scan_win2167; scan_win2169 <= scan_win2168; scan_win2170 <= scan_win2169; scan_win2171 <= scan_win2170; scan_win2172 <= scan_win2171; scan_win2173 <= scan_win2172; scan_win2174 <= scan_win2173; scan_win2175 <= scan_win2174; scan_win2176 <= scan_win2175; scan_win2177 <= scan_win2176; scan_win2178 <= scan_win2177; scan_win2179 <= scan_win2178; scan_win2180 <= scan_win2179; scan_win2181 <= scan_win2180; scan_win2182 <= scan_win2181; scan_win2183 <= scan_win2182; scan_win2184 <= scan_win2183; scan_win2185 <= scan_win2184; scan_win2186 <= scan_win2185; scan_win2187 <= scan_win2186; scan_win2188 <= scan_win2187; scan_win2189 <= scan_win2188; scan_win2190 <= scan_win2189; scan_win2191 <= scan_win2190; scan_win2192 <= scan_win2191; scan_win2193 <= scan_win2192; scan_win2194 <= scan_win2193; scan_win2195 <= scan_win2194; scan_win2196 <= scan_win2195; scan_win2197 <= scan_win2196; scan_win2198 <= scan_win2197; scan_win2199 <= scan_win2198; scan_win2200 <= scan_win2199; 
      scan_win2201 <= scan_win2200; scan_win2202 <= scan_win2201; scan_win2203 <= scan_win2202; scan_win2204 <= scan_win2203; scan_win2205 <= scan_win2204; scan_win2206 <= scan_win2205; scan_win2207 <= scan_win2206; scan_win2208 <= scan_win2207; scan_win2209 <= scan_win2208; scan_win2210 <= scan_win2209; scan_win2211 <= scan_win2210; scan_win2212 <= scan_win2211; scan_win2213 <= scan_win2212; scan_win2214 <= scan_win2213; scan_win2215 <= scan_win2214; scan_win2216 <= scan_win2215; scan_win2217 <= scan_win2216; scan_win2218 <= scan_win2217; scan_win2219 <= scan_win2218; scan_win2220 <= scan_win2219; scan_win2221 <= scan_win2220; scan_win2222 <= scan_win2221; scan_win2223 <= scan_win2222; scan_win2224 <= scan_win2223; scan_win2225 <= scan_win2224; scan_win2226 <= scan_win2225; scan_win2227 <= scan_win2226; scan_win2228 <= scan_win2227; scan_win2229 <= scan_win2228; scan_win2230 <= scan_win2229; scan_win2231 <= scan_win2230; scan_win2232 <= scan_win2231; scan_win2233 <= scan_win2232; scan_win2234 <= scan_win2233; scan_win2235 <= scan_win2234; scan_win2236 <= scan_win2235; scan_win2237 <= scan_win2236; scan_win2238 <= scan_win2237; scan_win2239 <= scan_win2238; scan_win2240 <= scan_win2239; scan_win2241 <= scan_win2240; scan_win2242 <= scan_win2241; scan_win2243 <= scan_win2242; scan_win2244 <= scan_win2243; scan_win2245 <= scan_win2244; scan_win2246 <= scan_win2245; scan_win2247 <= scan_win2246; scan_win2248 <= scan_win2247; scan_win2249 <= scan_win2248; scan_win2250 <= scan_win2249; scan_win2251 <= scan_win2250; scan_win2252 <= scan_win2251; scan_win2253 <= scan_win2252; scan_win2254 <= scan_win2253; scan_win2255 <= scan_win2254; scan_win2256 <= scan_win2255; scan_win2257 <= scan_win2256; scan_win2258 <= scan_win2257; scan_win2259 <= scan_win2258; scan_win2260 <= scan_win2259; scan_win2261 <= scan_win2260; scan_win2262 <= scan_win2261; scan_win2263 <= scan_win2262; scan_win2264 <= scan_win2263; scan_win2265 <= scan_win2264; scan_win2266 <= scan_win2265; scan_win2267 <= scan_win2266; scan_win2268 <= scan_win2267; scan_win2269 <= scan_win2268; scan_win2270 <= scan_win2269; scan_win2271 <= scan_win2270; scan_win2272 <= scan_win2271; scan_win2273 <= scan_win2272; scan_win2274 <= scan_win2273; scan_win2275 <= scan_win2274; scan_win2276 <= scan_win2275; scan_win2277 <= scan_win2276; scan_win2278 <= scan_win2277; scan_win2279 <= scan_win2278; scan_win2280 <= scan_win2279; scan_win2281 <= scan_win2280; scan_win2282 <= scan_win2281; scan_win2283 <= scan_win2282; scan_win2284 <= scan_win2283; scan_win2285 <= scan_win2284; scan_win2286 <= scan_win2285; scan_win2287 <= scan_win2286; scan_win2288 <= scan_win2287; scan_win2289 <= scan_win2288; scan_win2290 <= scan_win2289; scan_win2291 <= scan_win2290; scan_win2292 <= scan_win2291; scan_win2293 <= scan_win2292; scan_win2294 <= scan_win2293; scan_win2295 <= scan_win2294; scan_win2296 <= scan_win2295; scan_win2297 <= scan_win2296; scan_win2298 <= scan_win2297; scan_win2299 <= scan_win2298; scan_win2300 <= scan_win2299; scan_win2301 <= scan_win2300; scan_win2302 <= scan_win2301; scan_win2303 <= scan_win2302; scan_win2304 <= scan_win2303; scan_win2305 <= scan_win2304; scan_win2306 <= scan_win2305; scan_win2307 <= scan_win2306; scan_win2308 <= scan_win2307; scan_win2309 <= scan_win2308; scan_win2310 <= scan_win2309; scan_win2311 <= scan_win2310; scan_win2312 <= scan_win2311; scan_win2313 <= scan_win2312; scan_win2314 <= scan_win2313; scan_win2315 <= scan_win2314; scan_win2316 <= scan_win2315; scan_win2317 <= scan_win2316; scan_win2318 <= scan_win2317; scan_win2319 <= scan_win2318; scan_win2320 <= scan_win2319; scan_win2321 <= scan_win2320; scan_win2322 <= scan_win2321; scan_win2323 <= scan_win2322; scan_win2324 <= scan_win2323; scan_win2325 <= scan_win2324; scan_win2326 <= scan_win2325; scan_win2327 <= scan_win2326; scan_win2328 <= scan_win2327; scan_win2329 <= scan_win2328; scan_win2330 <= scan_win2329; scan_win2331 <= scan_win2330; scan_win2332 <= scan_win2331; scan_win2333 <= scan_win2332; scan_win2334 <= scan_win2333; scan_win2335 <= scan_win2334; scan_win2336 <= scan_win2335; scan_win2337 <= scan_win2336; scan_win2338 <= scan_win2337; scan_win2339 <= scan_win2338; scan_win2340 <= scan_win2339; scan_win2341 <= scan_win2340; scan_win2342 <= scan_win2341; scan_win2343 <= scan_win2342; scan_win2344 <= scan_win2343; scan_win2345 <= scan_win2344; scan_win2346 <= scan_win2345; scan_win2347 <= scan_win2346; scan_win2348 <= scan_win2347; scan_win2349 <= scan_win2348; scan_win2350 <= scan_win2349; scan_win2351 <= scan_win2350; scan_win2352 <= scan_win2351; scan_win2353 <= scan_win2352; scan_win2354 <= scan_win2353; scan_win2355 <= scan_win2354; scan_win2356 <= scan_win2355; scan_win2357 <= scan_win2356; scan_win2358 <= scan_win2357; scan_win2359 <= scan_win2358; scan_win2360 <= scan_win2359; scan_win2361 <= scan_win2360; scan_win2362 <= scan_win2361; scan_win2363 <= scan_win2362; scan_win2364 <= scan_win2363; scan_win2365 <= scan_win2364; scan_win2366 <= scan_win2365; scan_win2367 <= scan_win2366; scan_win2368 <= scan_win2367; scan_win2369 <= scan_win2368; scan_win2370 <= scan_win2369; scan_win2371 <= scan_win2370; scan_win2372 <= scan_win2371; scan_win2373 <= scan_win2372; scan_win2374 <= scan_win2373; scan_win2375 <= scan_win2374; scan_win2376 <= scan_win2375; scan_win2377 <= scan_win2376; scan_win2378 <= scan_win2377; scan_win2379 <= scan_win2378; scan_win2380 <= scan_win2379; scan_win2381 <= scan_win2380; scan_win2382 <= scan_win2381; scan_win2383 <= scan_win2382; scan_win2384 <= scan_win2383; scan_win2385 <= scan_win2384; scan_win2386 <= scan_win2385; scan_win2387 <= scan_win2386; scan_win2388 <= scan_win2387; scan_win2389 <= scan_win2388; scan_win2390 <= scan_win2389; scan_win2391 <= scan_win2390; scan_win2392 <= scan_win2391; scan_win2393 <= scan_win2392; scan_win2394 <= scan_win2393; scan_win2395 <= scan_win2394; scan_win2396 <= scan_win2395; scan_win2397 <= scan_win2396; scan_win2398 <= scan_win2397; scan_win2399 <= scan_win2398; scan_win2400 <= scan_win2399; 
      scan_win2401 <= scan_win2400; scan_win2402 <= scan_win2401; scan_win2403 <= scan_win2402; scan_win2404 <= scan_win2403; scan_win2405 <= scan_win2404; scan_win2406 <= scan_win2405; scan_win2407 <= scan_win2406; scan_win2408 <= scan_win2407; scan_win2409 <= scan_win2408; scan_win2410 <= scan_win2409; scan_win2411 <= scan_win2410; scan_win2412 <= scan_win2411; scan_win2413 <= scan_win2412; scan_win2414 <= scan_win2413; scan_win2415 <= scan_win2414; scan_win2416 <= scan_win2415; scan_win2417 <= scan_win2416; scan_win2418 <= scan_win2417; scan_win2419 <= scan_win2418; scan_win2420 <= scan_win2419; scan_win2421 <= scan_win2420; scan_win2422 <= scan_win2421; scan_win2423 <= scan_win2422; scan_win2424 <= scan_win2423; scan_win2425 <= scan_win2424; scan_win2426 <= scan_win2425; scan_win2427 <= scan_win2426; scan_win2428 <= scan_win2427; scan_win2429 <= scan_win2428; scan_win2430 <= scan_win2429; scan_win2431 <= scan_win2430; scan_win2432 <= scan_win2431; scan_win2433 <= scan_win2432; scan_win2434 <= scan_win2433; scan_win2435 <= scan_win2434; scan_win2436 <= scan_win2435; scan_win2437 <= scan_win2436; scan_win2438 <= scan_win2437; scan_win2439 <= scan_win2438; scan_win2440 <= scan_win2439; scan_win2441 <= scan_win2440; scan_win2442 <= scan_win2441; scan_win2443 <= scan_win2442; scan_win2444 <= scan_win2443; scan_win2445 <= scan_win2444; scan_win2446 <= scan_win2445; scan_win2447 <= scan_win2446; scan_win2448 <= scan_win2447; scan_win2449 <= scan_win2448; scan_win2450 <= scan_win2449; scan_win2451 <= scan_win2450; scan_win2452 <= scan_win2451; scan_win2453 <= scan_win2452; scan_win2454 <= scan_win2453; scan_win2455 <= scan_win2454; scan_win2456 <= scan_win2455; scan_win2457 <= scan_win2456; scan_win2458 <= scan_win2457; scan_win2459 <= scan_win2458; scan_win2460 <= scan_win2459; scan_win2461 <= scan_win2460; scan_win2462 <= scan_win2461; scan_win2463 <= scan_win2462; scan_win2464 <= scan_win2463; scan_win2465 <= scan_win2464; scan_win2466 <= scan_win2465; scan_win2467 <= scan_win2466; scan_win2468 <= scan_win2467; scan_win2469 <= scan_win2468; scan_win2470 <= scan_win2469; scan_win2471 <= scan_win2470; scan_win2472 <= scan_win2471; scan_win2473 <= scan_win2472; scan_win2474 <= scan_win2473; scan_win2475 <= scan_win2474; scan_win2476 <= scan_win2475; scan_win2477 <= scan_win2476; scan_win2478 <= scan_win2477; scan_win2479 <= scan_win2478; scan_win2480 <= scan_win2479; scan_win2481 <= scan_win2480; scan_win2482 <= scan_win2481; scan_win2483 <= scan_win2482; scan_win2484 <= scan_win2483; scan_win2485 <= scan_win2484; scan_win2486 <= scan_win2485; scan_win2487 <= scan_win2486; scan_win2488 <= scan_win2487; scan_win2489 <= scan_win2488; scan_win2490 <= scan_win2489; scan_win2491 <= scan_win2490; scan_win2492 <= scan_win2491; scan_win2493 <= scan_win2492; scan_win2494 <= scan_win2493; scan_win2495 <= scan_win2494; scan_win2496 <= scan_win2495; scan_win2497 <= scan_win2496; scan_win2498 <= scan_win2497; scan_win2499 <= scan_win2498; scan_win2500 <= scan_win2499; scan_win2501 <= scan_win2500; scan_win2502 <= scan_win2501; scan_win2503 <= scan_win2502; scan_win2504 <= scan_win2503; scan_win2505 <= scan_win2504; scan_win2506 <= scan_win2505; scan_win2507 <= scan_win2506; scan_win2508 <= scan_win2507; scan_win2509 <= scan_win2508; scan_win2510 <= scan_win2509; scan_win2511 <= scan_win2510; scan_win2512 <= scan_win2511; scan_win2513 <= scan_win2512; scan_win2514 <= scan_win2513; scan_win2515 <= scan_win2514; scan_win2516 <= scan_win2515; scan_win2517 <= scan_win2516; scan_win2518 <= scan_win2517; scan_win2519 <= scan_win2518; scan_win2520 <= scan_win2519; scan_win2521 <= scan_win2520; scan_win2522 <= scan_win2521; scan_win2523 <= scan_win2522; scan_win2524 <= scan_win2523; scan_win2525 <= scan_win2524; scan_win2526 <= scan_win2525; scan_win2527 <= scan_win2526; scan_win2528 <= scan_win2527; scan_win2529 <= scan_win2528; scan_win2530 <= scan_win2529; scan_win2531 <= scan_win2530; scan_win2532 <= scan_win2531; scan_win2533 <= scan_win2532; scan_win2534 <= scan_win2533; scan_win2535 <= scan_win2534; scan_win2536 <= scan_win2535; scan_win2537 <= scan_win2536; scan_win2538 <= scan_win2537; scan_win2539 <= scan_win2538; scan_win2540 <= scan_win2539; scan_win2541 <= scan_win2540; scan_win2542 <= scan_win2541; scan_win2543 <= scan_win2542; scan_win2544 <= scan_win2543; scan_win2545 <= scan_win2544; scan_win2546 <= scan_win2545; scan_win2547 <= scan_win2546; scan_win2548 <= scan_win2547; scan_win2549 <= scan_win2548; scan_win2550 <= scan_win2549; scan_win2551 <= scan_win2550; scan_win2552 <= scan_win2551; scan_win2553 <= scan_win2552; scan_win2554 <= scan_win2553; scan_win2555 <= scan_win2554; scan_win2556 <= scan_win2555; scan_win2557 <= scan_win2556; scan_win2558 <= scan_win2557; scan_win2559 <= scan_win2558; scan_win2560 <= scan_win2559; scan_win2561 <= scan_win2560; scan_win2562 <= scan_win2561; scan_win2563 <= scan_win2562; scan_win2564 <= scan_win2563; scan_win2565 <= scan_win2564; scan_win2566 <= scan_win2565; scan_win2567 <= scan_win2566; scan_win2568 <= scan_win2567; scan_win2569 <= scan_win2568; scan_win2570 <= scan_win2569; scan_win2571 <= scan_win2570; scan_win2572 <= scan_win2571; scan_win2573 <= scan_win2572; scan_win2574 <= scan_win2573; scan_win2575 <= scan_win2574; scan_win2576 <= scan_win2575; scan_win2577 <= scan_win2576; scan_win2578 <= scan_win2577; scan_win2579 <= scan_win2578; scan_win2580 <= scan_win2579; scan_win2581 <= scan_win2580; scan_win2582 <= scan_win2581; scan_win2583 <= scan_win2582; scan_win2584 <= scan_win2583; scan_win2585 <= scan_win2584; scan_win2586 <= scan_win2585; scan_win2587 <= scan_win2586; scan_win2588 <= scan_win2587; scan_win2589 <= scan_win2588; scan_win2590 <= scan_win2589; scan_win2591 <= scan_win2590; scan_win2592 <= scan_win2591; scan_win2593 <= scan_win2592; scan_win2594 <= scan_win2593; scan_win2595 <= scan_win2594; scan_win2596 <= scan_win2595; scan_win2597 <= scan_win2596; scan_win2598 <= scan_win2597; scan_win2599 <= scan_win2598; scan_win2600 <= scan_win2599; 
      scan_win2601 <= scan_win2600; scan_win2602 <= scan_win2601; scan_win2603 <= scan_win2602; scan_win2604 <= scan_win2603; scan_win2605 <= scan_win2604; scan_win2606 <= scan_win2605; scan_win2607 <= scan_win2606; scan_win2608 <= scan_win2607; scan_win2609 <= scan_win2608; scan_win2610 <= scan_win2609; scan_win2611 <= scan_win2610; scan_win2612 <= scan_win2611; scan_win2613 <= scan_win2612; scan_win2614 <= scan_win2613; scan_win2615 <= scan_win2614; scan_win2616 <= scan_win2615; scan_win2617 <= scan_win2616; scan_win2618 <= scan_win2617; scan_win2619 <= scan_win2618; scan_win2620 <= scan_win2619; scan_win2621 <= scan_win2620; scan_win2622 <= scan_win2621; scan_win2623 <= scan_win2622; scan_win2624 <= scan_win2623; scan_win2625 <= scan_win2624; scan_win2626 <= scan_win2625; scan_win2627 <= scan_win2626; scan_win2628 <= scan_win2627; scan_win2629 <= scan_win2628; scan_win2630 <= scan_win2629; scan_win2631 <= scan_win2630; scan_win2632 <= scan_win2631; scan_win2633 <= scan_win2632; scan_win2634 <= scan_win2633; scan_win2635 <= scan_win2634; scan_win2636 <= scan_win2635; scan_win2637 <= scan_win2636; scan_win2638 <= scan_win2637; scan_win2639 <= scan_win2638; scan_win2640 <= scan_win2639; scan_win2641 <= scan_win2640; scan_win2642 <= scan_win2641; scan_win2643 <= scan_win2642; scan_win2644 <= scan_win2643; scan_win2645 <= scan_win2644; scan_win2646 <= scan_win2645; scan_win2647 <= scan_win2646; scan_win2648 <= scan_win2647; scan_win2649 <= scan_win2648; scan_win2650 <= scan_win2649; scan_win2651 <= scan_win2650; scan_win2652 <= scan_win2651; scan_win2653 <= scan_win2652; scan_win2654 <= scan_win2653; scan_win2655 <= scan_win2654; scan_win2656 <= scan_win2655; scan_win2657 <= scan_win2656; scan_win2658 <= scan_win2657; scan_win2659 <= scan_win2658; scan_win2660 <= scan_win2659; scan_win2661 <= scan_win2660; scan_win2662 <= scan_win2661; scan_win2663 <= scan_win2662; scan_win2664 <= scan_win2663; scan_win2665 <= scan_win2664; scan_win2666 <= scan_win2665; scan_win2667 <= scan_win2666; scan_win2668 <= scan_win2667; scan_win2669 <= scan_win2668; scan_win2670 <= scan_win2669; scan_win2671 <= scan_win2670; scan_win2672 <= scan_win2671; scan_win2673 <= scan_win2672; scan_win2674 <= scan_win2673; scan_win2675 <= scan_win2674; scan_win2676 <= scan_win2675; scan_win2677 <= scan_win2676; scan_win2678 <= scan_win2677; scan_win2679 <= scan_win2678; scan_win2680 <= scan_win2679; scan_win2681 <= scan_win2680; scan_win2682 <= scan_win2681; scan_win2683 <= scan_win2682; scan_win2684 <= scan_win2683; scan_win2685 <= scan_win2684; scan_win2686 <= scan_win2685; scan_win2687 <= scan_win2686; scan_win2688 <= scan_win2687; scan_win2689 <= scan_win2688; scan_win2690 <= scan_win2689; scan_win2691 <= scan_win2690; scan_win2692 <= scan_win2691; scan_win2693 <= scan_win2692; scan_win2694 <= scan_win2693; scan_win2695 <= scan_win2694; scan_win2696 <= scan_win2695; scan_win2697 <= scan_win2696; scan_win2698 <= scan_win2697; scan_win2699 <= scan_win2698; scan_win2700 <= scan_win2699; scan_win2701 <= scan_win2700; scan_win2702 <= scan_win2701; scan_win2703 <= scan_win2702; scan_win2704 <= scan_win2703; scan_win2705 <= scan_win2704; scan_win2706 <= scan_win2705; scan_win2707 <= scan_win2706; scan_win2708 <= scan_win2707; scan_win2709 <= scan_win2708; scan_win2710 <= scan_win2709; scan_win2711 <= scan_win2710; scan_win2712 <= scan_win2711; scan_win2713 <= scan_win2712; scan_win2714 <= scan_win2713; scan_win2715 <= scan_win2714; scan_win2716 <= scan_win2715; scan_win2717 <= scan_win2716; scan_win2718 <= scan_win2717; scan_win2719 <= scan_win2718; scan_win2720 <= scan_win2719; scan_win2721 <= scan_win2720; scan_win2722 <= scan_win2721; scan_win2723 <= scan_win2722; scan_win2724 <= scan_win2723; scan_win2725 <= scan_win2724; scan_win2726 <= scan_win2725; scan_win2727 <= scan_win2726; scan_win2728 <= scan_win2727; scan_win2729 <= scan_win2728; scan_win2730 <= scan_win2729; scan_win2731 <= scan_win2730; scan_win2732 <= scan_win2731; scan_win2733 <= scan_win2732; scan_win2734 <= scan_win2733; scan_win2735 <= scan_win2734; scan_win2736 <= scan_win2735; scan_win2737 <= scan_win2736; scan_win2738 <= scan_win2737; scan_win2739 <= scan_win2738; scan_win2740 <= scan_win2739; scan_win2741 <= scan_win2740; scan_win2742 <= scan_win2741; scan_win2743 <= scan_win2742; scan_win2744 <= scan_win2743; scan_win2745 <= scan_win2744; scan_win2746 <= scan_win2745; scan_win2747 <= scan_win2746; scan_win2748 <= scan_win2747; scan_win2749 <= scan_win2748; scan_win2750 <= scan_win2749; scan_win2751 <= scan_win2750; scan_win2752 <= scan_win2751; scan_win2753 <= scan_win2752; scan_win2754 <= scan_win2753; scan_win2755 <= scan_win2754; scan_win2756 <= scan_win2755; scan_win2757 <= scan_win2756; scan_win2758 <= scan_win2757; scan_win2759 <= scan_win2758; scan_win2760 <= scan_win2759; scan_win2761 <= scan_win2760; scan_win2762 <= scan_win2761; scan_win2763 <= scan_win2762; scan_win2764 <= scan_win2763; scan_win2765 <= scan_win2764; scan_win2766 <= scan_win2765; scan_win2767 <= scan_win2766; scan_win2768 <= scan_win2767; scan_win2769 <= scan_win2768; scan_win2770 <= scan_win2769; scan_win2771 <= scan_win2770; scan_win2772 <= scan_win2771; scan_win2773 <= scan_win2772; scan_win2774 <= scan_win2773; scan_win2775 <= scan_win2774; scan_win2776 <= scan_win2775; scan_win2777 <= scan_win2776; scan_win2778 <= scan_win2777; scan_win2779 <= scan_win2778; scan_win2780 <= scan_win2779; scan_win2781 <= scan_win2780; scan_win2782 <= scan_win2781; scan_win2783 <= scan_win2782; scan_win2784 <= scan_win2783; scan_win2785 <= scan_win2784; scan_win2786 <= scan_win2785; scan_win2787 <= scan_win2786; scan_win2788 <= scan_win2787; scan_win2789 <= scan_win2788; scan_win2790 <= scan_win2789; scan_win2791 <= scan_win2790; scan_win2792 <= scan_win2791; scan_win2793 <= scan_win2792; scan_win2794 <= scan_win2793; scan_win2795 <= scan_win2794; scan_win2796 <= scan_win2795; scan_win2797 <= scan_win2796; scan_win2798 <= scan_win2797; scan_win2799 <= scan_win2798; scan_win2800 <= scan_win2799; 
      scan_win2801 <= scan_win2800; scan_win2802 <= scan_win2801; scan_win2803 <= scan_win2802; scan_win2804 <= scan_win2803; scan_win2805 <= scan_win2804; scan_win2806 <= scan_win2805; scan_win2807 <= scan_win2806; scan_win2808 <= scan_win2807; scan_win2809 <= scan_win2808; scan_win2810 <= scan_win2809; scan_win2811 <= scan_win2810; scan_win2812 <= scan_win2811; scan_win2813 <= scan_win2812; scan_win2814 <= scan_win2813; scan_win2815 <= scan_win2814; scan_win2816 <= scan_win2815; scan_win2817 <= scan_win2816; scan_win2818 <= scan_win2817; scan_win2819 <= scan_win2818; scan_win2820 <= scan_win2819; scan_win2821 <= scan_win2820; scan_win2822 <= scan_win2821; scan_win2823 <= scan_win2822; scan_win2824 <= scan_win2823; scan_win2825 <= scan_win2824; scan_win2826 <= scan_win2825; scan_win2827 <= scan_win2826; scan_win2828 <= scan_win2827; scan_win2829 <= scan_win2828; scan_win2830 <= scan_win2829; scan_win2831 <= scan_win2830; scan_win2832 <= scan_win2831; scan_win2833 <= scan_win2832; scan_win2834 <= scan_win2833; scan_win2835 <= scan_win2834; scan_win2836 <= scan_win2835; scan_win2837 <= scan_win2836; scan_win2838 <= scan_win2837; scan_win2839 <= scan_win2838; scan_win2840 <= scan_win2839; scan_win2841 <= scan_win2840; scan_win2842 <= scan_win2841; scan_win2843 <= scan_win2842; scan_win2844 <= scan_win2843; scan_win2845 <= scan_win2844; scan_win2846 <= scan_win2845; scan_win2847 <= scan_win2846; scan_win2848 <= scan_win2847; scan_win2849 <= scan_win2848; scan_win2850 <= scan_win2849; scan_win2851 <= scan_win2850; scan_win2852 <= scan_win2851; scan_win2853 <= scan_win2852; scan_win2854 <= scan_win2853; scan_win2855 <= scan_win2854; scan_win2856 <= scan_win2855; scan_win2857 <= scan_win2856; scan_win2858 <= scan_win2857; scan_win2859 <= scan_win2858; scan_win2860 <= scan_win2859; scan_win2861 <= scan_win2860; scan_win2862 <= scan_win2861; scan_win2863 <= scan_win2862; scan_win2864 <= scan_win2863; scan_win2865 <= scan_win2864; scan_win2866 <= scan_win2865; scan_win2867 <= scan_win2866; scan_win2868 <= scan_win2867; scan_win2869 <= scan_win2868; scan_win2870 <= scan_win2869; scan_win2871 <= scan_win2870; scan_win2872 <= scan_win2871; scan_win2873 <= scan_win2872; scan_win2874 <= scan_win2873; scan_win2875 <= scan_win2874; scan_win2876 <= scan_win2875; scan_win2877 <= scan_win2876; scan_win2878 <= scan_win2877; scan_win2879 <= scan_win2878; scan_win2880 <= scan_win2879; scan_win2881 <= scan_win2880; scan_win2882 <= scan_win2881; scan_win2883 <= scan_win2882; scan_win2884 <= scan_win2883; scan_win2885 <= scan_win2884; scan_win2886 <= scan_win2885; scan_win2887 <= scan_win2886; scan_win2888 <= scan_win2887; scan_win2889 <= scan_win2888; scan_win2890 <= scan_win2889; scan_win2891 <= scan_win2890; scan_win2892 <= scan_win2891; scan_win2893 <= scan_win2892; scan_win2894 <= scan_win2893; scan_win2895 <= scan_win2894; scan_win2896 <= scan_win2895; scan_win2897 <= scan_win2896; scan_win2898 <= scan_win2897; scan_win2899 <= scan_win2898; scan_win2900 <= scan_win2899; scan_win2901 <= scan_win2900; scan_win2902 <= scan_win2901; scan_win2903 <= scan_win2902; scan_win2904 <= scan_win2903; scan_win2905 <= scan_win2904; scan_win2906 <= scan_win2905; scan_win2907 <= scan_win2906; scan_win2908 <= scan_win2907; scan_win2909 <= scan_win2908; scan_win2910 <= scan_win2909; scan_win2911 <= scan_win2910; scan_win2912 <= scan_win2911; 
    end
  end

  accum_calculator #(.RECT1_X(rectangle1_xs[0]), .RECT1_Y(rectangle1_ys[0]), .RECT1_WIDTH(rectangle1_widths[0]), .RECT1_HEIGHT(rectangle1_heights[0]), .RECT1_WEIGHT(rectangle1_weights[0]), .RECT2_X(rectangle2_xs[0]), .RECT2_Y(rectangle2_ys[0]), .RECT2_WIDTH(rectangle2_widths[0]), .RECT2_HEIGHT(rectangle2_heights[0]), .RECT2_WEIGHT(rectangle2_weights[0]), .RECT3_X(rectangle3_xs[0]), .RECT3_Y(rectangle3_ys[0]), .RECT3_WIDTH(rectangle3_widths[0]), .RECT3_HEIGHT(rectangle3_heights[0]), .RECT3_WEIGHT(rectangle3_weights[0]), .FEAT_THRES(feature_thresholds[0]), .FEAT_ABOVE(feature_aboves[0]), .FEAT_BELOW(feature_belows[0])) ac0(.scan_win(scan_win0), .scan_win_std_dev(scan_win_std_dev[0]), .feature_accum(feature_accums[0]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1]), .RECT1_Y(rectangle1_ys[1]), .RECT1_WIDTH(rectangle1_widths[1]), .RECT1_HEIGHT(rectangle1_heights[1]), .RECT1_WEIGHT(rectangle1_weights[1]), .RECT2_X(rectangle2_xs[1]), .RECT2_Y(rectangle2_ys[1]), .RECT2_WIDTH(rectangle2_widths[1]), .RECT2_HEIGHT(rectangle2_heights[1]), .RECT2_WEIGHT(rectangle2_weights[1]), .RECT3_X(rectangle3_xs[1]), .RECT3_Y(rectangle3_ys[1]), .RECT3_WIDTH(rectangle3_widths[1]), .RECT3_HEIGHT(rectangle3_heights[1]), .RECT3_WEIGHT(rectangle3_weights[1]), .FEAT_THRES(feature_thresholds[1]), .FEAT_ABOVE(feature_aboves[1]), .FEAT_BELOW(feature_belows[1])) ac1(.scan_win(scan_win1), .scan_win_std_dev(scan_win_std_dev[1]), .feature_accum(feature_accums[1]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2]), .RECT1_Y(rectangle1_ys[2]), .RECT1_WIDTH(rectangle1_widths[2]), .RECT1_HEIGHT(rectangle1_heights[2]), .RECT1_WEIGHT(rectangle1_weights[2]), .RECT2_X(rectangle2_xs[2]), .RECT2_Y(rectangle2_ys[2]), .RECT2_WIDTH(rectangle2_widths[2]), .RECT2_HEIGHT(rectangle2_heights[2]), .RECT2_WEIGHT(rectangle2_weights[2]), .RECT3_X(rectangle3_xs[2]), .RECT3_Y(rectangle3_ys[2]), .RECT3_WIDTH(rectangle3_widths[2]), .RECT3_HEIGHT(rectangle3_heights[2]), .RECT3_WEIGHT(rectangle3_weights[2]), .FEAT_THRES(feature_thresholds[2]), .FEAT_ABOVE(feature_aboves[2]), .FEAT_BELOW(feature_belows[2])) ac2(.scan_win(scan_win2), .scan_win_std_dev(scan_win_std_dev[2]), .feature_accum(feature_accums[2]));
  accum_calculator #(.RECT1_X(rectangle1_xs[3]), .RECT1_Y(rectangle1_ys[3]), .RECT1_WIDTH(rectangle1_widths[3]), .RECT1_HEIGHT(rectangle1_heights[3]), .RECT1_WEIGHT(rectangle1_weights[3]), .RECT2_X(rectangle2_xs[3]), .RECT2_Y(rectangle2_ys[3]), .RECT2_WIDTH(rectangle2_widths[3]), .RECT2_HEIGHT(rectangle2_heights[3]), .RECT2_WEIGHT(rectangle2_weights[3]), .RECT3_X(rectangle3_xs[3]), .RECT3_Y(rectangle3_ys[3]), .RECT3_WIDTH(rectangle3_widths[3]), .RECT3_HEIGHT(rectangle3_heights[3]), .RECT3_WEIGHT(rectangle3_weights[3]), .FEAT_THRES(feature_thresholds[3]), .FEAT_ABOVE(feature_aboves[3]), .FEAT_BELOW(feature_belows[3])) ac3(.scan_win(scan_win3), .scan_win_std_dev(scan_win_std_dev[3]), .feature_accum(feature_accums[3]));
  accum_calculator #(.RECT1_X(rectangle1_xs[4]), .RECT1_Y(rectangle1_ys[4]), .RECT1_WIDTH(rectangle1_widths[4]), .RECT1_HEIGHT(rectangle1_heights[4]), .RECT1_WEIGHT(rectangle1_weights[4]), .RECT2_X(rectangle2_xs[4]), .RECT2_Y(rectangle2_ys[4]), .RECT2_WIDTH(rectangle2_widths[4]), .RECT2_HEIGHT(rectangle2_heights[4]), .RECT2_WEIGHT(rectangle2_weights[4]), .RECT3_X(rectangle3_xs[4]), .RECT3_Y(rectangle3_ys[4]), .RECT3_WIDTH(rectangle3_widths[4]), .RECT3_HEIGHT(rectangle3_heights[4]), .RECT3_WEIGHT(rectangle3_weights[4]), .FEAT_THRES(feature_thresholds[4]), .FEAT_ABOVE(feature_aboves[4]), .FEAT_BELOW(feature_belows[4])) ac4(.scan_win(scan_win4), .scan_win_std_dev(scan_win_std_dev[4]), .feature_accum(feature_accums[4]));
  accum_calculator #(.RECT1_X(rectangle1_xs[5]), .RECT1_Y(rectangle1_ys[5]), .RECT1_WIDTH(rectangle1_widths[5]), .RECT1_HEIGHT(rectangle1_heights[5]), .RECT1_WEIGHT(rectangle1_weights[5]), .RECT2_X(rectangle2_xs[5]), .RECT2_Y(rectangle2_ys[5]), .RECT2_WIDTH(rectangle2_widths[5]), .RECT2_HEIGHT(rectangle2_heights[5]), .RECT2_WEIGHT(rectangle2_weights[5]), .RECT3_X(rectangle3_xs[5]), .RECT3_Y(rectangle3_ys[5]), .RECT3_WIDTH(rectangle3_widths[5]), .RECT3_HEIGHT(rectangle3_heights[5]), .RECT3_WEIGHT(rectangle3_weights[5]), .FEAT_THRES(feature_thresholds[5]), .FEAT_ABOVE(feature_aboves[5]), .FEAT_BELOW(feature_belows[5])) ac5(.scan_win(scan_win5), .scan_win_std_dev(scan_win_std_dev[5]), .feature_accum(feature_accums[5]));
  accum_calculator #(.RECT1_X(rectangle1_xs[6]), .RECT1_Y(rectangle1_ys[6]), .RECT1_WIDTH(rectangle1_widths[6]), .RECT1_HEIGHT(rectangle1_heights[6]), .RECT1_WEIGHT(rectangle1_weights[6]), .RECT2_X(rectangle2_xs[6]), .RECT2_Y(rectangle2_ys[6]), .RECT2_WIDTH(rectangle2_widths[6]), .RECT2_HEIGHT(rectangle2_heights[6]), .RECT2_WEIGHT(rectangle2_weights[6]), .RECT3_X(rectangle3_xs[6]), .RECT3_Y(rectangle3_ys[6]), .RECT3_WIDTH(rectangle3_widths[6]), .RECT3_HEIGHT(rectangle3_heights[6]), .RECT3_WEIGHT(rectangle3_weights[6]), .FEAT_THRES(feature_thresholds[6]), .FEAT_ABOVE(feature_aboves[6]), .FEAT_BELOW(feature_belows[6])) ac6(.scan_win(scan_win6), .scan_win_std_dev(scan_win_std_dev[6]), .feature_accum(feature_accums[6]));
  accum_calculator #(.RECT1_X(rectangle1_xs[7]), .RECT1_Y(rectangle1_ys[7]), .RECT1_WIDTH(rectangle1_widths[7]), .RECT1_HEIGHT(rectangle1_heights[7]), .RECT1_WEIGHT(rectangle1_weights[7]), .RECT2_X(rectangle2_xs[7]), .RECT2_Y(rectangle2_ys[7]), .RECT2_WIDTH(rectangle2_widths[7]), .RECT2_HEIGHT(rectangle2_heights[7]), .RECT2_WEIGHT(rectangle2_weights[7]), .RECT3_X(rectangle3_xs[7]), .RECT3_Y(rectangle3_ys[7]), .RECT3_WIDTH(rectangle3_widths[7]), .RECT3_HEIGHT(rectangle3_heights[7]), .RECT3_WEIGHT(rectangle3_weights[7]), .FEAT_THRES(feature_thresholds[7]), .FEAT_ABOVE(feature_aboves[7]), .FEAT_BELOW(feature_belows[7])) ac7(.scan_win(scan_win7), .scan_win_std_dev(scan_win_std_dev[7]), .feature_accum(feature_accums[7]));
  accum_calculator #(.RECT1_X(rectangle1_xs[8]), .RECT1_Y(rectangle1_ys[8]), .RECT1_WIDTH(rectangle1_widths[8]), .RECT1_HEIGHT(rectangle1_heights[8]), .RECT1_WEIGHT(rectangle1_weights[8]), .RECT2_X(rectangle2_xs[8]), .RECT2_Y(rectangle2_ys[8]), .RECT2_WIDTH(rectangle2_widths[8]), .RECT2_HEIGHT(rectangle2_heights[8]), .RECT2_WEIGHT(rectangle2_weights[8]), .RECT3_X(rectangle3_xs[8]), .RECT3_Y(rectangle3_ys[8]), .RECT3_WIDTH(rectangle3_widths[8]), .RECT3_HEIGHT(rectangle3_heights[8]), .RECT3_WEIGHT(rectangle3_weights[8]), .FEAT_THRES(feature_thresholds[8]), .FEAT_ABOVE(feature_aboves[8]), .FEAT_BELOW(feature_belows[8])) ac8(.scan_win(scan_win8), .scan_win_std_dev(scan_win_std_dev[8]), .feature_accum(feature_accums[8]));
  accum_calculator #(.RECT1_X(rectangle1_xs[9]), .RECT1_Y(rectangle1_ys[9]), .RECT1_WIDTH(rectangle1_widths[9]), .RECT1_HEIGHT(rectangle1_heights[9]), .RECT1_WEIGHT(rectangle1_weights[9]), .RECT2_X(rectangle2_xs[9]), .RECT2_Y(rectangle2_ys[9]), .RECT2_WIDTH(rectangle2_widths[9]), .RECT2_HEIGHT(rectangle2_heights[9]), .RECT2_WEIGHT(rectangle2_weights[9]), .RECT3_X(rectangle3_xs[9]), .RECT3_Y(rectangle3_ys[9]), .RECT3_WIDTH(rectangle3_widths[9]), .RECT3_HEIGHT(rectangle3_heights[9]), .RECT3_WEIGHT(rectangle3_weights[9]), .FEAT_THRES(feature_thresholds[9]), .FEAT_ABOVE(feature_aboves[9]), .FEAT_BELOW(feature_belows[9])) ac9(.scan_win(scan_win9), .scan_win_std_dev(scan_win_std_dev[9]), .feature_accum(feature_accums[9]));
  accum_calculator #(.RECT1_X(rectangle1_xs[10]), .RECT1_Y(rectangle1_ys[10]), .RECT1_WIDTH(rectangle1_widths[10]), .RECT1_HEIGHT(rectangle1_heights[10]), .RECT1_WEIGHT(rectangle1_weights[10]), .RECT2_X(rectangle2_xs[10]), .RECT2_Y(rectangle2_ys[10]), .RECT2_WIDTH(rectangle2_widths[10]), .RECT2_HEIGHT(rectangle2_heights[10]), .RECT2_WEIGHT(rectangle2_weights[10]), .RECT3_X(rectangle3_xs[10]), .RECT3_Y(rectangle3_ys[10]), .RECT3_WIDTH(rectangle3_widths[10]), .RECT3_HEIGHT(rectangle3_heights[10]), .RECT3_WEIGHT(rectangle3_weights[10]), .FEAT_THRES(feature_thresholds[10]), .FEAT_ABOVE(feature_aboves[10]), .FEAT_BELOW(feature_belows[10])) ac10(.scan_win(scan_win10), .scan_win_std_dev(scan_win_std_dev[10]), .feature_accum(feature_accums[10]));
  accum_calculator #(.RECT1_X(rectangle1_xs[11]), .RECT1_Y(rectangle1_ys[11]), .RECT1_WIDTH(rectangle1_widths[11]), .RECT1_HEIGHT(rectangle1_heights[11]), .RECT1_WEIGHT(rectangle1_weights[11]), .RECT2_X(rectangle2_xs[11]), .RECT2_Y(rectangle2_ys[11]), .RECT2_WIDTH(rectangle2_widths[11]), .RECT2_HEIGHT(rectangle2_heights[11]), .RECT2_WEIGHT(rectangle2_weights[11]), .RECT3_X(rectangle3_xs[11]), .RECT3_Y(rectangle3_ys[11]), .RECT3_WIDTH(rectangle3_widths[11]), .RECT3_HEIGHT(rectangle3_heights[11]), .RECT3_WEIGHT(rectangle3_weights[11]), .FEAT_THRES(feature_thresholds[11]), .FEAT_ABOVE(feature_aboves[11]), .FEAT_BELOW(feature_belows[11])) ac11(.scan_win(scan_win11), .scan_win_std_dev(scan_win_std_dev[11]), .feature_accum(feature_accums[11]));
  accum_calculator #(.RECT1_X(rectangle1_xs[12]), .RECT1_Y(rectangle1_ys[12]), .RECT1_WIDTH(rectangle1_widths[12]), .RECT1_HEIGHT(rectangle1_heights[12]), .RECT1_WEIGHT(rectangle1_weights[12]), .RECT2_X(rectangle2_xs[12]), .RECT2_Y(rectangle2_ys[12]), .RECT2_WIDTH(rectangle2_widths[12]), .RECT2_HEIGHT(rectangle2_heights[12]), .RECT2_WEIGHT(rectangle2_weights[12]), .RECT3_X(rectangle3_xs[12]), .RECT3_Y(rectangle3_ys[12]), .RECT3_WIDTH(rectangle3_widths[12]), .RECT3_HEIGHT(rectangle3_heights[12]), .RECT3_WEIGHT(rectangle3_weights[12]), .FEAT_THRES(feature_thresholds[12]), .FEAT_ABOVE(feature_aboves[12]), .FEAT_BELOW(feature_belows[12])) ac12(.scan_win(scan_win12), .scan_win_std_dev(scan_win_std_dev[12]), .feature_accum(feature_accums[12]));
  accum_calculator #(.RECT1_X(rectangle1_xs[13]), .RECT1_Y(rectangle1_ys[13]), .RECT1_WIDTH(rectangle1_widths[13]), .RECT1_HEIGHT(rectangle1_heights[13]), .RECT1_WEIGHT(rectangle1_weights[13]), .RECT2_X(rectangle2_xs[13]), .RECT2_Y(rectangle2_ys[13]), .RECT2_WIDTH(rectangle2_widths[13]), .RECT2_HEIGHT(rectangle2_heights[13]), .RECT2_WEIGHT(rectangle2_weights[13]), .RECT3_X(rectangle3_xs[13]), .RECT3_Y(rectangle3_ys[13]), .RECT3_WIDTH(rectangle3_widths[13]), .RECT3_HEIGHT(rectangle3_heights[13]), .RECT3_WEIGHT(rectangle3_weights[13]), .FEAT_THRES(feature_thresholds[13]), .FEAT_ABOVE(feature_aboves[13]), .FEAT_BELOW(feature_belows[13])) ac13(.scan_win(scan_win13), .scan_win_std_dev(scan_win_std_dev[13]), .feature_accum(feature_accums[13]));
  accum_calculator #(.RECT1_X(rectangle1_xs[14]), .RECT1_Y(rectangle1_ys[14]), .RECT1_WIDTH(rectangle1_widths[14]), .RECT1_HEIGHT(rectangle1_heights[14]), .RECT1_WEIGHT(rectangle1_weights[14]), .RECT2_X(rectangle2_xs[14]), .RECT2_Y(rectangle2_ys[14]), .RECT2_WIDTH(rectangle2_widths[14]), .RECT2_HEIGHT(rectangle2_heights[14]), .RECT2_WEIGHT(rectangle2_weights[14]), .RECT3_X(rectangle3_xs[14]), .RECT3_Y(rectangle3_ys[14]), .RECT3_WIDTH(rectangle3_widths[14]), .RECT3_HEIGHT(rectangle3_heights[14]), .RECT3_WEIGHT(rectangle3_weights[14]), .FEAT_THRES(feature_thresholds[14]), .FEAT_ABOVE(feature_aboves[14]), .FEAT_BELOW(feature_belows[14])) ac14(.scan_win(scan_win14), .scan_win_std_dev(scan_win_std_dev[14]), .feature_accum(feature_accums[14]));
  accum_calculator #(.RECT1_X(rectangle1_xs[15]), .RECT1_Y(rectangle1_ys[15]), .RECT1_WIDTH(rectangle1_widths[15]), .RECT1_HEIGHT(rectangle1_heights[15]), .RECT1_WEIGHT(rectangle1_weights[15]), .RECT2_X(rectangle2_xs[15]), .RECT2_Y(rectangle2_ys[15]), .RECT2_WIDTH(rectangle2_widths[15]), .RECT2_HEIGHT(rectangle2_heights[15]), .RECT2_WEIGHT(rectangle2_weights[15]), .RECT3_X(rectangle3_xs[15]), .RECT3_Y(rectangle3_ys[15]), .RECT3_WIDTH(rectangle3_widths[15]), .RECT3_HEIGHT(rectangle3_heights[15]), .RECT3_WEIGHT(rectangle3_weights[15]), .FEAT_THRES(feature_thresholds[15]), .FEAT_ABOVE(feature_aboves[15]), .FEAT_BELOW(feature_belows[15])) ac15(.scan_win(scan_win15), .scan_win_std_dev(scan_win_std_dev[15]), .feature_accum(feature_accums[15]));
  accum_calculator #(.RECT1_X(rectangle1_xs[16]), .RECT1_Y(rectangle1_ys[16]), .RECT1_WIDTH(rectangle1_widths[16]), .RECT1_HEIGHT(rectangle1_heights[16]), .RECT1_WEIGHT(rectangle1_weights[16]), .RECT2_X(rectangle2_xs[16]), .RECT2_Y(rectangle2_ys[16]), .RECT2_WIDTH(rectangle2_widths[16]), .RECT2_HEIGHT(rectangle2_heights[16]), .RECT2_WEIGHT(rectangle2_weights[16]), .RECT3_X(rectangle3_xs[16]), .RECT3_Y(rectangle3_ys[16]), .RECT3_WIDTH(rectangle3_widths[16]), .RECT3_HEIGHT(rectangle3_heights[16]), .RECT3_WEIGHT(rectangle3_weights[16]), .FEAT_THRES(feature_thresholds[16]), .FEAT_ABOVE(feature_aboves[16]), .FEAT_BELOW(feature_belows[16])) ac16(.scan_win(scan_win16), .scan_win_std_dev(scan_win_std_dev[16]), .feature_accum(feature_accums[16]));
  accum_calculator #(.RECT1_X(rectangle1_xs[17]), .RECT1_Y(rectangle1_ys[17]), .RECT1_WIDTH(rectangle1_widths[17]), .RECT1_HEIGHT(rectangle1_heights[17]), .RECT1_WEIGHT(rectangle1_weights[17]), .RECT2_X(rectangle2_xs[17]), .RECT2_Y(rectangle2_ys[17]), .RECT2_WIDTH(rectangle2_widths[17]), .RECT2_HEIGHT(rectangle2_heights[17]), .RECT2_WEIGHT(rectangle2_weights[17]), .RECT3_X(rectangle3_xs[17]), .RECT3_Y(rectangle3_ys[17]), .RECT3_WIDTH(rectangle3_widths[17]), .RECT3_HEIGHT(rectangle3_heights[17]), .RECT3_WEIGHT(rectangle3_weights[17]), .FEAT_THRES(feature_thresholds[17]), .FEAT_ABOVE(feature_aboves[17]), .FEAT_BELOW(feature_belows[17])) ac17(.scan_win(scan_win17), .scan_win_std_dev(scan_win_std_dev[17]), .feature_accum(feature_accums[17]));
  accum_calculator #(.RECT1_X(rectangle1_xs[18]), .RECT1_Y(rectangle1_ys[18]), .RECT1_WIDTH(rectangle1_widths[18]), .RECT1_HEIGHT(rectangle1_heights[18]), .RECT1_WEIGHT(rectangle1_weights[18]), .RECT2_X(rectangle2_xs[18]), .RECT2_Y(rectangle2_ys[18]), .RECT2_WIDTH(rectangle2_widths[18]), .RECT2_HEIGHT(rectangle2_heights[18]), .RECT2_WEIGHT(rectangle2_weights[18]), .RECT3_X(rectangle3_xs[18]), .RECT3_Y(rectangle3_ys[18]), .RECT3_WIDTH(rectangle3_widths[18]), .RECT3_HEIGHT(rectangle3_heights[18]), .RECT3_WEIGHT(rectangle3_weights[18]), .FEAT_THRES(feature_thresholds[18]), .FEAT_ABOVE(feature_aboves[18]), .FEAT_BELOW(feature_belows[18])) ac18(.scan_win(scan_win18), .scan_win_std_dev(scan_win_std_dev[18]), .feature_accum(feature_accums[18]));
  accum_calculator #(.RECT1_X(rectangle1_xs[19]), .RECT1_Y(rectangle1_ys[19]), .RECT1_WIDTH(rectangle1_widths[19]), .RECT1_HEIGHT(rectangle1_heights[19]), .RECT1_WEIGHT(rectangle1_weights[19]), .RECT2_X(rectangle2_xs[19]), .RECT2_Y(rectangle2_ys[19]), .RECT2_WIDTH(rectangle2_widths[19]), .RECT2_HEIGHT(rectangle2_heights[19]), .RECT2_WEIGHT(rectangle2_weights[19]), .RECT3_X(rectangle3_xs[19]), .RECT3_Y(rectangle3_ys[19]), .RECT3_WIDTH(rectangle3_widths[19]), .RECT3_HEIGHT(rectangle3_heights[19]), .RECT3_WEIGHT(rectangle3_weights[19]), .FEAT_THRES(feature_thresholds[19]), .FEAT_ABOVE(feature_aboves[19]), .FEAT_BELOW(feature_belows[19])) ac19(.scan_win(scan_win19), .scan_win_std_dev(scan_win_std_dev[19]), .feature_accum(feature_accums[19]));
  accum_calculator #(.RECT1_X(rectangle1_xs[20]), .RECT1_Y(rectangle1_ys[20]), .RECT1_WIDTH(rectangle1_widths[20]), .RECT1_HEIGHT(rectangle1_heights[20]), .RECT1_WEIGHT(rectangle1_weights[20]), .RECT2_X(rectangle2_xs[20]), .RECT2_Y(rectangle2_ys[20]), .RECT2_WIDTH(rectangle2_widths[20]), .RECT2_HEIGHT(rectangle2_heights[20]), .RECT2_WEIGHT(rectangle2_weights[20]), .RECT3_X(rectangle3_xs[20]), .RECT3_Y(rectangle3_ys[20]), .RECT3_WIDTH(rectangle3_widths[20]), .RECT3_HEIGHT(rectangle3_heights[20]), .RECT3_WEIGHT(rectangle3_weights[20]), .FEAT_THRES(feature_thresholds[20]), .FEAT_ABOVE(feature_aboves[20]), .FEAT_BELOW(feature_belows[20])) ac20(.scan_win(scan_win20), .scan_win_std_dev(scan_win_std_dev[20]), .feature_accum(feature_accums[20]));
  accum_calculator #(.RECT1_X(rectangle1_xs[21]), .RECT1_Y(rectangle1_ys[21]), .RECT1_WIDTH(rectangle1_widths[21]), .RECT1_HEIGHT(rectangle1_heights[21]), .RECT1_WEIGHT(rectangle1_weights[21]), .RECT2_X(rectangle2_xs[21]), .RECT2_Y(rectangle2_ys[21]), .RECT2_WIDTH(rectangle2_widths[21]), .RECT2_HEIGHT(rectangle2_heights[21]), .RECT2_WEIGHT(rectangle2_weights[21]), .RECT3_X(rectangle3_xs[21]), .RECT3_Y(rectangle3_ys[21]), .RECT3_WIDTH(rectangle3_widths[21]), .RECT3_HEIGHT(rectangle3_heights[21]), .RECT3_WEIGHT(rectangle3_weights[21]), .FEAT_THRES(feature_thresholds[21]), .FEAT_ABOVE(feature_aboves[21]), .FEAT_BELOW(feature_belows[21])) ac21(.scan_win(scan_win21), .scan_win_std_dev(scan_win_std_dev[21]), .feature_accum(feature_accums[21]));
  accum_calculator #(.RECT1_X(rectangle1_xs[22]), .RECT1_Y(rectangle1_ys[22]), .RECT1_WIDTH(rectangle1_widths[22]), .RECT1_HEIGHT(rectangle1_heights[22]), .RECT1_WEIGHT(rectangle1_weights[22]), .RECT2_X(rectangle2_xs[22]), .RECT2_Y(rectangle2_ys[22]), .RECT2_WIDTH(rectangle2_widths[22]), .RECT2_HEIGHT(rectangle2_heights[22]), .RECT2_WEIGHT(rectangle2_weights[22]), .RECT3_X(rectangle3_xs[22]), .RECT3_Y(rectangle3_ys[22]), .RECT3_WIDTH(rectangle3_widths[22]), .RECT3_HEIGHT(rectangle3_heights[22]), .RECT3_WEIGHT(rectangle3_weights[22]), .FEAT_THRES(feature_thresholds[22]), .FEAT_ABOVE(feature_aboves[22]), .FEAT_BELOW(feature_belows[22])) ac22(.scan_win(scan_win22), .scan_win_std_dev(scan_win_std_dev[22]), .feature_accum(feature_accums[22]));
  accum_calculator #(.RECT1_X(rectangle1_xs[23]), .RECT1_Y(rectangle1_ys[23]), .RECT1_WIDTH(rectangle1_widths[23]), .RECT1_HEIGHT(rectangle1_heights[23]), .RECT1_WEIGHT(rectangle1_weights[23]), .RECT2_X(rectangle2_xs[23]), .RECT2_Y(rectangle2_ys[23]), .RECT2_WIDTH(rectangle2_widths[23]), .RECT2_HEIGHT(rectangle2_heights[23]), .RECT2_WEIGHT(rectangle2_weights[23]), .RECT3_X(rectangle3_xs[23]), .RECT3_Y(rectangle3_ys[23]), .RECT3_WIDTH(rectangle3_widths[23]), .RECT3_HEIGHT(rectangle3_heights[23]), .RECT3_WEIGHT(rectangle3_weights[23]), .FEAT_THRES(feature_thresholds[23]), .FEAT_ABOVE(feature_aboves[23]), .FEAT_BELOW(feature_belows[23])) ac23(.scan_win(scan_win23), .scan_win_std_dev(scan_win_std_dev[23]), .feature_accum(feature_accums[23]));
  accum_calculator #(.RECT1_X(rectangle1_xs[24]), .RECT1_Y(rectangle1_ys[24]), .RECT1_WIDTH(rectangle1_widths[24]), .RECT1_HEIGHT(rectangle1_heights[24]), .RECT1_WEIGHT(rectangle1_weights[24]), .RECT2_X(rectangle2_xs[24]), .RECT2_Y(rectangle2_ys[24]), .RECT2_WIDTH(rectangle2_widths[24]), .RECT2_HEIGHT(rectangle2_heights[24]), .RECT2_WEIGHT(rectangle2_weights[24]), .RECT3_X(rectangle3_xs[24]), .RECT3_Y(rectangle3_ys[24]), .RECT3_WIDTH(rectangle3_widths[24]), .RECT3_HEIGHT(rectangle3_heights[24]), .RECT3_WEIGHT(rectangle3_weights[24]), .FEAT_THRES(feature_thresholds[24]), .FEAT_ABOVE(feature_aboves[24]), .FEAT_BELOW(feature_belows[24])) ac24(.scan_win(scan_win24), .scan_win_std_dev(scan_win_std_dev[24]), .feature_accum(feature_accums[24]));
  accum_calculator #(.RECT1_X(rectangle1_xs[25]), .RECT1_Y(rectangle1_ys[25]), .RECT1_WIDTH(rectangle1_widths[25]), .RECT1_HEIGHT(rectangle1_heights[25]), .RECT1_WEIGHT(rectangle1_weights[25]), .RECT2_X(rectangle2_xs[25]), .RECT2_Y(rectangle2_ys[25]), .RECT2_WIDTH(rectangle2_widths[25]), .RECT2_HEIGHT(rectangle2_heights[25]), .RECT2_WEIGHT(rectangle2_weights[25]), .RECT3_X(rectangle3_xs[25]), .RECT3_Y(rectangle3_ys[25]), .RECT3_WIDTH(rectangle3_widths[25]), .RECT3_HEIGHT(rectangle3_heights[25]), .RECT3_WEIGHT(rectangle3_weights[25]), .FEAT_THRES(feature_thresholds[25]), .FEAT_ABOVE(feature_aboves[25]), .FEAT_BELOW(feature_belows[25])) ac25(.scan_win(scan_win25), .scan_win_std_dev(scan_win_std_dev[25]), .feature_accum(feature_accums[25]));
  accum_calculator #(.RECT1_X(rectangle1_xs[26]), .RECT1_Y(rectangle1_ys[26]), .RECT1_WIDTH(rectangle1_widths[26]), .RECT1_HEIGHT(rectangle1_heights[26]), .RECT1_WEIGHT(rectangle1_weights[26]), .RECT2_X(rectangle2_xs[26]), .RECT2_Y(rectangle2_ys[26]), .RECT2_WIDTH(rectangle2_widths[26]), .RECT2_HEIGHT(rectangle2_heights[26]), .RECT2_WEIGHT(rectangle2_weights[26]), .RECT3_X(rectangle3_xs[26]), .RECT3_Y(rectangle3_ys[26]), .RECT3_WIDTH(rectangle3_widths[26]), .RECT3_HEIGHT(rectangle3_heights[26]), .RECT3_WEIGHT(rectangle3_weights[26]), .FEAT_THRES(feature_thresholds[26]), .FEAT_ABOVE(feature_aboves[26]), .FEAT_BELOW(feature_belows[26])) ac26(.scan_win(scan_win26), .scan_win_std_dev(scan_win_std_dev[26]), .feature_accum(feature_accums[26]));
  accum_calculator #(.RECT1_X(rectangle1_xs[27]), .RECT1_Y(rectangle1_ys[27]), .RECT1_WIDTH(rectangle1_widths[27]), .RECT1_HEIGHT(rectangle1_heights[27]), .RECT1_WEIGHT(rectangle1_weights[27]), .RECT2_X(rectangle2_xs[27]), .RECT2_Y(rectangle2_ys[27]), .RECT2_WIDTH(rectangle2_widths[27]), .RECT2_HEIGHT(rectangle2_heights[27]), .RECT2_WEIGHT(rectangle2_weights[27]), .RECT3_X(rectangle3_xs[27]), .RECT3_Y(rectangle3_ys[27]), .RECT3_WIDTH(rectangle3_widths[27]), .RECT3_HEIGHT(rectangle3_heights[27]), .RECT3_WEIGHT(rectangle3_weights[27]), .FEAT_THRES(feature_thresholds[27]), .FEAT_ABOVE(feature_aboves[27]), .FEAT_BELOW(feature_belows[27])) ac27(.scan_win(scan_win27), .scan_win_std_dev(scan_win_std_dev[27]), .feature_accum(feature_accums[27]));
  accum_calculator #(.RECT1_X(rectangle1_xs[28]), .RECT1_Y(rectangle1_ys[28]), .RECT1_WIDTH(rectangle1_widths[28]), .RECT1_HEIGHT(rectangle1_heights[28]), .RECT1_WEIGHT(rectangle1_weights[28]), .RECT2_X(rectangle2_xs[28]), .RECT2_Y(rectangle2_ys[28]), .RECT2_WIDTH(rectangle2_widths[28]), .RECT2_HEIGHT(rectangle2_heights[28]), .RECT2_WEIGHT(rectangle2_weights[28]), .RECT3_X(rectangle3_xs[28]), .RECT3_Y(rectangle3_ys[28]), .RECT3_WIDTH(rectangle3_widths[28]), .RECT3_HEIGHT(rectangle3_heights[28]), .RECT3_WEIGHT(rectangle3_weights[28]), .FEAT_THRES(feature_thresholds[28]), .FEAT_ABOVE(feature_aboves[28]), .FEAT_BELOW(feature_belows[28])) ac28(.scan_win(scan_win28), .scan_win_std_dev(scan_win_std_dev[28]), .feature_accum(feature_accums[28]));
  accum_calculator #(.RECT1_X(rectangle1_xs[29]), .RECT1_Y(rectangle1_ys[29]), .RECT1_WIDTH(rectangle1_widths[29]), .RECT1_HEIGHT(rectangle1_heights[29]), .RECT1_WEIGHT(rectangle1_weights[29]), .RECT2_X(rectangle2_xs[29]), .RECT2_Y(rectangle2_ys[29]), .RECT2_WIDTH(rectangle2_widths[29]), .RECT2_HEIGHT(rectangle2_heights[29]), .RECT2_WEIGHT(rectangle2_weights[29]), .RECT3_X(rectangle3_xs[29]), .RECT3_Y(rectangle3_ys[29]), .RECT3_WIDTH(rectangle3_widths[29]), .RECT3_HEIGHT(rectangle3_heights[29]), .RECT3_WEIGHT(rectangle3_weights[29]), .FEAT_THRES(feature_thresholds[29]), .FEAT_ABOVE(feature_aboves[29]), .FEAT_BELOW(feature_belows[29])) ac29(.scan_win(scan_win29), .scan_win_std_dev(scan_win_std_dev[29]), .feature_accum(feature_accums[29]));
  accum_calculator #(.RECT1_X(rectangle1_xs[30]), .RECT1_Y(rectangle1_ys[30]), .RECT1_WIDTH(rectangle1_widths[30]), .RECT1_HEIGHT(rectangle1_heights[30]), .RECT1_WEIGHT(rectangle1_weights[30]), .RECT2_X(rectangle2_xs[30]), .RECT2_Y(rectangle2_ys[30]), .RECT2_WIDTH(rectangle2_widths[30]), .RECT2_HEIGHT(rectangle2_heights[30]), .RECT2_WEIGHT(rectangle2_weights[30]), .RECT3_X(rectangle3_xs[30]), .RECT3_Y(rectangle3_ys[30]), .RECT3_WIDTH(rectangle3_widths[30]), .RECT3_HEIGHT(rectangle3_heights[30]), .RECT3_WEIGHT(rectangle3_weights[30]), .FEAT_THRES(feature_thresholds[30]), .FEAT_ABOVE(feature_aboves[30]), .FEAT_BELOW(feature_belows[30])) ac30(.scan_win(scan_win30), .scan_win_std_dev(scan_win_std_dev[30]), .feature_accum(feature_accums[30]));
  accum_calculator #(.RECT1_X(rectangle1_xs[31]), .RECT1_Y(rectangle1_ys[31]), .RECT1_WIDTH(rectangle1_widths[31]), .RECT1_HEIGHT(rectangle1_heights[31]), .RECT1_WEIGHT(rectangle1_weights[31]), .RECT2_X(rectangle2_xs[31]), .RECT2_Y(rectangle2_ys[31]), .RECT2_WIDTH(rectangle2_widths[31]), .RECT2_HEIGHT(rectangle2_heights[31]), .RECT2_WEIGHT(rectangle2_weights[31]), .RECT3_X(rectangle3_xs[31]), .RECT3_Y(rectangle3_ys[31]), .RECT3_WIDTH(rectangle3_widths[31]), .RECT3_HEIGHT(rectangle3_heights[31]), .RECT3_WEIGHT(rectangle3_weights[31]), .FEAT_THRES(feature_thresholds[31]), .FEAT_ABOVE(feature_aboves[31]), .FEAT_BELOW(feature_belows[31])) ac31(.scan_win(scan_win31), .scan_win_std_dev(scan_win_std_dev[31]), .feature_accum(feature_accums[31]));
  accum_calculator #(.RECT1_X(rectangle1_xs[32]), .RECT1_Y(rectangle1_ys[32]), .RECT1_WIDTH(rectangle1_widths[32]), .RECT1_HEIGHT(rectangle1_heights[32]), .RECT1_WEIGHT(rectangle1_weights[32]), .RECT2_X(rectangle2_xs[32]), .RECT2_Y(rectangle2_ys[32]), .RECT2_WIDTH(rectangle2_widths[32]), .RECT2_HEIGHT(rectangle2_heights[32]), .RECT2_WEIGHT(rectangle2_weights[32]), .RECT3_X(rectangle3_xs[32]), .RECT3_Y(rectangle3_ys[32]), .RECT3_WIDTH(rectangle3_widths[32]), .RECT3_HEIGHT(rectangle3_heights[32]), .RECT3_WEIGHT(rectangle3_weights[32]), .FEAT_THRES(feature_thresholds[32]), .FEAT_ABOVE(feature_aboves[32]), .FEAT_BELOW(feature_belows[32])) ac32(.scan_win(scan_win32), .scan_win_std_dev(scan_win_std_dev[32]), .feature_accum(feature_accums[32]));
  accum_calculator #(.RECT1_X(rectangle1_xs[33]), .RECT1_Y(rectangle1_ys[33]), .RECT1_WIDTH(rectangle1_widths[33]), .RECT1_HEIGHT(rectangle1_heights[33]), .RECT1_WEIGHT(rectangle1_weights[33]), .RECT2_X(rectangle2_xs[33]), .RECT2_Y(rectangle2_ys[33]), .RECT2_WIDTH(rectangle2_widths[33]), .RECT2_HEIGHT(rectangle2_heights[33]), .RECT2_WEIGHT(rectangle2_weights[33]), .RECT3_X(rectangle3_xs[33]), .RECT3_Y(rectangle3_ys[33]), .RECT3_WIDTH(rectangle3_widths[33]), .RECT3_HEIGHT(rectangle3_heights[33]), .RECT3_WEIGHT(rectangle3_weights[33]), .FEAT_THRES(feature_thresholds[33]), .FEAT_ABOVE(feature_aboves[33]), .FEAT_BELOW(feature_belows[33])) ac33(.scan_win(scan_win33), .scan_win_std_dev(scan_win_std_dev[33]), .feature_accum(feature_accums[33]));
  accum_calculator #(.RECT1_X(rectangle1_xs[34]), .RECT1_Y(rectangle1_ys[34]), .RECT1_WIDTH(rectangle1_widths[34]), .RECT1_HEIGHT(rectangle1_heights[34]), .RECT1_WEIGHT(rectangle1_weights[34]), .RECT2_X(rectangle2_xs[34]), .RECT2_Y(rectangle2_ys[34]), .RECT2_WIDTH(rectangle2_widths[34]), .RECT2_HEIGHT(rectangle2_heights[34]), .RECT2_WEIGHT(rectangle2_weights[34]), .RECT3_X(rectangle3_xs[34]), .RECT3_Y(rectangle3_ys[34]), .RECT3_WIDTH(rectangle3_widths[34]), .RECT3_HEIGHT(rectangle3_heights[34]), .RECT3_WEIGHT(rectangle3_weights[34]), .FEAT_THRES(feature_thresholds[34]), .FEAT_ABOVE(feature_aboves[34]), .FEAT_BELOW(feature_belows[34])) ac34(.scan_win(scan_win34), .scan_win_std_dev(scan_win_std_dev[34]), .feature_accum(feature_accums[34]));
  accum_calculator #(.RECT1_X(rectangle1_xs[35]), .RECT1_Y(rectangle1_ys[35]), .RECT1_WIDTH(rectangle1_widths[35]), .RECT1_HEIGHT(rectangle1_heights[35]), .RECT1_WEIGHT(rectangle1_weights[35]), .RECT2_X(rectangle2_xs[35]), .RECT2_Y(rectangle2_ys[35]), .RECT2_WIDTH(rectangle2_widths[35]), .RECT2_HEIGHT(rectangle2_heights[35]), .RECT2_WEIGHT(rectangle2_weights[35]), .RECT3_X(rectangle3_xs[35]), .RECT3_Y(rectangle3_ys[35]), .RECT3_WIDTH(rectangle3_widths[35]), .RECT3_HEIGHT(rectangle3_heights[35]), .RECT3_WEIGHT(rectangle3_weights[35]), .FEAT_THRES(feature_thresholds[35]), .FEAT_ABOVE(feature_aboves[35]), .FEAT_BELOW(feature_belows[35])) ac35(.scan_win(scan_win35), .scan_win_std_dev(scan_win_std_dev[35]), .feature_accum(feature_accums[35]));
  accum_calculator #(.RECT1_X(rectangle1_xs[36]), .RECT1_Y(rectangle1_ys[36]), .RECT1_WIDTH(rectangle1_widths[36]), .RECT1_HEIGHT(rectangle1_heights[36]), .RECT1_WEIGHT(rectangle1_weights[36]), .RECT2_X(rectangle2_xs[36]), .RECT2_Y(rectangle2_ys[36]), .RECT2_WIDTH(rectangle2_widths[36]), .RECT2_HEIGHT(rectangle2_heights[36]), .RECT2_WEIGHT(rectangle2_weights[36]), .RECT3_X(rectangle3_xs[36]), .RECT3_Y(rectangle3_ys[36]), .RECT3_WIDTH(rectangle3_widths[36]), .RECT3_HEIGHT(rectangle3_heights[36]), .RECT3_WEIGHT(rectangle3_weights[36]), .FEAT_THRES(feature_thresholds[36]), .FEAT_ABOVE(feature_aboves[36]), .FEAT_BELOW(feature_belows[36])) ac36(.scan_win(scan_win36), .scan_win_std_dev(scan_win_std_dev[36]), .feature_accum(feature_accums[36]));
  accum_calculator #(.RECT1_X(rectangle1_xs[37]), .RECT1_Y(rectangle1_ys[37]), .RECT1_WIDTH(rectangle1_widths[37]), .RECT1_HEIGHT(rectangle1_heights[37]), .RECT1_WEIGHT(rectangle1_weights[37]), .RECT2_X(rectangle2_xs[37]), .RECT2_Y(rectangle2_ys[37]), .RECT2_WIDTH(rectangle2_widths[37]), .RECT2_HEIGHT(rectangle2_heights[37]), .RECT2_WEIGHT(rectangle2_weights[37]), .RECT3_X(rectangle3_xs[37]), .RECT3_Y(rectangle3_ys[37]), .RECT3_WIDTH(rectangle3_widths[37]), .RECT3_HEIGHT(rectangle3_heights[37]), .RECT3_WEIGHT(rectangle3_weights[37]), .FEAT_THRES(feature_thresholds[37]), .FEAT_ABOVE(feature_aboves[37]), .FEAT_BELOW(feature_belows[37])) ac37(.scan_win(scan_win37), .scan_win_std_dev(scan_win_std_dev[37]), .feature_accum(feature_accums[37]));
  accum_calculator #(.RECT1_X(rectangle1_xs[38]), .RECT1_Y(rectangle1_ys[38]), .RECT1_WIDTH(rectangle1_widths[38]), .RECT1_HEIGHT(rectangle1_heights[38]), .RECT1_WEIGHT(rectangle1_weights[38]), .RECT2_X(rectangle2_xs[38]), .RECT2_Y(rectangle2_ys[38]), .RECT2_WIDTH(rectangle2_widths[38]), .RECT2_HEIGHT(rectangle2_heights[38]), .RECT2_WEIGHT(rectangle2_weights[38]), .RECT3_X(rectangle3_xs[38]), .RECT3_Y(rectangle3_ys[38]), .RECT3_WIDTH(rectangle3_widths[38]), .RECT3_HEIGHT(rectangle3_heights[38]), .RECT3_WEIGHT(rectangle3_weights[38]), .FEAT_THRES(feature_thresholds[38]), .FEAT_ABOVE(feature_aboves[38]), .FEAT_BELOW(feature_belows[38])) ac38(.scan_win(scan_win38), .scan_win_std_dev(scan_win_std_dev[38]), .feature_accum(feature_accums[38]));
  accum_calculator #(.RECT1_X(rectangle1_xs[39]), .RECT1_Y(rectangle1_ys[39]), .RECT1_WIDTH(rectangle1_widths[39]), .RECT1_HEIGHT(rectangle1_heights[39]), .RECT1_WEIGHT(rectangle1_weights[39]), .RECT2_X(rectangle2_xs[39]), .RECT2_Y(rectangle2_ys[39]), .RECT2_WIDTH(rectangle2_widths[39]), .RECT2_HEIGHT(rectangle2_heights[39]), .RECT2_WEIGHT(rectangle2_weights[39]), .RECT3_X(rectangle3_xs[39]), .RECT3_Y(rectangle3_ys[39]), .RECT3_WIDTH(rectangle3_widths[39]), .RECT3_HEIGHT(rectangle3_heights[39]), .RECT3_WEIGHT(rectangle3_weights[39]), .FEAT_THRES(feature_thresholds[39]), .FEAT_ABOVE(feature_aboves[39]), .FEAT_BELOW(feature_belows[39])) ac39(.scan_win(scan_win39), .scan_win_std_dev(scan_win_std_dev[39]), .feature_accum(feature_accums[39]));
  accum_calculator #(.RECT1_X(rectangle1_xs[40]), .RECT1_Y(rectangle1_ys[40]), .RECT1_WIDTH(rectangle1_widths[40]), .RECT1_HEIGHT(rectangle1_heights[40]), .RECT1_WEIGHT(rectangle1_weights[40]), .RECT2_X(rectangle2_xs[40]), .RECT2_Y(rectangle2_ys[40]), .RECT2_WIDTH(rectangle2_widths[40]), .RECT2_HEIGHT(rectangle2_heights[40]), .RECT2_WEIGHT(rectangle2_weights[40]), .RECT3_X(rectangle3_xs[40]), .RECT3_Y(rectangle3_ys[40]), .RECT3_WIDTH(rectangle3_widths[40]), .RECT3_HEIGHT(rectangle3_heights[40]), .RECT3_WEIGHT(rectangle3_weights[40]), .FEAT_THRES(feature_thresholds[40]), .FEAT_ABOVE(feature_aboves[40]), .FEAT_BELOW(feature_belows[40])) ac40(.scan_win(scan_win40), .scan_win_std_dev(scan_win_std_dev[40]), .feature_accum(feature_accums[40]));
  accum_calculator #(.RECT1_X(rectangle1_xs[41]), .RECT1_Y(rectangle1_ys[41]), .RECT1_WIDTH(rectangle1_widths[41]), .RECT1_HEIGHT(rectangle1_heights[41]), .RECT1_WEIGHT(rectangle1_weights[41]), .RECT2_X(rectangle2_xs[41]), .RECT2_Y(rectangle2_ys[41]), .RECT2_WIDTH(rectangle2_widths[41]), .RECT2_HEIGHT(rectangle2_heights[41]), .RECT2_WEIGHT(rectangle2_weights[41]), .RECT3_X(rectangle3_xs[41]), .RECT3_Y(rectangle3_ys[41]), .RECT3_WIDTH(rectangle3_widths[41]), .RECT3_HEIGHT(rectangle3_heights[41]), .RECT3_WEIGHT(rectangle3_weights[41]), .FEAT_THRES(feature_thresholds[41]), .FEAT_ABOVE(feature_aboves[41]), .FEAT_BELOW(feature_belows[41])) ac41(.scan_win(scan_win41), .scan_win_std_dev(scan_win_std_dev[41]), .feature_accum(feature_accums[41]));
  accum_calculator #(.RECT1_X(rectangle1_xs[42]), .RECT1_Y(rectangle1_ys[42]), .RECT1_WIDTH(rectangle1_widths[42]), .RECT1_HEIGHT(rectangle1_heights[42]), .RECT1_WEIGHT(rectangle1_weights[42]), .RECT2_X(rectangle2_xs[42]), .RECT2_Y(rectangle2_ys[42]), .RECT2_WIDTH(rectangle2_widths[42]), .RECT2_HEIGHT(rectangle2_heights[42]), .RECT2_WEIGHT(rectangle2_weights[42]), .RECT3_X(rectangle3_xs[42]), .RECT3_Y(rectangle3_ys[42]), .RECT3_WIDTH(rectangle3_widths[42]), .RECT3_HEIGHT(rectangle3_heights[42]), .RECT3_WEIGHT(rectangle3_weights[42]), .FEAT_THRES(feature_thresholds[42]), .FEAT_ABOVE(feature_aboves[42]), .FEAT_BELOW(feature_belows[42])) ac42(.scan_win(scan_win42), .scan_win_std_dev(scan_win_std_dev[42]), .feature_accum(feature_accums[42]));
  accum_calculator #(.RECT1_X(rectangle1_xs[43]), .RECT1_Y(rectangle1_ys[43]), .RECT1_WIDTH(rectangle1_widths[43]), .RECT1_HEIGHT(rectangle1_heights[43]), .RECT1_WEIGHT(rectangle1_weights[43]), .RECT2_X(rectangle2_xs[43]), .RECT2_Y(rectangle2_ys[43]), .RECT2_WIDTH(rectangle2_widths[43]), .RECT2_HEIGHT(rectangle2_heights[43]), .RECT2_WEIGHT(rectangle2_weights[43]), .RECT3_X(rectangle3_xs[43]), .RECT3_Y(rectangle3_ys[43]), .RECT3_WIDTH(rectangle3_widths[43]), .RECT3_HEIGHT(rectangle3_heights[43]), .RECT3_WEIGHT(rectangle3_weights[43]), .FEAT_THRES(feature_thresholds[43]), .FEAT_ABOVE(feature_aboves[43]), .FEAT_BELOW(feature_belows[43])) ac43(.scan_win(scan_win43), .scan_win_std_dev(scan_win_std_dev[43]), .feature_accum(feature_accums[43]));
  accum_calculator #(.RECT1_X(rectangle1_xs[44]), .RECT1_Y(rectangle1_ys[44]), .RECT1_WIDTH(rectangle1_widths[44]), .RECT1_HEIGHT(rectangle1_heights[44]), .RECT1_WEIGHT(rectangle1_weights[44]), .RECT2_X(rectangle2_xs[44]), .RECT2_Y(rectangle2_ys[44]), .RECT2_WIDTH(rectangle2_widths[44]), .RECT2_HEIGHT(rectangle2_heights[44]), .RECT2_WEIGHT(rectangle2_weights[44]), .RECT3_X(rectangle3_xs[44]), .RECT3_Y(rectangle3_ys[44]), .RECT3_WIDTH(rectangle3_widths[44]), .RECT3_HEIGHT(rectangle3_heights[44]), .RECT3_WEIGHT(rectangle3_weights[44]), .FEAT_THRES(feature_thresholds[44]), .FEAT_ABOVE(feature_aboves[44]), .FEAT_BELOW(feature_belows[44])) ac44(.scan_win(scan_win44), .scan_win_std_dev(scan_win_std_dev[44]), .feature_accum(feature_accums[44]));
  accum_calculator #(.RECT1_X(rectangle1_xs[45]), .RECT1_Y(rectangle1_ys[45]), .RECT1_WIDTH(rectangle1_widths[45]), .RECT1_HEIGHT(rectangle1_heights[45]), .RECT1_WEIGHT(rectangle1_weights[45]), .RECT2_X(rectangle2_xs[45]), .RECT2_Y(rectangle2_ys[45]), .RECT2_WIDTH(rectangle2_widths[45]), .RECT2_HEIGHT(rectangle2_heights[45]), .RECT2_WEIGHT(rectangle2_weights[45]), .RECT3_X(rectangle3_xs[45]), .RECT3_Y(rectangle3_ys[45]), .RECT3_WIDTH(rectangle3_widths[45]), .RECT3_HEIGHT(rectangle3_heights[45]), .RECT3_WEIGHT(rectangle3_weights[45]), .FEAT_THRES(feature_thresholds[45]), .FEAT_ABOVE(feature_aboves[45]), .FEAT_BELOW(feature_belows[45])) ac45(.scan_win(scan_win45), .scan_win_std_dev(scan_win_std_dev[45]), .feature_accum(feature_accums[45]));
  accum_calculator #(.RECT1_X(rectangle1_xs[46]), .RECT1_Y(rectangle1_ys[46]), .RECT1_WIDTH(rectangle1_widths[46]), .RECT1_HEIGHT(rectangle1_heights[46]), .RECT1_WEIGHT(rectangle1_weights[46]), .RECT2_X(rectangle2_xs[46]), .RECT2_Y(rectangle2_ys[46]), .RECT2_WIDTH(rectangle2_widths[46]), .RECT2_HEIGHT(rectangle2_heights[46]), .RECT2_WEIGHT(rectangle2_weights[46]), .RECT3_X(rectangle3_xs[46]), .RECT3_Y(rectangle3_ys[46]), .RECT3_WIDTH(rectangle3_widths[46]), .RECT3_HEIGHT(rectangle3_heights[46]), .RECT3_WEIGHT(rectangle3_weights[46]), .FEAT_THRES(feature_thresholds[46]), .FEAT_ABOVE(feature_aboves[46]), .FEAT_BELOW(feature_belows[46])) ac46(.scan_win(scan_win46), .scan_win_std_dev(scan_win_std_dev[46]), .feature_accum(feature_accums[46]));
  accum_calculator #(.RECT1_X(rectangle1_xs[47]), .RECT1_Y(rectangle1_ys[47]), .RECT1_WIDTH(rectangle1_widths[47]), .RECT1_HEIGHT(rectangle1_heights[47]), .RECT1_WEIGHT(rectangle1_weights[47]), .RECT2_X(rectangle2_xs[47]), .RECT2_Y(rectangle2_ys[47]), .RECT2_WIDTH(rectangle2_widths[47]), .RECT2_HEIGHT(rectangle2_heights[47]), .RECT2_WEIGHT(rectangle2_weights[47]), .RECT3_X(rectangle3_xs[47]), .RECT3_Y(rectangle3_ys[47]), .RECT3_WIDTH(rectangle3_widths[47]), .RECT3_HEIGHT(rectangle3_heights[47]), .RECT3_WEIGHT(rectangle3_weights[47]), .FEAT_THRES(feature_thresholds[47]), .FEAT_ABOVE(feature_aboves[47]), .FEAT_BELOW(feature_belows[47])) ac47(.scan_win(scan_win47), .scan_win_std_dev(scan_win_std_dev[47]), .feature_accum(feature_accums[47]));
  accum_calculator #(.RECT1_X(rectangle1_xs[48]), .RECT1_Y(rectangle1_ys[48]), .RECT1_WIDTH(rectangle1_widths[48]), .RECT1_HEIGHT(rectangle1_heights[48]), .RECT1_WEIGHT(rectangle1_weights[48]), .RECT2_X(rectangle2_xs[48]), .RECT2_Y(rectangle2_ys[48]), .RECT2_WIDTH(rectangle2_widths[48]), .RECT2_HEIGHT(rectangle2_heights[48]), .RECT2_WEIGHT(rectangle2_weights[48]), .RECT3_X(rectangle3_xs[48]), .RECT3_Y(rectangle3_ys[48]), .RECT3_WIDTH(rectangle3_widths[48]), .RECT3_HEIGHT(rectangle3_heights[48]), .RECT3_WEIGHT(rectangle3_weights[48]), .FEAT_THRES(feature_thresholds[48]), .FEAT_ABOVE(feature_aboves[48]), .FEAT_BELOW(feature_belows[48])) ac48(.scan_win(scan_win48), .scan_win_std_dev(scan_win_std_dev[48]), .feature_accum(feature_accums[48]));
  accum_calculator #(.RECT1_X(rectangle1_xs[49]), .RECT1_Y(rectangle1_ys[49]), .RECT1_WIDTH(rectangle1_widths[49]), .RECT1_HEIGHT(rectangle1_heights[49]), .RECT1_WEIGHT(rectangle1_weights[49]), .RECT2_X(rectangle2_xs[49]), .RECT2_Y(rectangle2_ys[49]), .RECT2_WIDTH(rectangle2_widths[49]), .RECT2_HEIGHT(rectangle2_heights[49]), .RECT2_WEIGHT(rectangle2_weights[49]), .RECT3_X(rectangle3_xs[49]), .RECT3_Y(rectangle3_ys[49]), .RECT3_WIDTH(rectangle3_widths[49]), .RECT3_HEIGHT(rectangle3_heights[49]), .RECT3_WEIGHT(rectangle3_weights[49]), .FEAT_THRES(feature_thresholds[49]), .FEAT_ABOVE(feature_aboves[49]), .FEAT_BELOW(feature_belows[49])) ac49(.scan_win(scan_win49), .scan_win_std_dev(scan_win_std_dev[49]), .feature_accum(feature_accums[49]));
  accum_calculator #(.RECT1_X(rectangle1_xs[50]), .RECT1_Y(rectangle1_ys[50]), .RECT1_WIDTH(rectangle1_widths[50]), .RECT1_HEIGHT(rectangle1_heights[50]), .RECT1_WEIGHT(rectangle1_weights[50]), .RECT2_X(rectangle2_xs[50]), .RECT2_Y(rectangle2_ys[50]), .RECT2_WIDTH(rectangle2_widths[50]), .RECT2_HEIGHT(rectangle2_heights[50]), .RECT2_WEIGHT(rectangle2_weights[50]), .RECT3_X(rectangle3_xs[50]), .RECT3_Y(rectangle3_ys[50]), .RECT3_WIDTH(rectangle3_widths[50]), .RECT3_HEIGHT(rectangle3_heights[50]), .RECT3_WEIGHT(rectangle3_weights[50]), .FEAT_THRES(feature_thresholds[50]), .FEAT_ABOVE(feature_aboves[50]), .FEAT_BELOW(feature_belows[50])) ac50(.scan_win(scan_win50), .scan_win_std_dev(scan_win_std_dev[50]), .feature_accum(feature_accums[50]));
  accum_calculator #(.RECT1_X(rectangle1_xs[51]), .RECT1_Y(rectangle1_ys[51]), .RECT1_WIDTH(rectangle1_widths[51]), .RECT1_HEIGHT(rectangle1_heights[51]), .RECT1_WEIGHT(rectangle1_weights[51]), .RECT2_X(rectangle2_xs[51]), .RECT2_Y(rectangle2_ys[51]), .RECT2_WIDTH(rectangle2_widths[51]), .RECT2_HEIGHT(rectangle2_heights[51]), .RECT2_WEIGHT(rectangle2_weights[51]), .RECT3_X(rectangle3_xs[51]), .RECT3_Y(rectangle3_ys[51]), .RECT3_WIDTH(rectangle3_widths[51]), .RECT3_HEIGHT(rectangle3_heights[51]), .RECT3_WEIGHT(rectangle3_weights[51]), .FEAT_THRES(feature_thresholds[51]), .FEAT_ABOVE(feature_aboves[51]), .FEAT_BELOW(feature_belows[51])) ac51(.scan_win(scan_win51), .scan_win_std_dev(scan_win_std_dev[51]), .feature_accum(feature_accums[51]));
  accum_calculator #(.RECT1_X(rectangle1_xs[52]), .RECT1_Y(rectangle1_ys[52]), .RECT1_WIDTH(rectangle1_widths[52]), .RECT1_HEIGHT(rectangle1_heights[52]), .RECT1_WEIGHT(rectangle1_weights[52]), .RECT2_X(rectangle2_xs[52]), .RECT2_Y(rectangle2_ys[52]), .RECT2_WIDTH(rectangle2_widths[52]), .RECT2_HEIGHT(rectangle2_heights[52]), .RECT2_WEIGHT(rectangle2_weights[52]), .RECT3_X(rectangle3_xs[52]), .RECT3_Y(rectangle3_ys[52]), .RECT3_WIDTH(rectangle3_widths[52]), .RECT3_HEIGHT(rectangle3_heights[52]), .RECT3_WEIGHT(rectangle3_weights[52]), .FEAT_THRES(feature_thresholds[52]), .FEAT_ABOVE(feature_aboves[52]), .FEAT_BELOW(feature_belows[52])) ac52(.scan_win(scan_win52), .scan_win_std_dev(scan_win_std_dev[52]), .feature_accum(feature_accums[52]));
  accum_calculator #(.RECT1_X(rectangle1_xs[53]), .RECT1_Y(rectangle1_ys[53]), .RECT1_WIDTH(rectangle1_widths[53]), .RECT1_HEIGHT(rectangle1_heights[53]), .RECT1_WEIGHT(rectangle1_weights[53]), .RECT2_X(rectangle2_xs[53]), .RECT2_Y(rectangle2_ys[53]), .RECT2_WIDTH(rectangle2_widths[53]), .RECT2_HEIGHT(rectangle2_heights[53]), .RECT2_WEIGHT(rectangle2_weights[53]), .RECT3_X(rectangle3_xs[53]), .RECT3_Y(rectangle3_ys[53]), .RECT3_WIDTH(rectangle3_widths[53]), .RECT3_HEIGHT(rectangle3_heights[53]), .RECT3_WEIGHT(rectangle3_weights[53]), .FEAT_THRES(feature_thresholds[53]), .FEAT_ABOVE(feature_aboves[53]), .FEAT_BELOW(feature_belows[53])) ac53(.scan_win(scan_win53), .scan_win_std_dev(scan_win_std_dev[53]), .feature_accum(feature_accums[53]));
  accum_calculator #(.RECT1_X(rectangle1_xs[54]), .RECT1_Y(rectangle1_ys[54]), .RECT1_WIDTH(rectangle1_widths[54]), .RECT1_HEIGHT(rectangle1_heights[54]), .RECT1_WEIGHT(rectangle1_weights[54]), .RECT2_X(rectangle2_xs[54]), .RECT2_Y(rectangle2_ys[54]), .RECT2_WIDTH(rectangle2_widths[54]), .RECT2_HEIGHT(rectangle2_heights[54]), .RECT2_WEIGHT(rectangle2_weights[54]), .RECT3_X(rectangle3_xs[54]), .RECT3_Y(rectangle3_ys[54]), .RECT3_WIDTH(rectangle3_widths[54]), .RECT3_HEIGHT(rectangle3_heights[54]), .RECT3_WEIGHT(rectangle3_weights[54]), .FEAT_THRES(feature_thresholds[54]), .FEAT_ABOVE(feature_aboves[54]), .FEAT_BELOW(feature_belows[54])) ac54(.scan_win(scan_win54), .scan_win_std_dev(scan_win_std_dev[54]), .feature_accum(feature_accums[54]));
  accum_calculator #(.RECT1_X(rectangle1_xs[55]), .RECT1_Y(rectangle1_ys[55]), .RECT1_WIDTH(rectangle1_widths[55]), .RECT1_HEIGHT(rectangle1_heights[55]), .RECT1_WEIGHT(rectangle1_weights[55]), .RECT2_X(rectangle2_xs[55]), .RECT2_Y(rectangle2_ys[55]), .RECT2_WIDTH(rectangle2_widths[55]), .RECT2_HEIGHT(rectangle2_heights[55]), .RECT2_WEIGHT(rectangle2_weights[55]), .RECT3_X(rectangle3_xs[55]), .RECT3_Y(rectangle3_ys[55]), .RECT3_WIDTH(rectangle3_widths[55]), .RECT3_HEIGHT(rectangle3_heights[55]), .RECT3_WEIGHT(rectangle3_weights[55]), .FEAT_THRES(feature_thresholds[55]), .FEAT_ABOVE(feature_aboves[55]), .FEAT_BELOW(feature_belows[55])) ac55(.scan_win(scan_win55), .scan_win_std_dev(scan_win_std_dev[55]), .feature_accum(feature_accums[55]));
  accum_calculator #(.RECT1_X(rectangle1_xs[56]), .RECT1_Y(rectangle1_ys[56]), .RECT1_WIDTH(rectangle1_widths[56]), .RECT1_HEIGHT(rectangle1_heights[56]), .RECT1_WEIGHT(rectangle1_weights[56]), .RECT2_X(rectangle2_xs[56]), .RECT2_Y(rectangle2_ys[56]), .RECT2_WIDTH(rectangle2_widths[56]), .RECT2_HEIGHT(rectangle2_heights[56]), .RECT2_WEIGHT(rectangle2_weights[56]), .RECT3_X(rectangle3_xs[56]), .RECT3_Y(rectangle3_ys[56]), .RECT3_WIDTH(rectangle3_widths[56]), .RECT3_HEIGHT(rectangle3_heights[56]), .RECT3_WEIGHT(rectangle3_weights[56]), .FEAT_THRES(feature_thresholds[56]), .FEAT_ABOVE(feature_aboves[56]), .FEAT_BELOW(feature_belows[56])) ac56(.scan_win(scan_win56), .scan_win_std_dev(scan_win_std_dev[56]), .feature_accum(feature_accums[56]));
  accum_calculator #(.RECT1_X(rectangle1_xs[57]), .RECT1_Y(rectangle1_ys[57]), .RECT1_WIDTH(rectangle1_widths[57]), .RECT1_HEIGHT(rectangle1_heights[57]), .RECT1_WEIGHT(rectangle1_weights[57]), .RECT2_X(rectangle2_xs[57]), .RECT2_Y(rectangle2_ys[57]), .RECT2_WIDTH(rectangle2_widths[57]), .RECT2_HEIGHT(rectangle2_heights[57]), .RECT2_WEIGHT(rectangle2_weights[57]), .RECT3_X(rectangle3_xs[57]), .RECT3_Y(rectangle3_ys[57]), .RECT3_WIDTH(rectangle3_widths[57]), .RECT3_HEIGHT(rectangle3_heights[57]), .RECT3_WEIGHT(rectangle3_weights[57]), .FEAT_THRES(feature_thresholds[57]), .FEAT_ABOVE(feature_aboves[57]), .FEAT_BELOW(feature_belows[57])) ac57(.scan_win(scan_win57), .scan_win_std_dev(scan_win_std_dev[57]), .feature_accum(feature_accums[57]));
  accum_calculator #(.RECT1_X(rectangle1_xs[58]), .RECT1_Y(rectangle1_ys[58]), .RECT1_WIDTH(rectangle1_widths[58]), .RECT1_HEIGHT(rectangle1_heights[58]), .RECT1_WEIGHT(rectangle1_weights[58]), .RECT2_X(rectangle2_xs[58]), .RECT2_Y(rectangle2_ys[58]), .RECT2_WIDTH(rectangle2_widths[58]), .RECT2_HEIGHT(rectangle2_heights[58]), .RECT2_WEIGHT(rectangle2_weights[58]), .RECT3_X(rectangle3_xs[58]), .RECT3_Y(rectangle3_ys[58]), .RECT3_WIDTH(rectangle3_widths[58]), .RECT3_HEIGHT(rectangle3_heights[58]), .RECT3_WEIGHT(rectangle3_weights[58]), .FEAT_THRES(feature_thresholds[58]), .FEAT_ABOVE(feature_aboves[58]), .FEAT_BELOW(feature_belows[58])) ac58(.scan_win(scan_win58), .scan_win_std_dev(scan_win_std_dev[58]), .feature_accum(feature_accums[58]));
  accum_calculator #(.RECT1_X(rectangle1_xs[59]), .RECT1_Y(rectangle1_ys[59]), .RECT1_WIDTH(rectangle1_widths[59]), .RECT1_HEIGHT(rectangle1_heights[59]), .RECT1_WEIGHT(rectangle1_weights[59]), .RECT2_X(rectangle2_xs[59]), .RECT2_Y(rectangle2_ys[59]), .RECT2_WIDTH(rectangle2_widths[59]), .RECT2_HEIGHT(rectangle2_heights[59]), .RECT2_WEIGHT(rectangle2_weights[59]), .RECT3_X(rectangle3_xs[59]), .RECT3_Y(rectangle3_ys[59]), .RECT3_WIDTH(rectangle3_widths[59]), .RECT3_HEIGHT(rectangle3_heights[59]), .RECT3_WEIGHT(rectangle3_weights[59]), .FEAT_THRES(feature_thresholds[59]), .FEAT_ABOVE(feature_aboves[59]), .FEAT_BELOW(feature_belows[59])) ac59(.scan_win(scan_win59), .scan_win_std_dev(scan_win_std_dev[59]), .feature_accum(feature_accums[59]));
  accum_calculator #(.RECT1_X(rectangle1_xs[60]), .RECT1_Y(rectangle1_ys[60]), .RECT1_WIDTH(rectangle1_widths[60]), .RECT1_HEIGHT(rectangle1_heights[60]), .RECT1_WEIGHT(rectangle1_weights[60]), .RECT2_X(rectangle2_xs[60]), .RECT2_Y(rectangle2_ys[60]), .RECT2_WIDTH(rectangle2_widths[60]), .RECT2_HEIGHT(rectangle2_heights[60]), .RECT2_WEIGHT(rectangle2_weights[60]), .RECT3_X(rectangle3_xs[60]), .RECT3_Y(rectangle3_ys[60]), .RECT3_WIDTH(rectangle3_widths[60]), .RECT3_HEIGHT(rectangle3_heights[60]), .RECT3_WEIGHT(rectangle3_weights[60]), .FEAT_THRES(feature_thresholds[60]), .FEAT_ABOVE(feature_aboves[60]), .FEAT_BELOW(feature_belows[60])) ac60(.scan_win(scan_win60), .scan_win_std_dev(scan_win_std_dev[60]), .feature_accum(feature_accums[60]));
  accum_calculator #(.RECT1_X(rectangle1_xs[61]), .RECT1_Y(rectangle1_ys[61]), .RECT1_WIDTH(rectangle1_widths[61]), .RECT1_HEIGHT(rectangle1_heights[61]), .RECT1_WEIGHT(rectangle1_weights[61]), .RECT2_X(rectangle2_xs[61]), .RECT2_Y(rectangle2_ys[61]), .RECT2_WIDTH(rectangle2_widths[61]), .RECT2_HEIGHT(rectangle2_heights[61]), .RECT2_WEIGHT(rectangle2_weights[61]), .RECT3_X(rectangle3_xs[61]), .RECT3_Y(rectangle3_ys[61]), .RECT3_WIDTH(rectangle3_widths[61]), .RECT3_HEIGHT(rectangle3_heights[61]), .RECT3_WEIGHT(rectangle3_weights[61]), .FEAT_THRES(feature_thresholds[61]), .FEAT_ABOVE(feature_aboves[61]), .FEAT_BELOW(feature_belows[61])) ac61(.scan_win(scan_win61), .scan_win_std_dev(scan_win_std_dev[61]), .feature_accum(feature_accums[61]));
  accum_calculator #(.RECT1_X(rectangle1_xs[62]), .RECT1_Y(rectangle1_ys[62]), .RECT1_WIDTH(rectangle1_widths[62]), .RECT1_HEIGHT(rectangle1_heights[62]), .RECT1_WEIGHT(rectangle1_weights[62]), .RECT2_X(rectangle2_xs[62]), .RECT2_Y(rectangle2_ys[62]), .RECT2_WIDTH(rectangle2_widths[62]), .RECT2_HEIGHT(rectangle2_heights[62]), .RECT2_WEIGHT(rectangle2_weights[62]), .RECT3_X(rectangle3_xs[62]), .RECT3_Y(rectangle3_ys[62]), .RECT3_WIDTH(rectangle3_widths[62]), .RECT3_HEIGHT(rectangle3_heights[62]), .RECT3_WEIGHT(rectangle3_weights[62]), .FEAT_THRES(feature_thresholds[62]), .FEAT_ABOVE(feature_aboves[62]), .FEAT_BELOW(feature_belows[62])) ac62(.scan_win(scan_win62), .scan_win_std_dev(scan_win_std_dev[62]), .feature_accum(feature_accums[62]));
  accum_calculator #(.RECT1_X(rectangle1_xs[63]), .RECT1_Y(rectangle1_ys[63]), .RECT1_WIDTH(rectangle1_widths[63]), .RECT1_HEIGHT(rectangle1_heights[63]), .RECT1_WEIGHT(rectangle1_weights[63]), .RECT2_X(rectangle2_xs[63]), .RECT2_Y(rectangle2_ys[63]), .RECT2_WIDTH(rectangle2_widths[63]), .RECT2_HEIGHT(rectangle2_heights[63]), .RECT2_WEIGHT(rectangle2_weights[63]), .RECT3_X(rectangle3_xs[63]), .RECT3_Y(rectangle3_ys[63]), .RECT3_WIDTH(rectangle3_widths[63]), .RECT3_HEIGHT(rectangle3_heights[63]), .RECT3_WEIGHT(rectangle3_weights[63]), .FEAT_THRES(feature_thresholds[63]), .FEAT_ABOVE(feature_aboves[63]), .FEAT_BELOW(feature_belows[63])) ac63(.scan_win(scan_win63), .scan_win_std_dev(scan_win_std_dev[63]), .feature_accum(feature_accums[63]));
  accum_calculator #(.RECT1_X(rectangle1_xs[64]), .RECT1_Y(rectangle1_ys[64]), .RECT1_WIDTH(rectangle1_widths[64]), .RECT1_HEIGHT(rectangle1_heights[64]), .RECT1_WEIGHT(rectangle1_weights[64]), .RECT2_X(rectangle2_xs[64]), .RECT2_Y(rectangle2_ys[64]), .RECT2_WIDTH(rectangle2_widths[64]), .RECT2_HEIGHT(rectangle2_heights[64]), .RECT2_WEIGHT(rectangle2_weights[64]), .RECT3_X(rectangle3_xs[64]), .RECT3_Y(rectangle3_ys[64]), .RECT3_WIDTH(rectangle3_widths[64]), .RECT3_HEIGHT(rectangle3_heights[64]), .RECT3_WEIGHT(rectangle3_weights[64]), .FEAT_THRES(feature_thresholds[64]), .FEAT_ABOVE(feature_aboves[64]), .FEAT_BELOW(feature_belows[64])) ac64(.scan_win(scan_win64), .scan_win_std_dev(scan_win_std_dev[64]), .feature_accum(feature_accums[64]));
  accum_calculator #(.RECT1_X(rectangle1_xs[65]), .RECT1_Y(rectangle1_ys[65]), .RECT1_WIDTH(rectangle1_widths[65]), .RECT1_HEIGHT(rectangle1_heights[65]), .RECT1_WEIGHT(rectangle1_weights[65]), .RECT2_X(rectangle2_xs[65]), .RECT2_Y(rectangle2_ys[65]), .RECT2_WIDTH(rectangle2_widths[65]), .RECT2_HEIGHT(rectangle2_heights[65]), .RECT2_WEIGHT(rectangle2_weights[65]), .RECT3_X(rectangle3_xs[65]), .RECT3_Y(rectangle3_ys[65]), .RECT3_WIDTH(rectangle3_widths[65]), .RECT3_HEIGHT(rectangle3_heights[65]), .RECT3_WEIGHT(rectangle3_weights[65]), .FEAT_THRES(feature_thresholds[65]), .FEAT_ABOVE(feature_aboves[65]), .FEAT_BELOW(feature_belows[65])) ac65(.scan_win(scan_win65), .scan_win_std_dev(scan_win_std_dev[65]), .feature_accum(feature_accums[65]));
  accum_calculator #(.RECT1_X(rectangle1_xs[66]), .RECT1_Y(rectangle1_ys[66]), .RECT1_WIDTH(rectangle1_widths[66]), .RECT1_HEIGHT(rectangle1_heights[66]), .RECT1_WEIGHT(rectangle1_weights[66]), .RECT2_X(rectangle2_xs[66]), .RECT2_Y(rectangle2_ys[66]), .RECT2_WIDTH(rectangle2_widths[66]), .RECT2_HEIGHT(rectangle2_heights[66]), .RECT2_WEIGHT(rectangle2_weights[66]), .RECT3_X(rectangle3_xs[66]), .RECT3_Y(rectangle3_ys[66]), .RECT3_WIDTH(rectangle3_widths[66]), .RECT3_HEIGHT(rectangle3_heights[66]), .RECT3_WEIGHT(rectangle3_weights[66]), .FEAT_THRES(feature_thresholds[66]), .FEAT_ABOVE(feature_aboves[66]), .FEAT_BELOW(feature_belows[66])) ac66(.scan_win(scan_win66), .scan_win_std_dev(scan_win_std_dev[66]), .feature_accum(feature_accums[66]));
  accum_calculator #(.RECT1_X(rectangle1_xs[67]), .RECT1_Y(rectangle1_ys[67]), .RECT1_WIDTH(rectangle1_widths[67]), .RECT1_HEIGHT(rectangle1_heights[67]), .RECT1_WEIGHT(rectangle1_weights[67]), .RECT2_X(rectangle2_xs[67]), .RECT2_Y(rectangle2_ys[67]), .RECT2_WIDTH(rectangle2_widths[67]), .RECT2_HEIGHT(rectangle2_heights[67]), .RECT2_WEIGHT(rectangle2_weights[67]), .RECT3_X(rectangle3_xs[67]), .RECT3_Y(rectangle3_ys[67]), .RECT3_WIDTH(rectangle3_widths[67]), .RECT3_HEIGHT(rectangle3_heights[67]), .RECT3_WEIGHT(rectangle3_weights[67]), .FEAT_THRES(feature_thresholds[67]), .FEAT_ABOVE(feature_aboves[67]), .FEAT_BELOW(feature_belows[67])) ac67(.scan_win(scan_win67), .scan_win_std_dev(scan_win_std_dev[67]), .feature_accum(feature_accums[67]));
  accum_calculator #(.RECT1_X(rectangle1_xs[68]), .RECT1_Y(rectangle1_ys[68]), .RECT1_WIDTH(rectangle1_widths[68]), .RECT1_HEIGHT(rectangle1_heights[68]), .RECT1_WEIGHT(rectangle1_weights[68]), .RECT2_X(rectangle2_xs[68]), .RECT2_Y(rectangle2_ys[68]), .RECT2_WIDTH(rectangle2_widths[68]), .RECT2_HEIGHT(rectangle2_heights[68]), .RECT2_WEIGHT(rectangle2_weights[68]), .RECT3_X(rectangle3_xs[68]), .RECT3_Y(rectangle3_ys[68]), .RECT3_WIDTH(rectangle3_widths[68]), .RECT3_HEIGHT(rectangle3_heights[68]), .RECT3_WEIGHT(rectangle3_weights[68]), .FEAT_THRES(feature_thresholds[68]), .FEAT_ABOVE(feature_aboves[68]), .FEAT_BELOW(feature_belows[68])) ac68(.scan_win(scan_win68), .scan_win_std_dev(scan_win_std_dev[68]), .feature_accum(feature_accums[68]));
  accum_calculator #(.RECT1_X(rectangle1_xs[69]), .RECT1_Y(rectangle1_ys[69]), .RECT1_WIDTH(rectangle1_widths[69]), .RECT1_HEIGHT(rectangle1_heights[69]), .RECT1_WEIGHT(rectangle1_weights[69]), .RECT2_X(rectangle2_xs[69]), .RECT2_Y(rectangle2_ys[69]), .RECT2_WIDTH(rectangle2_widths[69]), .RECT2_HEIGHT(rectangle2_heights[69]), .RECT2_WEIGHT(rectangle2_weights[69]), .RECT3_X(rectangle3_xs[69]), .RECT3_Y(rectangle3_ys[69]), .RECT3_WIDTH(rectangle3_widths[69]), .RECT3_HEIGHT(rectangle3_heights[69]), .RECT3_WEIGHT(rectangle3_weights[69]), .FEAT_THRES(feature_thresholds[69]), .FEAT_ABOVE(feature_aboves[69]), .FEAT_BELOW(feature_belows[69])) ac69(.scan_win(scan_win69), .scan_win_std_dev(scan_win_std_dev[69]), .feature_accum(feature_accums[69]));
  accum_calculator #(.RECT1_X(rectangle1_xs[70]), .RECT1_Y(rectangle1_ys[70]), .RECT1_WIDTH(rectangle1_widths[70]), .RECT1_HEIGHT(rectangle1_heights[70]), .RECT1_WEIGHT(rectangle1_weights[70]), .RECT2_X(rectangle2_xs[70]), .RECT2_Y(rectangle2_ys[70]), .RECT2_WIDTH(rectangle2_widths[70]), .RECT2_HEIGHT(rectangle2_heights[70]), .RECT2_WEIGHT(rectangle2_weights[70]), .RECT3_X(rectangle3_xs[70]), .RECT3_Y(rectangle3_ys[70]), .RECT3_WIDTH(rectangle3_widths[70]), .RECT3_HEIGHT(rectangle3_heights[70]), .RECT3_WEIGHT(rectangle3_weights[70]), .FEAT_THRES(feature_thresholds[70]), .FEAT_ABOVE(feature_aboves[70]), .FEAT_BELOW(feature_belows[70])) ac70(.scan_win(scan_win70), .scan_win_std_dev(scan_win_std_dev[70]), .feature_accum(feature_accums[70]));
  accum_calculator #(.RECT1_X(rectangle1_xs[71]), .RECT1_Y(rectangle1_ys[71]), .RECT1_WIDTH(rectangle1_widths[71]), .RECT1_HEIGHT(rectangle1_heights[71]), .RECT1_WEIGHT(rectangle1_weights[71]), .RECT2_X(rectangle2_xs[71]), .RECT2_Y(rectangle2_ys[71]), .RECT2_WIDTH(rectangle2_widths[71]), .RECT2_HEIGHT(rectangle2_heights[71]), .RECT2_WEIGHT(rectangle2_weights[71]), .RECT3_X(rectangle3_xs[71]), .RECT3_Y(rectangle3_ys[71]), .RECT3_WIDTH(rectangle3_widths[71]), .RECT3_HEIGHT(rectangle3_heights[71]), .RECT3_WEIGHT(rectangle3_weights[71]), .FEAT_THRES(feature_thresholds[71]), .FEAT_ABOVE(feature_aboves[71]), .FEAT_BELOW(feature_belows[71])) ac71(.scan_win(scan_win71), .scan_win_std_dev(scan_win_std_dev[71]), .feature_accum(feature_accums[71]));
  accum_calculator #(.RECT1_X(rectangle1_xs[72]), .RECT1_Y(rectangle1_ys[72]), .RECT1_WIDTH(rectangle1_widths[72]), .RECT1_HEIGHT(rectangle1_heights[72]), .RECT1_WEIGHT(rectangle1_weights[72]), .RECT2_X(rectangle2_xs[72]), .RECT2_Y(rectangle2_ys[72]), .RECT2_WIDTH(rectangle2_widths[72]), .RECT2_HEIGHT(rectangle2_heights[72]), .RECT2_WEIGHT(rectangle2_weights[72]), .RECT3_X(rectangle3_xs[72]), .RECT3_Y(rectangle3_ys[72]), .RECT3_WIDTH(rectangle3_widths[72]), .RECT3_HEIGHT(rectangle3_heights[72]), .RECT3_WEIGHT(rectangle3_weights[72]), .FEAT_THRES(feature_thresholds[72]), .FEAT_ABOVE(feature_aboves[72]), .FEAT_BELOW(feature_belows[72])) ac72(.scan_win(scan_win72), .scan_win_std_dev(scan_win_std_dev[72]), .feature_accum(feature_accums[72]));
  accum_calculator #(.RECT1_X(rectangle1_xs[73]), .RECT1_Y(rectangle1_ys[73]), .RECT1_WIDTH(rectangle1_widths[73]), .RECT1_HEIGHT(rectangle1_heights[73]), .RECT1_WEIGHT(rectangle1_weights[73]), .RECT2_X(rectangle2_xs[73]), .RECT2_Y(rectangle2_ys[73]), .RECT2_WIDTH(rectangle2_widths[73]), .RECT2_HEIGHT(rectangle2_heights[73]), .RECT2_WEIGHT(rectangle2_weights[73]), .RECT3_X(rectangle3_xs[73]), .RECT3_Y(rectangle3_ys[73]), .RECT3_WIDTH(rectangle3_widths[73]), .RECT3_HEIGHT(rectangle3_heights[73]), .RECT3_WEIGHT(rectangle3_weights[73]), .FEAT_THRES(feature_thresholds[73]), .FEAT_ABOVE(feature_aboves[73]), .FEAT_BELOW(feature_belows[73])) ac73(.scan_win(scan_win73), .scan_win_std_dev(scan_win_std_dev[73]), .feature_accum(feature_accums[73]));
  accum_calculator #(.RECT1_X(rectangle1_xs[74]), .RECT1_Y(rectangle1_ys[74]), .RECT1_WIDTH(rectangle1_widths[74]), .RECT1_HEIGHT(rectangle1_heights[74]), .RECT1_WEIGHT(rectangle1_weights[74]), .RECT2_X(rectangle2_xs[74]), .RECT2_Y(rectangle2_ys[74]), .RECT2_WIDTH(rectangle2_widths[74]), .RECT2_HEIGHT(rectangle2_heights[74]), .RECT2_WEIGHT(rectangle2_weights[74]), .RECT3_X(rectangle3_xs[74]), .RECT3_Y(rectangle3_ys[74]), .RECT3_WIDTH(rectangle3_widths[74]), .RECT3_HEIGHT(rectangle3_heights[74]), .RECT3_WEIGHT(rectangle3_weights[74]), .FEAT_THRES(feature_thresholds[74]), .FEAT_ABOVE(feature_aboves[74]), .FEAT_BELOW(feature_belows[74])) ac74(.scan_win(scan_win74), .scan_win_std_dev(scan_win_std_dev[74]), .feature_accum(feature_accums[74]));
  accum_calculator #(.RECT1_X(rectangle1_xs[75]), .RECT1_Y(rectangle1_ys[75]), .RECT1_WIDTH(rectangle1_widths[75]), .RECT1_HEIGHT(rectangle1_heights[75]), .RECT1_WEIGHT(rectangle1_weights[75]), .RECT2_X(rectangle2_xs[75]), .RECT2_Y(rectangle2_ys[75]), .RECT2_WIDTH(rectangle2_widths[75]), .RECT2_HEIGHT(rectangle2_heights[75]), .RECT2_WEIGHT(rectangle2_weights[75]), .RECT3_X(rectangle3_xs[75]), .RECT3_Y(rectangle3_ys[75]), .RECT3_WIDTH(rectangle3_widths[75]), .RECT3_HEIGHT(rectangle3_heights[75]), .RECT3_WEIGHT(rectangle3_weights[75]), .FEAT_THRES(feature_thresholds[75]), .FEAT_ABOVE(feature_aboves[75]), .FEAT_BELOW(feature_belows[75])) ac75(.scan_win(scan_win75), .scan_win_std_dev(scan_win_std_dev[75]), .feature_accum(feature_accums[75]));
  accum_calculator #(.RECT1_X(rectangle1_xs[76]), .RECT1_Y(rectangle1_ys[76]), .RECT1_WIDTH(rectangle1_widths[76]), .RECT1_HEIGHT(rectangle1_heights[76]), .RECT1_WEIGHT(rectangle1_weights[76]), .RECT2_X(rectangle2_xs[76]), .RECT2_Y(rectangle2_ys[76]), .RECT2_WIDTH(rectangle2_widths[76]), .RECT2_HEIGHT(rectangle2_heights[76]), .RECT2_WEIGHT(rectangle2_weights[76]), .RECT3_X(rectangle3_xs[76]), .RECT3_Y(rectangle3_ys[76]), .RECT3_WIDTH(rectangle3_widths[76]), .RECT3_HEIGHT(rectangle3_heights[76]), .RECT3_WEIGHT(rectangle3_weights[76]), .FEAT_THRES(feature_thresholds[76]), .FEAT_ABOVE(feature_aboves[76]), .FEAT_BELOW(feature_belows[76])) ac76(.scan_win(scan_win76), .scan_win_std_dev(scan_win_std_dev[76]), .feature_accum(feature_accums[76]));
  accum_calculator #(.RECT1_X(rectangle1_xs[77]), .RECT1_Y(rectangle1_ys[77]), .RECT1_WIDTH(rectangle1_widths[77]), .RECT1_HEIGHT(rectangle1_heights[77]), .RECT1_WEIGHT(rectangle1_weights[77]), .RECT2_X(rectangle2_xs[77]), .RECT2_Y(rectangle2_ys[77]), .RECT2_WIDTH(rectangle2_widths[77]), .RECT2_HEIGHT(rectangle2_heights[77]), .RECT2_WEIGHT(rectangle2_weights[77]), .RECT3_X(rectangle3_xs[77]), .RECT3_Y(rectangle3_ys[77]), .RECT3_WIDTH(rectangle3_widths[77]), .RECT3_HEIGHT(rectangle3_heights[77]), .RECT3_WEIGHT(rectangle3_weights[77]), .FEAT_THRES(feature_thresholds[77]), .FEAT_ABOVE(feature_aboves[77]), .FEAT_BELOW(feature_belows[77])) ac77(.scan_win(scan_win77), .scan_win_std_dev(scan_win_std_dev[77]), .feature_accum(feature_accums[77]));
  accum_calculator #(.RECT1_X(rectangle1_xs[78]), .RECT1_Y(rectangle1_ys[78]), .RECT1_WIDTH(rectangle1_widths[78]), .RECT1_HEIGHT(rectangle1_heights[78]), .RECT1_WEIGHT(rectangle1_weights[78]), .RECT2_X(rectangle2_xs[78]), .RECT2_Y(rectangle2_ys[78]), .RECT2_WIDTH(rectangle2_widths[78]), .RECT2_HEIGHT(rectangle2_heights[78]), .RECT2_WEIGHT(rectangle2_weights[78]), .RECT3_X(rectangle3_xs[78]), .RECT3_Y(rectangle3_ys[78]), .RECT3_WIDTH(rectangle3_widths[78]), .RECT3_HEIGHT(rectangle3_heights[78]), .RECT3_WEIGHT(rectangle3_weights[78]), .FEAT_THRES(feature_thresholds[78]), .FEAT_ABOVE(feature_aboves[78]), .FEAT_BELOW(feature_belows[78])) ac78(.scan_win(scan_win78), .scan_win_std_dev(scan_win_std_dev[78]), .feature_accum(feature_accums[78]));
  accum_calculator #(.RECT1_X(rectangle1_xs[79]), .RECT1_Y(rectangle1_ys[79]), .RECT1_WIDTH(rectangle1_widths[79]), .RECT1_HEIGHT(rectangle1_heights[79]), .RECT1_WEIGHT(rectangle1_weights[79]), .RECT2_X(rectangle2_xs[79]), .RECT2_Y(rectangle2_ys[79]), .RECT2_WIDTH(rectangle2_widths[79]), .RECT2_HEIGHT(rectangle2_heights[79]), .RECT2_WEIGHT(rectangle2_weights[79]), .RECT3_X(rectangle3_xs[79]), .RECT3_Y(rectangle3_ys[79]), .RECT3_WIDTH(rectangle3_widths[79]), .RECT3_HEIGHT(rectangle3_heights[79]), .RECT3_WEIGHT(rectangle3_weights[79]), .FEAT_THRES(feature_thresholds[79]), .FEAT_ABOVE(feature_aboves[79]), .FEAT_BELOW(feature_belows[79])) ac79(.scan_win(scan_win79), .scan_win_std_dev(scan_win_std_dev[79]), .feature_accum(feature_accums[79]));
  accum_calculator #(.RECT1_X(rectangle1_xs[80]), .RECT1_Y(rectangle1_ys[80]), .RECT1_WIDTH(rectangle1_widths[80]), .RECT1_HEIGHT(rectangle1_heights[80]), .RECT1_WEIGHT(rectangle1_weights[80]), .RECT2_X(rectangle2_xs[80]), .RECT2_Y(rectangle2_ys[80]), .RECT2_WIDTH(rectangle2_widths[80]), .RECT2_HEIGHT(rectangle2_heights[80]), .RECT2_WEIGHT(rectangle2_weights[80]), .RECT3_X(rectangle3_xs[80]), .RECT3_Y(rectangle3_ys[80]), .RECT3_WIDTH(rectangle3_widths[80]), .RECT3_HEIGHT(rectangle3_heights[80]), .RECT3_WEIGHT(rectangle3_weights[80]), .FEAT_THRES(feature_thresholds[80]), .FEAT_ABOVE(feature_aboves[80]), .FEAT_BELOW(feature_belows[80])) ac80(.scan_win(scan_win80), .scan_win_std_dev(scan_win_std_dev[80]), .feature_accum(feature_accums[80]));
  accum_calculator #(.RECT1_X(rectangle1_xs[81]), .RECT1_Y(rectangle1_ys[81]), .RECT1_WIDTH(rectangle1_widths[81]), .RECT1_HEIGHT(rectangle1_heights[81]), .RECT1_WEIGHT(rectangle1_weights[81]), .RECT2_X(rectangle2_xs[81]), .RECT2_Y(rectangle2_ys[81]), .RECT2_WIDTH(rectangle2_widths[81]), .RECT2_HEIGHT(rectangle2_heights[81]), .RECT2_WEIGHT(rectangle2_weights[81]), .RECT3_X(rectangle3_xs[81]), .RECT3_Y(rectangle3_ys[81]), .RECT3_WIDTH(rectangle3_widths[81]), .RECT3_HEIGHT(rectangle3_heights[81]), .RECT3_WEIGHT(rectangle3_weights[81]), .FEAT_THRES(feature_thresholds[81]), .FEAT_ABOVE(feature_aboves[81]), .FEAT_BELOW(feature_belows[81])) ac81(.scan_win(scan_win81), .scan_win_std_dev(scan_win_std_dev[81]), .feature_accum(feature_accums[81]));
  accum_calculator #(.RECT1_X(rectangle1_xs[82]), .RECT1_Y(rectangle1_ys[82]), .RECT1_WIDTH(rectangle1_widths[82]), .RECT1_HEIGHT(rectangle1_heights[82]), .RECT1_WEIGHT(rectangle1_weights[82]), .RECT2_X(rectangle2_xs[82]), .RECT2_Y(rectangle2_ys[82]), .RECT2_WIDTH(rectangle2_widths[82]), .RECT2_HEIGHT(rectangle2_heights[82]), .RECT2_WEIGHT(rectangle2_weights[82]), .RECT3_X(rectangle3_xs[82]), .RECT3_Y(rectangle3_ys[82]), .RECT3_WIDTH(rectangle3_widths[82]), .RECT3_HEIGHT(rectangle3_heights[82]), .RECT3_WEIGHT(rectangle3_weights[82]), .FEAT_THRES(feature_thresholds[82]), .FEAT_ABOVE(feature_aboves[82]), .FEAT_BELOW(feature_belows[82])) ac82(.scan_win(scan_win82), .scan_win_std_dev(scan_win_std_dev[82]), .feature_accum(feature_accums[82]));
  accum_calculator #(.RECT1_X(rectangle1_xs[83]), .RECT1_Y(rectangle1_ys[83]), .RECT1_WIDTH(rectangle1_widths[83]), .RECT1_HEIGHT(rectangle1_heights[83]), .RECT1_WEIGHT(rectangle1_weights[83]), .RECT2_X(rectangle2_xs[83]), .RECT2_Y(rectangle2_ys[83]), .RECT2_WIDTH(rectangle2_widths[83]), .RECT2_HEIGHT(rectangle2_heights[83]), .RECT2_WEIGHT(rectangle2_weights[83]), .RECT3_X(rectangle3_xs[83]), .RECT3_Y(rectangle3_ys[83]), .RECT3_WIDTH(rectangle3_widths[83]), .RECT3_HEIGHT(rectangle3_heights[83]), .RECT3_WEIGHT(rectangle3_weights[83]), .FEAT_THRES(feature_thresholds[83]), .FEAT_ABOVE(feature_aboves[83]), .FEAT_BELOW(feature_belows[83])) ac83(.scan_win(scan_win83), .scan_win_std_dev(scan_win_std_dev[83]), .feature_accum(feature_accums[83]));
  accum_calculator #(.RECT1_X(rectangle1_xs[84]), .RECT1_Y(rectangle1_ys[84]), .RECT1_WIDTH(rectangle1_widths[84]), .RECT1_HEIGHT(rectangle1_heights[84]), .RECT1_WEIGHT(rectangle1_weights[84]), .RECT2_X(rectangle2_xs[84]), .RECT2_Y(rectangle2_ys[84]), .RECT2_WIDTH(rectangle2_widths[84]), .RECT2_HEIGHT(rectangle2_heights[84]), .RECT2_WEIGHT(rectangle2_weights[84]), .RECT3_X(rectangle3_xs[84]), .RECT3_Y(rectangle3_ys[84]), .RECT3_WIDTH(rectangle3_widths[84]), .RECT3_HEIGHT(rectangle3_heights[84]), .RECT3_WEIGHT(rectangle3_weights[84]), .FEAT_THRES(feature_thresholds[84]), .FEAT_ABOVE(feature_aboves[84]), .FEAT_BELOW(feature_belows[84])) ac84(.scan_win(scan_win84), .scan_win_std_dev(scan_win_std_dev[84]), .feature_accum(feature_accums[84]));
  accum_calculator #(.RECT1_X(rectangle1_xs[85]), .RECT1_Y(rectangle1_ys[85]), .RECT1_WIDTH(rectangle1_widths[85]), .RECT1_HEIGHT(rectangle1_heights[85]), .RECT1_WEIGHT(rectangle1_weights[85]), .RECT2_X(rectangle2_xs[85]), .RECT2_Y(rectangle2_ys[85]), .RECT2_WIDTH(rectangle2_widths[85]), .RECT2_HEIGHT(rectangle2_heights[85]), .RECT2_WEIGHT(rectangle2_weights[85]), .RECT3_X(rectangle3_xs[85]), .RECT3_Y(rectangle3_ys[85]), .RECT3_WIDTH(rectangle3_widths[85]), .RECT3_HEIGHT(rectangle3_heights[85]), .RECT3_WEIGHT(rectangle3_weights[85]), .FEAT_THRES(feature_thresholds[85]), .FEAT_ABOVE(feature_aboves[85]), .FEAT_BELOW(feature_belows[85])) ac85(.scan_win(scan_win85), .scan_win_std_dev(scan_win_std_dev[85]), .feature_accum(feature_accums[85]));
  accum_calculator #(.RECT1_X(rectangle1_xs[86]), .RECT1_Y(rectangle1_ys[86]), .RECT1_WIDTH(rectangle1_widths[86]), .RECT1_HEIGHT(rectangle1_heights[86]), .RECT1_WEIGHT(rectangle1_weights[86]), .RECT2_X(rectangle2_xs[86]), .RECT2_Y(rectangle2_ys[86]), .RECT2_WIDTH(rectangle2_widths[86]), .RECT2_HEIGHT(rectangle2_heights[86]), .RECT2_WEIGHT(rectangle2_weights[86]), .RECT3_X(rectangle3_xs[86]), .RECT3_Y(rectangle3_ys[86]), .RECT3_WIDTH(rectangle3_widths[86]), .RECT3_HEIGHT(rectangle3_heights[86]), .RECT3_WEIGHT(rectangle3_weights[86]), .FEAT_THRES(feature_thresholds[86]), .FEAT_ABOVE(feature_aboves[86]), .FEAT_BELOW(feature_belows[86])) ac86(.scan_win(scan_win86), .scan_win_std_dev(scan_win_std_dev[86]), .feature_accum(feature_accums[86]));
  accum_calculator #(.RECT1_X(rectangle1_xs[87]), .RECT1_Y(rectangle1_ys[87]), .RECT1_WIDTH(rectangle1_widths[87]), .RECT1_HEIGHT(rectangle1_heights[87]), .RECT1_WEIGHT(rectangle1_weights[87]), .RECT2_X(rectangle2_xs[87]), .RECT2_Y(rectangle2_ys[87]), .RECT2_WIDTH(rectangle2_widths[87]), .RECT2_HEIGHT(rectangle2_heights[87]), .RECT2_WEIGHT(rectangle2_weights[87]), .RECT3_X(rectangle3_xs[87]), .RECT3_Y(rectangle3_ys[87]), .RECT3_WIDTH(rectangle3_widths[87]), .RECT3_HEIGHT(rectangle3_heights[87]), .RECT3_WEIGHT(rectangle3_weights[87]), .FEAT_THRES(feature_thresholds[87]), .FEAT_ABOVE(feature_aboves[87]), .FEAT_BELOW(feature_belows[87])) ac87(.scan_win(scan_win87), .scan_win_std_dev(scan_win_std_dev[87]), .feature_accum(feature_accums[87]));
  accum_calculator #(.RECT1_X(rectangle1_xs[88]), .RECT1_Y(rectangle1_ys[88]), .RECT1_WIDTH(rectangle1_widths[88]), .RECT1_HEIGHT(rectangle1_heights[88]), .RECT1_WEIGHT(rectangle1_weights[88]), .RECT2_X(rectangle2_xs[88]), .RECT2_Y(rectangle2_ys[88]), .RECT2_WIDTH(rectangle2_widths[88]), .RECT2_HEIGHT(rectangle2_heights[88]), .RECT2_WEIGHT(rectangle2_weights[88]), .RECT3_X(rectangle3_xs[88]), .RECT3_Y(rectangle3_ys[88]), .RECT3_WIDTH(rectangle3_widths[88]), .RECT3_HEIGHT(rectangle3_heights[88]), .RECT3_WEIGHT(rectangle3_weights[88]), .FEAT_THRES(feature_thresholds[88]), .FEAT_ABOVE(feature_aboves[88]), .FEAT_BELOW(feature_belows[88])) ac88(.scan_win(scan_win88), .scan_win_std_dev(scan_win_std_dev[88]), .feature_accum(feature_accums[88]));
  accum_calculator #(.RECT1_X(rectangle1_xs[89]), .RECT1_Y(rectangle1_ys[89]), .RECT1_WIDTH(rectangle1_widths[89]), .RECT1_HEIGHT(rectangle1_heights[89]), .RECT1_WEIGHT(rectangle1_weights[89]), .RECT2_X(rectangle2_xs[89]), .RECT2_Y(rectangle2_ys[89]), .RECT2_WIDTH(rectangle2_widths[89]), .RECT2_HEIGHT(rectangle2_heights[89]), .RECT2_WEIGHT(rectangle2_weights[89]), .RECT3_X(rectangle3_xs[89]), .RECT3_Y(rectangle3_ys[89]), .RECT3_WIDTH(rectangle3_widths[89]), .RECT3_HEIGHT(rectangle3_heights[89]), .RECT3_WEIGHT(rectangle3_weights[89]), .FEAT_THRES(feature_thresholds[89]), .FEAT_ABOVE(feature_aboves[89]), .FEAT_BELOW(feature_belows[89])) ac89(.scan_win(scan_win89), .scan_win_std_dev(scan_win_std_dev[89]), .feature_accum(feature_accums[89]));
  accum_calculator #(.RECT1_X(rectangle1_xs[90]), .RECT1_Y(rectangle1_ys[90]), .RECT1_WIDTH(rectangle1_widths[90]), .RECT1_HEIGHT(rectangle1_heights[90]), .RECT1_WEIGHT(rectangle1_weights[90]), .RECT2_X(rectangle2_xs[90]), .RECT2_Y(rectangle2_ys[90]), .RECT2_WIDTH(rectangle2_widths[90]), .RECT2_HEIGHT(rectangle2_heights[90]), .RECT2_WEIGHT(rectangle2_weights[90]), .RECT3_X(rectangle3_xs[90]), .RECT3_Y(rectangle3_ys[90]), .RECT3_WIDTH(rectangle3_widths[90]), .RECT3_HEIGHT(rectangle3_heights[90]), .RECT3_WEIGHT(rectangle3_weights[90]), .FEAT_THRES(feature_thresholds[90]), .FEAT_ABOVE(feature_aboves[90]), .FEAT_BELOW(feature_belows[90])) ac90(.scan_win(scan_win90), .scan_win_std_dev(scan_win_std_dev[90]), .feature_accum(feature_accums[90]));
  accum_calculator #(.RECT1_X(rectangle1_xs[91]), .RECT1_Y(rectangle1_ys[91]), .RECT1_WIDTH(rectangle1_widths[91]), .RECT1_HEIGHT(rectangle1_heights[91]), .RECT1_WEIGHT(rectangle1_weights[91]), .RECT2_X(rectangle2_xs[91]), .RECT2_Y(rectangle2_ys[91]), .RECT2_WIDTH(rectangle2_widths[91]), .RECT2_HEIGHT(rectangle2_heights[91]), .RECT2_WEIGHT(rectangle2_weights[91]), .RECT3_X(rectangle3_xs[91]), .RECT3_Y(rectangle3_ys[91]), .RECT3_WIDTH(rectangle3_widths[91]), .RECT3_HEIGHT(rectangle3_heights[91]), .RECT3_WEIGHT(rectangle3_weights[91]), .FEAT_THRES(feature_thresholds[91]), .FEAT_ABOVE(feature_aboves[91]), .FEAT_BELOW(feature_belows[91])) ac91(.scan_win(scan_win91), .scan_win_std_dev(scan_win_std_dev[91]), .feature_accum(feature_accums[91]));
  accum_calculator #(.RECT1_X(rectangle1_xs[92]), .RECT1_Y(rectangle1_ys[92]), .RECT1_WIDTH(rectangle1_widths[92]), .RECT1_HEIGHT(rectangle1_heights[92]), .RECT1_WEIGHT(rectangle1_weights[92]), .RECT2_X(rectangle2_xs[92]), .RECT2_Y(rectangle2_ys[92]), .RECT2_WIDTH(rectangle2_widths[92]), .RECT2_HEIGHT(rectangle2_heights[92]), .RECT2_WEIGHT(rectangle2_weights[92]), .RECT3_X(rectangle3_xs[92]), .RECT3_Y(rectangle3_ys[92]), .RECT3_WIDTH(rectangle3_widths[92]), .RECT3_HEIGHT(rectangle3_heights[92]), .RECT3_WEIGHT(rectangle3_weights[92]), .FEAT_THRES(feature_thresholds[92]), .FEAT_ABOVE(feature_aboves[92]), .FEAT_BELOW(feature_belows[92])) ac92(.scan_win(scan_win92), .scan_win_std_dev(scan_win_std_dev[92]), .feature_accum(feature_accums[92]));
  accum_calculator #(.RECT1_X(rectangle1_xs[93]), .RECT1_Y(rectangle1_ys[93]), .RECT1_WIDTH(rectangle1_widths[93]), .RECT1_HEIGHT(rectangle1_heights[93]), .RECT1_WEIGHT(rectangle1_weights[93]), .RECT2_X(rectangle2_xs[93]), .RECT2_Y(rectangle2_ys[93]), .RECT2_WIDTH(rectangle2_widths[93]), .RECT2_HEIGHT(rectangle2_heights[93]), .RECT2_WEIGHT(rectangle2_weights[93]), .RECT3_X(rectangle3_xs[93]), .RECT3_Y(rectangle3_ys[93]), .RECT3_WIDTH(rectangle3_widths[93]), .RECT3_HEIGHT(rectangle3_heights[93]), .RECT3_WEIGHT(rectangle3_weights[93]), .FEAT_THRES(feature_thresholds[93]), .FEAT_ABOVE(feature_aboves[93]), .FEAT_BELOW(feature_belows[93])) ac93(.scan_win(scan_win93), .scan_win_std_dev(scan_win_std_dev[93]), .feature_accum(feature_accums[93]));
  accum_calculator #(.RECT1_X(rectangle1_xs[94]), .RECT1_Y(rectangle1_ys[94]), .RECT1_WIDTH(rectangle1_widths[94]), .RECT1_HEIGHT(rectangle1_heights[94]), .RECT1_WEIGHT(rectangle1_weights[94]), .RECT2_X(rectangle2_xs[94]), .RECT2_Y(rectangle2_ys[94]), .RECT2_WIDTH(rectangle2_widths[94]), .RECT2_HEIGHT(rectangle2_heights[94]), .RECT2_WEIGHT(rectangle2_weights[94]), .RECT3_X(rectangle3_xs[94]), .RECT3_Y(rectangle3_ys[94]), .RECT3_WIDTH(rectangle3_widths[94]), .RECT3_HEIGHT(rectangle3_heights[94]), .RECT3_WEIGHT(rectangle3_weights[94]), .FEAT_THRES(feature_thresholds[94]), .FEAT_ABOVE(feature_aboves[94]), .FEAT_BELOW(feature_belows[94])) ac94(.scan_win(scan_win94), .scan_win_std_dev(scan_win_std_dev[94]), .feature_accum(feature_accums[94]));
  accum_calculator #(.RECT1_X(rectangle1_xs[95]), .RECT1_Y(rectangle1_ys[95]), .RECT1_WIDTH(rectangle1_widths[95]), .RECT1_HEIGHT(rectangle1_heights[95]), .RECT1_WEIGHT(rectangle1_weights[95]), .RECT2_X(rectangle2_xs[95]), .RECT2_Y(rectangle2_ys[95]), .RECT2_WIDTH(rectangle2_widths[95]), .RECT2_HEIGHT(rectangle2_heights[95]), .RECT2_WEIGHT(rectangle2_weights[95]), .RECT3_X(rectangle3_xs[95]), .RECT3_Y(rectangle3_ys[95]), .RECT3_WIDTH(rectangle3_widths[95]), .RECT3_HEIGHT(rectangle3_heights[95]), .RECT3_WEIGHT(rectangle3_weights[95]), .FEAT_THRES(feature_thresholds[95]), .FEAT_ABOVE(feature_aboves[95]), .FEAT_BELOW(feature_belows[95])) ac95(.scan_win(scan_win95), .scan_win_std_dev(scan_win_std_dev[95]), .feature_accum(feature_accums[95]));
  accum_calculator #(.RECT1_X(rectangle1_xs[96]), .RECT1_Y(rectangle1_ys[96]), .RECT1_WIDTH(rectangle1_widths[96]), .RECT1_HEIGHT(rectangle1_heights[96]), .RECT1_WEIGHT(rectangle1_weights[96]), .RECT2_X(rectangle2_xs[96]), .RECT2_Y(rectangle2_ys[96]), .RECT2_WIDTH(rectangle2_widths[96]), .RECT2_HEIGHT(rectangle2_heights[96]), .RECT2_WEIGHT(rectangle2_weights[96]), .RECT3_X(rectangle3_xs[96]), .RECT3_Y(rectangle3_ys[96]), .RECT3_WIDTH(rectangle3_widths[96]), .RECT3_HEIGHT(rectangle3_heights[96]), .RECT3_WEIGHT(rectangle3_weights[96]), .FEAT_THRES(feature_thresholds[96]), .FEAT_ABOVE(feature_aboves[96]), .FEAT_BELOW(feature_belows[96])) ac96(.scan_win(scan_win96), .scan_win_std_dev(scan_win_std_dev[96]), .feature_accum(feature_accums[96]));
  accum_calculator #(.RECT1_X(rectangle1_xs[97]), .RECT1_Y(rectangle1_ys[97]), .RECT1_WIDTH(rectangle1_widths[97]), .RECT1_HEIGHT(rectangle1_heights[97]), .RECT1_WEIGHT(rectangle1_weights[97]), .RECT2_X(rectangle2_xs[97]), .RECT2_Y(rectangle2_ys[97]), .RECT2_WIDTH(rectangle2_widths[97]), .RECT2_HEIGHT(rectangle2_heights[97]), .RECT2_WEIGHT(rectangle2_weights[97]), .RECT3_X(rectangle3_xs[97]), .RECT3_Y(rectangle3_ys[97]), .RECT3_WIDTH(rectangle3_widths[97]), .RECT3_HEIGHT(rectangle3_heights[97]), .RECT3_WEIGHT(rectangle3_weights[97]), .FEAT_THRES(feature_thresholds[97]), .FEAT_ABOVE(feature_aboves[97]), .FEAT_BELOW(feature_belows[97])) ac97(.scan_win(scan_win97), .scan_win_std_dev(scan_win_std_dev[97]), .feature_accum(feature_accums[97]));
  accum_calculator #(.RECT1_X(rectangle1_xs[98]), .RECT1_Y(rectangle1_ys[98]), .RECT1_WIDTH(rectangle1_widths[98]), .RECT1_HEIGHT(rectangle1_heights[98]), .RECT1_WEIGHT(rectangle1_weights[98]), .RECT2_X(rectangle2_xs[98]), .RECT2_Y(rectangle2_ys[98]), .RECT2_WIDTH(rectangle2_widths[98]), .RECT2_HEIGHT(rectangle2_heights[98]), .RECT2_WEIGHT(rectangle2_weights[98]), .RECT3_X(rectangle3_xs[98]), .RECT3_Y(rectangle3_ys[98]), .RECT3_WIDTH(rectangle3_widths[98]), .RECT3_HEIGHT(rectangle3_heights[98]), .RECT3_WEIGHT(rectangle3_weights[98]), .FEAT_THRES(feature_thresholds[98]), .FEAT_ABOVE(feature_aboves[98]), .FEAT_BELOW(feature_belows[98])) ac98(.scan_win(scan_win98), .scan_win_std_dev(scan_win_std_dev[98]), .feature_accum(feature_accums[98]));
  accum_calculator #(.RECT1_X(rectangle1_xs[99]), .RECT1_Y(rectangle1_ys[99]), .RECT1_WIDTH(rectangle1_widths[99]), .RECT1_HEIGHT(rectangle1_heights[99]), .RECT1_WEIGHT(rectangle1_weights[99]), .RECT2_X(rectangle2_xs[99]), .RECT2_Y(rectangle2_ys[99]), .RECT2_WIDTH(rectangle2_widths[99]), .RECT2_HEIGHT(rectangle2_heights[99]), .RECT2_WEIGHT(rectangle2_weights[99]), .RECT3_X(rectangle3_xs[99]), .RECT3_Y(rectangle3_ys[99]), .RECT3_WIDTH(rectangle3_widths[99]), .RECT3_HEIGHT(rectangle3_heights[99]), .RECT3_WEIGHT(rectangle3_weights[99]), .FEAT_THRES(feature_thresholds[99]), .FEAT_ABOVE(feature_aboves[99]), .FEAT_BELOW(feature_belows[99])) ac99(.scan_win(scan_win99), .scan_win_std_dev(scan_win_std_dev[99]), .feature_accum(feature_accums[99]));
  accum_calculator #(.RECT1_X(rectangle1_xs[100]), .RECT1_Y(rectangle1_ys[100]), .RECT1_WIDTH(rectangle1_widths[100]), .RECT1_HEIGHT(rectangle1_heights[100]), .RECT1_WEIGHT(rectangle1_weights[100]), .RECT2_X(rectangle2_xs[100]), .RECT2_Y(rectangle2_ys[100]), .RECT2_WIDTH(rectangle2_widths[100]), .RECT2_HEIGHT(rectangle2_heights[100]), .RECT2_WEIGHT(rectangle2_weights[100]), .RECT3_X(rectangle3_xs[100]), .RECT3_Y(rectangle3_ys[100]), .RECT3_WIDTH(rectangle3_widths[100]), .RECT3_HEIGHT(rectangle3_heights[100]), .RECT3_WEIGHT(rectangle3_weights[100]), .FEAT_THRES(feature_thresholds[100]), .FEAT_ABOVE(feature_aboves[100]), .FEAT_BELOW(feature_belows[100])) ac100(.scan_win(scan_win100), .scan_win_std_dev(scan_win_std_dev[100]), .feature_accum(feature_accums[100]));
  accum_calculator #(.RECT1_X(rectangle1_xs[101]), .RECT1_Y(rectangle1_ys[101]), .RECT1_WIDTH(rectangle1_widths[101]), .RECT1_HEIGHT(rectangle1_heights[101]), .RECT1_WEIGHT(rectangle1_weights[101]), .RECT2_X(rectangle2_xs[101]), .RECT2_Y(rectangle2_ys[101]), .RECT2_WIDTH(rectangle2_widths[101]), .RECT2_HEIGHT(rectangle2_heights[101]), .RECT2_WEIGHT(rectangle2_weights[101]), .RECT3_X(rectangle3_xs[101]), .RECT3_Y(rectangle3_ys[101]), .RECT3_WIDTH(rectangle3_widths[101]), .RECT3_HEIGHT(rectangle3_heights[101]), .RECT3_WEIGHT(rectangle3_weights[101]), .FEAT_THRES(feature_thresholds[101]), .FEAT_ABOVE(feature_aboves[101]), .FEAT_BELOW(feature_belows[101])) ac101(.scan_win(scan_win101), .scan_win_std_dev(scan_win_std_dev[101]), .feature_accum(feature_accums[101]));
  accum_calculator #(.RECT1_X(rectangle1_xs[102]), .RECT1_Y(rectangle1_ys[102]), .RECT1_WIDTH(rectangle1_widths[102]), .RECT1_HEIGHT(rectangle1_heights[102]), .RECT1_WEIGHT(rectangle1_weights[102]), .RECT2_X(rectangle2_xs[102]), .RECT2_Y(rectangle2_ys[102]), .RECT2_WIDTH(rectangle2_widths[102]), .RECT2_HEIGHT(rectangle2_heights[102]), .RECT2_WEIGHT(rectangle2_weights[102]), .RECT3_X(rectangle3_xs[102]), .RECT3_Y(rectangle3_ys[102]), .RECT3_WIDTH(rectangle3_widths[102]), .RECT3_HEIGHT(rectangle3_heights[102]), .RECT3_WEIGHT(rectangle3_weights[102]), .FEAT_THRES(feature_thresholds[102]), .FEAT_ABOVE(feature_aboves[102]), .FEAT_BELOW(feature_belows[102])) ac102(.scan_win(scan_win102), .scan_win_std_dev(scan_win_std_dev[102]), .feature_accum(feature_accums[102]));
  accum_calculator #(.RECT1_X(rectangle1_xs[103]), .RECT1_Y(rectangle1_ys[103]), .RECT1_WIDTH(rectangle1_widths[103]), .RECT1_HEIGHT(rectangle1_heights[103]), .RECT1_WEIGHT(rectangle1_weights[103]), .RECT2_X(rectangle2_xs[103]), .RECT2_Y(rectangle2_ys[103]), .RECT2_WIDTH(rectangle2_widths[103]), .RECT2_HEIGHT(rectangle2_heights[103]), .RECT2_WEIGHT(rectangle2_weights[103]), .RECT3_X(rectangle3_xs[103]), .RECT3_Y(rectangle3_ys[103]), .RECT3_WIDTH(rectangle3_widths[103]), .RECT3_HEIGHT(rectangle3_heights[103]), .RECT3_WEIGHT(rectangle3_weights[103]), .FEAT_THRES(feature_thresholds[103]), .FEAT_ABOVE(feature_aboves[103]), .FEAT_BELOW(feature_belows[103])) ac103(.scan_win(scan_win103), .scan_win_std_dev(scan_win_std_dev[103]), .feature_accum(feature_accums[103]));
  accum_calculator #(.RECT1_X(rectangle1_xs[104]), .RECT1_Y(rectangle1_ys[104]), .RECT1_WIDTH(rectangle1_widths[104]), .RECT1_HEIGHT(rectangle1_heights[104]), .RECT1_WEIGHT(rectangle1_weights[104]), .RECT2_X(rectangle2_xs[104]), .RECT2_Y(rectangle2_ys[104]), .RECT2_WIDTH(rectangle2_widths[104]), .RECT2_HEIGHT(rectangle2_heights[104]), .RECT2_WEIGHT(rectangle2_weights[104]), .RECT3_X(rectangle3_xs[104]), .RECT3_Y(rectangle3_ys[104]), .RECT3_WIDTH(rectangle3_widths[104]), .RECT3_HEIGHT(rectangle3_heights[104]), .RECT3_WEIGHT(rectangle3_weights[104]), .FEAT_THRES(feature_thresholds[104]), .FEAT_ABOVE(feature_aboves[104]), .FEAT_BELOW(feature_belows[104])) ac104(.scan_win(scan_win104), .scan_win_std_dev(scan_win_std_dev[104]), .feature_accum(feature_accums[104]));
  accum_calculator #(.RECT1_X(rectangle1_xs[105]), .RECT1_Y(rectangle1_ys[105]), .RECT1_WIDTH(rectangle1_widths[105]), .RECT1_HEIGHT(rectangle1_heights[105]), .RECT1_WEIGHT(rectangle1_weights[105]), .RECT2_X(rectangle2_xs[105]), .RECT2_Y(rectangle2_ys[105]), .RECT2_WIDTH(rectangle2_widths[105]), .RECT2_HEIGHT(rectangle2_heights[105]), .RECT2_WEIGHT(rectangle2_weights[105]), .RECT3_X(rectangle3_xs[105]), .RECT3_Y(rectangle3_ys[105]), .RECT3_WIDTH(rectangle3_widths[105]), .RECT3_HEIGHT(rectangle3_heights[105]), .RECT3_WEIGHT(rectangle3_weights[105]), .FEAT_THRES(feature_thresholds[105]), .FEAT_ABOVE(feature_aboves[105]), .FEAT_BELOW(feature_belows[105])) ac105(.scan_win(scan_win105), .scan_win_std_dev(scan_win_std_dev[105]), .feature_accum(feature_accums[105]));
  accum_calculator #(.RECT1_X(rectangle1_xs[106]), .RECT1_Y(rectangle1_ys[106]), .RECT1_WIDTH(rectangle1_widths[106]), .RECT1_HEIGHT(rectangle1_heights[106]), .RECT1_WEIGHT(rectangle1_weights[106]), .RECT2_X(rectangle2_xs[106]), .RECT2_Y(rectangle2_ys[106]), .RECT2_WIDTH(rectangle2_widths[106]), .RECT2_HEIGHT(rectangle2_heights[106]), .RECT2_WEIGHT(rectangle2_weights[106]), .RECT3_X(rectangle3_xs[106]), .RECT3_Y(rectangle3_ys[106]), .RECT3_WIDTH(rectangle3_widths[106]), .RECT3_HEIGHT(rectangle3_heights[106]), .RECT3_WEIGHT(rectangle3_weights[106]), .FEAT_THRES(feature_thresholds[106]), .FEAT_ABOVE(feature_aboves[106]), .FEAT_BELOW(feature_belows[106])) ac106(.scan_win(scan_win106), .scan_win_std_dev(scan_win_std_dev[106]), .feature_accum(feature_accums[106]));
  accum_calculator #(.RECT1_X(rectangle1_xs[107]), .RECT1_Y(rectangle1_ys[107]), .RECT1_WIDTH(rectangle1_widths[107]), .RECT1_HEIGHT(rectangle1_heights[107]), .RECT1_WEIGHT(rectangle1_weights[107]), .RECT2_X(rectangle2_xs[107]), .RECT2_Y(rectangle2_ys[107]), .RECT2_WIDTH(rectangle2_widths[107]), .RECT2_HEIGHT(rectangle2_heights[107]), .RECT2_WEIGHT(rectangle2_weights[107]), .RECT3_X(rectangle3_xs[107]), .RECT3_Y(rectangle3_ys[107]), .RECT3_WIDTH(rectangle3_widths[107]), .RECT3_HEIGHT(rectangle3_heights[107]), .RECT3_WEIGHT(rectangle3_weights[107]), .FEAT_THRES(feature_thresholds[107]), .FEAT_ABOVE(feature_aboves[107]), .FEAT_BELOW(feature_belows[107])) ac107(.scan_win(scan_win107), .scan_win_std_dev(scan_win_std_dev[107]), .feature_accum(feature_accums[107]));
  accum_calculator #(.RECT1_X(rectangle1_xs[108]), .RECT1_Y(rectangle1_ys[108]), .RECT1_WIDTH(rectangle1_widths[108]), .RECT1_HEIGHT(rectangle1_heights[108]), .RECT1_WEIGHT(rectangle1_weights[108]), .RECT2_X(rectangle2_xs[108]), .RECT2_Y(rectangle2_ys[108]), .RECT2_WIDTH(rectangle2_widths[108]), .RECT2_HEIGHT(rectangle2_heights[108]), .RECT2_WEIGHT(rectangle2_weights[108]), .RECT3_X(rectangle3_xs[108]), .RECT3_Y(rectangle3_ys[108]), .RECT3_WIDTH(rectangle3_widths[108]), .RECT3_HEIGHT(rectangle3_heights[108]), .RECT3_WEIGHT(rectangle3_weights[108]), .FEAT_THRES(feature_thresholds[108]), .FEAT_ABOVE(feature_aboves[108]), .FEAT_BELOW(feature_belows[108])) ac108(.scan_win(scan_win108), .scan_win_std_dev(scan_win_std_dev[108]), .feature_accum(feature_accums[108]));
  accum_calculator #(.RECT1_X(rectangle1_xs[109]), .RECT1_Y(rectangle1_ys[109]), .RECT1_WIDTH(rectangle1_widths[109]), .RECT1_HEIGHT(rectangle1_heights[109]), .RECT1_WEIGHT(rectangle1_weights[109]), .RECT2_X(rectangle2_xs[109]), .RECT2_Y(rectangle2_ys[109]), .RECT2_WIDTH(rectangle2_widths[109]), .RECT2_HEIGHT(rectangle2_heights[109]), .RECT2_WEIGHT(rectangle2_weights[109]), .RECT3_X(rectangle3_xs[109]), .RECT3_Y(rectangle3_ys[109]), .RECT3_WIDTH(rectangle3_widths[109]), .RECT3_HEIGHT(rectangle3_heights[109]), .RECT3_WEIGHT(rectangle3_weights[109]), .FEAT_THRES(feature_thresholds[109]), .FEAT_ABOVE(feature_aboves[109]), .FEAT_BELOW(feature_belows[109])) ac109(.scan_win(scan_win109), .scan_win_std_dev(scan_win_std_dev[109]), .feature_accum(feature_accums[109]));
  accum_calculator #(.RECT1_X(rectangle1_xs[110]), .RECT1_Y(rectangle1_ys[110]), .RECT1_WIDTH(rectangle1_widths[110]), .RECT1_HEIGHT(rectangle1_heights[110]), .RECT1_WEIGHT(rectangle1_weights[110]), .RECT2_X(rectangle2_xs[110]), .RECT2_Y(rectangle2_ys[110]), .RECT2_WIDTH(rectangle2_widths[110]), .RECT2_HEIGHT(rectangle2_heights[110]), .RECT2_WEIGHT(rectangle2_weights[110]), .RECT3_X(rectangle3_xs[110]), .RECT3_Y(rectangle3_ys[110]), .RECT3_WIDTH(rectangle3_widths[110]), .RECT3_HEIGHT(rectangle3_heights[110]), .RECT3_WEIGHT(rectangle3_weights[110]), .FEAT_THRES(feature_thresholds[110]), .FEAT_ABOVE(feature_aboves[110]), .FEAT_BELOW(feature_belows[110])) ac110(.scan_win(scan_win110), .scan_win_std_dev(scan_win_std_dev[110]), .feature_accum(feature_accums[110]));
  accum_calculator #(.RECT1_X(rectangle1_xs[111]), .RECT1_Y(rectangle1_ys[111]), .RECT1_WIDTH(rectangle1_widths[111]), .RECT1_HEIGHT(rectangle1_heights[111]), .RECT1_WEIGHT(rectangle1_weights[111]), .RECT2_X(rectangle2_xs[111]), .RECT2_Y(rectangle2_ys[111]), .RECT2_WIDTH(rectangle2_widths[111]), .RECT2_HEIGHT(rectangle2_heights[111]), .RECT2_WEIGHT(rectangle2_weights[111]), .RECT3_X(rectangle3_xs[111]), .RECT3_Y(rectangle3_ys[111]), .RECT3_WIDTH(rectangle3_widths[111]), .RECT3_HEIGHT(rectangle3_heights[111]), .RECT3_WEIGHT(rectangle3_weights[111]), .FEAT_THRES(feature_thresholds[111]), .FEAT_ABOVE(feature_aboves[111]), .FEAT_BELOW(feature_belows[111])) ac111(.scan_win(scan_win111), .scan_win_std_dev(scan_win_std_dev[111]), .feature_accum(feature_accums[111]));
  accum_calculator #(.RECT1_X(rectangle1_xs[112]), .RECT1_Y(rectangle1_ys[112]), .RECT1_WIDTH(rectangle1_widths[112]), .RECT1_HEIGHT(rectangle1_heights[112]), .RECT1_WEIGHT(rectangle1_weights[112]), .RECT2_X(rectangle2_xs[112]), .RECT2_Y(rectangle2_ys[112]), .RECT2_WIDTH(rectangle2_widths[112]), .RECT2_HEIGHT(rectangle2_heights[112]), .RECT2_WEIGHT(rectangle2_weights[112]), .RECT3_X(rectangle3_xs[112]), .RECT3_Y(rectangle3_ys[112]), .RECT3_WIDTH(rectangle3_widths[112]), .RECT3_HEIGHT(rectangle3_heights[112]), .RECT3_WEIGHT(rectangle3_weights[112]), .FEAT_THRES(feature_thresholds[112]), .FEAT_ABOVE(feature_aboves[112]), .FEAT_BELOW(feature_belows[112])) ac112(.scan_win(scan_win112), .scan_win_std_dev(scan_win_std_dev[112]), .feature_accum(feature_accums[112]));
  accum_calculator #(.RECT1_X(rectangle1_xs[113]), .RECT1_Y(rectangle1_ys[113]), .RECT1_WIDTH(rectangle1_widths[113]), .RECT1_HEIGHT(rectangle1_heights[113]), .RECT1_WEIGHT(rectangle1_weights[113]), .RECT2_X(rectangle2_xs[113]), .RECT2_Y(rectangle2_ys[113]), .RECT2_WIDTH(rectangle2_widths[113]), .RECT2_HEIGHT(rectangle2_heights[113]), .RECT2_WEIGHT(rectangle2_weights[113]), .RECT3_X(rectangle3_xs[113]), .RECT3_Y(rectangle3_ys[113]), .RECT3_WIDTH(rectangle3_widths[113]), .RECT3_HEIGHT(rectangle3_heights[113]), .RECT3_WEIGHT(rectangle3_weights[113]), .FEAT_THRES(feature_thresholds[113]), .FEAT_ABOVE(feature_aboves[113]), .FEAT_BELOW(feature_belows[113])) ac113(.scan_win(scan_win113), .scan_win_std_dev(scan_win_std_dev[113]), .feature_accum(feature_accums[113]));
  accum_calculator #(.RECT1_X(rectangle1_xs[114]), .RECT1_Y(rectangle1_ys[114]), .RECT1_WIDTH(rectangle1_widths[114]), .RECT1_HEIGHT(rectangle1_heights[114]), .RECT1_WEIGHT(rectangle1_weights[114]), .RECT2_X(rectangle2_xs[114]), .RECT2_Y(rectangle2_ys[114]), .RECT2_WIDTH(rectangle2_widths[114]), .RECT2_HEIGHT(rectangle2_heights[114]), .RECT2_WEIGHT(rectangle2_weights[114]), .RECT3_X(rectangle3_xs[114]), .RECT3_Y(rectangle3_ys[114]), .RECT3_WIDTH(rectangle3_widths[114]), .RECT3_HEIGHT(rectangle3_heights[114]), .RECT3_WEIGHT(rectangle3_weights[114]), .FEAT_THRES(feature_thresholds[114]), .FEAT_ABOVE(feature_aboves[114]), .FEAT_BELOW(feature_belows[114])) ac114(.scan_win(scan_win114), .scan_win_std_dev(scan_win_std_dev[114]), .feature_accum(feature_accums[114]));
  accum_calculator #(.RECT1_X(rectangle1_xs[115]), .RECT1_Y(rectangle1_ys[115]), .RECT1_WIDTH(rectangle1_widths[115]), .RECT1_HEIGHT(rectangle1_heights[115]), .RECT1_WEIGHT(rectangle1_weights[115]), .RECT2_X(rectangle2_xs[115]), .RECT2_Y(rectangle2_ys[115]), .RECT2_WIDTH(rectangle2_widths[115]), .RECT2_HEIGHT(rectangle2_heights[115]), .RECT2_WEIGHT(rectangle2_weights[115]), .RECT3_X(rectangle3_xs[115]), .RECT3_Y(rectangle3_ys[115]), .RECT3_WIDTH(rectangle3_widths[115]), .RECT3_HEIGHT(rectangle3_heights[115]), .RECT3_WEIGHT(rectangle3_weights[115]), .FEAT_THRES(feature_thresholds[115]), .FEAT_ABOVE(feature_aboves[115]), .FEAT_BELOW(feature_belows[115])) ac115(.scan_win(scan_win115), .scan_win_std_dev(scan_win_std_dev[115]), .feature_accum(feature_accums[115]));
  accum_calculator #(.RECT1_X(rectangle1_xs[116]), .RECT1_Y(rectangle1_ys[116]), .RECT1_WIDTH(rectangle1_widths[116]), .RECT1_HEIGHT(rectangle1_heights[116]), .RECT1_WEIGHT(rectangle1_weights[116]), .RECT2_X(rectangle2_xs[116]), .RECT2_Y(rectangle2_ys[116]), .RECT2_WIDTH(rectangle2_widths[116]), .RECT2_HEIGHT(rectangle2_heights[116]), .RECT2_WEIGHT(rectangle2_weights[116]), .RECT3_X(rectangle3_xs[116]), .RECT3_Y(rectangle3_ys[116]), .RECT3_WIDTH(rectangle3_widths[116]), .RECT3_HEIGHT(rectangle3_heights[116]), .RECT3_WEIGHT(rectangle3_weights[116]), .FEAT_THRES(feature_thresholds[116]), .FEAT_ABOVE(feature_aboves[116]), .FEAT_BELOW(feature_belows[116])) ac116(.scan_win(scan_win116), .scan_win_std_dev(scan_win_std_dev[116]), .feature_accum(feature_accums[116]));
  accum_calculator #(.RECT1_X(rectangle1_xs[117]), .RECT1_Y(rectangle1_ys[117]), .RECT1_WIDTH(rectangle1_widths[117]), .RECT1_HEIGHT(rectangle1_heights[117]), .RECT1_WEIGHT(rectangle1_weights[117]), .RECT2_X(rectangle2_xs[117]), .RECT2_Y(rectangle2_ys[117]), .RECT2_WIDTH(rectangle2_widths[117]), .RECT2_HEIGHT(rectangle2_heights[117]), .RECT2_WEIGHT(rectangle2_weights[117]), .RECT3_X(rectangle3_xs[117]), .RECT3_Y(rectangle3_ys[117]), .RECT3_WIDTH(rectangle3_widths[117]), .RECT3_HEIGHT(rectangle3_heights[117]), .RECT3_WEIGHT(rectangle3_weights[117]), .FEAT_THRES(feature_thresholds[117]), .FEAT_ABOVE(feature_aboves[117]), .FEAT_BELOW(feature_belows[117])) ac117(.scan_win(scan_win117), .scan_win_std_dev(scan_win_std_dev[117]), .feature_accum(feature_accums[117]));
  accum_calculator #(.RECT1_X(rectangle1_xs[118]), .RECT1_Y(rectangle1_ys[118]), .RECT1_WIDTH(rectangle1_widths[118]), .RECT1_HEIGHT(rectangle1_heights[118]), .RECT1_WEIGHT(rectangle1_weights[118]), .RECT2_X(rectangle2_xs[118]), .RECT2_Y(rectangle2_ys[118]), .RECT2_WIDTH(rectangle2_widths[118]), .RECT2_HEIGHT(rectangle2_heights[118]), .RECT2_WEIGHT(rectangle2_weights[118]), .RECT3_X(rectangle3_xs[118]), .RECT3_Y(rectangle3_ys[118]), .RECT3_WIDTH(rectangle3_widths[118]), .RECT3_HEIGHT(rectangle3_heights[118]), .RECT3_WEIGHT(rectangle3_weights[118]), .FEAT_THRES(feature_thresholds[118]), .FEAT_ABOVE(feature_aboves[118]), .FEAT_BELOW(feature_belows[118])) ac118(.scan_win(scan_win118), .scan_win_std_dev(scan_win_std_dev[118]), .feature_accum(feature_accums[118]));
  accum_calculator #(.RECT1_X(rectangle1_xs[119]), .RECT1_Y(rectangle1_ys[119]), .RECT1_WIDTH(rectangle1_widths[119]), .RECT1_HEIGHT(rectangle1_heights[119]), .RECT1_WEIGHT(rectangle1_weights[119]), .RECT2_X(rectangle2_xs[119]), .RECT2_Y(rectangle2_ys[119]), .RECT2_WIDTH(rectangle2_widths[119]), .RECT2_HEIGHT(rectangle2_heights[119]), .RECT2_WEIGHT(rectangle2_weights[119]), .RECT3_X(rectangle3_xs[119]), .RECT3_Y(rectangle3_ys[119]), .RECT3_WIDTH(rectangle3_widths[119]), .RECT3_HEIGHT(rectangle3_heights[119]), .RECT3_WEIGHT(rectangle3_weights[119]), .FEAT_THRES(feature_thresholds[119]), .FEAT_ABOVE(feature_aboves[119]), .FEAT_BELOW(feature_belows[119])) ac119(.scan_win(scan_win119), .scan_win_std_dev(scan_win_std_dev[119]), .feature_accum(feature_accums[119]));
  accum_calculator #(.RECT1_X(rectangle1_xs[120]), .RECT1_Y(rectangle1_ys[120]), .RECT1_WIDTH(rectangle1_widths[120]), .RECT1_HEIGHT(rectangle1_heights[120]), .RECT1_WEIGHT(rectangle1_weights[120]), .RECT2_X(rectangle2_xs[120]), .RECT2_Y(rectangle2_ys[120]), .RECT2_WIDTH(rectangle2_widths[120]), .RECT2_HEIGHT(rectangle2_heights[120]), .RECT2_WEIGHT(rectangle2_weights[120]), .RECT3_X(rectangle3_xs[120]), .RECT3_Y(rectangle3_ys[120]), .RECT3_WIDTH(rectangle3_widths[120]), .RECT3_HEIGHT(rectangle3_heights[120]), .RECT3_WEIGHT(rectangle3_weights[120]), .FEAT_THRES(feature_thresholds[120]), .FEAT_ABOVE(feature_aboves[120]), .FEAT_BELOW(feature_belows[120])) ac120(.scan_win(scan_win120), .scan_win_std_dev(scan_win_std_dev[120]), .feature_accum(feature_accums[120]));
  accum_calculator #(.RECT1_X(rectangle1_xs[121]), .RECT1_Y(rectangle1_ys[121]), .RECT1_WIDTH(rectangle1_widths[121]), .RECT1_HEIGHT(rectangle1_heights[121]), .RECT1_WEIGHT(rectangle1_weights[121]), .RECT2_X(rectangle2_xs[121]), .RECT2_Y(rectangle2_ys[121]), .RECT2_WIDTH(rectangle2_widths[121]), .RECT2_HEIGHT(rectangle2_heights[121]), .RECT2_WEIGHT(rectangle2_weights[121]), .RECT3_X(rectangle3_xs[121]), .RECT3_Y(rectangle3_ys[121]), .RECT3_WIDTH(rectangle3_widths[121]), .RECT3_HEIGHT(rectangle3_heights[121]), .RECT3_WEIGHT(rectangle3_weights[121]), .FEAT_THRES(feature_thresholds[121]), .FEAT_ABOVE(feature_aboves[121]), .FEAT_BELOW(feature_belows[121])) ac121(.scan_win(scan_win121), .scan_win_std_dev(scan_win_std_dev[121]), .feature_accum(feature_accums[121]));
  accum_calculator #(.RECT1_X(rectangle1_xs[122]), .RECT1_Y(rectangle1_ys[122]), .RECT1_WIDTH(rectangle1_widths[122]), .RECT1_HEIGHT(rectangle1_heights[122]), .RECT1_WEIGHT(rectangle1_weights[122]), .RECT2_X(rectangle2_xs[122]), .RECT2_Y(rectangle2_ys[122]), .RECT2_WIDTH(rectangle2_widths[122]), .RECT2_HEIGHT(rectangle2_heights[122]), .RECT2_WEIGHT(rectangle2_weights[122]), .RECT3_X(rectangle3_xs[122]), .RECT3_Y(rectangle3_ys[122]), .RECT3_WIDTH(rectangle3_widths[122]), .RECT3_HEIGHT(rectangle3_heights[122]), .RECT3_WEIGHT(rectangle3_weights[122]), .FEAT_THRES(feature_thresholds[122]), .FEAT_ABOVE(feature_aboves[122]), .FEAT_BELOW(feature_belows[122])) ac122(.scan_win(scan_win122), .scan_win_std_dev(scan_win_std_dev[122]), .feature_accum(feature_accums[122]));
  accum_calculator #(.RECT1_X(rectangle1_xs[123]), .RECT1_Y(rectangle1_ys[123]), .RECT1_WIDTH(rectangle1_widths[123]), .RECT1_HEIGHT(rectangle1_heights[123]), .RECT1_WEIGHT(rectangle1_weights[123]), .RECT2_X(rectangle2_xs[123]), .RECT2_Y(rectangle2_ys[123]), .RECT2_WIDTH(rectangle2_widths[123]), .RECT2_HEIGHT(rectangle2_heights[123]), .RECT2_WEIGHT(rectangle2_weights[123]), .RECT3_X(rectangle3_xs[123]), .RECT3_Y(rectangle3_ys[123]), .RECT3_WIDTH(rectangle3_widths[123]), .RECT3_HEIGHT(rectangle3_heights[123]), .RECT3_WEIGHT(rectangle3_weights[123]), .FEAT_THRES(feature_thresholds[123]), .FEAT_ABOVE(feature_aboves[123]), .FEAT_BELOW(feature_belows[123])) ac123(.scan_win(scan_win123), .scan_win_std_dev(scan_win_std_dev[123]), .feature_accum(feature_accums[123]));
  accum_calculator #(.RECT1_X(rectangle1_xs[124]), .RECT1_Y(rectangle1_ys[124]), .RECT1_WIDTH(rectangle1_widths[124]), .RECT1_HEIGHT(rectangle1_heights[124]), .RECT1_WEIGHT(rectangle1_weights[124]), .RECT2_X(rectangle2_xs[124]), .RECT2_Y(rectangle2_ys[124]), .RECT2_WIDTH(rectangle2_widths[124]), .RECT2_HEIGHT(rectangle2_heights[124]), .RECT2_WEIGHT(rectangle2_weights[124]), .RECT3_X(rectangle3_xs[124]), .RECT3_Y(rectangle3_ys[124]), .RECT3_WIDTH(rectangle3_widths[124]), .RECT3_HEIGHT(rectangle3_heights[124]), .RECT3_WEIGHT(rectangle3_weights[124]), .FEAT_THRES(feature_thresholds[124]), .FEAT_ABOVE(feature_aboves[124]), .FEAT_BELOW(feature_belows[124])) ac124(.scan_win(scan_win124), .scan_win_std_dev(scan_win_std_dev[124]), .feature_accum(feature_accums[124]));
  accum_calculator #(.RECT1_X(rectangle1_xs[125]), .RECT1_Y(rectangle1_ys[125]), .RECT1_WIDTH(rectangle1_widths[125]), .RECT1_HEIGHT(rectangle1_heights[125]), .RECT1_WEIGHT(rectangle1_weights[125]), .RECT2_X(rectangle2_xs[125]), .RECT2_Y(rectangle2_ys[125]), .RECT2_WIDTH(rectangle2_widths[125]), .RECT2_HEIGHT(rectangle2_heights[125]), .RECT2_WEIGHT(rectangle2_weights[125]), .RECT3_X(rectangle3_xs[125]), .RECT3_Y(rectangle3_ys[125]), .RECT3_WIDTH(rectangle3_widths[125]), .RECT3_HEIGHT(rectangle3_heights[125]), .RECT3_WEIGHT(rectangle3_weights[125]), .FEAT_THRES(feature_thresholds[125]), .FEAT_ABOVE(feature_aboves[125]), .FEAT_BELOW(feature_belows[125])) ac125(.scan_win(scan_win125), .scan_win_std_dev(scan_win_std_dev[125]), .feature_accum(feature_accums[125]));
  accum_calculator #(.RECT1_X(rectangle1_xs[126]), .RECT1_Y(rectangle1_ys[126]), .RECT1_WIDTH(rectangle1_widths[126]), .RECT1_HEIGHT(rectangle1_heights[126]), .RECT1_WEIGHT(rectangle1_weights[126]), .RECT2_X(rectangle2_xs[126]), .RECT2_Y(rectangle2_ys[126]), .RECT2_WIDTH(rectangle2_widths[126]), .RECT2_HEIGHT(rectangle2_heights[126]), .RECT2_WEIGHT(rectangle2_weights[126]), .RECT3_X(rectangle3_xs[126]), .RECT3_Y(rectangle3_ys[126]), .RECT3_WIDTH(rectangle3_widths[126]), .RECT3_HEIGHT(rectangle3_heights[126]), .RECT3_WEIGHT(rectangle3_weights[126]), .FEAT_THRES(feature_thresholds[126]), .FEAT_ABOVE(feature_aboves[126]), .FEAT_BELOW(feature_belows[126])) ac126(.scan_win(scan_win126), .scan_win_std_dev(scan_win_std_dev[126]), .feature_accum(feature_accums[126]));
  accum_calculator #(.RECT1_X(rectangle1_xs[127]), .RECT1_Y(rectangle1_ys[127]), .RECT1_WIDTH(rectangle1_widths[127]), .RECT1_HEIGHT(rectangle1_heights[127]), .RECT1_WEIGHT(rectangle1_weights[127]), .RECT2_X(rectangle2_xs[127]), .RECT2_Y(rectangle2_ys[127]), .RECT2_WIDTH(rectangle2_widths[127]), .RECT2_HEIGHT(rectangle2_heights[127]), .RECT2_WEIGHT(rectangle2_weights[127]), .RECT3_X(rectangle3_xs[127]), .RECT3_Y(rectangle3_ys[127]), .RECT3_WIDTH(rectangle3_widths[127]), .RECT3_HEIGHT(rectangle3_heights[127]), .RECT3_WEIGHT(rectangle3_weights[127]), .FEAT_THRES(feature_thresholds[127]), .FEAT_ABOVE(feature_aboves[127]), .FEAT_BELOW(feature_belows[127])) ac127(.scan_win(scan_win127), .scan_win_std_dev(scan_win_std_dev[127]), .feature_accum(feature_accums[127]));
  accum_calculator #(.RECT1_X(rectangle1_xs[128]), .RECT1_Y(rectangle1_ys[128]), .RECT1_WIDTH(rectangle1_widths[128]), .RECT1_HEIGHT(rectangle1_heights[128]), .RECT1_WEIGHT(rectangle1_weights[128]), .RECT2_X(rectangle2_xs[128]), .RECT2_Y(rectangle2_ys[128]), .RECT2_WIDTH(rectangle2_widths[128]), .RECT2_HEIGHT(rectangle2_heights[128]), .RECT2_WEIGHT(rectangle2_weights[128]), .RECT3_X(rectangle3_xs[128]), .RECT3_Y(rectangle3_ys[128]), .RECT3_WIDTH(rectangle3_widths[128]), .RECT3_HEIGHT(rectangle3_heights[128]), .RECT3_WEIGHT(rectangle3_weights[128]), .FEAT_THRES(feature_thresholds[128]), .FEAT_ABOVE(feature_aboves[128]), .FEAT_BELOW(feature_belows[128])) ac128(.scan_win(scan_win128), .scan_win_std_dev(scan_win_std_dev[128]), .feature_accum(feature_accums[128]));
  accum_calculator #(.RECT1_X(rectangle1_xs[129]), .RECT1_Y(rectangle1_ys[129]), .RECT1_WIDTH(rectangle1_widths[129]), .RECT1_HEIGHT(rectangle1_heights[129]), .RECT1_WEIGHT(rectangle1_weights[129]), .RECT2_X(rectangle2_xs[129]), .RECT2_Y(rectangle2_ys[129]), .RECT2_WIDTH(rectangle2_widths[129]), .RECT2_HEIGHT(rectangle2_heights[129]), .RECT2_WEIGHT(rectangle2_weights[129]), .RECT3_X(rectangle3_xs[129]), .RECT3_Y(rectangle3_ys[129]), .RECT3_WIDTH(rectangle3_widths[129]), .RECT3_HEIGHT(rectangle3_heights[129]), .RECT3_WEIGHT(rectangle3_weights[129]), .FEAT_THRES(feature_thresholds[129]), .FEAT_ABOVE(feature_aboves[129]), .FEAT_BELOW(feature_belows[129])) ac129(.scan_win(scan_win129), .scan_win_std_dev(scan_win_std_dev[129]), .feature_accum(feature_accums[129]));
  accum_calculator #(.RECT1_X(rectangle1_xs[130]), .RECT1_Y(rectangle1_ys[130]), .RECT1_WIDTH(rectangle1_widths[130]), .RECT1_HEIGHT(rectangle1_heights[130]), .RECT1_WEIGHT(rectangle1_weights[130]), .RECT2_X(rectangle2_xs[130]), .RECT2_Y(rectangle2_ys[130]), .RECT2_WIDTH(rectangle2_widths[130]), .RECT2_HEIGHT(rectangle2_heights[130]), .RECT2_WEIGHT(rectangle2_weights[130]), .RECT3_X(rectangle3_xs[130]), .RECT3_Y(rectangle3_ys[130]), .RECT3_WIDTH(rectangle3_widths[130]), .RECT3_HEIGHT(rectangle3_heights[130]), .RECT3_WEIGHT(rectangle3_weights[130]), .FEAT_THRES(feature_thresholds[130]), .FEAT_ABOVE(feature_aboves[130]), .FEAT_BELOW(feature_belows[130])) ac130(.scan_win(scan_win130), .scan_win_std_dev(scan_win_std_dev[130]), .feature_accum(feature_accums[130]));
  accum_calculator #(.RECT1_X(rectangle1_xs[131]), .RECT1_Y(rectangle1_ys[131]), .RECT1_WIDTH(rectangle1_widths[131]), .RECT1_HEIGHT(rectangle1_heights[131]), .RECT1_WEIGHT(rectangle1_weights[131]), .RECT2_X(rectangle2_xs[131]), .RECT2_Y(rectangle2_ys[131]), .RECT2_WIDTH(rectangle2_widths[131]), .RECT2_HEIGHT(rectangle2_heights[131]), .RECT2_WEIGHT(rectangle2_weights[131]), .RECT3_X(rectangle3_xs[131]), .RECT3_Y(rectangle3_ys[131]), .RECT3_WIDTH(rectangle3_widths[131]), .RECT3_HEIGHT(rectangle3_heights[131]), .RECT3_WEIGHT(rectangle3_weights[131]), .FEAT_THRES(feature_thresholds[131]), .FEAT_ABOVE(feature_aboves[131]), .FEAT_BELOW(feature_belows[131])) ac131(.scan_win(scan_win131), .scan_win_std_dev(scan_win_std_dev[131]), .feature_accum(feature_accums[131]));
  accum_calculator #(.RECT1_X(rectangle1_xs[132]), .RECT1_Y(rectangle1_ys[132]), .RECT1_WIDTH(rectangle1_widths[132]), .RECT1_HEIGHT(rectangle1_heights[132]), .RECT1_WEIGHT(rectangle1_weights[132]), .RECT2_X(rectangle2_xs[132]), .RECT2_Y(rectangle2_ys[132]), .RECT2_WIDTH(rectangle2_widths[132]), .RECT2_HEIGHT(rectangle2_heights[132]), .RECT2_WEIGHT(rectangle2_weights[132]), .RECT3_X(rectangle3_xs[132]), .RECT3_Y(rectangle3_ys[132]), .RECT3_WIDTH(rectangle3_widths[132]), .RECT3_HEIGHT(rectangle3_heights[132]), .RECT3_WEIGHT(rectangle3_weights[132]), .FEAT_THRES(feature_thresholds[132]), .FEAT_ABOVE(feature_aboves[132]), .FEAT_BELOW(feature_belows[132])) ac132(.scan_win(scan_win132), .scan_win_std_dev(scan_win_std_dev[132]), .feature_accum(feature_accums[132]));
  accum_calculator #(.RECT1_X(rectangle1_xs[133]), .RECT1_Y(rectangle1_ys[133]), .RECT1_WIDTH(rectangle1_widths[133]), .RECT1_HEIGHT(rectangle1_heights[133]), .RECT1_WEIGHT(rectangle1_weights[133]), .RECT2_X(rectangle2_xs[133]), .RECT2_Y(rectangle2_ys[133]), .RECT2_WIDTH(rectangle2_widths[133]), .RECT2_HEIGHT(rectangle2_heights[133]), .RECT2_WEIGHT(rectangle2_weights[133]), .RECT3_X(rectangle3_xs[133]), .RECT3_Y(rectangle3_ys[133]), .RECT3_WIDTH(rectangle3_widths[133]), .RECT3_HEIGHT(rectangle3_heights[133]), .RECT3_WEIGHT(rectangle3_weights[133]), .FEAT_THRES(feature_thresholds[133]), .FEAT_ABOVE(feature_aboves[133]), .FEAT_BELOW(feature_belows[133])) ac133(.scan_win(scan_win133), .scan_win_std_dev(scan_win_std_dev[133]), .feature_accum(feature_accums[133]));
  accum_calculator #(.RECT1_X(rectangle1_xs[134]), .RECT1_Y(rectangle1_ys[134]), .RECT1_WIDTH(rectangle1_widths[134]), .RECT1_HEIGHT(rectangle1_heights[134]), .RECT1_WEIGHT(rectangle1_weights[134]), .RECT2_X(rectangle2_xs[134]), .RECT2_Y(rectangle2_ys[134]), .RECT2_WIDTH(rectangle2_widths[134]), .RECT2_HEIGHT(rectangle2_heights[134]), .RECT2_WEIGHT(rectangle2_weights[134]), .RECT3_X(rectangle3_xs[134]), .RECT3_Y(rectangle3_ys[134]), .RECT3_WIDTH(rectangle3_widths[134]), .RECT3_HEIGHT(rectangle3_heights[134]), .RECT3_WEIGHT(rectangle3_weights[134]), .FEAT_THRES(feature_thresholds[134]), .FEAT_ABOVE(feature_aboves[134]), .FEAT_BELOW(feature_belows[134])) ac134(.scan_win(scan_win134), .scan_win_std_dev(scan_win_std_dev[134]), .feature_accum(feature_accums[134]));
  accum_calculator #(.RECT1_X(rectangle1_xs[135]), .RECT1_Y(rectangle1_ys[135]), .RECT1_WIDTH(rectangle1_widths[135]), .RECT1_HEIGHT(rectangle1_heights[135]), .RECT1_WEIGHT(rectangle1_weights[135]), .RECT2_X(rectangle2_xs[135]), .RECT2_Y(rectangle2_ys[135]), .RECT2_WIDTH(rectangle2_widths[135]), .RECT2_HEIGHT(rectangle2_heights[135]), .RECT2_WEIGHT(rectangle2_weights[135]), .RECT3_X(rectangle3_xs[135]), .RECT3_Y(rectangle3_ys[135]), .RECT3_WIDTH(rectangle3_widths[135]), .RECT3_HEIGHT(rectangle3_heights[135]), .RECT3_WEIGHT(rectangle3_weights[135]), .FEAT_THRES(feature_thresholds[135]), .FEAT_ABOVE(feature_aboves[135]), .FEAT_BELOW(feature_belows[135])) ac135(.scan_win(scan_win135), .scan_win_std_dev(scan_win_std_dev[135]), .feature_accum(feature_accums[135]));
  accum_calculator #(.RECT1_X(rectangle1_xs[136]), .RECT1_Y(rectangle1_ys[136]), .RECT1_WIDTH(rectangle1_widths[136]), .RECT1_HEIGHT(rectangle1_heights[136]), .RECT1_WEIGHT(rectangle1_weights[136]), .RECT2_X(rectangle2_xs[136]), .RECT2_Y(rectangle2_ys[136]), .RECT2_WIDTH(rectangle2_widths[136]), .RECT2_HEIGHT(rectangle2_heights[136]), .RECT2_WEIGHT(rectangle2_weights[136]), .RECT3_X(rectangle3_xs[136]), .RECT3_Y(rectangle3_ys[136]), .RECT3_WIDTH(rectangle3_widths[136]), .RECT3_HEIGHT(rectangle3_heights[136]), .RECT3_WEIGHT(rectangle3_weights[136]), .FEAT_THRES(feature_thresholds[136]), .FEAT_ABOVE(feature_aboves[136]), .FEAT_BELOW(feature_belows[136])) ac136(.scan_win(scan_win136), .scan_win_std_dev(scan_win_std_dev[136]), .feature_accum(feature_accums[136]));
  accum_calculator #(.RECT1_X(rectangle1_xs[137]), .RECT1_Y(rectangle1_ys[137]), .RECT1_WIDTH(rectangle1_widths[137]), .RECT1_HEIGHT(rectangle1_heights[137]), .RECT1_WEIGHT(rectangle1_weights[137]), .RECT2_X(rectangle2_xs[137]), .RECT2_Y(rectangle2_ys[137]), .RECT2_WIDTH(rectangle2_widths[137]), .RECT2_HEIGHT(rectangle2_heights[137]), .RECT2_WEIGHT(rectangle2_weights[137]), .RECT3_X(rectangle3_xs[137]), .RECT3_Y(rectangle3_ys[137]), .RECT3_WIDTH(rectangle3_widths[137]), .RECT3_HEIGHT(rectangle3_heights[137]), .RECT3_WEIGHT(rectangle3_weights[137]), .FEAT_THRES(feature_thresholds[137]), .FEAT_ABOVE(feature_aboves[137]), .FEAT_BELOW(feature_belows[137])) ac137(.scan_win(scan_win137), .scan_win_std_dev(scan_win_std_dev[137]), .feature_accum(feature_accums[137]));
  accum_calculator #(.RECT1_X(rectangle1_xs[138]), .RECT1_Y(rectangle1_ys[138]), .RECT1_WIDTH(rectangle1_widths[138]), .RECT1_HEIGHT(rectangle1_heights[138]), .RECT1_WEIGHT(rectangle1_weights[138]), .RECT2_X(rectangle2_xs[138]), .RECT2_Y(rectangle2_ys[138]), .RECT2_WIDTH(rectangle2_widths[138]), .RECT2_HEIGHT(rectangle2_heights[138]), .RECT2_WEIGHT(rectangle2_weights[138]), .RECT3_X(rectangle3_xs[138]), .RECT3_Y(rectangle3_ys[138]), .RECT3_WIDTH(rectangle3_widths[138]), .RECT3_HEIGHT(rectangle3_heights[138]), .RECT3_WEIGHT(rectangle3_weights[138]), .FEAT_THRES(feature_thresholds[138]), .FEAT_ABOVE(feature_aboves[138]), .FEAT_BELOW(feature_belows[138])) ac138(.scan_win(scan_win138), .scan_win_std_dev(scan_win_std_dev[138]), .feature_accum(feature_accums[138]));
  accum_calculator #(.RECT1_X(rectangle1_xs[139]), .RECT1_Y(rectangle1_ys[139]), .RECT1_WIDTH(rectangle1_widths[139]), .RECT1_HEIGHT(rectangle1_heights[139]), .RECT1_WEIGHT(rectangle1_weights[139]), .RECT2_X(rectangle2_xs[139]), .RECT2_Y(rectangle2_ys[139]), .RECT2_WIDTH(rectangle2_widths[139]), .RECT2_HEIGHT(rectangle2_heights[139]), .RECT2_WEIGHT(rectangle2_weights[139]), .RECT3_X(rectangle3_xs[139]), .RECT3_Y(rectangle3_ys[139]), .RECT3_WIDTH(rectangle3_widths[139]), .RECT3_HEIGHT(rectangle3_heights[139]), .RECT3_WEIGHT(rectangle3_weights[139]), .FEAT_THRES(feature_thresholds[139]), .FEAT_ABOVE(feature_aboves[139]), .FEAT_BELOW(feature_belows[139])) ac139(.scan_win(scan_win139), .scan_win_std_dev(scan_win_std_dev[139]), .feature_accum(feature_accums[139]));
  accum_calculator #(.RECT1_X(rectangle1_xs[140]), .RECT1_Y(rectangle1_ys[140]), .RECT1_WIDTH(rectangle1_widths[140]), .RECT1_HEIGHT(rectangle1_heights[140]), .RECT1_WEIGHT(rectangle1_weights[140]), .RECT2_X(rectangle2_xs[140]), .RECT2_Y(rectangle2_ys[140]), .RECT2_WIDTH(rectangle2_widths[140]), .RECT2_HEIGHT(rectangle2_heights[140]), .RECT2_WEIGHT(rectangle2_weights[140]), .RECT3_X(rectangle3_xs[140]), .RECT3_Y(rectangle3_ys[140]), .RECT3_WIDTH(rectangle3_widths[140]), .RECT3_HEIGHT(rectangle3_heights[140]), .RECT3_WEIGHT(rectangle3_weights[140]), .FEAT_THRES(feature_thresholds[140]), .FEAT_ABOVE(feature_aboves[140]), .FEAT_BELOW(feature_belows[140])) ac140(.scan_win(scan_win140), .scan_win_std_dev(scan_win_std_dev[140]), .feature_accum(feature_accums[140]));
  accum_calculator #(.RECT1_X(rectangle1_xs[141]), .RECT1_Y(rectangle1_ys[141]), .RECT1_WIDTH(rectangle1_widths[141]), .RECT1_HEIGHT(rectangle1_heights[141]), .RECT1_WEIGHT(rectangle1_weights[141]), .RECT2_X(rectangle2_xs[141]), .RECT2_Y(rectangle2_ys[141]), .RECT2_WIDTH(rectangle2_widths[141]), .RECT2_HEIGHT(rectangle2_heights[141]), .RECT2_WEIGHT(rectangle2_weights[141]), .RECT3_X(rectangle3_xs[141]), .RECT3_Y(rectangle3_ys[141]), .RECT3_WIDTH(rectangle3_widths[141]), .RECT3_HEIGHT(rectangle3_heights[141]), .RECT3_WEIGHT(rectangle3_weights[141]), .FEAT_THRES(feature_thresholds[141]), .FEAT_ABOVE(feature_aboves[141]), .FEAT_BELOW(feature_belows[141])) ac141(.scan_win(scan_win141), .scan_win_std_dev(scan_win_std_dev[141]), .feature_accum(feature_accums[141]));
  accum_calculator #(.RECT1_X(rectangle1_xs[142]), .RECT1_Y(rectangle1_ys[142]), .RECT1_WIDTH(rectangle1_widths[142]), .RECT1_HEIGHT(rectangle1_heights[142]), .RECT1_WEIGHT(rectangle1_weights[142]), .RECT2_X(rectangle2_xs[142]), .RECT2_Y(rectangle2_ys[142]), .RECT2_WIDTH(rectangle2_widths[142]), .RECT2_HEIGHT(rectangle2_heights[142]), .RECT2_WEIGHT(rectangle2_weights[142]), .RECT3_X(rectangle3_xs[142]), .RECT3_Y(rectangle3_ys[142]), .RECT3_WIDTH(rectangle3_widths[142]), .RECT3_HEIGHT(rectangle3_heights[142]), .RECT3_WEIGHT(rectangle3_weights[142]), .FEAT_THRES(feature_thresholds[142]), .FEAT_ABOVE(feature_aboves[142]), .FEAT_BELOW(feature_belows[142])) ac142(.scan_win(scan_win142), .scan_win_std_dev(scan_win_std_dev[142]), .feature_accum(feature_accums[142]));
  accum_calculator #(.RECT1_X(rectangle1_xs[143]), .RECT1_Y(rectangle1_ys[143]), .RECT1_WIDTH(rectangle1_widths[143]), .RECT1_HEIGHT(rectangle1_heights[143]), .RECT1_WEIGHT(rectangle1_weights[143]), .RECT2_X(rectangle2_xs[143]), .RECT2_Y(rectangle2_ys[143]), .RECT2_WIDTH(rectangle2_widths[143]), .RECT2_HEIGHT(rectangle2_heights[143]), .RECT2_WEIGHT(rectangle2_weights[143]), .RECT3_X(rectangle3_xs[143]), .RECT3_Y(rectangle3_ys[143]), .RECT3_WIDTH(rectangle3_widths[143]), .RECT3_HEIGHT(rectangle3_heights[143]), .RECT3_WEIGHT(rectangle3_weights[143]), .FEAT_THRES(feature_thresholds[143]), .FEAT_ABOVE(feature_aboves[143]), .FEAT_BELOW(feature_belows[143])) ac143(.scan_win(scan_win143), .scan_win_std_dev(scan_win_std_dev[143]), .feature_accum(feature_accums[143]));
  accum_calculator #(.RECT1_X(rectangle1_xs[144]), .RECT1_Y(rectangle1_ys[144]), .RECT1_WIDTH(rectangle1_widths[144]), .RECT1_HEIGHT(rectangle1_heights[144]), .RECT1_WEIGHT(rectangle1_weights[144]), .RECT2_X(rectangle2_xs[144]), .RECT2_Y(rectangle2_ys[144]), .RECT2_WIDTH(rectangle2_widths[144]), .RECT2_HEIGHT(rectangle2_heights[144]), .RECT2_WEIGHT(rectangle2_weights[144]), .RECT3_X(rectangle3_xs[144]), .RECT3_Y(rectangle3_ys[144]), .RECT3_WIDTH(rectangle3_widths[144]), .RECT3_HEIGHT(rectangle3_heights[144]), .RECT3_WEIGHT(rectangle3_weights[144]), .FEAT_THRES(feature_thresholds[144]), .FEAT_ABOVE(feature_aboves[144]), .FEAT_BELOW(feature_belows[144])) ac144(.scan_win(scan_win144), .scan_win_std_dev(scan_win_std_dev[144]), .feature_accum(feature_accums[144]));
  accum_calculator #(.RECT1_X(rectangle1_xs[145]), .RECT1_Y(rectangle1_ys[145]), .RECT1_WIDTH(rectangle1_widths[145]), .RECT1_HEIGHT(rectangle1_heights[145]), .RECT1_WEIGHT(rectangle1_weights[145]), .RECT2_X(rectangle2_xs[145]), .RECT2_Y(rectangle2_ys[145]), .RECT2_WIDTH(rectangle2_widths[145]), .RECT2_HEIGHT(rectangle2_heights[145]), .RECT2_WEIGHT(rectangle2_weights[145]), .RECT3_X(rectangle3_xs[145]), .RECT3_Y(rectangle3_ys[145]), .RECT3_WIDTH(rectangle3_widths[145]), .RECT3_HEIGHT(rectangle3_heights[145]), .RECT3_WEIGHT(rectangle3_weights[145]), .FEAT_THRES(feature_thresholds[145]), .FEAT_ABOVE(feature_aboves[145]), .FEAT_BELOW(feature_belows[145])) ac145(.scan_win(scan_win145), .scan_win_std_dev(scan_win_std_dev[145]), .feature_accum(feature_accums[145]));
  accum_calculator #(.RECT1_X(rectangle1_xs[146]), .RECT1_Y(rectangle1_ys[146]), .RECT1_WIDTH(rectangle1_widths[146]), .RECT1_HEIGHT(rectangle1_heights[146]), .RECT1_WEIGHT(rectangle1_weights[146]), .RECT2_X(rectangle2_xs[146]), .RECT2_Y(rectangle2_ys[146]), .RECT2_WIDTH(rectangle2_widths[146]), .RECT2_HEIGHT(rectangle2_heights[146]), .RECT2_WEIGHT(rectangle2_weights[146]), .RECT3_X(rectangle3_xs[146]), .RECT3_Y(rectangle3_ys[146]), .RECT3_WIDTH(rectangle3_widths[146]), .RECT3_HEIGHT(rectangle3_heights[146]), .RECT3_WEIGHT(rectangle3_weights[146]), .FEAT_THRES(feature_thresholds[146]), .FEAT_ABOVE(feature_aboves[146]), .FEAT_BELOW(feature_belows[146])) ac146(.scan_win(scan_win146), .scan_win_std_dev(scan_win_std_dev[146]), .feature_accum(feature_accums[146]));
  accum_calculator #(.RECT1_X(rectangle1_xs[147]), .RECT1_Y(rectangle1_ys[147]), .RECT1_WIDTH(rectangle1_widths[147]), .RECT1_HEIGHT(rectangle1_heights[147]), .RECT1_WEIGHT(rectangle1_weights[147]), .RECT2_X(rectangle2_xs[147]), .RECT2_Y(rectangle2_ys[147]), .RECT2_WIDTH(rectangle2_widths[147]), .RECT2_HEIGHT(rectangle2_heights[147]), .RECT2_WEIGHT(rectangle2_weights[147]), .RECT3_X(rectangle3_xs[147]), .RECT3_Y(rectangle3_ys[147]), .RECT3_WIDTH(rectangle3_widths[147]), .RECT3_HEIGHT(rectangle3_heights[147]), .RECT3_WEIGHT(rectangle3_weights[147]), .FEAT_THRES(feature_thresholds[147]), .FEAT_ABOVE(feature_aboves[147]), .FEAT_BELOW(feature_belows[147])) ac147(.scan_win(scan_win147), .scan_win_std_dev(scan_win_std_dev[147]), .feature_accum(feature_accums[147]));
  accum_calculator #(.RECT1_X(rectangle1_xs[148]), .RECT1_Y(rectangle1_ys[148]), .RECT1_WIDTH(rectangle1_widths[148]), .RECT1_HEIGHT(rectangle1_heights[148]), .RECT1_WEIGHT(rectangle1_weights[148]), .RECT2_X(rectangle2_xs[148]), .RECT2_Y(rectangle2_ys[148]), .RECT2_WIDTH(rectangle2_widths[148]), .RECT2_HEIGHT(rectangle2_heights[148]), .RECT2_WEIGHT(rectangle2_weights[148]), .RECT3_X(rectangle3_xs[148]), .RECT3_Y(rectangle3_ys[148]), .RECT3_WIDTH(rectangle3_widths[148]), .RECT3_HEIGHT(rectangle3_heights[148]), .RECT3_WEIGHT(rectangle3_weights[148]), .FEAT_THRES(feature_thresholds[148]), .FEAT_ABOVE(feature_aboves[148]), .FEAT_BELOW(feature_belows[148])) ac148(.scan_win(scan_win148), .scan_win_std_dev(scan_win_std_dev[148]), .feature_accum(feature_accums[148]));
  accum_calculator #(.RECT1_X(rectangle1_xs[149]), .RECT1_Y(rectangle1_ys[149]), .RECT1_WIDTH(rectangle1_widths[149]), .RECT1_HEIGHT(rectangle1_heights[149]), .RECT1_WEIGHT(rectangle1_weights[149]), .RECT2_X(rectangle2_xs[149]), .RECT2_Y(rectangle2_ys[149]), .RECT2_WIDTH(rectangle2_widths[149]), .RECT2_HEIGHT(rectangle2_heights[149]), .RECT2_WEIGHT(rectangle2_weights[149]), .RECT3_X(rectangle3_xs[149]), .RECT3_Y(rectangle3_ys[149]), .RECT3_WIDTH(rectangle3_widths[149]), .RECT3_HEIGHT(rectangle3_heights[149]), .RECT3_WEIGHT(rectangle3_weights[149]), .FEAT_THRES(feature_thresholds[149]), .FEAT_ABOVE(feature_aboves[149]), .FEAT_BELOW(feature_belows[149])) ac149(.scan_win(scan_win149), .scan_win_std_dev(scan_win_std_dev[149]), .feature_accum(feature_accums[149]));
  accum_calculator #(.RECT1_X(rectangle1_xs[150]), .RECT1_Y(rectangle1_ys[150]), .RECT1_WIDTH(rectangle1_widths[150]), .RECT1_HEIGHT(rectangle1_heights[150]), .RECT1_WEIGHT(rectangle1_weights[150]), .RECT2_X(rectangle2_xs[150]), .RECT2_Y(rectangle2_ys[150]), .RECT2_WIDTH(rectangle2_widths[150]), .RECT2_HEIGHT(rectangle2_heights[150]), .RECT2_WEIGHT(rectangle2_weights[150]), .RECT3_X(rectangle3_xs[150]), .RECT3_Y(rectangle3_ys[150]), .RECT3_WIDTH(rectangle3_widths[150]), .RECT3_HEIGHT(rectangle3_heights[150]), .RECT3_WEIGHT(rectangle3_weights[150]), .FEAT_THRES(feature_thresholds[150]), .FEAT_ABOVE(feature_aboves[150]), .FEAT_BELOW(feature_belows[150])) ac150(.scan_win(scan_win150), .scan_win_std_dev(scan_win_std_dev[150]), .feature_accum(feature_accums[150]));
  accum_calculator #(.RECT1_X(rectangle1_xs[151]), .RECT1_Y(rectangle1_ys[151]), .RECT1_WIDTH(rectangle1_widths[151]), .RECT1_HEIGHT(rectangle1_heights[151]), .RECT1_WEIGHT(rectangle1_weights[151]), .RECT2_X(rectangle2_xs[151]), .RECT2_Y(rectangle2_ys[151]), .RECT2_WIDTH(rectangle2_widths[151]), .RECT2_HEIGHT(rectangle2_heights[151]), .RECT2_WEIGHT(rectangle2_weights[151]), .RECT3_X(rectangle3_xs[151]), .RECT3_Y(rectangle3_ys[151]), .RECT3_WIDTH(rectangle3_widths[151]), .RECT3_HEIGHT(rectangle3_heights[151]), .RECT3_WEIGHT(rectangle3_weights[151]), .FEAT_THRES(feature_thresholds[151]), .FEAT_ABOVE(feature_aboves[151]), .FEAT_BELOW(feature_belows[151])) ac151(.scan_win(scan_win151), .scan_win_std_dev(scan_win_std_dev[151]), .feature_accum(feature_accums[151]));
  accum_calculator #(.RECT1_X(rectangle1_xs[152]), .RECT1_Y(rectangle1_ys[152]), .RECT1_WIDTH(rectangle1_widths[152]), .RECT1_HEIGHT(rectangle1_heights[152]), .RECT1_WEIGHT(rectangle1_weights[152]), .RECT2_X(rectangle2_xs[152]), .RECT2_Y(rectangle2_ys[152]), .RECT2_WIDTH(rectangle2_widths[152]), .RECT2_HEIGHT(rectangle2_heights[152]), .RECT2_WEIGHT(rectangle2_weights[152]), .RECT3_X(rectangle3_xs[152]), .RECT3_Y(rectangle3_ys[152]), .RECT3_WIDTH(rectangle3_widths[152]), .RECT3_HEIGHT(rectangle3_heights[152]), .RECT3_WEIGHT(rectangle3_weights[152]), .FEAT_THRES(feature_thresholds[152]), .FEAT_ABOVE(feature_aboves[152]), .FEAT_BELOW(feature_belows[152])) ac152(.scan_win(scan_win152), .scan_win_std_dev(scan_win_std_dev[152]), .feature_accum(feature_accums[152]));
  accum_calculator #(.RECT1_X(rectangle1_xs[153]), .RECT1_Y(rectangle1_ys[153]), .RECT1_WIDTH(rectangle1_widths[153]), .RECT1_HEIGHT(rectangle1_heights[153]), .RECT1_WEIGHT(rectangle1_weights[153]), .RECT2_X(rectangle2_xs[153]), .RECT2_Y(rectangle2_ys[153]), .RECT2_WIDTH(rectangle2_widths[153]), .RECT2_HEIGHT(rectangle2_heights[153]), .RECT2_WEIGHT(rectangle2_weights[153]), .RECT3_X(rectangle3_xs[153]), .RECT3_Y(rectangle3_ys[153]), .RECT3_WIDTH(rectangle3_widths[153]), .RECT3_HEIGHT(rectangle3_heights[153]), .RECT3_WEIGHT(rectangle3_weights[153]), .FEAT_THRES(feature_thresholds[153]), .FEAT_ABOVE(feature_aboves[153]), .FEAT_BELOW(feature_belows[153])) ac153(.scan_win(scan_win153), .scan_win_std_dev(scan_win_std_dev[153]), .feature_accum(feature_accums[153]));
  accum_calculator #(.RECT1_X(rectangle1_xs[154]), .RECT1_Y(rectangle1_ys[154]), .RECT1_WIDTH(rectangle1_widths[154]), .RECT1_HEIGHT(rectangle1_heights[154]), .RECT1_WEIGHT(rectangle1_weights[154]), .RECT2_X(rectangle2_xs[154]), .RECT2_Y(rectangle2_ys[154]), .RECT2_WIDTH(rectangle2_widths[154]), .RECT2_HEIGHT(rectangle2_heights[154]), .RECT2_WEIGHT(rectangle2_weights[154]), .RECT3_X(rectangle3_xs[154]), .RECT3_Y(rectangle3_ys[154]), .RECT3_WIDTH(rectangle3_widths[154]), .RECT3_HEIGHT(rectangle3_heights[154]), .RECT3_WEIGHT(rectangle3_weights[154]), .FEAT_THRES(feature_thresholds[154]), .FEAT_ABOVE(feature_aboves[154]), .FEAT_BELOW(feature_belows[154])) ac154(.scan_win(scan_win154), .scan_win_std_dev(scan_win_std_dev[154]), .feature_accum(feature_accums[154]));
  accum_calculator #(.RECT1_X(rectangle1_xs[155]), .RECT1_Y(rectangle1_ys[155]), .RECT1_WIDTH(rectangle1_widths[155]), .RECT1_HEIGHT(rectangle1_heights[155]), .RECT1_WEIGHT(rectangle1_weights[155]), .RECT2_X(rectangle2_xs[155]), .RECT2_Y(rectangle2_ys[155]), .RECT2_WIDTH(rectangle2_widths[155]), .RECT2_HEIGHT(rectangle2_heights[155]), .RECT2_WEIGHT(rectangle2_weights[155]), .RECT3_X(rectangle3_xs[155]), .RECT3_Y(rectangle3_ys[155]), .RECT3_WIDTH(rectangle3_widths[155]), .RECT3_HEIGHT(rectangle3_heights[155]), .RECT3_WEIGHT(rectangle3_weights[155]), .FEAT_THRES(feature_thresholds[155]), .FEAT_ABOVE(feature_aboves[155]), .FEAT_BELOW(feature_belows[155])) ac155(.scan_win(scan_win155), .scan_win_std_dev(scan_win_std_dev[155]), .feature_accum(feature_accums[155]));
  accum_calculator #(.RECT1_X(rectangle1_xs[156]), .RECT1_Y(rectangle1_ys[156]), .RECT1_WIDTH(rectangle1_widths[156]), .RECT1_HEIGHT(rectangle1_heights[156]), .RECT1_WEIGHT(rectangle1_weights[156]), .RECT2_X(rectangle2_xs[156]), .RECT2_Y(rectangle2_ys[156]), .RECT2_WIDTH(rectangle2_widths[156]), .RECT2_HEIGHT(rectangle2_heights[156]), .RECT2_WEIGHT(rectangle2_weights[156]), .RECT3_X(rectangle3_xs[156]), .RECT3_Y(rectangle3_ys[156]), .RECT3_WIDTH(rectangle3_widths[156]), .RECT3_HEIGHT(rectangle3_heights[156]), .RECT3_WEIGHT(rectangle3_weights[156]), .FEAT_THRES(feature_thresholds[156]), .FEAT_ABOVE(feature_aboves[156]), .FEAT_BELOW(feature_belows[156])) ac156(.scan_win(scan_win156), .scan_win_std_dev(scan_win_std_dev[156]), .feature_accum(feature_accums[156]));
  accum_calculator #(.RECT1_X(rectangle1_xs[157]), .RECT1_Y(rectangle1_ys[157]), .RECT1_WIDTH(rectangle1_widths[157]), .RECT1_HEIGHT(rectangle1_heights[157]), .RECT1_WEIGHT(rectangle1_weights[157]), .RECT2_X(rectangle2_xs[157]), .RECT2_Y(rectangle2_ys[157]), .RECT2_WIDTH(rectangle2_widths[157]), .RECT2_HEIGHT(rectangle2_heights[157]), .RECT2_WEIGHT(rectangle2_weights[157]), .RECT3_X(rectangle3_xs[157]), .RECT3_Y(rectangle3_ys[157]), .RECT3_WIDTH(rectangle3_widths[157]), .RECT3_HEIGHT(rectangle3_heights[157]), .RECT3_WEIGHT(rectangle3_weights[157]), .FEAT_THRES(feature_thresholds[157]), .FEAT_ABOVE(feature_aboves[157]), .FEAT_BELOW(feature_belows[157])) ac157(.scan_win(scan_win157), .scan_win_std_dev(scan_win_std_dev[157]), .feature_accum(feature_accums[157]));
  accum_calculator #(.RECT1_X(rectangle1_xs[158]), .RECT1_Y(rectangle1_ys[158]), .RECT1_WIDTH(rectangle1_widths[158]), .RECT1_HEIGHT(rectangle1_heights[158]), .RECT1_WEIGHT(rectangle1_weights[158]), .RECT2_X(rectangle2_xs[158]), .RECT2_Y(rectangle2_ys[158]), .RECT2_WIDTH(rectangle2_widths[158]), .RECT2_HEIGHT(rectangle2_heights[158]), .RECT2_WEIGHT(rectangle2_weights[158]), .RECT3_X(rectangle3_xs[158]), .RECT3_Y(rectangle3_ys[158]), .RECT3_WIDTH(rectangle3_widths[158]), .RECT3_HEIGHT(rectangle3_heights[158]), .RECT3_WEIGHT(rectangle3_weights[158]), .FEAT_THRES(feature_thresholds[158]), .FEAT_ABOVE(feature_aboves[158]), .FEAT_BELOW(feature_belows[158])) ac158(.scan_win(scan_win158), .scan_win_std_dev(scan_win_std_dev[158]), .feature_accum(feature_accums[158]));
  accum_calculator #(.RECT1_X(rectangle1_xs[159]), .RECT1_Y(rectangle1_ys[159]), .RECT1_WIDTH(rectangle1_widths[159]), .RECT1_HEIGHT(rectangle1_heights[159]), .RECT1_WEIGHT(rectangle1_weights[159]), .RECT2_X(rectangle2_xs[159]), .RECT2_Y(rectangle2_ys[159]), .RECT2_WIDTH(rectangle2_widths[159]), .RECT2_HEIGHT(rectangle2_heights[159]), .RECT2_WEIGHT(rectangle2_weights[159]), .RECT3_X(rectangle3_xs[159]), .RECT3_Y(rectangle3_ys[159]), .RECT3_WIDTH(rectangle3_widths[159]), .RECT3_HEIGHT(rectangle3_heights[159]), .RECT3_WEIGHT(rectangle3_weights[159]), .FEAT_THRES(feature_thresholds[159]), .FEAT_ABOVE(feature_aboves[159]), .FEAT_BELOW(feature_belows[159])) ac159(.scan_win(scan_win159), .scan_win_std_dev(scan_win_std_dev[159]), .feature_accum(feature_accums[159]));
  accum_calculator #(.RECT1_X(rectangle1_xs[160]), .RECT1_Y(rectangle1_ys[160]), .RECT1_WIDTH(rectangle1_widths[160]), .RECT1_HEIGHT(rectangle1_heights[160]), .RECT1_WEIGHT(rectangle1_weights[160]), .RECT2_X(rectangle2_xs[160]), .RECT2_Y(rectangle2_ys[160]), .RECT2_WIDTH(rectangle2_widths[160]), .RECT2_HEIGHT(rectangle2_heights[160]), .RECT2_WEIGHT(rectangle2_weights[160]), .RECT3_X(rectangle3_xs[160]), .RECT3_Y(rectangle3_ys[160]), .RECT3_WIDTH(rectangle3_widths[160]), .RECT3_HEIGHT(rectangle3_heights[160]), .RECT3_WEIGHT(rectangle3_weights[160]), .FEAT_THRES(feature_thresholds[160]), .FEAT_ABOVE(feature_aboves[160]), .FEAT_BELOW(feature_belows[160])) ac160(.scan_win(scan_win160), .scan_win_std_dev(scan_win_std_dev[160]), .feature_accum(feature_accums[160]));
  accum_calculator #(.RECT1_X(rectangle1_xs[161]), .RECT1_Y(rectangle1_ys[161]), .RECT1_WIDTH(rectangle1_widths[161]), .RECT1_HEIGHT(rectangle1_heights[161]), .RECT1_WEIGHT(rectangle1_weights[161]), .RECT2_X(rectangle2_xs[161]), .RECT2_Y(rectangle2_ys[161]), .RECT2_WIDTH(rectangle2_widths[161]), .RECT2_HEIGHT(rectangle2_heights[161]), .RECT2_WEIGHT(rectangle2_weights[161]), .RECT3_X(rectangle3_xs[161]), .RECT3_Y(rectangle3_ys[161]), .RECT3_WIDTH(rectangle3_widths[161]), .RECT3_HEIGHT(rectangle3_heights[161]), .RECT3_WEIGHT(rectangle3_weights[161]), .FEAT_THRES(feature_thresholds[161]), .FEAT_ABOVE(feature_aboves[161]), .FEAT_BELOW(feature_belows[161])) ac161(.scan_win(scan_win161), .scan_win_std_dev(scan_win_std_dev[161]), .feature_accum(feature_accums[161]));
  accum_calculator #(.RECT1_X(rectangle1_xs[162]), .RECT1_Y(rectangle1_ys[162]), .RECT1_WIDTH(rectangle1_widths[162]), .RECT1_HEIGHT(rectangle1_heights[162]), .RECT1_WEIGHT(rectangle1_weights[162]), .RECT2_X(rectangle2_xs[162]), .RECT2_Y(rectangle2_ys[162]), .RECT2_WIDTH(rectangle2_widths[162]), .RECT2_HEIGHT(rectangle2_heights[162]), .RECT2_WEIGHT(rectangle2_weights[162]), .RECT3_X(rectangle3_xs[162]), .RECT3_Y(rectangle3_ys[162]), .RECT3_WIDTH(rectangle3_widths[162]), .RECT3_HEIGHT(rectangle3_heights[162]), .RECT3_WEIGHT(rectangle3_weights[162]), .FEAT_THRES(feature_thresholds[162]), .FEAT_ABOVE(feature_aboves[162]), .FEAT_BELOW(feature_belows[162])) ac162(.scan_win(scan_win162), .scan_win_std_dev(scan_win_std_dev[162]), .feature_accum(feature_accums[162]));
  accum_calculator #(.RECT1_X(rectangle1_xs[163]), .RECT1_Y(rectangle1_ys[163]), .RECT1_WIDTH(rectangle1_widths[163]), .RECT1_HEIGHT(rectangle1_heights[163]), .RECT1_WEIGHT(rectangle1_weights[163]), .RECT2_X(rectangle2_xs[163]), .RECT2_Y(rectangle2_ys[163]), .RECT2_WIDTH(rectangle2_widths[163]), .RECT2_HEIGHT(rectangle2_heights[163]), .RECT2_WEIGHT(rectangle2_weights[163]), .RECT3_X(rectangle3_xs[163]), .RECT3_Y(rectangle3_ys[163]), .RECT3_WIDTH(rectangle3_widths[163]), .RECT3_HEIGHT(rectangle3_heights[163]), .RECT3_WEIGHT(rectangle3_weights[163]), .FEAT_THRES(feature_thresholds[163]), .FEAT_ABOVE(feature_aboves[163]), .FEAT_BELOW(feature_belows[163])) ac163(.scan_win(scan_win163), .scan_win_std_dev(scan_win_std_dev[163]), .feature_accum(feature_accums[163]));
  accum_calculator #(.RECT1_X(rectangle1_xs[164]), .RECT1_Y(rectangle1_ys[164]), .RECT1_WIDTH(rectangle1_widths[164]), .RECT1_HEIGHT(rectangle1_heights[164]), .RECT1_WEIGHT(rectangle1_weights[164]), .RECT2_X(rectangle2_xs[164]), .RECT2_Y(rectangle2_ys[164]), .RECT2_WIDTH(rectangle2_widths[164]), .RECT2_HEIGHT(rectangle2_heights[164]), .RECT2_WEIGHT(rectangle2_weights[164]), .RECT3_X(rectangle3_xs[164]), .RECT3_Y(rectangle3_ys[164]), .RECT3_WIDTH(rectangle3_widths[164]), .RECT3_HEIGHT(rectangle3_heights[164]), .RECT3_WEIGHT(rectangle3_weights[164]), .FEAT_THRES(feature_thresholds[164]), .FEAT_ABOVE(feature_aboves[164]), .FEAT_BELOW(feature_belows[164])) ac164(.scan_win(scan_win164), .scan_win_std_dev(scan_win_std_dev[164]), .feature_accum(feature_accums[164]));
  accum_calculator #(.RECT1_X(rectangle1_xs[165]), .RECT1_Y(rectangle1_ys[165]), .RECT1_WIDTH(rectangle1_widths[165]), .RECT1_HEIGHT(rectangle1_heights[165]), .RECT1_WEIGHT(rectangle1_weights[165]), .RECT2_X(rectangle2_xs[165]), .RECT2_Y(rectangle2_ys[165]), .RECT2_WIDTH(rectangle2_widths[165]), .RECT2_HEIGHT(rectangle2_heights[165]), .RECT2_WEIGHT(rectangle2_weights[165]), .RECT3_X(rectangle3_xs[165]), .RECT3_Y(rectangle3_ys[165]), .RECT3_WIDTH(rectangle3_widths[165]), .RECT3_HEIGHT(rectangle3_heights[165]), .RECT3_WEIGHT(rectangle3_weights[165]), .FEAT_THRES(feature_thresholds[165]), .FEAT_ABOVE(feature_aboves[165]), .FEAT_BELOW(feature_belows[165])) ac165(.scan_win(scan_win165), .scan_win_std_dev(scan_win_std_dev[165]), .feature_accum(feature_accums[165]));
  accum_calculator #(.RECT1_X(rectangle1_xs[166]), .RECT1_Y(rectangle1_ys[166]), .RECT1_WIDTH(rectangle1_widths[166]), .RECT1_HEIGHT(rectangle1_heights[166]), .RECT1_WEIGHT(rectangle1_weights[166]), .RECT2_X(rectangle2_xs[166]), .RECT2_Y(rectangle2_ys[166]), .RECT2_WIDTH(rectangle2_widths[166]), .RECT2_HEIGHT(rectangle2_heights[166]), .RECT2_WEIGHT(rectangle2_weights[166]), .RECT3_X(rectangle3_xs[166]), .RECT3_Y(rectangle3_ys[166]), .RECT3_WIDTH(rectangle3_widths[166]), .RECT3_HEIGHT(rectangle3_heights[166]), .RECT3_WEIGHT(rectangle3_weights[166]), .FEAT_THRES(feature_thresholds[166]), .FEAT_ABOVE(feature_aboves[166]), .FEAT_BELOW(feature_belows[166])) ac166(.scan_win(scan_win166), .scan_win_std_dev(scan_win_std_dev[166]), .feature_accum(feature_accums[166]));
  accum_calculator #(.RECT1_X(rectangle1_xs[167]), .RECT1_Y(rectangle1_ys[167]), .RECT1_WIDTH(rectangle1_widths[167]), .RECT1_HEIGHT(rectangle1_heights[167]), .RECT1_WEIGHT(rectangle1_weights[167]), .RECT2_X(rectangle2_xs[167]), .RECT2_Y(rectangle2_ys[167]), .RECT2_WIDTH(rectangle2_widths[167]), .RECT2_HEIGHT(rectangle2_heights[167]), .RECT2_WEIGHT(rectangle2_weights[167]), .RECT3_X(rectangle3_xs[167]), .RECT3_Y(rectangle3_ys[167]), .RECT3_WIDTH(rectangle3_widths[167]), .RECT3_HEIGHT(rectangle3_heights[167]), .RECT3_WEIGHT(rectangle3_weights[167]), .FEAT_THRES(feature_thresholds[167]), .FEAT_ABOVE(feature_aboves[167]), .FEAT_BELOW(feature_belows[167])) ac167(.scan_win(scan_win167), .scan_win_std_dev(scan_win_std_dev[167]), .feature_accum(feature_accums[167]));
  accum_calculator #(.RECT1_X(rectangle1_xs[168]), .RECT1_Y(rectangle1_ys[168]), .RECT1_WIDTH(rectangle1_widths[168]), .RECT1_HEIGHT(rectangle1_heights[168]), .RECT1_WEIGHT(rectangle1_weights[168]), .RECT2_X(rectangle2_xs[168]), .RECT2_Y(rectangle2_ys[168]), .RECT2_WIDTH(rectangle2_widths[168]), .RECT2_HEIGHT(rectangle2_heights[168]), .RECT2_WEIGHT(rectangle2_weights[168]), .RECT3_X(rectangle3_xs[168]), .RECT3_Y(rectangle3_ys[168]), .RECT3_WIDTH(rectangle3_widths[168]), .RECT3_HEIGHT(rectangle3_heights[168]), .RECT3_WEIGHT(rectangle3_weights[168]), .FEAT_THRES(feature_thresholds[168]), .FEAT_ABOVE(feature_aboves[168]), .FEAT_BELOW(feature_belows[168])) ac168(.scan_win(scan_win168), .scan_win_std_dev(scan_win_std_dev[168]), .feature_accum(feature_accums[168]));
  accum_calculator #(.RECT1_X(rectangle1_xs[169]), .RECT1_Y(rectangle1_ys[169]), .RECT1_WIDTH(rectangle1_widths[169]), .RECT1_HEIGHT(rectangle1_heights[169]), .RECT1_WEIGHT(rectangle1_weights[169]), .RECT2_X(rectangle2_xs[169]), .RECT2_Y(rectangle2_ys[169]), .RECT2_WIDTH(rectangle2_widths[169]), .RECT2_HEIGHT(rectangle2_heights[169]), .RECT2_WEIGHT(rectangle2_weights[169]), .RECT3_X(rectangle3_xs[169]), .RECT3_Y(rectangle3_ys[169]), .RECT3_WIDTH(rectangle3_widths[169]), .RECT3_HEIGHT(rectangle3_heights[169]), .RECT3_WEIGHT(rectangle3_weights[169]), .FEAT_THRES(feature_thresholds[169]), .FEAT_ABOVE(feature_aboves[169]), .FEAT_BELOW(feature_belows[169])) ac169(.scan_win(scan_win169), .scan_win_std_dev(scan_win_std_dev[169]), .feature_accum(feature_accums[169]));
  accum_calculator #(.RECT1_X(rectangle1_xs[170]), .RECT1_Y(rectangle1_ys[170]), .RECT1_WIDTH(rectangle1_widths[170]), .RECT1_HEIGHT(rectangle1_heights[170]), .RECT1_WEIGHT(rectangle1_weights[170]), .RECT2_X(rectangle2_xs[170]), .RECT2_Y(rectangle2_ys[170]), .RECT2_WIDTH(rectangle2_widths[170]), .RECT2_HEIGHT(rectangle2_heights[170]), .RECT2_WEIGHT(rectangle2_weights[170]), .RECT3_X(rectangle3_xs[170]), .RECT3_Y(rectangle3_ys[170]), .RECT3_WIDTH(rectangle3_widths[170]), .RECT3_HEIGHT(rectangle3_heights[170]), .RECT3_WEIGHT(rectangle3_weights[170]), .FEAT_THRES(feature_thresholds[170]), .FEAT_ABOVE(feature_aboves[170]), .FEAT_BELOW(feature_belows[170])) ac170(.scan_win(scan_win170), .scan_win_std_dev(scan_win_std_dev[170]), .feature_accum(feature_accums[170]));
  accum_calculator #(.RECT1_X(rectangle1_xs[171]), .RECT1_Y(rectangle1_ys[171]), .RECT1_WIDTH(rectangle1_widths[171]), .RECT1_HEIGHT(rectangle1_heights[171]), .RECT1_WEIGHT(rectangle1_weights[171]), .RECT2_X(rectangle2_xs[171]), .RECT2_Y(rectangle2_ys[171]), .RECT2_WIDTH(rectangle2_widths[171]), .RECT2_HEIGHT(rectangle2_heights[171]), .RECT2_WEIGHT(rectangle2_weights[171]), .RECT3_X(rectangle3_xs[171]), .RECT3_Y(rectangle3_ys[171]), .RECT3_WIDTH(rectangle3_widths[171]), .RECT3_HEIGHT(rectangle3_heights[171]), .RECT3_WEIGHT(rectangle3_weights[171]), .FEAT_THRES(feature_thresholds[171]), .FEAT_ABOVE(feature_aboves[171]), .FEAT_BELOW(feature_belows[171])) ac171(.scan_win(scan_win171), .scan_win_std_dev(scan_win_std_dev[171]), .feature_accum(feature_accums[171]));
  accum_calculator #(.RECT1_X(rectangle1_xs[172]), .RECT1_Y(rectangle1_ys[172]), .RECT1_WIDTH(rectangle1_widths[172]), .RECT1_HEIGHT(rectangle1_heights[172]), .RECT1_WEIGHT(rectangle1_weights[172]), .RECT2_X(rectangle2_xs[172]), .RECT2_Y(rectangle2_ys[172]), .RECT2_WIDTH(rectangle2_widths[172]), .RECT2_HEIGHT(rectangle2_heights[172]), .RECT2_WEIGHT(rectangle2_weights[172]), .RECT3_X(rectangle3_xs[172]), .RECT3_Y(rectangle3_ys[172]), .RECT3_WIDTH(rectangle3_widths[172]), .RECT3_HEIGHT(rectangle3_heights[172]), .RECT3_WEIGHT(rectangle3_weights[172]), .FEAT_THRES(feature_thresholds[172]), .FEAT_ABOVE(feature_aboves[172]), .FEAT_BELOW(feature_belows[172])) ac172(.scan_win(scan_win172), .scan_win_std_dev(scan_win_std_dev[172]), .feature_accum(feature_accums[172]));
  accum_calculator #(.RECT1_X(rectangle1_xs[173]), .RECT1_Y(rectangle1_ys[173]), .RECT1_WIDTH(rectangle1_widths[173]), .RECT1_HEIGHT(rectangle1_heights[173]), .RECT1_WEIGHT(rectangle1_weights[173]), .RECT2_X(rectangle2_xs[173]), .RECT2_Y(rectangle2_ys[173]), .RECT2_WIDTH(rectangle2_widths[173]), .RECT2_HEIGHT(rectangle2_heights[173]), .RECT2_WEIGHT(rectangle2_weights[173]), .RECT3_X(rectangle3_xs[173]), .RECT3_Y(rectangle3_ys[173]), .RECT3_WIDTH(rectangle3_widths[173]), .RECT3_HEIGHT(rectangle3_heights[173]), .RECT3_WEIGHT(rectangle3_weights[173]), .FEAT_THRES(feature_thresholds[173]), .FEAT_ABOVE(feature_aboves[173]), .FEAT_BELOW(feature_belows[173])) ac173(.scan_win(scan_win173), .scan_win_std_dev(scan_win_std_dev[173]), .feature_accum(feature_accums[173]));
  accum_calculator #(.RECT1_X(rectangle1_xs[174]), .RECT1_Y(rectangle1_ys[174]), .RECT1_WIDTH(rectangle1_widths[174]), .RECT1_HEIGHT(rectangle1_heights[174]), .RECT1_WEIGHT(rectangle1_weights[174]), .RECT2_X(rectangle2_xs[174]), .RECT2_Y(rectangle2_ys[174]), .RECT2_WIDTH(rectangle2_widths[174]), .RECT2_HEIGHT(rectangle2_heights[174]), .RECT2_WEIGHT(rectangle2_weights[174]), .RECT3_X(rectangle3_xs[174]), .RECT3_Y(rectangle3_ys[174]), .RECT3_WIDTH(rectangle3_widths[174]), .RECT3_HEIGHT(rectangle3_heights[174]), .RECT3_WEIGHT(rectangle3_weights[174]), .FEAT_THRES(feature_thresholds[174]), .FEAT_ABOVE(feature_aboves[174]), .FEAT_BELOW(feature_belows[174])) ac174(.scan_win(scan_win174), .scan_win_std_dev(scan_win_std_dev[174]), .feature_accum(feature_accums[174]));
  accum_calculator #(.RECT1_X(rectangle1_xs[175]), .RECT1_Y(rectangle1_ys[175]), .RECT1_WIDTH(rectangle1_widths[175]), .RECT1_HEIGHT(rectangle1_heights[175]), .RECT1_WEIGHT(rectangle1_weights[175]), .RECT2_X(rectangle2_xs[175]), .RECT2_Y(rectangle2_ys[175]), .RECT2_WIDTH(rectangle2_widths[175]), .RECT2_HEIGHT(rectangle2_heights[175]), .RECT2_WEIGHT(rectangle2_weights[175]), .RECT3_X(rectangle3_xs[175]), .RECT3_Y(rectangle3_ys[175]), .RECT3_WIDTH(rectangle3_widths[175]), .RECT3_HEIGHT(rectangle3_heights[175]), .RECT3_WEIGHT(rectangle3_weights[175]), .FEAT_THRES(feature_thresholds[175]), .FEAT_ABOVE(feature_aboves[175]), .FEAT_BELOW(feature_belows[175])) ac175(.scan_win(scan_win175), .scan_win_std_dev(scan_win_std_dev[175]), .feature_accum(feature_accums[175]));
  accum_calculator #(.RECT1_X(rectangle1_xs[176]), .RECT1_Y(rectangle1_ys[176]), .RECT1_WIDTH(rectangle1_widths[176]), .RECT1_HEIGHT(rectangle1_heights[176]), .RECT1_WEIGHT(rectangle1_weights[176]), .RECT2_X(rectangle2_xs[176]), .RECT2_Y(rectangle2_ys[176]), .RECT2_WIDTH(rectangle2_widths[176]), .RECT2_HEIGHT(rectangle2_heights[176]), .RECT2_WEIGHT(rectangle2_weights[176]), .RECT3_X(rectangle3_xs[176]), .RECT3_Y(rectangle3_ys[176]), .RECT3_WIDTH(rectangle3_widths[176]), .RECT3_HEIGHT(rectangle3_heights[176]), .RECT3_WEIGHT(rectangle3_weights[176]), .FEAT_THRES(feature_thresholds[176]), .FEAT_ABOVE(feature_aboves[176]), .FEAT_BELOW(feature_belows[176])) ac176(.scan_win(scan_win176), .scan_win_std_dev(scan_win_std_dev[176]), .feature_accum(feature_accums[176]));
  accum_calculator #(.RECT1_X(rectangle1_xs[177]), .RECT1_Y(rectangle1_ys[177]), .RECT1_WIDTH(rectangle1_widths[177]), .RECT1_HEIGHT(rectangle1_heights[177]), .RECT1_WEIGHT(rectangle1_weights[177]), .RECT2_X(rectangle2_xs[177]), .RECT2_Y(rectangle2_ys[177]), .RECT2_WIDTH(rectangle2_widths[177]), .RECT2_HEIGHT(rectangle2_heights[177]), .RECT2_WEIGHT(rectangle2_weights[177]), .RECT3_X(rectangle3_xs[177]), .RECT3_Y(rectangle3_ys[177]), .RECT3_WIDTH(rectangle3_widths[177]), .RECT3_HEIGHT(rectangle3_heights[177]), .RECT3_WEIGHT(rectangle3_weights[177]), .FEAT_THRES(feature_thresholds[177]), .FEAT_ABOVE(feature_aboves[177]), .FEAT_BELOW(feature_belows[177])) ac177(.scan_win(scan_win177), .scan_win_std_dev(scan_win_std_dev[177]), .feature_accum(feature_accums[177]));
  accum_calculator #(.RECT1_X(rectangle1_xs[178]), .RECT1_Y(rectangle1_ys[178]), .RECT1_WIDTH(rectangle1_widths[178]), .RECT1_HEIGHT(rectangle1_heights[178]), .RECT1_WEIGHT(rectangle1_weights[178]), .RECT2_X(rectangle2_xs[178]), .RECT2_Y(rectangle2_ys[178]), .RECT2_WIDTH(rectangle2_widths[178]), .RECT2_HEIGHT(rectangle2_heights[178]), .RECT2_WEIGHT(rectangle2_weights[178]), .RECT3_X(rectangle3_xs[178]), .RECT3_Y(rectangle3_ys[178]), .RECT3_WIDTH(rectangle3_widths[178]), .RECT3_HEIGHT(rectangle3_heights[178]), .RECT3_WEIGHT(rectangle3_weights[178]), .FEAT_THRES(feature_thresholds[178]), .FEAT_ABOVE(feature_aboves[178]), .FEAT_BELOW(feature_belows[178])) ac178(.scan_win(scan_win178), .scan_win_std_dev(scan_win_std_dev[178]), .feature_accum(feature_accums[178]));
  accum_calculator #(.RECT1_X(rectangle1_xs[179]), .RECT1_Y(rectangle1_ys[179]), .RECT1_WIDTH(rectangle1_widths[179]), .RECT1_HEIGHT(rectangle1_heights[179]), .RECT1_WEIGHT(rectangle1_weights[179]), .RECT2_X(rectangle2_xs[179]), .RECT2_Y(rectangle2_ys[179]), .RECT2_WIDTH(rectangle2_widths[179]), .RECT2_HEIGHT(rectangle2_heights[179]), .RECT2_WEIGHT(rectangle2_weights[179]), .RECT3_X(rectangle3_xs[179]), .RECT3_Y(rectangle3_ys[179]), .RECT3_WIDTH(rectangle3_widths[179]), .RECT3_HEIGHT(rectangle3_heights[179]), .RECT3_WEIGHT(rectangle3_weights[179]), .FEAT_THRES(feature_thresholds[179]), .FEAT_ABOVE(feature_aboves[179]), .FEAT_BELOW(feature_belows[179])) ac179(.scan_win(scan_win179), .scan_win_std_dev(scan_win_std_dev[179]), .feature_accum(feature_accums[179]));
  accum_calculator #(.RECT1_X(rectangle1_xs[180]), .RECT1_Y(rectangle1_ys[180]), .RECT1_WIDTH(rectangle1_widths[180]), .RECT1_HEIGHT(rectangle1_heights[180]), .RECT1_WEIGHT(rectangle1_weights[180]), .RECT2_X(rectangle2_xs[180]), .RECT2_Y(rectangle2_ys[180]), .RECT2_WIDTH(rectangle2_widths[180]), .RECT2_HEIGHT(rectangle2_heights[180]), .RECT2_WEIGHT(rectangle2_weights[180]), .RECT3_X(rectangle3_xs[180]), .RECT3_Y(rectangle3_ys[180]), .RECT3_WIDTH(rectangle3_widths[180]), .RECT3_HEIGHT(rectangle3_heights[180]), .RECT3_WEIGHT(rectangle3_weights[180]), .FEAT_THRES(feature_thresholds[180]), .FEAT_ABOVE(feature_aboves[180]), .FEAT_BELOW(feature_belows[180])) ac180(.scan_win(scan_win180), .scan_win_std_dev(scan_win_std_dev[180]), .feature_accum(feature_accums[180]));
  accum_calculator #(.RECT1_X(rectangle1_xs[181]), .RECT1_Y(rectangle1_ys[181]), .RECT1_WIDTH(rectangle1_widths[181]), .RECT1_HEIGHT(rectangle1_heights[181]), .RECT1_WEIGHT(rectangle1_weights[181]), .RECT2_X(rectangle2_xs[181]), .RECT2_Y(rectangle2_ys[181]), .RECT2_WIDTH(rectangle2_widths[181]), .RECT2_HEIGHT(rectangle2_heights[181]), .RECT2_WEIGHT(rectangle2_weights[181]), .RECT3_X(rectangle3_xs[181]), .RECT3_Y(rectangle3_ys[181]), .RECT3_WIDTH(rectangle3_widths[181]), .RECT3_HEIGHT(rectangle3_heights[181]), .RECT3_WEIGHT(rectangle3_weights[181]), .FEAT_THRES(feature_thresholds[181]), .FEAT_ABOVE(feature_aboves[181]), .FEAT_BELOW(feature_belows[181])) ac181(.scan_win(scan_win181), .scan_win_std_dev(scan_win_std_dev[181]), .feature_accum(feature_accums[181]));
  accum_calculator #(.RECT1_X(rectangle1_xs[182]), .RECT1_Y(rectangle1_ys[182]), .RECT1_WIDTH(rectangle1_widths[182]), .RECT1_HEIGHT(rectangle1_heights[182]), .RECT1_WEIGHT(rectangle1_weights[182]), .RECT2_X(rectangle2_xs[182]), .RECT2_Y(rectangle2_ys[182]), .RECT2_WIDTH(rectangle2_widths[182]), .RECT2_HEIGHT(rectangle2_heights[182]), .RECT2_WEIGHT(rectangle2_weights[182]), .RECT3_X(rectangle3_xs[182]), .RECT3_Y(rectangle3_ys[182]), .RECT3_WIDTH(rectangle3_widths[182]), .RECT3_HEIGHT(rectangle3_heights[182]), .RECT3_WEIGHT(rectangle3_weights[182]), .FEAT_THRES(feature_thresholds[182]), .FEAT_ABOVE(feature_aboves[182]), .FEAT_BELOW(feature_belows[182])) ac182(.scan_win(scan_win182), .scan_win_std_dev(scan_win_std_dev[182]), .feature_accum(feature_accums[182]));
  accum_calculator #(.RECT1_X(rectangle1_xs[183]), .RECT1_Y(rectangle1_ys[183]), .RECT1_WIDTH(rectangle1_widths[183]), .RECT1_HEIGHT(rectangle1_heights[183]), .RECT1_WEIGHT(rectangle1_weights[183]), .RECT2_X(rectangle2_xs[183]), .RECT2_Y(rectangle2_ys[183]), .RECT2_WIDTH(rectangle2_widths[183]), .RECT2_HEIGHT(rectangle2_heights[183]), .RECT2_WEIGHT(rectangle2_weights[183]), .RECT3_X(rectangle3_xs[183]), .RECT3_Y(rectangle3_ys[183]), .RECT3_WIDTH(rectangle3_widths[183]), .RECT3_HEIGHT(rectangle3_heights[183]), .RECT3_WEIGHT(rectangle3_weights[183]), .FEAT_THRES(feature_thresholds[183]), .FEAT_ABOVE(feature_aboves[183]), .FEAT_BELOW(feature_belows[183])) ac183(.scan_win(scan_win183), .scan_win_std_dev(scan_win_std_dev[183]), .feature_accum(feature_accums[183]));
  accum_calculator #(.RECT1_X(rectangle1_xs[184]), .RECT1_Y(rectangle1_ys[184]), .RECT1_WIDTH(rectangle1_widths[184]), .RECT1_HEIGHT(rectangle1_heights[184]), .RECT1_WEIGHT(rectangle1_weights[184]), .RECT2_X(rectangle2_xs[184]), .RECT2_Y(rectangle2_ys[184]), .RECT2_WIDTH(rectangle2_widths[184]), .RECT2_HEIGHT(rectangle2_heights[184]), .RECT2_WEIGHT(rectangle2_weights[184]), .RECT3_X(rectangle3_xs[184]), .RECT3_Y(rectangle3_ys[184]), .RECT3_WIDTH(rectangle3_widths[184]), .RECT3_HEIGHT(rectangle3_heights[184]), .RECT3_WEIGHT(rectangle3_weights[184]), .FEAT_THRES(feature_thresholds[184]), .FEAT_ABOVE(feature_aboves[184]), .FEAT_BELOW(feature_belows[184])) ac184(.scan_win(scan_win184), .scan_win_std_dev(scan_win_std_dev[184]), .feature_accum(feature_accums[184]));
  accum_calculator #(.RECT1_X(rectangle1_xs[185]), .RECT1_Y(rectangle1_ys[185]), .RECT1_WIDTH(rectangle1_widths[185]), .RECT1_HEIGHT(rectangle1_heights[185]), .RECT1_WEIGHT(rectangle1_weights[185]), .RECT2_X(rectangle2_xs[185]), .RECT2_Y(rectangle2_ys[185]), .RECT2_WIDTH(rectangle2_widths[185]), .RECT2_HEIGHT(rectangle2_heights[185]), .RECT2_WEIGHT(rectangle2_weights[185]), .RECT3_X(rectangle3_xs[185]), .RECT3_Y(rectangle3_ys[185]), .RECT3_WIDTH(rectangle3_widths[185]), .RECT3_HEIGHT(rectangle3_heights[185]), .RECT3_WEIGHT(rectangle3_weights[185]), .FEAT_THRES(feature_thresholds[185]), .FEAT_ABOVE(feature_aboves[185]), .FEAT_BELOW(feature_belows[185])) ac185(.scan_win(scan_win185), .scan_win_std_dev(scan_win_std_dev[185]), .feature_accum(feature_accums[185]));
  accum_calculator #(.RECT1_X(rectangle1_xs[186]), .RECT1_Y(rectangle1_ys[186]), .RECT1_WIDTH(rectangle1_widths[186]), .RECT1_HEIGHT(rectangle1_heights[186]), .RECT1_WEIGHT(rectangle1_weights[186]), .RECT2_X(rectangle2_xs[186]), .RECT2_Y(rectangle2_ys[186]), .RECT2_WIDTH(rectangle2_widths[186]), .RECT2_HEIGHT(rectangle2_heights[186]), .RECT2_WEIGHT(rectangle2_weights[186]), .RECT3_X(rectangle3_xs[186]), .RECT3_Y(rectangle3_ys[186]), .RECT3_WIDTH(rectangle3_widths[186]), .RECT3_HEIGHT(rectangle3_heights[186]), .RECT3_WEIGHT(rectangle3_weights[186]), .FEAT_THRES(feature_thresholds[186]), .FEAT_ABOVE(feature_aboves[186]), .FEAT_BELOW(feature_belows[186])) ac186(.scan_win(scan_win186), .scan_win_std_dev(scan_win_std_dev[186]), .feature_accum(feature_accums[186]));
  accum_calculator #(.RECT1_X(rectangle1_xs[187]), .RECT1_Y(rectangle1_ys[187]), .RECT1_WIDTH(rectangle1_widths[187]), .RECT1_HEIGHT(rectangle1_heights[187]), .RECT1_WEIGHT(rectangle1_weights[187]), .RECT2_X(rectangle2_xs[187]), .RECT2_Y(rectangle2_ys[187]), .RECT2_WIDTH(rectangle2_widths[187]), .RECT2_HEIGHT(rectangle2_heights[187]), .RECT2_WEIGHT(rectangle2_weights[187]), .RECT3_X(rectangle3_xs[187]), .RECT3_Y(rectangle3_ys[187]), .RECT3_WIDTH(rectangle3_widths[187]), .RECT3_HEIGHT(rectangle3_heights[187]), .RECT3_WEIGHT(rectangle3_weights[187]), .FEAT_THRES(feature_thresholds[187]), .FEAT_ABOVE(feature_aboves[187]), .FEAT_BELOW(feature_belows[187])) ac187(.scan_win(scan_win187), .scan_win_std_dev(scan_win_std_dev[187]), .feature_accum(feature_accums[187]));
  accum_calculator #(.RECT1_X(rectangle1_xs[188]), .RECT1_Y(rectangle1_ys[188]), .RECT1_WIDTH(rectangle1_widths[188]), .RECT1_HEIGHT(rectangle1_heights[188]), .RECT1_WEIGHT(rectangle1_weights[188]), .RECT2_X(rectangle2_xs[188]), .RECT2_Y(rectangle2_ys[188]), .RECT2_WIDTH(rectangle2_widths[188]), .RECT2_HEIGHT(rectangle2_heights[188]), .RECT2_WEIGHT(rectangle2_weights[188]), .RECT3_X(rectangle3_xs[188]), .RECT3_Y(rectangle3_ys[188]), .RECT3_WIDTH(rectangle3_widths[188]), .RECT3_HEIGHT(rectangle3_heights[188]), .RECT3_WEIGHT(rectangle3_weights[188]), .FEAT_THRES(feature_thresholds[188]), .FEAT_ABOVE(feature_aboves[188]), .FEAT_BELOW(feature_belows[188])) ac188(.scan_win(scan_win188), .scan_win_std_dev(scan_win_std_dev[188]), .feature_accum(feature_accums[188]));
  accum_calculator #(.RECT1_X(rectangle1_xs[189]), .RECT1_Y(rectangle1_ys[189]), .RECT1_WIDTH(rectangle1_widths[189]), .RECT1_HEIGHT(rectangle1_heights[189]), .RECT1_WEIGHT(rectangle1_weights[189]), .RECT2_X(rectangle2_xs[189]), .RECT2_Y(rectangle2_ys[189]), .RECT2_WIDTH(rectangle2_widths[189]), .RECT2_HEIGHT(rectangle2_heights[189]), .RECT2_WEIGHT(rectangle2_weights[189]), .RECT3_X(rectangle3_xs[189]), .RECT3_Y(rectangle3_ys[189]), .RECT3_WIDTH(rectangle3_widths[189]), .RECT3_HEIGHT(rectangle3_heights[189]), .RECT3_WEIGHT(rectangle3_weights[189]), .FEAT_THRES(feature_thresholds[189]), .FEAT_ABOVE(feature_aboves[189]), .FEAT_BELOW(feature_belows[189])) ac189(.scan_win(scan_win189), .scan_win_std_dev(scan_win_std_dev[189]), .feature_accum(feature_accums[189]));
  accum_calculator #(.RECT1_X(rectangle1_xs[190]), .RECT1_Y(rectangle1_ys[190]), .RECT1_WIDTH(rectangle1_widths[190]), .RECT1_HEIGHT(rectangle1_heights[190]), .RECT1_WEIGHT(rectangle1_weights[190]), .RECT2_X(rectangle2_xs[190]), .RECT2_Y(rectangle2_ys[190]), .RECT2_WIDTH(rectangle2_widths[190]), .RECT2_HEIGHT(rectangle2_heights[190]), .RECT2_WEIGHT(rectangle2_weights[190]), .RECT3_X(rectangle3_xs[190]), .RECT3_Y(rectangle3_ys[190]), .RECT3_WIDTH(rectangle3_widths[190]), .RECT3_HEIGHT(rectangle3_heights[190]), .RECT3_WEIGHT(rectangle3_weights[190]), .FEAT_THRES(feature_thresholds[190]), .FEAT_ABOVE(feature_aboves[190]), .FEAT_BELOW(feature_belows[190])) ac190(.scan_win(scan_win190), .scan_win_std_dev(scan_win_std_dev[190]), .feature_accum(feature_accums[190]));
  accum_calculator #(.RECT1_X(rectangle1_xs[191]), .RECT1_Y(rectangle1_ys[191]), .RECT1_WIDTH(rectangle1_widths[191]), .RECT1_HEIGHT(rectangle1_heights[191]), .RECT1_WEIGHT(rectangle1_weights[191]), .RECT2_X(rectangle2_xs[191]), .RECT2_Y(rectangle2_ys[191]), .RECT2_WIDTH(rectangle2_widths[191]), .RECT2_HEIGHT(rectangle2_heights[191]), .RECT2_WEIGHT(rectangle2_weights[191]), .RECT3_X(rectangle3_xs[191]), .RECT3_Y(rectangle3_ys[191]), .RECT3_WIDTH(rectangle3_widths[191]), .RECT3_HEIGHT(rectangle3_heights[191]), .RECT3_WEIGHT(rectangle3_weights[191]), .FEAT_THRES(feature_thresholds[191]), .FEAT_ABOVE(feature_aboves[191]), .FEAT_BELOW(feature_belows[191])) ac191(.scan_win(scan_win191), .scan_win_std_dev(scan_win_std_dev[191]), .feature_accum(feature_accums[191]));
  accum_calculator #(.RECT1_X(rectangle1_xs[192]), .RECT1_Y(rectangle1_ys[192]), .RECT1_WIDTH(rectangle1_widths[192]), .RECT1_HEIGHT(rectangle1_heights[192]), .RECT1_WEIGHT(rectangle1_weights[192]), .RECT2_X(rectangle2_xs[192]), .RECT2_Y(rectangle2_ys[192]), .RECT2_WIDTH(rectangle2_widths[192]), .RECT2_HEIGHT(rectangle2_heights[192]), .RECT2_WEIGHT(rectangle2_weights[192]), .RECT3_X(rectangle3_xs[192]), .RECT3_Y(rectangle3_ys[192]), .RECT3_WIDTH(rectangle3_widths[192]), .RECT3_HEIGHT(rectangle3_heights[192]), .RECT3_WEIGHT(rectangle3_weights[192]), .FEAT_THRES(feature_thresholds[192]), .FEAT_ABOVE(feature_aboves[192]), .FEAT_BELOW(feature_belows[192])) ac192(.scan_win(scan_win192), .scan_win_std_dev(scan_win_std_dev[192]), .feature_accum(feature_accums[192]));
  accum_calculator #(.RECT1_X(rectangle1_xs[193]), .RECT1_Y(rectangle1_ys[193]), .RECT1_WIDTH(rectangle1_widths[193]), .RECT1_HEIGHT(rectangle1_heights[193]), .RECT1_WEIGHT(rectangle1_weights[193]), .RECT2_X(rectangle2_xs[193]), .RECT2_Y(rectangle2_ys[193]), .RECT2_WIDTH(rectangle2_widths[193]), .RECT2_HEIGHT(rectangle2_heights[193]), .RECT2_WEIGHT(rectangle2_weights[193]), .RECT3_X(rectangle3_xs[193]), .RECT3_Y(rectangle3_ys[193]), .RECT3_WIDTH(rectangle3_widths[193]), .RECT3_HEIGHT(rectangle3_heights[193]), .RECT3_WEIGHT(rectangle3_weights[193]), .FEAT_THRES(feature_thresholds[193]), .FEAT_ABOVE(feature_aboves[193]), .FEAT_BELOW(feature_belows[193])) ac193(.scan_win(scan_win193), .scan_win_std_dev(scan_win_std_dev[193]), .feature_accum(feature_accums[193]));
  accum_calculator #(.RECT1_X(rectangle1_xs[194]), .RECT1_Y(rectangle1_ys[194]), .RECT1_WIDTH(rectangle1_widths[194]), .RECT1_HEIGHT(rectangle1_heights[194]), .RECT1_WEIGHT(rectangle1_weights[194]), .RECT2_X(rectangle2_xs[194]), .RECT2_Y(rectangle2_ys[194]), .RECT2_WIDTH(rectangle2_widths[194]), .RECT2_HEIGHT(rectangle2_heights[194]), .RECT2_WEIGHT(rectangle2_weights[194]), .RECT3_X(rectangle3_xs[194]), .RECT3_Y(rectangle3_ys[194]), .RECT3_WIDTH(rectangle3_widths[194]), .RECT3_HEIGHT(rectangle3_heights[194]), .RECT3_WEIGHT(rectangle3_weights[194]), .FEAT_THRES(feature_thresholds[194]), .FEAT_ABOVE(feature_aboves[194]), .FEAT_BELOW(feature_belows[194])) ac194(.scan_win(scan_win194), .scan_win_std_dev(scan_win_std_dev[194]), .feature_accum(feature_accums[194]));
  accum_calculator #(.RECT1_X(rectangle1_xs[195]), .RECT1_Y(rectangle1_ys[195]), .RECT1_WIDTH(rectangle1_widths[195]), .RECT1_HEIGHT(rectangle1_heights[195]), .RECT1_WEIGHT(rectangle1_weights[195]), .RECT2_X(rectangle2_xs[195]), .RECT2_Y(rectangle2_ys[195]), .RECT2_WIDTH(rectangle2_widths[195]), .RECT2_HEIGHT(rectangle2_heights[195]), .RECT2_WEIGHT(rectangle2_weights[195]), .RECT3_X(rectangle3_xs[195]), .RECT3_Y(rectangle3_ys[195]), .RECT3_WIDTH(rectangle3_widths[195]), .RECT3_HEIGHT(rectangle3_heights[195]), .RECT3_WEIGHT(rectangle3_weights[195]), .FEAT_THRES(feature_thresholds[195]), .FEAT_ABOVE(feature_aboves[195]), .FEAT_BELOW(feature_belows[195])) ac195(.scan_win(scan_win195), .scan_win_std_dev(scan_win_std_dev[195]), .feature_accum(feature_accums[195]));
  accum_calculator #(.RECT1_X(rectangle1_xs[196]), .RECT1_Y(rectangle1_ys[196]), .RECT1_WIDTH(rectangle1_widths[196]), .RECT1_HEIGHT(rectangle1_heights[196]), .RECT1_WEIGHT(rectangle1_weights[196]), .RECT2_X(rectangle2_xs[196]), .RECT2_Y(rectangle2_ys[196]), .RECT2_WIDTH(rectangle2_widths[196]), .RECT2_HEIGHT(rectangle2_heights[196]), .RECT2_WEIGHT(rectangle2_weights[196]), .RECT3_X(rectangle3_xs[196]), .RECT3_Y(rectangle3_ys[196]), .RECT3_WIDTH(rectangle3_widths[196]), .RECT3_HEIGHT(rectangle3_heights[196]), .RECT3_WEIGHT(rectangle3_weights[196]), .FEAT_THRES(feature_thresholds[196]), .FEAT_ABOVE(feature_aboves[196]), .FEAT_BELOW(feature_belows[196])) ac196(.scan_win(scan_win196), .scan_win_std_dev(scan_win_std_dev[196]), .feature_accum(feature_accums[196]));
  accum_calculator #(.RECT1_X(rectangle1_xs[197]), .RECT1_Y(rectangle1_ys[197]), .RECT1_WIDTH(rectangle1_widths[197]), .RECT1_HEIGHT(rectangle1_heights[197]), .RECT1_WEIGHT(rectangle1_weights[197]), .RECT2_X(rectangle2_xs[197]), .RECT2_Y(rectangle2_ys[197]), .RECT2_WIDTH(rectangle2_widths[197]), .RECT2_HEIGHT(rectangle2_heights[197]), .RECT2_WEIGHT(rectangle2_weights[197]), .RECT3_X(rectangle3_xs[197]), .RECT3_Y(rectangle3_ys[197]), .RECT3_WIDTH(rectangle3_widths[197]), .RECT3_HEIGHT(rectangle3_heights[197]), .RECT3_WEIGHT(rectangle3_weights[197]), .FEAT_THRES(feature_thresholds[197]), .FEAT_ABOVE(feature_aboves[197]), .FEAT_BELOW(feature_belows[197])) ac197(.scan_win(scan_win197), .scan_win_std_dev(scan_win_std_dev[197]), .feature_accum(feature_accums[197]));
  accum_calculator #(.RECT1_X(rectangle1_xs[198]), .RECT1_Y(rectangle1_ys[198]), .RECT1_WIDTH(rectangle1_widths[198]), .RECT1_HEIGHT(rectangle1_heights[198]), .RECT1_WEIGHT(rectangle1_weights[198]), .RECT2_X(rectangle2_xs[198]), .RECT2_Y(rectangle2_ys[198]), .RECT2_WIDTH(rectangle2_widths[198]), .RECT2_HEIGHT(rectangle2_heights[198]), .RECT2_WEIGHT(rectangle2_weights[198]), .RECT3_X(rectangle3_xs[198]), .RECT3_Y(rectangle3_ys[198]), .RECT3_WIDTH(rectangle3_widths[198]), .RECT3_HEIGHT(rectangle3_heights[198]), .RECT3_WEIGHT(rectangle3_weights[198]), .FEAT_THRES(feature_thresholds[198]), .FEAT_ABOVE(feature_aboves[198]), .FEAT_BELOW(feature_belows[198])) ac198(.scan_win(scan_win198), .scan_win_std_dev(scan_win_std_dev[198]), .feature_accum(feature_accums[198]));
  accum_calculator #(.RECT1_X(rectangle1_xs[199]), .RECT1_Y(rectangle1_ys[199]), .RECT1_WIDTH(rectangle1_widths[199]), .RECT1_HEIGHT(rectangle1_heights[199]), .RECT1_WEIGHT(rectangle1_weights[199]), .RECT2_X(rectangle2_xs[199]), .RECT2_Y(rectangle2_ys[199]), .RECT2_WIDTH(rectangle2_widths[199]), .RECT2_HEIGHT(rectangle2_heights[199]), .RECT2_WEIGHT(rectangle2_weights[199]), .RECT3_X(rectangle3_xs[199]), .RECT3_Y(rectangle3_ys[199]), .RECT3_WIDTH(rectangle3_widths[199]), .RECT3_HEIGHT(rectangle3_heights[199]), .RECT3_WEIGHT(rectangle3_weights[199]), .FEAT_THRES(feature_thresholds[199]), .FEAT_ABOVE(feature_aboves[199]), .FEAT_BELOW(feature_belows[199])) ac199(.scan_win(scan_win199), .scan_win_std_dev(scan_win_std_dev[199]), .feature_accum(feature_accums[199]));
  accum_calculator #(.RECT1_X(rectangle1_xs[200]), .RECT1_Y(rectangle1_ys[200]), .RECT1_WIDTH(rectangle1_widths[200]), .RECT1_HEIGHT(rectangle1_heights[200]), .RECT1_WEIGHT(rectangle1_weights[200]), .RECT2_X(rectangle2_xs[200]), .RECT2_Y(rectangle2_ys[200]), .RECT2_WIDTH(rectangle2_widths[200]), .RECT2_HEIGHT(rectangle2_heights[200]), .RECT2_WEIGHT(rectangle2_weights[200]), .RECT3_X(rectangle3_xs[200]), .RECT3_Y(rectangle3_ys[200]), .RECT3_WIDTH(rectangle3_widths[200]), .RECT3_HEIGHT(rectangle3_heights[200]), .RECT3_WEIGHT(rectangle3_weights[200]), .FEAT_THRES(feature_thresholds[200]), .FEAT_ABOVE(feature_aboves[200]), .FEAT_BELOW(feature_belows[200])) ac200(.scan_win(scan_win200), .scan_win_std_dev(scan_win_std_dev[200]), .feature_accum(feature_accums[200]));
  accum_calculator #(.RECT1_X(rectangle1_xs[201]), .RECT1_Y(rectangle1_ys[201]), .RECT1_WIDTH(rectangle1_widths[201]), .RECT1_HEIGHT(rectangle1_heights[201]), .RECT1_WEIGHT(rectangle1_weights[201]), .RECT2_X(rectangle2_xs[201]), .RECT2_Y(rectangle2_ys[201]), .RECT2_WIDTH(rectangle2_widths[201]), .RECT2_HEIGHT(rectangle2_heights[201]), .RECT2_WEIGHT(rectangle2_weights[201]), .RECT3_X(rectangle3_xs[201]), .RECT3_Y(rectangle3_ys[201]), .RECT3_WIDTH(rectangle3_widths[201]), .RECT3_HEIGHT(rectangle3_heights[201]), .RECT3_WEIGHT(rectangle3_weights[201]), .FEAT_THRES(feature_thresholds[201]), .FEAT_ABOVE(feature_aboves[201]), .FEAT_BELOW(feature_belows[201])) ac201(.scan_win(scan_win201), .scan_win_std_dev(scan_win_std_dev[201]), .feature_accum(feature_accums[201]));
  accum_calculator #(.RECT1_X(rectangle1_xs[202]), .RECT1_Y(rectangle1_ys[202]), .RECT1_WIDTH(rectangle1_widths[202]), .RECT1_HEIGHT(rectangle1_heights[202]), .RECT1_WEIGHT(rectangle1_weights[202]), .RECT2_X(rectangle2_xs[202]), .RECT2_Y(rectangle2_ys[202]), .RECT2_WIDTH(rectangle2_widths[202]), .RECT2_HEIGHT(rectangle2_heights[202]), .RECT2_WEIGHT(rectangle2_weights[202]), .RECT3_X(rectangle3_xs[202]), .RECT3_Y(rectangle3_ys[202]), .RECT3_WIDTH(rectangle3_widths[202]), .RECT3_HEIGHT(rectangle3_heights[202]), .RECT3_WEIGHT(rectangle3_weights[202]), .FEAT_THRES(feature_thresholds[202]), .FEAT_ABOVE(feature_aboves[202]), .FEAT_BELOW(feature_belows[202])) ac202(.scan_win(scan_win202), .scan_win_std_dev(scan_win_std_dev[202]), .feature_accum(feature_accums[202]));
  accum_calculator #(.RECT1_X(rectangle1_xs[203]), .RECT1_Y(rectangle1_ys[203]), .RECT1_WIDTH(rectangle1_widths[203]), .RECT1_HEIGHT(rectangle1_heights[203]), .RECT1_WEIGHT(rectangle1_weights[203]), .RECT2_X(rectangle2_xs[203]), .RECT2_Y(rectangle2_ys[203]), .RECT2_WIDTH(rectangle2_widths[203]), .RECT2_HEIGHT(rectangle2_heights[203]), .RECT2_WEIGHT(rectangle2_weights[203]), .RECT3_X(rectangle3_xs[203]), .RECT3_Y(rectangle3_ys[203]), .RECT3_WIDTH(rectangle3_widths[203]), .RECT3_HEIGHT(rectangle3_heights[203]), .RECT3_WEIGHT(rectangle3_weights[203]), .FEAT_THRES(feature_thresholds[203]), .FEAT_ABOVE(feature_aboves[203]), .FEAT_BELOW(feature_belows[203])) ac203(.scan_win(scan_win203), .scan_win_std_dev(scan_win_std_dev[203]), .feature_accum(feature_accums[203]));
  accum_calculator #(.RECT1_X(rectangle1_xs[204]), .RECT1_Y(rectangle1_ys[204]), .RECT1_WIDTH(rectangle1_widths[204]), .RECT1_HEIGHT(rectangle1_heights[204]), .RECT1_WEIGHT(rectangle1_weights[204]), .RECT2_X(rectangle2_xs[204]), .RECT2_Y(rectangle2_ys[204]), .RECT2_WIDTH(rectangle2_widths[204]), .RECT2_HEIGHT(rectangle2_heights[204]), .RECT2_WEIGHT(rectangle2_weights[204]), .RECT3_X(rectangle3_xs[204]), .RECT3_Y(rectangle3_ys[204]), .RECT3_WIDTH(rectangle3_widths[204]), .RECT3_HEIGHT(rectangle3_heights[204]), .RECT3_WEIGHT(rectangle3_weights[204]), .FEAT_THRES(feature_thresholds[204]), .FEAT_ABOVE(feature_aboves[204]), .FEAT_BELOW(feature_belows[204])) ac204(.scan_win(scan_win204), .scan_win_std_dev(scan_win_std_dev[204]), .feature_accum(feature_accums[204]));
  accum_calculator #(.RECT1_X(rectangle1_xs[205]), .RECT1_Y(rectangle1_ys[205]), .RECT1_WIDTH(rectangle1_widths[205]), .RECT1_HEIGHT(rectangle1_heights[205]), .RECT1_WEIGHT(rectangle1_weights[205]), .RECT2_X(rectangle2_xs[205]), .RECT2_Y(rectangle2_ys[205]), .RECT2_WIDTH(rectangle2_widths[205]), .RECT2_HEIGHT(rectangle2_heights[205]), .RECT2_WEIGHT(rectangle2_weights[205]), .RECT3_X(rectangle3_xs[205]), .RECT3_Y(rectangle3_ys[205]), .RECT3_WIDTH(rectangle3_widths[205]), .RECT3_HEIGHT(rectangle3_heights[205]), .RECT3_WEIGHT(rectangle3_weights[205]), .FEAT_THRES(feature_thresholds[205]), .FEAT_ABOVE(feature_aboves[205]), .FEAT_BELOW(feature_belows[205])) ac205(.scan_win(scan_win205), .scan_win_std_dev(scan_win_std_dev[205]), .feature_accum(feature_accums[205]));
  accum_calculator #(.RECT1_X(rectangle1_xs[206]), .RECT1_Y(rectangle1_ys[206]), .RECT1_WIDTH(rectangle1_widths[206]), .RECT1_HEIGHT(rectangle1_heights[206]), .RECT1_WEIGHT(rectangle1_weights[206]), .RECT2_X(rectangle2_xs[206]), .RECT2_Y(rectangle2_ys[206]), .RECT2_WIDTH(rectangle2_widths[206]), .RECT2_HEIGHT(rectangle2_heights[206]), .RECT2_WEIGHT(rectangle2_weights[206]), .RECT3_X(rectangle3_xs[206]), .RECT3_Y(rectangle3_ys[206]), .RECT3_WIDTH(rectangle3_widths[206]), .RECT3_HEIGHT(rectangle3_heights[206]), .RECT3_WEIGHT(rectangle3_weights[206]), .FEAT_THRES(feature_thresholds[206]), .FEAT_ABOVE(feature_aboves[206]), .FEAT_BELOW(feature_belows[206])) ac206(.scan_win(scan_win206), .scan_win_std_dev(scan_win_std_dev[206]), .feature_accum(feature_accums[206]));
  accum_calculator #(.RECT1_X(rectangle1_xs[207]), .RECT1_Y(rectangle1_ys[207]), .RECT1_WIDTH(rectangle1_widths[207]), .RECT1_HEIGHT(rectangle1_heights[207]), .RECT1_WEIGHT(rectangle1_weights[207]), .RECT2_X(rectangle2_xs[207]), .RECT2_Y(rectangle2_ys[207]), .RECT2_WIDTH(rectangle2_widths[207]), .RECT2_HEIGHT(rectangle2_heights[207]), .RECT2_WEIGHT(rectangle2_weights[207]), .RECT3_X(rectangle3_xs[207]), .RECT3_Y(rectangle3_ys[207]), .RECT3_WIDTH(rectangle3_widths[207]), .RECT3_HEIGHT(rectangle3_heights[207]), .RECT3_WEIGHT(rectangle3_weights[207]), .FEAT_THRES(feature_thresholds[207]), .FEAT_ABOVE(feature_aboves[207]), .FEAT_BELOW(feature_belows[207])) ac207(.scan_win(scan_win207), .scan_win_std_dev(scan_win_std_dev[207]), .feature_accum(feature_accums[207]));
  accum_calculator #(.RECT1_X(rectangle1_xs[208]), .RECT1_Y(rectangle1_ys[208]), .RECT1_WIDTH(rectangle1_widths[208]), .RECT1_HEIGHT(rectangle1_heights[208]), .RECT1_WEIGHT(rectangle1_weights[208]), .RECT2_X(rectangle2_xs[208]), .RECT2_Y(rectangle2_ys[208]), .RECT2_WIDTH(rectangle2_widths[208]), .RECT2_HEIGHT(rectangle2_heights[208]), .RECT2_WEIGHT(rectangle2_weights[208]), .RECT3_X(rectangle3_xs[208]), .RECT3_Y(rectangle3_ys[208]), .RECT3_WIDTH(rectangle3_widths[208]), .RECT3_HEIGHT(rectangle3_heights[208]), .RECT3_WEIGHT(rectangle3_weights[208]), .FEAT_THRES(feature_thresholds[208]), .FEAT_ABOVE(feature_aboves[208]), .FEAT_BELOW(feature_belows[208])) ac208(.scan_win(scan_win208), .scan_win_std_dev(scan_win_std_dev[208]), .feature_accum(feature_accums[208]));
  accum_calculator #(.RECT1_X(rectangle1_xs[209]), .RECT1_Y(rectangle1_ys[209]), .RECT1_WIDTH(rectangle1_widths[209]), .RECT1_HEIGHT(rectangle1_heights[209]), .RECT1_WEIGHT(rectangle1_weights[209]), .RECT2_X(rectangle2_xs[209]), .RECT2_Y(rectangle2_ys[209]), .RECT2_WIDTH(rectangle2_widths[209]), .RECT2_HEIGHT(rectangle2_heights[209]), .RECT2_WEIGHT(rectangle2_weights[209]), .RECT3_X(rectangle3_xs[209]), .RECT3_Y(rectangle3_ys[209]), .RECT3_WIDTH(rectangle3_widths[209]), .RECT3_HEIGHT(rectangle3_heights[209]), .RECT3_WEIGHT(rectangle3_weights[209]), .FEAT_THRES(feature_thresholds[209]), .FEAT_ABOVE(feature_aboves[209]), .FEAT_BELOW(feature_belows[209])) ac209(.scan_win(scan_win209), .scan_win_std_dev(scan_win_std_dev[209]), .feature_accum(feature_accums[209]));
  accum_calculator #(.RECT1_X(rectangle1_xs[210]), .RECT1_Y(rectangle1_ys[210]), .RECT1_WIDTH(rectangle1_widths[210]), .RECT1_HEIGHT(rectangle1_heights[210]), .RECT1_WEIGHT(rectangle1_weights[210]), .RECT2_X(rectangle2_xs[210]), .RECT2_Y(rectangle2_ys[210]), .RECT2_WIDTH(rectangle2_widths[210]), .RECT2_HEIGHT(rectangle2_heights[210]), .RECT2_WEIGHT(rectangle2_weights[210]), .RECT3_X(rectangle3_xs[210]), .RECT3_Y(rectangle3_ys[210]), .RECT3_WIDTH(rectangle3_widths[210]), .RECT3_HEIGHT(rectangle3_heights[210]), .RECT3_WEIGHT(rectangle3_weights[210]), .FEAT_THRES(feature_thresholds[210]), .FEAT_ABOVE(feature_aboves[210]), .FEAT_BELOW(feature_belows[210])) ac210(.scan_win(scan_win210), .scan_win_std_dev(scan_win_std_dev[210]), .feature_accum(feature_accums[210]));
  accum_calculator #(.RECT1_X(rectangle1_xs[211]), .RECT1_Y(rectangle1_ys[211]), .RECT1_WIDTH(rectangle1_widths[211]), .RECT1_HEIGHT(rectangle1_heights[211]), .RECT1_WEIGHT(rectangle1_weights[211]), .RECT2_X(rectangle2_xs[211]), .RECT2_Y(rectangle2_ys[211]), .RECT2_WIDTH(rectangle2_widths[211]), .RECT2_HEIGHT(rectangle2_heights[211]), .RECT2_WEIGHT(rectangle2_weights[211]), .RECT3_X(rectangle3_xs[211]), .RECT3_Y(rectangle3_ys[211]), .RECT3_WIDTH(rectangle3_widths[211]), .RECT3_HEIGHT(rectangle3_heights[211]), .RECT3_WEIGHT(rectangle3_weights[211]), .FEAT_THRES(feature_thresholds[211]), .FEAT_ABOVE(feature_aboves[211]), .FEAT_BELOW(feature_belows[211])) ac211(.scan_win(scan_win211), .scan_win_std_dev(scan_win_std_dev[211]), .feature_accum(feature_accums[211]));
  accum_calculator #(.RECT1_X(rectangle1_xs[212]), .RECT1_Y(rectangle1_ys[212]), .RECT1_WIDTH(rectangle1_widths[212]), .RECT1_HEIGHT(rectangle1_heights[212]), .RECT1_WEIGHT(rectangle1_weights[212]), .RECT2_X(rectangle2_xs[212]), .RECT2_Y(rectangle2_ys[212]), .RECT2_WIDTH(rectangle2_widths[212]), .RECT2_HEIGHT(rectangle2_heights[212]), .RECT2_WEIGHT(rectangle2_weights[212]), .RECT3_X(rectangle3_xs[212]), .RECT3_Y(rectangle3_ys[212]), .RECT3_WIDTH(rectangle3_widths[212]), .RECT3_HEIGHT(rectangle3_heights[212]), .RECT3_WEIGHT(rectangle3_weights[212]), .FEAT_THRES(feature_thresholds[212]), .FEAT_ABOVE(feature_aboves[212]), .FEAT_BELOW(feature_belows[212])) ac212(.scan_win(scan_win212), .scan_win_std_dev(scan_win_std_dev[212]), .feature_accum(feature_accums[212]));
  accum_calculator #(.RECT1_X(rectangle1_xs[213]), .RECT1_Y(rectangle1_ys[213]), .RECT1_WIDTH(rectangle1_widths[213]), .RECT1_HEIGHT(rectangle1_heights[213]), .RECT1_WEIGHT(rectangle1_weights[213]), .RECT2_X(rectangle2_xs[213]), .RECT2_Y(rectangle2_ys[213]), .RECT2_WIDTH(rectangle2_widths[213]), .RECT2_HEIGHT(rectangle2_heights[213]), .RECT2_WEIGHT(rectangle2_weights[213]), .RECT3_X(rectangle3_xs[213]), .RECT3_Y(rectangle3_ys[213]), .RECT3_WIDTH(rectangle3_widths[213]), .RECT3_HEIGHT(rectangle3_heights[213]), .RECT3_WEIGHT(rectangle3_weights[213]), .FEAT_THRES(feature_thresholds[213]), .FEAT_ABOVE(feature_aboves[213]), .FEAT_BELOW(feature_belows[213])) ac213(.scan_win(scan_win213), .scan_win_std_dev(scan_win_std_dev[213]), .feature_accum(feature_accums[213]));
  accum_calculator #(.RECT1_X(rectangle1_xs[214]), .RECT1_Y(rectangle1_ys[214]), .RECT1_WIDTH(rectangle1_widths[214]), .RECT1_HEIGHT(rectangle1_heights[214]), .RECT1_WEIGHT(rectangle1_weights[214]), .RECT2_X(rectangle2_xs[214]), .RECT2_Y(rectangle2_ys[214]), .RECT2_WIDTH(rectangle2_widths[214]), .RECT2_HEIGHT(rectangle2_heights[214]), .RECT2_WEIGHT(rectangle2_weights[214]), .RECT3_X(rectangle3_xs[214]), .RECT3_Y(rectangle3_ys[214]), .RECT3_WIDTH(rectangle3_widths[214]), .RECT3_HEIGHT(rectangle3_heights[214]), .RECT3_WEIGHT(rectangle3_weights[214]), .FEAT_THRES(feature_thresholds[214]), .FEAT_ABOVE(feature_aboves[214]), .FEAT_BELOW(feature_belows[214])) ac214(.scan_win(scan_win214), .scan_win_std_dev(scan_win_std_dev[214]), .feature_accum(feature_accums[214]));
  accum_calculator #(.RECT1_X(rectangle1_xs[215]), .RECT1_Y(rectangle1_ys[215]), .RECT1_WIDTH(rectangle1_widths[215]), .RECT1_HEIGHT(rectangle1_heights[215]), .RECT1_WEIGHT(rectangle1_weights[215]), .RECT2_X(rectangle2_xs[215]), .RECT2_Y(rectangle2_ys[215]), .RECT2_WIDTH(rectangle2_widths[215]), .RECT2_HEIGHT(rectangle2_heights[215]), .RECT2_WEIGHT(rectangle2_weights[215]), .RECT3_X(rectangle3_xs[215]), .RECT3_Y(rectangle3_ys[215]), .RECT3_WIDTH(rectangle3_widths[215]), .RECT3_HEIGHT(rectangle3_heights[215]), .RECT3_WEIGHT(rectangle3_weights[215]), .FEAT_THRES(feature_thresholds[215]), .FEAT_ABOVE(feature_aboves[215]), .FEAT_BELOW(feature_belows[215])) ac215(.scan_win(scan_win215), .scan_win_std_dev(scan_win_std_dev[215]), .feature_accum(feature_accums[215]));
  accum_calculator #(.RECT1_X(rectangle1_xs[216]), .RECT1_Y(rectangle1_ys[216]), .RECT1_WIDTH(rectangle1_widths[216]), .RECT1_HEIGHT(rectangle1_heights[216]), .RECT1_WEIGHT(rectangle1_weights[216]), .RECT2_X(rectangle2_xs[216]), .RECT2_Y(rectangle2_ys[216]), .RECT2_WIDTH(rectangle2_widths[216]), .RECT2_HEIGHT(rectangle2_heights[216]), .RECT2_WEIGHT(rectangle2_weights[216]), .RECT3_X(rectangle3_xs[216]), .RECT3_Y(rectangle3_ys[216]), .RECT3_WIDTH(rectangle3_widths[216]), .RECT3_HEIGHT(rectangle3_heights[216]), .RECT3_WEIGHT(rectangle3_weights[216]), .FEAT_THRES(feature_thresholds[216]), .FEAT_ABOVE(feature_aboves[216]), .FEAT_BELOW(feature_belows[216])) ac216(.scan_win(scan_win216), .scan_win_std_dev(scan_win_std_dev[216]), .feature_accum(feature_accums[216]));
  accum_calculator #(.RECT1_X(rectangle1_xs[217]), .RECT1_Y(rectangle1_ys[217]), .RECT1_WIDTH(rectangle1_widths[217]), .RECT1_HEIGHT(rectangle1_heights[217]), .RECT1_WEIGHT(rectangle1_weights[217]), .RECT2_X(rectangle2_xs[217]), .RECT2_Y(rectangle2_ys[217]), .RECT2_WIDTH(rectangle2_widths[217]), .RECT2_HEIGHT(rectangle2_heights[217]), .RECT2_WEIGHT(rectangle2_weights[217]), .RECT3_X(rectangle3_xs[217]), .RECT3_Y(rectangle3_ys[217]), .RECT3_WIDTH(rectangle3_widths[217]), .RECT3_HEIGHT(rectangle3_heights[217]), .RECT3_WEIGHT(rectangle3_weights[217]), .FEAT_THRES(feature_thresholds[217]), .FEAT_ABOVE(feature_aboves[217]), .FEAT_BELOW(feature_belows[217])) ac217(.scan_win(scan_win217), .scan_win_std_dev(scan_win_std_dev[217]), .feature_accum(feature_accums[217]));
  accum_calculator #(.RECT1_X(rectangle1_xs[218]), .RECT1_Y(rectangle1_ys[218]), .RECT1_WIDTH(rectangle1_widths[218]), .RECT1_HEIGHT(rectangle1_heights[218]), .RECT1_WEIGHT(rectangle1_weights[218]), .RECT2_X(rectangle2_xs[218]), .RECT2_Y(rectangle2_ys[218]), .RECT2_WIDTH(rectangle2_widths[218]), .RECT2_HEIGHT(rectangle2_heights[218]), .RECT2_WEIGHT(rectangle2_weights[218]), .RECT3_X(rectangle3_xs[218]), .RECT3_Y(rectangle3_ys[218]), .RECT3_WIDTH(rectangle3_widths[218]), .RECT3_HEIGHT(rectangle3_heights[218]), .RECT3_WEIGHT(rectangle3_weights[218]), .FEAT_THRES(feature_thresholds[218]), .FEAT_ABOVE(feature_aboves[218]), .FEAT_BELOW(feature_belows[218])) ac218(.scan_win(scan_win218), .scan_win_std_dev(scan_win_std_dev[218]), .feature_accum(feature_accums[218]));
  accum_calculator #(.RECT1_X(rectangle1_xs[219]), .RECT1_Y(rectangle1_ys[219]), .RECT1_WIDTH(rectangle1_widths[219]), .RECT1_HEIGHT(rectangle1_heights[219]), .RECT1_WEIGHT(rectangle1_weights[219]), .RECT2_X(rectangle2_xs[219]), .RECT2_Y(rectangle2_ys[219]), .RECT2_WIDTH(rectangle2_widths[219]), .RECT2_HEIGHT(rectangle2_heights[219]), .RECT2_WEIGHT(rectangle2_weights[219]), .RECT3_X(rectangle3_xs[219]), .RECT3_Y(rectangle3_ys[219]), .RECT3_WIDTH(rectangle3_widths[219]), .RECT3_HEIGHT(rectangle3_heights[219]), .RECT3_WEIGHT(rectangle3_weights[219]), .FEAT_THRES(feature_thresholds[219]), .FEAT_ABOVE(feature_aboves[219]), .FEAT_BELOW(feature_belows[219])) ac219(.scan_win(scan_win219), .scan_win_std_dev(scan_win_std_dev[219]), .feature_accum(feature_accums[219]));
  accum_calculator #(.RECT1_X(rectangle1_xs[220]), .RECT1_Y(rectangle1_ys[220]), .RECT1_WIDTH(rectangle1_widths[220]), .RECT1_HEIGHT(rectangle1_heights[220]), .RECT1_WEIGHT(rectangle1_weights[220]), .RECT2_X(rectangle2_xs[220]), .RECT2_Y(rectangle2_ys[220]), .RECT2_WIDTH(rectangle2_widths[220]), .RECT2_HEIGHT(rectangle2_heights[220]), .RECT2_WEIGHT(rectangle2_weights[220]), .RECT3_X(rectangle3_xs[220]), .RECT3_Y(rectangle3_ys[220]), .RECT3_WIDTH(rectangle3_widths[220]), .RECT3_HEIGHT(rectangle3_heights[220]), .RECT3_WEIGHT(rectangle3_weights[220]), .FEAT_THRES(feature_thresholds[220]), .FEAT_ABOVE(feature_aboves[220]), .FEAT_BELOW(feature_belows[220])) ac220(.scan_win(scan_win220), .scan_win_std_dev(scan_win_std_dev[220]), .feature_accum(feature_accums[220]));
  accum_calculator #(.RECT1_X(rectangle1_xs[221]), .RECT1_Y(rectangle1_ys[221]), .RECT1_WIDTH(rectangle1_widths[221]), .RECT1_HEIGHT(rectangle1_heights[221]), .RECT1_WEIGHT(rectangle1_weights[221]), .RECT2_X(rectangle2_xs[221]), .RECT2_Y(rectangle2_ys[221]), .RECT2_WIDTH(rectangle2_widths[221]), .RECT2_HEIGHT(rectangle2_heights[221]), .RECT2_WEIGHT(rectangle2_weights[221]), .RECT3_X(rectangle3_xs[221]), .RECT3_Y(rectangle3_ys[221]), .RECT3_WIDTH(rectangle3_widths[221]), .RECT3_HEIGHT(rectangle3_heights[221]), .RECT3_WEIGHT(rectangle3_weights[221]), .FEAT_THRES(feature_thresholds[221]), .FEAT_ABOVE(feature_aboves[221]), .FEAT_BELOW(feature_belows[221])) ac221(.scan_win(scan_win221), .scan_win_std_dev(scan_win_std_dev[221]), .feature_accum(feature_accums[221]));
  accum_calculator #(.RECT1_X(rectangle1_xs[222]), .RECT1_Y(rectangle1_ys[222]), .RECT1_WIDTH(rectangle1_widths[222]), .RECT1_HEIGHT(rectangle1_heights[222]), .RECT1_WEIGHT(rectangle1_weights[222]), .RECT2_X(rectangle2_xs[222]), .RECT2_Y(rectangle2_ys[222]), .RECT2_WIDTH(rectangle2_widths[222]), .RECT2_HEIGHT(rectangle2_heights[222]), .RECT2_WEIGHT(rectangle2_weights[222]), .RECT3_X(rectangle3_xs[222]), .RECT3_Y(rectangle3_ys[222]), .RECT3_WIDTH(rectangle3_widths[222]), .RECT3_HEIGHT(rectangle3_heights[222]), .RECT3_WEIGHT(rectangle3_weights[222]), .FEAT_THRES(feature_thresholds[222]), .FEAT_ABOVE(feature_aboves[222]), .FEAT_BELOW(feature_belows[222])) ac222(.scan_win(scan_win222), .scan_win_std_dev(scan_win_std_dev[222]), .feature_accum(feature_accums[222]));
  accum_calculator #(.RECT1_X(rectangle1_xs[223]), .RECT1_Y(rectangle1_ys[223]), .RECT1_WIDTH(rectangle1_widths[223]), .RECT1_HEIGHT(rectangle1_heights[223]), .RECT1_WEIGHT(rectangle1_weights[223]), .RECT2_X(rectangle2_xs[223]), .RECT2_Y(rectangle2_ys[223]), .RECT2_WIDTH(rectangle2_widths[223]), .RECT2_HEIGHT(rectangle2_heights[223]), .RECT2_WEIGHT(rectangle2_weights[223]), .RECT3_X(rectangle3_xs[223]), .RECT3_Y(rectangle3_ys[223]), .RECT3_WIDTH(rectangle3_widths[223]), .RECT3_HEIGHT(rectangle3_heights[223]), .RECT3_WEIGHT(rectangle3_weights[223]), .FEAT_THRES(feature_thresholds[223]), .FEAT_ABOVE(feature_aboves[223]), .FEAT_BELOW(feature_belows[223])) ac223(.scan_win(scan_win223), .scan_win_std_dev(scan_win_std_dev[223]), .feature_accum(feature_accums[223]));
  accum_calculator #(.RECT1_X(rectangle1_xs[224]), .RECT1_Y(rectangle1_ys[224]), .RECT1_WIDTH(rectangle1_widths[224]), .RECT1_HEIGHT(rectangle1_heights[224]), .RECT1_WEIGHT(rectangle1_weights[224]), .RECT2_X(rectangle2_xs[224]), .RECT2_Y(rectangle2_ys[224]), .RECT2_WIDTH(rectangle2_widths[224]), .RECT2_HEIGHT(rectangle2_heights[224]), .RECT2_WEIGHT(rectangle2_weights[224]), .RECT3_X(rectangle3_xs[224]), .RECT3_Y(rectangle3_ys[224]), .RECT3_WIDTH(rectangle3_widths[224]), .RECT3_HEIGHT(rectangle3_heights[224]), .RECT3_WEIGHT(rectangle3_weights[224]), .FEAT_THRES(feature_thresholds[224]), .FEAT_ABOVE(feature_aboves[224]), .FEAT_BELOW(feature_belows[224])) ac224(.scan_win(scan_win224), .scan_win_std_dev(scan_win_std_dev[224]), .feature_accum(feature_accums[224]));
  accum_calculator #(.RECT1_X(rectangle1_xs[225]), .RECT1_Y(rectangle1_ys[225]), .RECT1_WIDTH(rectangle1_widths[225]), .RECT1_HEIGHT(rectangle1_heights[225]), .RECT1_WEIGHT(rectangle1_weights[225]), .RECT2_X(rectangle2_xs[225]), .RECT2_Y(rectangle2_ys[225]), .RECT2_WIDTH(rectangle2_widths[225]), .RECT2_HEIGHT(rectangle2_heights[225]), .RECT2_WEIGHT(rectangle2_weights[225]), .RECT3_X(rectangle3_xs[225]), .RECT3_Y(rectangle3_ys[225]), .RECT3_WIDTH(rectangle3_widths[225]), .RECT3_HEIGHT(rectangle3_heights[225]), .RECT3_WEIGHT(rectangle3_weights[225]), .FEAT_THRES(feature_thresholds[225]), .FEAT_ABOVE(feature_aboves[225]), .FEAT_BELOW(feature_belows[225])) ac225(.scan_win(scan_win225), .scan_win_std_dev(scan_win_std_dev[225]), .feature_accum(feature_accums[225]));
  accum_calculator #(.RECT1_X(rectangle1_xs[226]), .RECT1_Y(rectangle1_ys[226]), .RECT1_WIDTH(rectangle1_widths[226]), .RECT1_HEIGHT(rectangle1_heights[226]), .RECT1_WEIGHT(rectangle1_weights[226]), .RECT2_X(rectangle2_xs[226]), .RECT2_Y(rectangle2_ys[226]), .RECT2_WIDTH(rectangle2_widths[226]), .RECT2_HEIGHT(rectangle2_heights[226]), .RECT2_WEIGHT(rectangle2_weights[226]), .RECT3_X(rectangle3_xs[226]), .RECT3_Y(rectangle3_ys[226]), .RECT3_WIDTH(rectangle3_widths[226]), .RECT3_HEIGHT(rectangle3_heights[226]), .RECT3_WEIGHT(rectangle3_weights[226]), .FEAT_THRES(feature_thresholds[226]), .FEAT_ABOVE(feature_aboves[226]), .FEAT_BELOW(feature_belows[226])) ac226(.scan_win(scan_win226), .scan_win_std_dev(scan_win_std_dev[226]), .feature_accum(feature_accums[226]));
  accum_calculator #(.RECT1_X(rectangle1_xs[227]), .RECT1_Y(rectangle1_ys[227]), .RECT1_WIDTH(rectangle1_widths[227]), .RECT1_HEIGHT(rectangle1_heights[227]), .RECT1_WEIGHT(rectangle1_weights[227]), .RECT2_X(rectangle2_xs[227]), .RECT2_Y(rectangle2_ys[227]), .RECT2_WIDTH(rectangle2_widths[227]), .RECT2_HEIGHT(rectangle2_heights[227]), .RECT2_WEIGHT(rectangle2_weights[227]), .RECT3_X(rectangle3_xs[227]), .RECT3_Y(rectangle3_ys[227]), .RECT3_WIDTH(rectangle3_widths[227]), .RECT3_HEIGHT(rectangle3_heights[227]), .RECT3_WEIGHT(rectangle3_weights[227]), .FEAT_THRES(feature_thresholds[227]), .FEAT_ABOVE(feature_aboves[227]), .FEAT_BELOW(feature_belows[227])) ac227(.scan_win(scan_win227), .scan_win_std_dev(scan_win_std_dev[227]), .feature_accum(feature_accums[227]));
  accum_calculator #(.RECT1_X(rectangle1_xs[228]), .RECT1_Y(rectangle1_ys[228]), .RECT1_WIDTH(rectangle1_widths[228]), .RECT1_HEIGHT(rectangle1_heights[228]), .RECT1_WEIGHT(rectangle1_weights[228]), .RECT2_X(rectangle2_xs[228]), .RECT2_Y(rectangle2_ys[228]), .RECT2_WIDTH(rectangle2_widths[228]), .RECT2_HEIGHT(rectangle2_heights[228]), .RECT2_WEIGHT(rectangle2_weights[228]), .RECT3_X(rectangle3_xs[228]), .RECT3_Y(rectangle3_ys[228]), .RECT3_WIDTH(rectangle3_widths[228]), .RECT3_HEIGHT(rectangle3_heights[228]), .RECT3_WEIGHT(rectangle3_weights[228]), .FEAT_THRES(feature_thresholds[228]), .FEAT_ABOVE(feature_aboves[228]), .FEAT_BELOW(feature_belows[228])) ac228(.scan_win(scan_win228), .scan_win_std_dev(scan_win_std_dev[228]), .feature_accum(feature_accums[228]));
  accum_calculator #(.RECT1_X(rectangle1_xs[229]), .RECT1_Y(rectangle1_ys[229]), .RECT1_WIDTH(rectangle1_widths[229]), .RECT1_HEIGHT(rectangle1_heights[229]), .RECT1_WEIGHT(rectangle1_weights[229]), .RECT2_X(rectangle2_xs[229]), .RECT2_Y(rectangle2_ys[229]), .RECT2_WIDTH(rectangle2_widths[229]), .RECT2_HEIGHT(rectangle2_heights[229]), .RECT2_WEIGHT(rectangle2_weights[229]), .RECT3_X(rectangle3_xs[229]), .RECT3_Y(rectangle3_ys[229]), .RECT3_WIDTH(rectangle3_widths[229]), .RECT3_HEIGHT(rectangle3_heights[229]), .RECT3_WEIGHT(rectangle3_weights[229]), .FEAT_THRES(feature_thresholds[229]), .FEAT_ABOVE(feature_aboves[229]), .FEAT_BELOW(feature_belows[229])) ac229(.scan_win(scan_win229), .scan_win_std_dev(scan_win_std_dev[229]), .feature_accum(feature_accums[229]));
  accum_calculator #(.RECT1_X(rectangle1_xs[230]), .RECT1_Y(rectangle1_ys[230]), .RECT1_WIDTH(rectangle1_widths[230]), .RECT1_HEIGHT(rectangle1_heights[230]), .RECT1_WEIGHT(rectangle1_weights[230]), .RECT2_X(rectangle2_xs[230]), .RECT2_Y(rectangle2_ys[230]), .RECT2_WIDTH(rectangle2_widths[230]), .RECT2_HEIGHT(rectangle2_heights[230]), .RECT2_WEIGHT(rectangle2_weights[230]), .RECT3_X(rectangle3_xs[230]), .RECT3_Y(rectangle3_ys[230]), .RECT3_WIDTH(rectangle3_widths[230]), .RECT3_HEIGHT(rectangle3_heights[230]), .RECT3_WEIGHT(rectangle3_weights[230]), .FEAT_THRES(feature_thresholds[230]), .FEAT_ABOVE(feature_aboves[230]), .FEAT_BELOW(feature_belows[230])) ac230(.scan_win(scan_win230), .scan_win_std_dev(scan_win_std_dev[230]), .feature_accum(feature_accums[230]));
  accum_calculator #(.RECT1_X(rectangle1_xs[231]), .RECT1_Y(rectangle1_ys[231]), .RECT1_WIDTH(rectangle1_widths[231]), .RECT1_HEIGHT(rectangle1_heights[231]), .RECT1_WEIGHT(rectangle1_weights[231]), .RECT2_X(rectangle2_xs[231]), .RECT2_Y(rectangle2_ys[231]), .RECT2_WIDTH(rectangle2_widths[231]), .RECT2_HEIGHT(rectangle2_heights[231]), .RECT2_WEIGHT(rectangle2_weights[231]), .RECT3_X(rectangle3_xs[231]), .RECT3_Y(rectangle3_ys[231]), .RECT3_WIDTH(rectangle3_widths[231]), .RECT3_HEIGHT(rectangle3_heights[231]), .RECT3_WEIGHT(rectangle3_weights[231]), .FEAT_THRES(feature_thresholds[231]), .FEAT_ABOVE(feature_aboves[231]), .FEAT_BELOW(feature_belows[231])) ac231(.scan_win(scan_win231), .scan_win_std_dev(scan_win_std_dev[231]), .feature_accum(feature_accums[231]));
  accum_calculator #(.RECT1_X(rectangle1_xs[232]), .RECT1_Y(rectangle1_ys[232]), .RECT1_WIDTH(rectangle1_widths[232]), .RECT1_HEIGHT(rectangle1_heights[232]), .RECT1_WEIGHT(rectangle1_weights[232]), .RECT2_X(rectangle2_xs[232]), .RECT2_Y(rectangle2_ys[232]), .RECT2_WIDTH(rectangle2_widths[232]), .RECT2_HEIGHT(rectangle2_heights[232]), .RECT2_WEIGHT(rectangle2_weights[232]), .RECT3_X(rectangle3_xs[232]), .RECT3_Y(rectangle3_ys[232]), .RECT3_WIDTH(rectangle3_widths[232]), .RECT3_HEIGHT(rectangle3_heights[232]), .RECT3_WEIGHT(rectangle3_weights[232]), .FEAT_THRES(feature_thresholds[232]), .FEAT_ABOVE(feature_aboves[232]), .FEAT_BELOW(feature_belows[232])) ac232(.scan_win(scan_win232), .scan_win_std_dev(scan_win_std_dev[232]), .feature_accum(feature_accums[232]));
  accum_calculator #(.RECT1_X(rectangle1_xs[233]), .RECT1_Y(rectangle1_ys[233]), .RECT1_WIDTH(rectangle1_widths[233]), .RECT1_HEIGHT(rectangle1_heights[233]), .RECT1_WEIGHT(rectangle1_weights[233]), .RECT2_X(rectangle2_xs[233]), .RECT2_Y(rectangle2_ys[233]), .RECT2_WIDTH(rectangle2_widths[233]), .RECT2_HEIGHT(rectangle2_heights[233]), .RECT2_WEIGHT(rectangle2_weights[233]), .RECT3_X(rectangle3_xs[233]), .RECT3_Y(rectangle3_ys[233]), .RECT3_WIDTH(rectangle3_widths[233]), .RECT3_HEIGHT(rectangle3_heights[233]), .RECT3_WEIGHT(rectangle3_weights[233]), .FEAT_THRES(feature_thresholds[233]), .FEAT_ABOVE(feature_aboves[233]), .FEAT_BELOW(feature_belows[233])) ac233(.scan_win(scan_win233), .scan_win_std_dev(scan_win_std_dev[233]), .feature_accum(feature_accums[233]));
  accum_calculator #(.RECT1_X(rectangle1_xs[234]), .RECT1_Y(rectangle1_ys[234]), .RECT1_WIDTH(rectangle1_widths[234]), .RECT1_HEIGHT(rectangle1_heights[234]), .RECT1_WEIGHT(rectangle1_weights[234]), .RECT2_X(rectangle2_xs[234]), .RECT2_Y(rectangle2_ys[234]), .RECT2_WIDTH(rectangle2_widths[234]), .RECT2_HEIGHT(rectangle2_heights[234]), .RECT2_WEIGHT(rectangle2_weights[234]), .RECT3_X(rectangle3_xs[234]), .RECT3_Y(rectangle3_ys[234]), .RECT3_WIDTH(rectangle3_widths[234]), .RECT3_HEIGHT(rectangle3_heights[234]), .RECT3_WEIGHT(rectangle3_weights[234]), .FEAT_THRES(feature_thresholds[234]), .FEAT_ABOVE(feature_aboves[234]), .FEAT_BELOW(feature_belows[234])) ac234(.scan_win(scan_win234), .scan_win_std_dev(scan_win_std_dev[234]), .feature_accum(feature_accums[234]));
  accum_calculator #(.RECT1_X(rectangle1_xs[235]), .RECT1_Y(rectangle1_ys[235]), .RECT1_WIDTH(rectangle1_widths[235]), .RECT1_HEIGHT(rectangle1_heights[235]), .RECT1_WEIGHT(rectangle1_weights[235]), .RECT2_X(rectangle2_xs[235]), .RECT2_Y(rectangle2_ys[235]), .RECT2_WIDTH(rectangle2_widths[235]), .RECT2_HEIGHT(rectangle2_heights[235]), .RECT2_WEIGHT(rectangle2_weights[235]), .RECT3_X(rectangle3_xs[235]), .RECT3_Y(rectangle3_ys[235]), .RECT3_WIDTH(rectangle3_widths[235]), .RECT3_HEIGHT(rectangle3_heights[235]), .RECT3_WEIGHT(rectangle3_weights[235]), .FEAT_THRES(feature_thresholds[235]), .FEAT_ABOVE(feature_aboves[235]), .FEAT_BELOW(feature_belows[235])) ac235(.scan_win(scan_win235), .scan_win_std_dev(scan_win_std_dev[235]), .feature_accum(feature_accums[235]));
  accum_calculator #(.RECT1_X(rectangle1_xs[236]), .RECT1_Y(rectangle1_ys[236]), .RECT1_WIDTH(rectangle1_widths[236]), .RECT1_HEIGHT(rectangle1_heights[236]), .RECT1_WEIGHT(rectangle1_weights[236]), .RECT2_X(rectangle2_xs[236]), .RECT2_Y(rectangle2_ys[236]), .RECT2_WIDTH(rectangle2_widths[236]), .RECT2_HEIGHT(rectangle2_heights[236]), .RECT2_WEIGHT(rectangle2_weights[236]), .RECT3_X(rectangle3_xs[236]), .RECT3_Y(rectangle3_ys[236]), .RECT3_WIDTH(rectangle3_widths[236]), .RECT3_HEIGHT(rectangle3_heights[236]), .RECT3_WEIGHT(rectangle3_weights[236]), .FEAT_THRES(feature_thresholds[236]), .FEAT_ABOVE(feature_aboves[236]), .FEAT_BELOW(feature_belows[236])) ac236(.scan_win(scan_win236), .scan_win_std_dev(scan_win_std_dev[236]), .feature_accum(feature_accums[236]));
  accum_calculator #(.RECT1_X(rectangle1_xs[237]), .RECT1_Y(rectangle1_ys[237]), .RECT1_WIDTH(rectangle1_widths[237]), .RECT1_HEIGHT(rectangle1_heights[237]), .RECT1_WEIGHT(rectangle1_weights[237]), .RECT2_X(rectangle2_xs[237]), .RECT2_Y(rectangle2_ys[237]), .RECT2_WIDTH(rectangle2_widths[237]), .RECT2_HEIGHT(rectangle2_heights[237]), .RECT2_WEIGHT(rectangle2_weights[237]), .RECT3_X(rectangle3_xs[237]), .RECT3_Y(rectangle3_ys[237]), .RECT3_WIDTH(rectangle3_widths[237]), .RECT3_HEIGHT(rectangle3_heights[237]), .RECT3_WEIGHT(rectangle3_weights[237]), .FEAT_THRES(feature_thresholds[237]), .FEAT_ABOVE(feature_aboves[237]), .FEAT_BELOW(feature_belows[237])) ac237(.scan_win(scan_win237), .scan_win_std_dev(scan_win_std_dev[237]), .feature_accum(feature_accums[237]));
  accum_calculator #(.RECT1_X(rectangle1_xs[238]), .RECT1_Y(rectangle1_ys[238]), .RECT1_WIDTH(rectangle1_widths[238]), .RECT1_HEIGHT(rectangle1_heights[238]), .RECT1_WEIGHT(rectangle1_weights[238]), .RECT2_X(rectangle2_xs[238]), .RECT2_Y(rectangle2_ys[238]), .RECT2_WIDTH(rectangle2_widths[238]), .RECT2_HEIGHT(rectangle2_heights[238]), .RECT2_WEIGHT(rectangle2_weights[238]), .RECT3_X(rectangle3_xs[238]), .RECT3_Y(rectangle3_ys[238]), .RECT3_WIDTH(rectangle3_widths[238]), .RECT3_HEIGHT(rectangle3_heights[238]), .RECT3_WEIGHT(rectangle3_weights[238]), .FEAT_THRES(feature_thresholds[238]), .FEAT_ABOVE(feature_aboves[238]), .FEAT_BELOW(feature_belows[238])) ac238(.scan_win(scan_win238), .scan_win_std_dev(scan_win_std_dev[238]), .feature_accum(feature_accums[238]));
  accum_calculator #(.RECT1_X(rectangle1_xs[239]), .RECT1_Y(rectangle1_ys[239]), .RECT1_WIDTH(rectangle1_widths[239]), .RECT1_HEIGHT(rectangle1_heights[239]), .RECT1_WEIGHT(rectangle1_weights[239]), .RECT2_X(rectangle2_xs[239]), .RECT2_Y(rectangle2_ys[239]), .RECT2_WIDTH(rectangle2_widths[239]), .RECT2_HEIGHT(rectangle2_heights[239]), .RECT2_WEIGHT(rectangle2_weights[239]), .RECT3_X(rectangle3_xs[239]), .RECT3_Y(rectangle3_ys[239]), .RECT3_WIDTH(rectangle3_widths[239]), .RECT3_HEIGHT(rectangle3_heights[239]), .RECT3_WEIGHT(rectangle3_weights[239]), .FEAT_THRES(feature_thresholds[239]), .FEAT_ABOVE(feature_aboves[239]), .FEAT_BELOW(feature_belows[239])) ac239(.scan_win(scan_win239), .scan_win_std_dev(scan_win_std_dev[239]), .feature_accum(feature_accums[239]));
  accum_calculator #(.RECT1_X(rectangle1_xs[240]), .RECT1_Y(rectangle1_ys[240]), .RECT1_WIDTH(rectangle1_widths[240]), .RECT1_HEIGHT(rectangle1_heights[240]), .RECT1_WEIGHT(rectangle1_weights[240]), .RECT2_X(rectangle2_xs[240]), .RECT2_Y(rectangle2_ys[240]), .RECT2_WIDTH(rectangle2_widths[240]), .RECT2_HEIGHT(rectangle2_heights[240]), .RECT2_WEIGHT(rectangle2_weights[240]), .RECT3_X(rectangle3_xs[240]), .RECT3_Y(rectangle3_ys[240]), .RECT3_WIDTH(rectangle3_widths[240]), .RECT3_HEIGHT(rectangle3_heights[240]), .RECT3_WEIGHT(rectangle3_weights[240]), .FEAT_THRES(feature_thresholds[240]), .FEAT_ABOVE(feature_aboves[240]), .FEAT_BELOW(feature_belows[240])) ac240(.scan_win(scan_win240), .scan_win_std_dev(scan_win_std_dev[240]), .feature_accum(feature_accums[240]));
  accum_calculator #(.RECT1_X(rectangle1_xs[241]), .RECT1_Y(rectangle1_ys[241]), .RECT1_WIDTH(rectangle1_widths[241]), .RECT1_HEIGHT(rectangle1_heights[241]), .RECT1_WEIGHT(rectangle1_weights[241]), .RECT2_X(rectangle2_xs[241]), .RECT2_Y(rectangle2_ys[241]), .RECT2_WIDTH(rectangle2_widths[241]), .RECT2_HEIGHT(rectangle2_heights[241]), .RECT2_WEIGHT(rectangle2_weights[241]), .RECT3_X(rectangle3_xs[241]), .RECT3_Y(rectangle3_ys[241]), .RECT3_WIDTH(rectangle3_widths[241]), .RECT3_HEIGHT(rectangle3_heights[241]), .RECT3_WEIGHT(rectangle3_weights[241]), .FEAT_THRES(feature_thresholds[241]), .FEAT_ABOVE(feature_aboves[241]), .FEAT_BELOW(feature_belows[241])) ac241(.scan_win(scan_win241), .scan_win_std_dev(scan_win_std_dev[241]), .feature_accum(feature_accums[241]));
  accum_calculator #(.RECT1_X(rectangle1_xs[242]), .RECT1_Y(rectangle1_ys[242]), .RECT1_WIDTH(rectangle1_widths[242]), .RECT1_HEIGHT(rectangle1_heights[242]), .RECT1_WEIGHT(rectangle1_weights[242]), .RECT2_X(rectangle2_xs[242]), .RECT2_Y(rectangle2_ys[242]), .RECT2_WIDTH(rectangle2_widths[242]), .RECT2_HEIGHT(rectangle2_heights[242]), .RECT2_WEIGHT(rectangle2_weights[242]), .RECT3_X(rectangle3_xs[242]), .RECT3_Y(rectangle3_ys[242]), .RECT3_WIDTH(rectangle3_widths[242]), .RECT3_HEIGHT(rectangle3_heights[242]), .RECT3_WEIGHT(rectangle3_weights[242]), .FEAT_THRES(feature_thresholds[242]), .FEAT_ABOVE(feature_aboves[242]), .FEAT_BELOW(feature_belows[242])) ac242(.scan_win(scan_win242), .scan_win_std_dev(scan_win_std_dev[242]), .feature_accum(feature_accums[242]));
  accum_calculator #(.RECT1_X(rectangle1_xs[243]), .RECT1_Y(rectangle1_ys[243]), .RECT1_WIDTH(rectangle1_widths[243]), .RECT1_HEIGHT(rectangle1_heights[243]), .RECT1_WEIGHT(rectangle1_weights[243]), .RECT2_X(rectangle2_xs[243]), .RECT2_Y(rectangle2_ys[243]), .RECT2_WIDTH(rectangle2_widths[243]), .RECT2_HEIGHT(rectangle2_heights[243]), .RECT2_WEIGHT(rectangle2_weights[243]), .RECT3_X(rectangle3_xs[243]), .RECT3_Y(rectangle3_ys[243]), .RECT3_WIDTH(rectangle3_widths[243]), .RECT3_HEIGHT(rectangle3_heights[243]), .RECT3_WEIGHT(rectangle3_weights[243]), .FEAT_THRES(feature_thresholds[243]), .FEAT_ABOVE(feature_aboves[243]), .FEAT_BELOW(feature_belows[243])) ac243(.scan_win(scan_win243), .scan_win_std_dev(scan_win_std_dev[243]), .feature_accum(feature_accums[243]));
  accum_calculator #(.RECT1_X(rectangle1_xs[244]), .RECT1_Y(rectangle1_ys[244]), .RECT1_WIDTH(rectangle1_widths[244]), .RECT1_HEIGHT(rectangle1_heights[244]), .RECT1_WEIGHT(rectangle1_weights[244]), .RECT2_X(rectangle2_xs[244]), .RECT2_Y(rectangle2_ys[244]), .RECT2_WIDTH(rectangle2_widths[244]), .RECT2_HEIGHT(rectangle2_heights[244]), .RECT2_WEIGHT(rectangle2_weights[244]), .RECT3_X(rectangle3_xs[244]), .RECT3_Y(rectangle3_ys[244]), .RECT3_WIDTH(rectangle3_widths[244]), .RECT3_HEIGHT(rectangle3_heights[244]), .RECT3_WEIGHT(rectangle3_weights[244]), .FEAT_THRES(feature_thresholds[244]), .FEAT_ABOVE(feature_aboves[244]), .FEAT_BELOW(feature_belows[244])) ac244(.scan_win(scan_win244), .scan_win_std_dev(scan_win_std_dev[244]), .feature_accum(feature_accums[244]));
  accum_calculator #(.RECT1_X(rectangle1_xs[245]), .RECT1_Y(rectangle1_ys[245]), .RECT1_WIDTH(rectangle1_widths[245]), .RECT1_HEIGHT(rectangle1_heights[245]), .RECT1_WEIGHT(rectangle1_weights[245]), .RECT2_X(rectangle2_xs[245]), .RECT2_Y(rectangle2_ys[245]), .RECT2_WIDTH(rectangle2_widths[245]), .RECT2_HEIGHT(rectangle2_heights[245]), .RECT2_WEIGHT(rectangle2_weights[245]), .RECT3_X(rectangle3_xs[245]), .RECT3_Y(rectangle3_ys[245]), .RECT3_WIDTH(rectangle3_widths[245]), .RECT3_HEIGHT(rectangle3_heights[245]), .RECT3_WEIGHT(rectangle3_weights[245]), .FEAT_THRES(feature_thresholds[245]), .FEAT_ABOVE(feature_aboves[245]), .FEAT_BELOW(feature_belows[245])) ac245(.scan_win(scan_win245), .scan_win_std_dev(scan_win_std_dev[245]), .feature_accum(feature_accums[245]));
  accum_calculator #(.RECT1_X(rectangle1_xs[246]), .RECT1_Y(rectangle1_ys[246]), .RECT1_WIDTH(rectangle1_widths[246]), .RECT1_HEIGHT(rectangle1_heights[246]), .RECT1_WEIGHT(rectangle1_weights[246]), .RECT2_X(rectangle2_xs[246]), .RECT2_Y(rectangle2_ys[246]), .RECT2_WIDTH(rectangle2_widths[246]), .RECT2_HEIGHT(rectangle2_heights[246]), .RECT2_WEIGHT(rectangle2_weights[246]), .RECT3_X(rectangle3_xs[246]), .RECT3_Y(rectangle3_ys[246]), .RECT3_WIDTH(rectangle3_widths[246]), .RECT3_HEIGHT(rectangle3_heights[246]), .RECT3_WEIGHT(rectangle3_weights[246]), .FEAT_THRES(feature_thresholds[246]), .FEAT_ABOVE(feature_aboves[246]), .FEAT_BELOW(feature_belows[246])) ac246(.scan_win(scan_win246), .scan_win_std_dev(scan_win_std_dev[246]), .feature_accum(feature_accums[246]));
  accum_calculator #(.RECT1_X(rectangle1_xs[247]), .RECT1_Y(rectangle1_ys[247]), .RECT1_WIDTH(rectangle1_widths[247]), .RECT1_HEIGHT(rectangle1_heights[247]), .RECT1_WEIGHT(rectangle1_weights[247]), .RECT2_X(rectangle2_xs[247]), .RECT2_Y(rectangle2_ys[247]), .RECT2_WIDTH(rectangle2_widths[247]), .RECT2_HEIGHT(rectangle2_heights[247]), .RECT2_WEIGHT(rectangle2_weights[247]), .RECT3_X(rectangle3_xs[247]), .RECT3_Y(rectangle3_ys[247]), .RECT3_WIDTH(rectangle3_widths[247]), .RECT3_HEIGHT(rectangle3_heights[247]), .RECT3_WEIGHT(rectangle3_weights[247]), .FEAT_THRES(feature_thresholds[247]), .FEAT_ABOVE(feature_aboves[247]), .FEAT_BELOW(feature_belows[247])) ac247(.scan_win(scan_win247), .scan_win_std_dev(scan_win_std_dev[247]), .feature_accum(feature_accums[247]));
  accum_calculator #(.RECT1_X(rectangle1_xs[248]), .RECT1_Y(rectangle1_ys[248]), .RECT1_WIDTH(rectangle1_widths[248]), .RECT1_HEIGHT(rectangle1_heights[248]), .RECT1_WEIGHT(rectangle1_weights[248]), .RECT2_X(rectangle2_xs[248]), .RECT2_Y(rectangle2_ys[248]), .RECT2_WIDTH(rectangle2_widths[248]), .RECT2_HEIGHT(rectangle2_heights[248]), .RECT2_WEIGHT(rectangle2_weights[248]), .RECT3_X(rectangle3_xs[248]), .RECT3_Y(rectangle3_ys[248]), .RECT3_WIDTH(rectangle3_widths[248]), .RECT3_HEIGHT(rectangle3_heights[248]), .RECT3_WEIGHT(rectangle3_weights[248]), .FEAT_THRES(feature_thresholds[248]), .FEAT_ABOVE(feature_aboves[248]), .FEAT_BELOW(feature_belows[248])) ac248(.scan_win(scan_win248), .scan_win_std_dev(scan_win_std_dev[248]), .feature_accum(feature_accums[248]));
  accum_calculator #(.RECT1_X(rectangle1_xs[249]), .RECT1_Y(rectangle1_ys[249]), .RECT1_WIDTH(rectangle1_widths[249]), .RECT1_HEIGHT(rectangle1_heights[249]), .RECT1_WEIGHT(rectangle1_weights[249]), .RECT2_X(rectangle2_xs[249]), .RECT2_Y(rectangle2_ys[249]), .RECT2_WIDTH(rectangle2_widths[249]), .RECT2_HEIGHT(rectangle2_heights[249]), .RECT2_WEIGHT(rectangle2_weights[249]), .RECT3_X(rectangle3_xs[249]), .RECT3_Y(rectangle3_ys[249]), .RECT3_WIDTH(rectangle3_widths[249]), .RECT3_HEIGHT(rectangle3_heights[249]), .RECT3_WEIGHT(rectangle3_weights[249]), .FEAT_THRES(feature_thresholds[249]), .FEAT_ABOVE(feature_aboves[249]), .FEAT_BELOW(feature_belows[249])) ac249(.scan_win(scan_win249), .scan_win_std_dev(scan_win_std_dev[249]), .feature_accum(feature_accums[249]));
  accum_calculator #(.RECT1_X(rectangle1_xs[250]), .RECT1_Y(rectangle1_ys[250]), .RECT1_WIDTH(rectangle1_widths[250]), .RECT1_HEIGHT(rectangle1_heights[250]), .RECT1_WEIGHT(rectangle1_weights[250]), .RECT2_X(rectangle2_xs[250]), .RECT2_Y(rectangle2_ys[250]), .RECT2_WIDTH(rectangle2_widths[250]), .RECT2_HEIGHT(rectangle2_heights[250]), .RECT2_WEIGHT(rectangle2_weights[250]), .RECT3_X(rectangle3_xs[250]), .RECT3_Y(rectangle3_ys[250]), .RECT3_WIDTH(rectangle3_widths[250]), .RECT3_HEIGHT(rectangle3_heights[250]), .RECT3_WEIGHT(rectangle3_weights[250]), .FEAT_THRES(feature_thresholds[250]), .FEAT_ABOVE(feature_aboves[250]), .FEAT_BELOW(feature_belows[250])) ac250(.scan_win(scan_win250), .scan_win_std_dev(scan_win_std_dev[250]), .feature_accum(feature_accums[250]));
  accum_calculator #(.RECT1_X(rectangle1_xs[251]), .RECT1_Y(rectangle1_ys[251]), .RECT1_WIDTH(rectangle1_widths[251]), .RECT1_HEIGHT(rectangle1_heights[251]), .RECT1_WEIGHT(rectangle1_weights[251]), .RECT2_X(rectangle2_xs[251]), .RECT2_Y(rectangle2_ys[251]), .RECT2_WIDTH(rectangle2_widths[251]), .RECT2_HEIGHT(rectangle2_heights[251]), .RECT2_WEIGHT(rectangle2_weights[251]), .RECT3_X(rectangle3_xs[251]), .RECT3_Y(rectangle3_ys[251]), .RECT3_WIDTH(rectangle3_widths[251]), .RECT3_HEIGHT(rectangle3_heights[251]), .RECT3_WEIGHT(rectangle3_weights[251]), .FEAT_THRES(feature_thresholds[251]), .FEAT_ABOVE(feature_aboves[251]), .FEAT_BELOW(feature_belows[251])) ac251(.scan_win(scan_win251), .scan_win_std_dev(scan_win_std_dev[251]), .feature_accum(feature_accums[251]));
  accum_calculator #(.RECT1_X(rectangle1_xs[252]), .RECT1_Y(rectangle1_ys[252]), .RECT1_WIDTH(rectangle1_widths[252]), .RECT1_HEIGHT(rectangle1_heights[252]), .RECT1_WEIGHT(rectangle1_weights[252]), .RECT2_X(rectangle2_xs[252]), .RECT2_Y(rectangle2_ys[252]), .RECT2_WIDTH(rectangle2_widths[252]), .RECT2_HEIGHT(rectangle2_heights[252]), .RECT2_WEIGHT(rectangle2_weights[252]), .RECT3_X(rectangle3_xs[252]), .RECT3_Y(rectangle3_ys[252]), .RECT3_WIDTH(rectangle3_widths[252]), .RECT3_HEIGHT(rectangle3_heights[252]), .RECT3_WEIGHT(rectangle3_weights[252]), .FEAT_THRES(feature_thresholds[252]), .FEAT_ABOVE(feature_aboves[252]), .FEAT_BELOW(feature_belows[252])) ac252(.scan_win(scan_win252), .scan_win_std_dev(scan_win_std_dev[252]), .feature_accum(feature_accums[252]));
  accum_calculator #(.RECT1_X(rectangle1_xs[253]), .RECT1_Y(rectangle1_ys[253]), .RECT1_WIDTH(rectangle1_widths[253]), .RECT1_HEIGHT(rectangle1_heights[253]), .RECT1_WEIGHT(rectangle1_weights[253]), .RECT2_X(rectangle2_xs[253]), .RECT2_Y(rectangle2_ys[253]), .RECT2_WIDTH(rectangle2_widths[253]), .RECT2_HEIGHT(rectangle2_heights[253]), .RECT2_WEIGHT(rectangle2_weights[253]), .RECT3_X(rectangle3_xs[253]), .RECT3_Y(rectangle3_ys[253]), .RECT3_WIDTH(rectangle3_widths[253]), .RECT3_HEIGHT(rectangle3_heights[253]), .RECT3_WEIGHT(rectangle3_weights[253]), .FEAT_THRES(feature_thresholds[253]), .FEAT_ABOVE(feature_aboves[253]), .FEAT_BELOW(feature_belows[253])) ac253(.scan_win(scan_win253), .scan_win_std_dev(scan_win_std_dev[253]), .feature_accum(feature_accums[253]));
  accum_calculator #(.RECT1_X(rectangle1_xs[254]), .RECT1_Y(rectangle1_ys[254]), .RECT1_WIDTH(rectangle1_widths[254]), .RECT1_HEIGHT(rectangle1_heights[254]), .RECT1_WEIGHT(rectangle1_weights[254]), .RECT2_X(rectangle2_xs[254]), .RECT2_Y(rectangle2_ys[254]), .RECT2_WIDTH(rectangle2_widths[254]), .RECT2_HEIGHT(rectangle2_heights[254]), .RECT2_WEIGHT(rectangle2_weights[254]), .RECT3_X(rectangle3_xs[254]), .RECT3_Y(rectangle3_ys[254]), .RECT3_WIDTH(rectangle3_widths[254]), .RECT3_HEIGHT(rectangle3_heights[254]), .RECT3_WEIGHT(rectangle3_weights[254]), .FEAT_THRES(feature_thresholds[254]), .FEAT_ABOVE(feature_aboves[254]), .FEAT_BELOW(feature_belows[254])) ac254(.scan_win(scan_win254), .scan_win_std_dev(scan_win_std_dev[254]), .feature_accum(feature_accums[254]));
  accum_calculator #(.RECT1_X(rectangle1_xs[255]), .RECT1_Y(rectangle1_ys[255]), .RECT1_WIDTH(rectangle1_widths[255]), .RECT1_HEIGHT(rectangle1_heights[255]), .RECT1_WEIGHT(rectangle1_weights[255]), .RECT2_X(rectangle2_xs[255]), .RECT2_Y(rectangle2_ys[255]), .RECT2_WIDTH(rectangle2_widths[255]), .RECT2_HEIGHT(rectangle2_heights[255]), .RECT2_WEIGHT(rectangle2_weights[255]), .RECT3_X(rectangle3_xs[255]), .RECT3_Y(rectangle3_ys[255]), .RECT3_WIDTH(rectangle3_widths[255]), .RECT3_HEIGHT(rectangle3_heights[255]), .RECT3_WEIGHT(rectangle3_weights[255]), .FEAT_THRES(feature_thresholds[255]), .FEAT_ABOVE(feature_aboves[255]), .FEAT_BELOW(feature_belows[255])) ac255(.scan_win(scan_win255), .scan_win_std_dev(scan_win_std_dev[255]), .feature_accum(feature_accums[255]));
  accum_calculator #(.RECT1_X(rectangle1_xs[256]), .RECT1_Y(rectangle1_ys[256]), .RECT1_WIDTH(rectangle1_widths[256]), .RECT1_HEIGHT(rectangle1_heights[256]), .RECT1_WEIGHT(rectangle1_weights[256]), .RECT2_X(rectangle2_xs[256]), .RECT2_Y(rectangle2_ys[256]), .RECT2_WIDTH(rectangle2_widths[256]), .RECT2_HEIGHT(rectangle2_heights[256]), .RECT2_WEIGHT(rectangle2_weights[256]), .RECT3_X(rectangle3_xs[256]), .RECT3_Y(rectangle3_ys[256]), .RECT3_WIDTH(rectangle3_widths[256]), .RECT3_HEIGHT(rectangle3_heights[256]), .RECT3_WEIGHT(rectangle3_weights[256]), .FEAT_THRES(feature_thresholds[256]), .FEAT_ABOVE(feature_aboves[256]), .FEAT_BELOW(feature_belows[256])) ac256(.scan_win(scan_win256), .scan_win_std_dev(scan_win_std_dev[256]), .feature_accum(feature_accums[256]));
  accum_calculator #(.RECT1_X(rectangle1_xs[257]), .RECT1_Y(rectangle1_ys[257]), .RECT1_WIDTH(rectangle1_widths[257]), .RECT1_HEIGHT(rectangle1_heights[257]), .RECT1_WEIGHT(rectangle1_weights[257]), .RECT2_X(rectangle2_xs[257]), .RECT2_Y(rectangle2_ys[257]), .RECT2_WIDTH(rectangle2_widths[257]), .RECT2_HEIGHT(rectangle2_heights[257]), .RECT2_WEIGHT(rectangle2_weights[257]), .RECT3_X(rectangle3_xs[257]), .RECT3_Y(rectangle3_ys[257]), .RECT3_WIDTH(rectangle3_widths[257]), .RECT3_HEIGHT(rectangle3_heights[257]), .RECT3_WEIGHT(rectangle3_weights[257]), .FEAT_THRES(feature_thresholds[257]), .FEAT_ABOVE(feature_aboves[257]), .FEAT_BELOW(feature_belows[257])) ac257(.scan_win(scan_win257), .scan_win_std_dev(scan_win_std_dev[257]), .feature_accum(feature_accums[257]));
  accum_calculator #(.RECT1_X(rectangle1_xs[258]), .RECT1_Y(rectangle1_ys[258]), .RECT1_WIDTH(rectangle1_widths[258]), .RECT1_HEIGHT(rectangle1_heights[258]), .RECT1_WEIGHT(rectangle1_weights[258]), .RECT2_X(rectangle2_xs[258]), .RECT2_Y(rectangle2_ys[258]), .RECT2_WIDTH(rectangle2_widths[258]), .RECT2_HEIGHT(rectangle2_heights[258]), .RECT2_WEIGHT(rectangle2_weights[258]), .RECT3_X(rectangle3_xs[258]), .RECT3_Y(rectangle3_ys[258]), .RECT3_WIDTH(rectangle3_widths[258]), .RECT3_HEIGHT(rectangle3_heights[258]), .RECT3_WEIGHT(rectangle3_weights[258]), .FEAT_THRES(feature_thresholds[258]), .FEAT_ABOVE(feature_aboves[258]), .FEAT_BELOW(feature_belows[258])) ac258(.scan_win(scan_win258), .scan_win_std_dev(scan_win_std_dev[258]), .feature_accum(feature_accums[258]));
  accum_calculator #(.RECT1_X(rectangle1_xs[259]), .RECT1_Y(rectangle1_ys[259]), .RECT1_WIDTH(rectangle1_widths[259]), .RECT1_HEIGHT(rectangle1_heights[259]), .RECT1_WEIGHT(rectangle1_weights[259]), .RECT2_X(rectangle2_xs[259]), .RECT2_Y(rectangle2_ys[259]), .RECT2_WIDTH(rectangle2_widths[259]), .RECT2_HEIGHT(rectangle2_heights[259]), .RECT2_WEIGHT(rectangle2_weights[259]), .RECT3_X(rectangle3_xs[259]), .RECT3_Y(rectangle3_ys[259]), .RECT3_WIDTH(rectangle3_widths[259]), .RECT3_HEIGHT(rectangle3_heights[259]), .RECT3_WEIGHT(rectangle3_weights[259]), .FEAT_THRES(feature_thresholds[259]), .FEAT_ABOVE(feature_aboves[259]), .FEAT_BELOW(feature_belows[259])) ac259(.scan_win(scan_win259), .scan_win_std_dev(scan_win_std_dev[259]), .feature_accum(feature_accums[259]));
  accum_calculator #(.RECT1_X(rectangle1_xs[260]), .RECT1_Y(rectangle1_ys[260]), .RECT1_WIDTH(rectangle1_widths[260]), .RECT1_HEIGHT(rectangle1_heights[260]), .RECT1_WEIGHT(rectangle1_weights[260]), .RECT2_X(rectangle2_xs[260]), .RECT2_Y(rectangle2_ys[260]), .RECT2_WIDTH(rectangle2_widths[260]), .RECT2_HEIGHT(rectangle2_heights[260]), .RECT2_WEIGHT(rectangle2_weights[260]), .RECT3_X(rectangle3_xs[260]), .RECT3_Y(rectangle3_ys[260]), .RECT3_WIDTH(rectangle3_widths[260]), .RECT3_HEIGHT(rectangle3_heights[260]), .RECT3_WEIGHT(rectangle3_weights[260]), .FEAT_THRES(feature_thresholds[260]), .FEAT_ABOVE(feature_aboves[260]), .FEAT_BELOW(feature_belows[260])) ac260(.scan_win(scan_win260), .scan_win_std_dev(scan_win_std_dev[260]), .feature_accum(feature_accums[260]));
  accum_calculator #(.RECT1_X(rectangle1_xs[261]), .RECT1_Y(rectangle1_ys[261]), .RECT1_WIDTH(rectangle1_widths[261]), .RECT1_HEIGHT(rectangle1_heights[261]), .RECT1_WEIGHT(rectangle1_weights[261]), .RECT2_X(rectangle2_xs[261]), .RECT2_Y(rectangle2_ys[261]), .RECT2_WIDTH(rectangle2_widths[261]), .RECT2_HEIGHT(rectangle2_heights[261]), .RECT2_WEIGHT(rectangle2_weights[261]), .RECT3_X(rectangle3_xs[261]), .RECT3_Y(rectangle3_ys[261]), .RECT3_WIDTH(rectangle3_widths[261]), .RECT3_HEIGHT(rectangle3_heights[261]), .RECT3_WEIGHT(rectangle3_weights[261]), .FEAT_THRES(feature_thresholds[261]), .FEAT_ABOVE(feature_aboves[261]), .FEAT_BELOW(feature_belows[261])) ac261(.scan_win(scan_win261), .scan_win_std_dev(scan_win_std_dev[261]), .feature_accum(feature_accums[261]));
  accum_calculator #(.RECT1_X(rectangle1_xs[262]), .RECT1_Y(rectangle1_ys[262]), .RECT1_WIDTH(rectangle1_widths[262]), .RECT1_HEIGHT(rectangle1_heights[262]), .RECT1_WEIGHT(rectangle1_weights[262]), .RECT2_X(rectangle2_xs[262]), .RECT2_Y(rectangle2_ys[262]), .RECT2_WIDTH(rectangle2_widths[262]), .RECT2_HEIGHT(rectangle2_heights[262]), .RECT2_WEIGHT(rectangle2_weights[262]), .RECT3_X(rectangle3_xs[262]), .RECT3_Y(rectangle3_ys[262]), .RECT3_WIDTH(rectangle3_widths[262]), .RECT3_HEIGHT(rectangle3_heights[262]), .RECT3_WEIGHT(rectangle3_weights[262]), .FEAT_THRES(feature_thresholds[262]), .FEAT_ABOVE(feature_aboves[262]), .FEAT_BELOW(feature_belows[262])) ac262(.scan_win(scan_win262), .scan_win_std_dev(scan_win_std_dev[262]), .feature_accum(feature_accums[262]));
  accum_calculator #(.RECT1_X(rectangle1_xs[263]), .RECT1_Y(rectangle1_ys[263]), .RECT1_WIDTH(rectangle1_widths[263]), .RECT1_HEIGHT(rectangle1_heights[263]), .RECT1_WEIGHT(rectangle1_weights[263]), .RECT2_X(rectangle2_xs[263]), .RECT2_Y(rectangle2_ys[263]), .RECT2_WIDTH(rectangle2_widths[263]), .RECT2_HEIGHT(rectangle2_heights[263]), .RECT2_WEIGHT(rectangle2_weights[263]), .RECT3_X(rectangle3_xs[263]), .RECT3_Y(rectangle3_ys[263]), .RECT3_WIDTH(rectangle3_widths[263]), .RECT3_HEIGHT(rectangle3_heights[263]), .RECT3_WEIGHT(rectangle3_weights[263]), .FEAT_THRES(feature_thresholds[263]), .FEAT_ABOVE(feature_aboves[263]), .FEAT_BELOW(feature_belows[263])) ac263(.scan_win(scan_win263), .scan_win_std_dev(scan_win_std_dev[263]), .feature_accum(feature_accums[263]));
  accum_calculator #(.RECT1_X(rectangle1_xs[264]), .RECT1_Y(rectangle1_ys[264]), .RECT1_WIDTH(rectangle1_widths[264]), .RECT1_HEIGHT(rectangle1_heights[264]), .RECT1_WEIGHT(rectangle1_weights[264]), .RECT2_X(rectangle2_xs[264]), .RECT2_Y(rectangle2_ys[264]), .RECT2_WIDTH(rectangle2_widths[264]), .RECT2_HEIGHT(rectangle2_heights[264]), .RECT2_WEIGHT(rectangle2_weights[264]), .RECT3_X(rectangle3_xs[264]), .RECT3_Y(rectangle3_ys[264]), .RECT3_WIDTH(rectangle3_widths[264]), .RECT3_HEIGHT(rectangle3_heights[264]), .RECT3_WEIGHT(rectangle3_weights[264]), .FEAT_THRES(feature_thresholds[264]), .FEAT_ABOVE(feature_aboves[264]), .FEAT_BELOW(feature_belows[264])) ac264(.scan_win(scan_win264), .scan_win_std_dev(scan_win_std_dev[264]), .feature_accum(feature_accums[264]));
  accum_calculator #(.RECT1_X(rectangle1_xs[265]), .RECT1_Y(rectangle1_ys[265]), .RECT1_WIDTH(rectangle1_widths[265]), .RECT1_HEIGHT(rectangle1_heights[265]), .RECT1_WEIGHT(rectangle1_weights[265]), .RECT2_X(rectangle2_xs[265]), .RECT2_Y(rectangle2_ys[265]), .RECT2_WIDTH(rectangle2_widths[265]), .RECT2_HEIGHT(rectangle2_heights[265]), .RECT2_WEIGHT(rectangle2_weights[265]), .RECT3_X(rectangle3_xs[265]), .RECT3_Y(rectangle3_ys[265]), .RECT3_WIDTH(rectangle3_widths[265]), .RECT3_HEIGHT(rectangle3_heights[265]), .RECT3_WEIGHT(rectangle3_weights[265]), .FEAT_THRES(feature_thresholds[265]), .FEAT_ABOVE(feature_aboves[265]), .FEAT_BELOW(feature_belows[265])) ac265(.scan_win(scan_win265), .scan_win_std_dev(scan_win_std_dev[265]), .feature_accum(feature_accums[265]));
  accum_calculator #(.RECT1_X(rectangle1_xs[266]), .RECT1_Y(rectangle1_ys[266]), .RECT1_WIDTH(rectangle1_widths[266]), .RECT1_HEIGHT(rectangle1_heights[266]), .RECT1_WEIGHT(rectangle1_weights[266]), .RECT2_X(rectangle2_xs[266]), .RECT2_Y(rectangle2_ys[266]), .RECT2_WIDTH(rectangle2_widths[266]), .RECT2_HEIGHT(rectangle2_heights[266]), .RECT2_WEIGHT(rectangle2_weights[266]), .RECT3_X(rectangle3_xs[266]), .RECT3_Y(rectangle3_ys[266]), .RECT3_WIDTH(rectangle3_widths[266]), .RECT3_HEIGHT(rectangle3_heights[266]), .RECT3_WEIGHT(rectangle3_weights[266]), .FEAT_THRES(feature_thresholds[266]), .FEAT_ABOVE(feature_aboves[266]), .FEAT_BELOW(feature_belows[266])) ac266(.scan_win(scan_win266), .scan_win_std_dev(scan_win_std_dev[266]), .feature_accum(feature_accums[266]));
  accum_calculator #(.RECT1_X(rectangle1_xs[267]), .RECT1_Y(rectangle1_ys[267]), .RECT1_WIDTH(rectangle1_widths[267]), .RECT1_HEIGHT(rectangle1_heights[267]), .RECT1_WEIGHT(rectangle1_weights[267]), .RECT2_X(rectangle2_xs[267]), .RECT2_Y(rectangle2_ys[267]), .RECT2_WIDTH(rectangle2_widths[267]), .RECT2_HEIGHT(rectangle2_heights[267]), .RECT2_WEIGHT(rectangle2_weights[267]), .RECT3_X(rectangle3_xs[267]), .RECT3_Y(rectangle3_ys[267]), .RECT3_WIDTH(rectangle3_widths[267]), .RECT3_HEIGHT(rectangle3_heights[267]), .RECT3_WEIGHT(rectangle3_weights[267]), .FEAT_THRES(feature_thresholds[267]), .FEAT_ABOVE(feature_aboves[267]), .FEAT_BELOW(feature_belows[267])) ac267(.scan_win(scan_win267), .scan_win_std_dev(scan_win_std_dev[267]), .feature_accum(feature_accums[267]));
  accum_calculator #(.RECT1_X(rectangle1_xs[268]), .RECT1_Y(rectangle1_ys[268]), .RECT1_WIDTH(rectangle1_widths[268]), .RECT1_HEIGHT(rectangle1_heights[268]), .RECT1_WEIGHT(rectangle1_weights[268]), .RECT2_X(rectangle2_xs[268]), .RECT2_Y(rectangle2_ys[268]), .RECT2_WIDTH(rectangle2_widths[268]), .RECT2_HEIGHT(rectangle2_heights[268]), .RECT2_WEIGHT(rectangle2_weights[268]), .RECT3_X(rectangle3_xs[268]), .RECT3_Y(rectangle3_ys[268]), .RECT3_WIDTH(rectangle3_widths[268]), .RECT3_HEIGHT(rectangle3_heights[268]), .RECT3_WEIGHT(rectangle3_weights[268]), .FEAT_THRES(feature_thresholds[268]), .FEAT_ABOVE(feature_aboves[268]), .FEAT_BELOW(feature_belows[268])) ac268(.scan_win(scan_win268), .scan_win_std_dev(scan_win_std_dev[268]), .feature_accum(feature_accums[268]));
  accum_calculator #(.RECT1_X(rectangle1_xs[269]), .RECT1_Y(rectangle1_ys[269]), .RECT1_WIDTH(rectangle1_widths[269]), .RECT1_HEIGHT(rectangle1_heights[269]), .RECT1_WEIGHT(rectangle1_weights[269]), .RECT2_X(rectangle2_xs[269]), .RECT2_Y(rectangle2_ys[269]), .RECT2_WIDTH(rectangle2_widths[269]), .RECT2_HEIGHT(rectangle2_heights[269]), .RECT2_WEIGHT(rectangle2_weights[269]), .RECT3_X(rectangle3_xs[269]), .RECT3_Y(rectangle3_ys[269]), .RECT3_WIDTH(rectangle3_widths[269]), .RECT3_HEIGHT(rectangle3_heights[269]), .RECT3_WEIGHT(rectangle3_weights[269]), .FEAT_THRES(feature_thresholds[269]), .FEAT_ABOVE(feature_aboves[269]), .FEAT_BELOW(feature_belows[269])) ac269(.scan_win(scan_win269), .scan_win_std_dev(scan_win_std_dev[269]), .feature_accum(feature_accums[269]));
  accum_calculator #(.RECT1_X(rectangle1_xs[270]), .RECT1_Y(rectangle1_ys[270]), .RECT1_WIDTH(rectangle1_widths[270]), .RECT1_HEIGHT(rectangle1_heights[270]), .RECT1_WEIGHT(rectangle1_weights[270]), .RECT2_X(rectangle2_xs[270]), .RECT2_Y(rectangle2_ys[270]), .RECT2_WIDTH(rectangle2_widths[270]), .RECT2_HEIGHT(rectangle2_heights[270]), .RECT2_WEIGHT(rectangle2_weights[270]), .RECT3_X(rectangle3_xs[270]), .RECT3_Y(rectangle3_ys[270]), .RECT3_WIDTH(rectangle3_widths[270]), .RECT3_HEIGHT(rectangle3_heights[270]), .RECT3_WEIGHT(rectangle3_weights[270]), .FEAT_THRES(feature_thresholds[270]), .FEAT_ABOVE(feature_aboves[270]), .FEAT_BELOW(feature_belows[270])) ac270(.scan_win(scan_win270), .scan_win_std_dev(scan_win_std_dev[270]), .feature_accum(feature_accums[270]));
  accum_calculator #(.RECT1_X(rectangle1_xs[271]), .RECT1_Y(rectangle1_ys[271]), .RECT1_WIDTH(rectangle1_widths[271]), .RECT1_HEIGHT(rectangle1_heights[271]), .RECT1_WEIGHT(rectangle1_weights[271]), .RECT2_X(rectangle2_xs[271]), .RECT2_Y(rectangle2_ys[271]), .RECT2_WIDTH(rectangle2_widths[271]), .RECT2_HEIGHT(rectangle2_heights[271]), .RECT2_WEIGHT(rectangle2_weights[271]), .RECT3_X(rectangle3_xs[271]), .RECT3_Y(rectangle3_ys[271]), .RECT3_WIDTH(rectangle3_widths[271]), .RECT3_HEIGHT(rectangle3_heights[271]), .RECT3_WEIGHT(rectangle3_weights[271]), .FEAT_THRES(feature_thresholds[271]), .FEAT_ABOVE(feature_aboves[271]), .FEAT_BELOW(feature_belows[271])) ac271(.scan_win(scan_win271), .scan_win_std_dev(scan_win_std_dev[271]), .feature_accum(feature_accums[271]));
  accum_calculator #(.RECT1_X(rectangle1_xs[272]), .RECT1_Y(rectangle1_ys[272]), .RECT1_WIDTH(rectangle1_widths[272]), .RECT1_HEIGHT(rectangle1_heights[272]), .RECT1_WEIGHT(rectangle1_weights[272]), .RECT2_X(rectangle2_xs[272]), .RECT2_Y(rectangle2_ys[272]), .RECT2_WIDTH(rectangle2_widths[272]), .RECT2_HEIGHT(rectangle2_heights[272]), .RECT2_WEIGHT(rectangle2_weights[272]), .RECT3_X(rectangle3_xs[272]), .RECT3_Y(rectangle3_ys[272]), .RECT3_WIDTH(rectangle3_widths[272]), .RECT3_HEIGHT(rectangle3_heights[272]), .RECT3_WEIGHT(rectangle3_weights[272]), .FEAT_THRES(feature_thresholds[272]), .FEAT_ABOVE(feature_aboves[272]), .FEAT_BELOW(feature_belows[272])) ac272(.scan_win(scan_win272), .scan_win_std_dev(scan_win_std_dev[272]), .feature_accum(feature_accums[272]));
  accum_calculator #(.RECT1_X(rectangle1_xs[273]), .RECT1_Y(rectangle1_ys[273]), .RECT1_WIDTH(rectangle1_widths[273]), .RECT1_HEIGHT(rectangle1_heights[273]), .RECT1_WEIGHT(rectangle1_weights[273]), .RECT2_X(rectangle2_xs[273]), .RECT2_Y(rectangle2_ys[273]), .RECT2_WIDTH(rectangle2_widths[273]), .RECT2_HEIGHT(rectangle2_heights[273]), .RECT2_WEIGHT(rectangle2_weights[273]), .RECT3_X(rectangle3_xs[273]), .RECT3_Y(rectangle3_ys[273]), .RECT3_WIDTH(rectangle3_widths[273]), .RECT3_HEIGHT(rectangle3_heights[273]), .RECT3_WEIGHT(rectangle3_weights[273]), .FEAT_THRES(feature_thresholds[273]), .FEAT_ABOVE(feature_aboves[273]), .FEAT_BELOW(feature_belows[273])) ac273(.scan_win(scan_win273), .scan_win_std_dev(scan_win_std_dev[273]), .feature_accum(feature_accums[273]));
  accum_calculator #(.RECT1_X(rectangle1_xs[274]), .RECT1_Y(rectangle1_ys[274]), .RECT1_WIDTH(rectangle1_widths[274]), .RECT1_HEIGHT(rectangle1_heights[274]), .RECT1_WEIGHT(rectangle1_weights[274]), .RECT2_X(rectangle2_xs[274]), .RECT2_Y(rectangle2_ys[274]), .RECT2_WIDTH(rectangle2_widths[274]), .RECT2_HEIGHT(rectangle2_heights[274]), .RECT2_WEIGHT(rectangle2_weights[274]), .RECT3_X(rectangle3_xs[274]), .RECT3_Y(rectangle3_ys[274]), .RECT3_WIDTH(rectangle3_widths[274]), .RECT3_HEIGHT(rectangle3_heights[274]), .RECT3_WEIGHT(rectangle3_weights[274]), .FEAT_THRES(feature_thresholds[274]), .FEAT_ABOVE(feature_aboves[274]), .FEAT_BELOW(feature_belows[274])) ac274(.scan_win(scan_win274), .scan_win_std_dev(scan_win_std_dev[274]), .feature_accum(feature_accums[274]));
  accum_calculator #(.RECT1_X(rectangle1_xs[275]), .RECT1_Y(rectangle1_ys[275]), .RECT1_WIDTH(rectangle1_widths[275]), .RECT1_HEIGHT(rectangle1_heights[275]), .RECT1_WEIGHT(rectangle1_weights[275]), .RECT2_X(rectangle2_xs[275]), .RECT2_Y(rectangle2_ys[275]), .RECT2_WIDTH(rectangle2_widths[275]), .RECT2_HEIGHT(rectangle2_heights[275]), .RECT2_WEIGHT(rectangle2_weights[275]), .RECT3_X(rectangle3_xs[275]), .RECT3_Y(rectangle3_ys[275]), .RECT3_WIDTH(rectangle3_widths[275]), .RECT3_HEIGHT(rectangle3_heights[275]), .RECT3_WEIGHT(rectangle3_weights[275]), .FEAT_THRES(feature_thresholds[275]), .FEAT_ABOVE(feature_aboves[275]), .FEAT_BELOW(feature_belows[275])) ac275(.scan_win(scan_win275), .scan_win_std_dev(scan_win_std_dev[275]), .feature_accum(feature_accums[275]));
  accum_calculator #(.RECT1_X(rectangle1_xs[276]), .RECT1_Y(rectangle1_ys[276]), .RECT1_WIDTH(rectangle1_widths[276]), .RECT1_HEIGHT(rectangle1_heights[276]), .RECT1_WEIGHT(rectangle1_weights[276]), .RECT2_X(rectangle2_xs[276]), .RECT2_Y(rectangle2_ys[276]), .RECT2_WIDTH(rectangle2_widths[276]), .RECT2_HEIGHT(rectangle2_heights[276]), .RECT2_WEIGHT(rectangle2_weights[276]), .RECT3_X(rectangle3_xs[276]), .RECT3_Y(rectangle3_ys[276]), .RECT3_WIDTH(rectangle3_widths[276]), .RECT3_HEIGHT(rectangle3_heights[276]), .RECT3_WEIGHT(rectangle3_weights[276]), .FEAT_THRES(feature_thresholds[276]), .FEAT_ABOVE(feature_aboves[276]), .FEAT_BELOW(feature_belows[276])) ac276(.scan_win(scan_win276), .scan_win_std_dev(scan_win_std_dev[276]), .feature_accum(feature_accums[276]));
  accum_calculator #(.RECT1_X(rectangle1_xs[277]), .RECT1_Y(rectangle1_ys[277]), .RECT1_WIDTH(rectangle1_widths[277]), .RECT1_HEIGHT(rectangle1_heights[277]), .RECT1_WEIGHT(rectangle1_weights[277]), .RECT2_X(rectangle2_xs[277]), .RECT2_Y(rectangle2_ys[277]), .RECT2_WIDTH(rectangle2_widths[277]), .RECT2_HEIGHT(rectangle2_heights[277]), .RECT2_WEIGHT(rectangle2_weights[277]), .RECT3_X(rectangle3_xs[277]), .RECT3_Y(rectangle3_ys[277]), .RECT3_WIDTH(rectangle3_widths[277]), .RECT3_HEIGHT(rectangle3_heights[277]), .RECT3_WEIGHT(rectangle3_weights[277]), .FEAT_THRES(feature_thresholds[277]), .FEAT_ABOVE(feature_aboves[277]), .FEAT_BELOW(feature_belows[277])) ac277(.scan_win(scan_win277), .scan_win_std_dev(scan_win_std_dev[277]), .feature_accum(feature_accums[277]));
  accum_calculator #(.RECT1_X(rectangle1_xs[278]), .RECT1_Y(rectangle1_ys[278]), .RECT1_WIDTH(rectangle1_widths[278]), .RECT1_HEIGHT(rectangle1_heights[278]), .RECT1_WEIGHT(rectangle1_weights[278]), .RECT2_X(rectangle2_xs[278]), .RECT2_Y(rectangle2_ys[278]), .RECT2_WIDTH(rectangle2_widths[278]), .RECT2_HEIGHT(rectangle2_heights[278]), .RECT2_WEIGHT(rectangle2_weights[278]), .RECT3_X(rectangle3_xs[278]), .RECT3_Y(rectangle3_ys[278]), .RECT3_WIDTH(rectangle3_widths[278]), .RECT3_HEIGHT(rectangle3_heights[278]), .RECT3_WEIGHT(rectangle3_weights[278]), .FEAT_THRES(feature_thresholds[278]), .FEAT_ABOVE(feature_aboves[278]), .FEAT_BELOW(feature_belows[278])) ac278(.scan_win(scan_win278), .scan_win_std_dev(scan_win_std_dev[278]), .feature_accum(feature_accums[278]));
  accum_calculator #(.RECT1_X(rectangle1_xs[279]), .RECT1_Y(rectangle1_ys[279]), .RECT1_WIDTH(rectangle1_widths[279]), .RECT1_HEIGHT(rectangle1_heights[279]), .RECT1_WEIGHT(rectangle1_weights[279]), .RECT2_X(rectangle2_xs[279]), .RECT2_Y(rectangle2_ys[279]), .RECT2_WIDTH(rectangle2_widths[279]), .RECT2_HEIGHT(rectangle2_heights[279]), .RECT2_WEIGHT(rectangle2_weights[279]), .RECT3_X(rectangle3_xs[279]), .RECT3_Y(rectangle3_ys[279]), .RECT3_WIDTH(rectangle3_widths[279]), .RECT3_HEIGHT(rectangle3_heights[279]), .RECT3_WEIGHT(rectangle3_weights[279]), .FEAT_THRES(feature_thresholds[279]), .FEAT_ABOVE(feature_aboves[279]), .FEAT_BELOW(feature_belows[279])) ac279(.scan_win(scan_win279), .scan_win_std_dev(scan_win_std_dev[279]), .feature_accum(feature_accums[279]));
  accum_calculator #(.RECT1_X(rectangle1_xs[280]), .RECT1_Y(rectangle1_ys[280]), .RECT1_WIDTH(rectangle1_widths[280]), .RECT1_HEIGHT(rectangle1_heights[280]), .RECT1_WEIGHT(rectangle1_weights[280]), .RECT2_X(rectangle2_xs[280]), .RECT2_Y(rectangle2_ys[280]), .RECT2_WIDTH(rectangle2_widths[280]), .RECT2_HEIGHT(rectangle2_heights[280]), .RECT2_WEIGHT(rectangle2_weights[280]), .RECT3_X(rectangle3_xs[280]), .RECT3_Y(rectangle3_ys[280]), .RECT3_WIDTH(rectangle3_widths[280]), .RECT3_HEIGHT(rectangle3_heights[280]), .RECT3_WEIGHT(rectangle3_weights[280]), .FEAT_THRES(feature_thresholds[280]), .FEAT_ABOVE(feature_aboves[280]), .FEAT_BELOW(feature_belows[280])) ac280(.scan_win(scan_win280), .scan_win_std_dev(scan_win_std_dev[280]), .feature_accum(feature_accums[280]));
  accum_calculator #(.RECT1_X(rectangle1_xs[281]), .RECT1_Y(rectangle1_ys[281]), .RECT1_WIDTH(rectangle1_widths[281]), .RECT1_HEIGHT(rectangle1_heights[281]), .RECT1_WEIGHT(rectangle1_weights[281]), .RECT2_X(rectangle2_xs[281]), .RECT2_Y(rectangle2_ys[281]), .RECT2_WIDTH(rectangle2_widths[281]), .RECT2_HEIGHT(rectangle2_heights[281]), .RECT2_WEIGHT(rectangle2_weights[281]), .RECT3_X(rectangle3_xs[281]), .RECT3_Y(rectangle3_ys[281]), .RECT3_WIDTH(rectangle3_widths[281]), .RECT3_HEIGHT(rectangle3_heights[281]), .RECT3_WEIGHT(rectangle3_weights[281]), .FEAT_THRES(feature_thresholds[281]), .FEAT_ABOVE(feature_aboves[281]), .FEAT_BELOW(feature_belows[281])) ac281(.scan_win(scan_win281), .scan_win_std_dev(scan_win_std_dev[281]), .feature_accum(feature_accums[281]));
  accum_calculator #(.RECT1_X(rectangle1_xs[282]), .RECT1_Y(rectangle1_ys[282]), .RECT1_WIDTH(rectangle1_widths[282]), .RECT1_HEIGHT(rectangle1_heights[282]), .RECT1_WEIGHT(rectangle1_weights[282]), .RECT2_X(rectangle2_xs[282]), .RECT2_Y(rectangle2_ys[282]), .RECT2_WIDTH(rectangle2_widths[282]), .RECT2_HEIGHT(rectangle2_heights[282]), .RECT2_WEIGHT(rectangle2_weights[282]), .RECT3_X(rectangle3_xs[282]), .RECT3_Y(rectangle3_ys[282]), .RECT3_WIDTH(rectangle3_widths[282]), .RECT3_HEIGHT(rectangle3_heights[282]), .RECT3_WEIGHT(rectangle3_weights[282]), .FEAT_THRES(feature_thresholds[282]), .FEAT_ABOVE(feature_aboves[282]), .FEAT_BELOW(feature_belows[282])) ac282(.scan_win(scan_win282), .scan_win_std_dev(scan_win_std_dev[282]), .feature_accum(feature_accums[282]));
  accum_calculator #(.RECT1_X(rectangle1_xs[283]), .RECT1_Y(rectangle1_ys[283]), .RECT1_WIDTH(rectangle1_widths[283]), .RECT1_HEIGHT(rectangle1_heights[283]), .RECT1_WEIGHT(rectangle1_weights[283]), .RECT2_X(rectangle2_xs[283]), .RECT2_Y(rectangle2_ys[283]), .RECT2_WIDTH(rectangle2_widths[283]), .RECT2_HEIGHT(rectangle2_heights[283]), .RECT2_WEIGHT(rectangle2_weights[283]), .RECT3_X(rectangle3_xs[283]), .RECT3_Y(rectangle3_ys[283]), .RECT3_WIDTH(rectangle3_widths[283]), .RECT3_HEIGHT(rectangle3_heights[283]), .RECT3_WEIGHT(rectangle3_weights[283]), .FEAT_THRES(feature_thresholds[283]), .FEAT_ABOVE(feature_aboves[283]), .FEAT_BELOW(feature_belows[283])) ac283(.scan_win(scan_win283), .scan_win_std_dev(scan_win_std_dev[283]), .feature_accum(feature_accums[283]));
  accum_calculator #(.RECT1_X(rectangle1_xs[284]), .RECT1_Y(rectangle1_ys[284]), .RECT1_WIDTH(rectangle1_widths[284]), .RECT1_HEIGHT(rectangle1_heights[284]), .RECT1_WEIGHT(rectangle1_weights[284]), .RECT2_X(rectangle2_xs[284]), .RECT2_Y(rectangle2_ys[284]), .RECT2_WIDTH(rectangle2_widths[284]), .RECT2_HEIGHT(rectangle2_heights[284]), .RECT2_WEIGHT(rectangle2_weights[284]), .RECT3_X(rectangle3_xs[284]), .RECT3_Y(rectangle3_ys[284]), .RECT3_WIDTH(rectangle3_widths[284]), .RECT3_HEIGHT(rectangle3_heights[284]), .RECT3_WEIGHT(rectangle3_weights[284]), .FEAT_THRES(feature_thresholds[284]), .FEAT_ABOVE(feature_aboves[284]), .FEAT_BELOW(feature_belows[284])) ac284(.scan_win(scan_win284), .scan_win_std_dev(scan_win_std_dev[284]), .feature_accum(feature_accums[284]));
  accum_calculator #(.RECT1_X(rectangle1_xs[285]), .RECT1_Y(rectangle1_ys[285]), .RECT1_WIDTH(rectangle1_widths[285]), .RECT1_HEIGHT(rectangle1_heights[285]), .RECT1_WEIGHT(rectangle1_weights[285]), .RECT2_X(rectangle2_xs[285]), .RECT2_Y(rectangle2_ys[285]), .RECT2_WIDTH(rectangle2_widths[285]), .RECT2_HEIGHT(rectangle2_heights[285]), .RECT2_WEIGHT(rectangle2_weights[285]), .RECT3_X(rectangle3_xs[285]), .RECT3_Y(rectangle3_ys[285]), .RECT3_WIDTH(rectangle3_widths[285]), .RECT3_HEIGHT(rectangle3_heights[285]), .RECT3_WEIGHT(rectangle3_weights[285]), .FEAT_THRES(feature_thresholds[285]), .FEAT_ABOVE(feature_aboves[285]), .FEAT_BELOW(feature_belows[285])) ac285(.scan_win(scan_win285), .scan_win_std_dev(scan_win_std_dev[285]), .feature_accum(feature_accums[285]));
  accum_calculator #(.RECT1_X(rectangle1_xs[286]), .RECT1_Y(rectangle1_ys[286]), .RECT1_WIDTH(rectangle1_widths[286]), .RECT1_HEIGHT(rectangle1_heights[286]), .RECT1_WEIGHT(rectangle1_weights[286]), .RECT2_X(rectangle2_xs[286]), .RECT2_Y(rectangle2_ys[286]), .RECT2_WIDTH(rectangle2_widths[286]), .RECT2_HEIGHT(rectangle2_heights[286]), .RECT2_WEIGHT(rectangle2_weights[286]), .RECT3_X(rectangle3_xs[286]), .RECT3_Y(rectangle3_ys[286]), .RECT3_WIDTH(rectangle3_widths[286]), .RECT3_HEIGHT(rectangle3_heights[286]), .RECT3_WEIGHT(rectangle3_weights[286]), .FEAT_THRES(feature_thresholds[286]), .FEAT_ABOVE(feature_aboves[286]), .FEAT_BELOW(feature_belows[286])) ac286(.scan_win(scan_win286), .scan_win_std_dev(scan_win_std_dev[286]), .feature_accum(feature_accums[286]));
  accum_calculator #(.RECT1_X(rectangle1_xs[287]), .RECT1_Y(rectangle1_ys[287]), .RECT1_WIDTH(rectangle1_widths[287]), .RECT1_HEIGHT(rectangle1_heights[287]), .RECT1_WEIGHT(rectangle1_weights[287]), .RECT2_X(rectangle2_xs[287]), .RECT2_Y(rectangle2_ys[287]), .RECT2_WIDTH(rectangle2_widths[287]), .RECT2_HEIGHT(rectangle2_heights[287]), .RECT2_WEIGHT(rectangle2_weights[287]), .RECT3_X(rectangle3_xs[287]), .RECT3_Y(rectangle3_ys[287]), .RECT3_WIDTH(rectangle3_widths[287]), .RECT3_HEIGHT(rectangle3_heights[287]), .RECT3_WEIGHT(rectangle3_weights[287]), .FEAT_THRES(feature_thresholds[287]), .FEAT_ABOVE(feature_aboves[287]), .FEAT_BELOW(feature_belows[287])) ac287(.scan_win(scan_win287), .scan_win_std_dev(scan_win_std_dev[287]), .feature_accum(feature_accums[287]));
  accum_calculator #(.RECT1_X(rectangle1_xs[288]), .RECT1_Y(rectangle1_ys[288]), .RECT1_WIDTH(rectangle1_widths[288]), .RECT1_HEIGHT(rectangle1_heights[288]), .RECT1_WEIGHT(rectangle1_weights[288]), .RECT2_X(rectangle2_xs[288]), .RECT2_Y(rectangle2_ys[288]), .RECT2_WIDTH(rectangle2_widths[288]), .RECT2_HEIGHT(rectangle2_heights[288]), .RECT2_WEIGHT(rectangle2_weights[288]), .RECT3_X(rectangle3_xs[288]), .RECT3_Y(rectangle3_ys[288]), .RECT3_WIDTH(rectangle3_widths[288]), .RECT3_HEIGHT(rectangle3_heights[288]), .RECT3_WEIGHT(rectangle3_weights[288]), .FEAT_THRES(feature_thresholds[288]), .FEAT_ABOVE(feature_aboves[288]), .FEAT_BELOW(feature_belows[288])) ac288(.scan_win(scan_win288), .scan_win_std_dev(scan_win_std_dev[288]), .feature_accum(feature_accums[288]));
  accum_calculator #(.RECT1_X(rectangle1_xs[289]), .RECT1_Y(rectangle1_ys[289]), .RECT1_WIDTH(rectangle1_widths[289]), .RECT1_HEIGHT(rectangle1_heights[289]), .RECT1_WEIGHT(rectangle1_weights[289]), .RECT2_X(rectangle2_xs[289]), .RECT2_Y(rectangle2_ys[289]), .RECT2_WIDTH(rectangle2_widths[289]), .RECT2_HEIGHT(rectangle2_heights[289]), .RECT2_WEIGHT(rectangle2_weights[289]), .RECT3_X(rectangle3_xs[289]), .RECT3_Y(rectangle3_ys[289]), .RECT3_WIDTH(rectangle3_widths[289]), .RECT3_HEIGHT(rectangle3_heights[289]), .RECT3_WEIGHT(rectangle3_weights[289]), .FEAT_THRES(feature_thresholds[289]), .FEAT_ABOVE(feature_aboves[289]), .FEAT_BELOW(feature_belows[289])) ac289(.scan_win(scan_win289), .scan_win_std_dev(scan_win_std_dev[289]), .feature_accum(feature_accums[289]));
  accum_calculator #(.RECT1_X(rectangle1_xs[290]), .RECT1_Y(rectangle1_ys[290]), .RECT1_WIDTH(rectangle1_widths[290]), .RECT1_HEIGHT(rectangle1_heights[290]), .RECT1_WEIGHT(rectangle1_weights[290]), .RECT2_X(rectangle2_xs[290]), .RECT2_Y(rectangle2_ys[290]), .RECT2_WIDTH(rectangle2_widths[290]), .RECT2_HEIGHT(rectangle2_heights[290]), .RECT2_WEIGHT(rectangle2_weights[290]), .RECT3_X(rectangle3_xs[290]), .RECT3_Y(rectangle3_ys[290]), .RECT3_WIDTH(rectangle3_widths[290]), .RECT3_HEIGHT(rectangle3_heights[290]), .RECT3_WEIGHT(rectangle3_weights[290]), .FEAT_THRES(feature_thresholds[290]), .FEAT_ABOVE(feature_aboves[290]), .FEAT_BELOW(feature_belows[290])) ac290(.scan_win(scan_win290), .scan_win_std_dev(scan_win_std_dev[290]), .feature_accum(feature_accums[290]));
  accum_calculator #(.RECT1_X(rectangle1_xs[291]), .RECT1_Y(rectangle1_ys[291]), .RECT1_WIDTH(rectangle1_widths[291]), .RECT1_HEIGHT(rectangle1_heights[291]), .RECT1_WEIGHT(rectangle1_weights[291]), .RECT2_X(rectangle2_xs[291]), .RECT2_Y(rectangle2_ys[291]), .RECT2_WIDTH(rectangle2_widths[291]), .RECT2_HEIGHT(rectangle2_heights[291]), .RECT2_WEIGHT(rectangle2_weights[291]), .RECT3_X(rectangle3_xs[291]), .RECT3_Y(rectangle3_ys[291]), .RECT3_WIDTH(rectangle3_widths[291]), .RECT3_HEIGHT(rectangle3_heights[291]), .RECT3_WEIGHT(rectangle3_weights[291]), .FEAT_THRES(feature_thresholds[291]), .FEAT_ABOVE(feature_aboves[291]), .FEAT_BELOW(feature_belows[291])) ac291(.scan_win(scan_win291), .scan_win_std_dev(scan_win_std_dev[291]), .feature_accum(feature_accums[291]));
  accum_calculator #(.RECT1_X(rectangle1_xs[292]), .RECT1_Y(rectangle1_ys[292]), .RECT1_WIDTH(rectangle1_widths[292]), .RECT1_HEIGHT(rectangle1_heights[292]), .RECT1_WEIGHT(rectangle1_weights[292]), .RECT2_X(rectangle2_xs[292]), .RECT2_Y(rectangle2_ys[292]), .RECT2_WIDTH(rectangle2_widths[292]), .RECT2_HEIGHT(rectangle2_heights[292]), .RECT2_WEIGHT(rectangle2_weights[292]), .RECT3_X(rectangle3_xs[292]), .RECT3_Y(rectangle3_ys[292]), .RECT3_WIDTH(rectangle3_widths[292]), .RECT3_HEIGHT(rectangle3_heights[292]), .RECT3_WEIGHT(rectangle3_weights[292]), .FEAT_THRES(feature_thresholds[292]), .FEAT_ABOVE(feature_aboves[292]), .FEAT_BELOW(feature_belows[292])) ac292(.scan_win(scan_win292), .scan_win_std_dev(scan_win_std_dev[292]), .feature_accum(feature_accums[292]));
  accum_calculator #(.RECT1_X(rectangle1_xs[293]), .RECT1_Y(rectangle1_ys[293]), .RECT1_WIDTH(rectangle1_widths[293]), .RECT1_HEIGHT(rectangle1_heights[293]), .RECT1_WEIGHT(rectangle1_weights[293]), .RECT2_X(rectangle2_xs[293]), .RECT2_Y(rectangle2_ys[293]), .RECT2_WIDTH(rectangle2_widths[293]), .RECT2_HEIGHT(rectangle2_heights[293]), .RECT2_WEIGHT(rectangle2_weights[293]), .RECT3_X(rectangle3_xs[293]), .RECT3_Y(rectangle3_ys[293]), .RECT3_WIDTH(rectangle3_widths[293]), .RECT3_HEIGHT(rectangle3_heights[293]), .RECT3_WEIGHT(rectangle3_weights[293]), .FEAT_THRES(feature_thresholds[293]), .FEAT_ABOVE(feature_aboves[293]), .FEAT_BELOW(feature_belows[293])) ac293(.scan_win(scan_win293), .scan_win_std_dev(scan_win_std_dev[293]), .feature_accum(feature_accums[293]));
  accum_calculator #(.RECT1_X(rectangle1_xs[294]), .RECT1_Y(rectangle1_ys[294]), .RECT1_WIDTH(rectangle1_widths[294]), .RECT1_HEIGHT(rectangle1_heights[294]), .RECT1_WEIGHT(rectangle1_weights[294]), .RECT2_X(rectangle2_xs[294]), .RECT2_Y(rectangle2_ys[294]), .RECT2_WIDTH(rectangle2_widths[294]), .RECT2_HEIGHT(rectangle2_heights[294]), .RECT2_WEIGHT(rectangle2_weights[294]), .RECT3_X(rectangle3_xs[294]), .RECT3_Y(rectangle3_ys[294]), .RECT3_WIDTH(rectangle3_widths[294]), .RECT3_HEIGHT(rectangle3_heights[294]), .RECT3_WEIGHT(rectangle3_weights[294]), .FEAT_THRES(feature_thresholds[294]), .FEAT_ABOVE(feature_aboves[294]), .FEAT_BELOW(feature_belows[294])) ac294(.scan_win(scan_win294), .scan_win_std_dev(scan_win_std_dev[294]), .feature_accum(feature_accums[294]));
  accum_calculator #(.RECT1_X(rectangle1_xs[295]), .RECT1_Y(rectangle1_ys[295]), .RECT1_WIDTH(rectangle1_widths[295]), .RECT1_HEIGHT(rectangle1_heights[295]), .RECT1_WEIGHT(rectangle1_weights[295]), .RECT2_X(rectangle2_xs[295]), .RECT2_Y(rectangle2_ys[295]), .RECT2_WIDTH(rectangle2_widths[295]), .RECT2_HEIGHT(rectangle2_heights[295]), .RECT2_WEIGHT(rectangle2_weights[295]), .RECT3_X(rectangle3_xs[295]), .RECT3_Y(rectangle3_ys[295]), .RECT3_WIDTH(rectangle3_widths[295]), .RECT3_HEIGHT(rectangle3_heights[295]), .RECT3_WEIGHT(rectangle3_weights[295]), .FEAT_THRES(feature_thresholds[295]), .FEAT_ABOVE(feature_aboves[295]), .FEAT_BELOW(feature_belows[295])) ac295(.scan_win(scan_win295), .scan_win_std_dev(scan_win_std_dev[295]), .feature_accum(feature_accums[295]));
  accum_calculator #(.RECT1_X(rectangle1_xs[296]), .RECT1_Y(rectangle1_ys[296]), .RECT1_WIDTH(rectangle1_widths[296]), .RECT1_HEIGHT(rectangle1_heights[296]), .RECT1_WEIGHT(rectangle1_weights[296]), .RECT2_X(rectangle2_xs[296]), .RECT2_Y(rectangle2_ys[296]), .RECT2_WIDTH(rectangle2_widths[296]), .RECT2_HEIGHT(rectangle2_heights[296]), .RECT2_WEIGHT(rectangle2_weights[296]), .RECT3_X(rectangle3_xs[296]), .RECT3_Y(rectangle3_ys[296]), .RECT3_WIDTH(rectangle3_widths[296]), .RECT3_HEIGHT(rectangle3_heights[296]), .RECT3_WEIGHT(rectangle3_weights[296]), .FEAT_THRES(feature_thresholds[296]), .FEAT_ABOVE(feature_aboves[296]), .FEAT_BELOW(feature_belows[296])) ac296(.scan_win(scan_win296), .scan_win_std_dev(scan_win_std_dev[296]), .feature_accum(feature_accums[296]));
  accum_calculator #(.RECT1_X(rectangle1_xs[297]), .RECT1_Y(rectangle1_ys[297]), .RECT1_WIDTH(rectangle1_widths[297]), .RECT1_HEIGHT(rectangle1_heights[297]), .RECT1_WEIGHT(rectangle1_weights[297]), .RECT2_X(rectangle2_xs[297]), .RECT2_Y(rectangle2_ys[297]), .RECT2_WIDTH(rectangle2_widths[297]), .RECT2_HEIGHT(rectangle2_heights[297]), .RECT2_WEIGHT(rectangle2_weights[297]), .RECT3_X(rectangle3_xs[297]), .RECT3_Y(rectangle3_ys[297]), .RECT3_WIDTH(rectangle3_widths[297]), .RECT3_HEIGHT(rectangle3_heights[297]), .RECT3_WEIGHT(rectangle3_weights[297]), .FEAT_THRES(feature_thresholds[297]), .FEAT_ABOVE(feature_aboves[297]), .FEAT_BELOW(feature_belows[297])) ac297(.scan_win(scan_win297), .scan_win_std_dev(scan_win_std_dev[297]), .feature_accum(feature_accums[297]));
  accum_calculator #(.RECT1_X(rectangle1_xs[298]), .RECT1_Y(rectangle1_ys[298]), .RECT1_WIDTH(rectangle1_widths[298]), .RECT1_HEIGHT(rectangle1_heights[298]), .RECT1_WEIGHT(rectangle1_weights[298]), .RECT2_X(rectangle2_xs[298]), .RECT2_Y(rectangle2_ys[298]), .RECT2_WIDTH(rectangle2_widths[298]), .RECT2_HEIGHT(rectangle2_heights[298]), .RECT2_WEIGHT(rectangle2_weights[298]), .RECT3_X(rectangle3_xs[298]), .RECT3_Y(rectangle3_ys[298]), .RECT3_WIDTH(rectangle3_widths[298]), .RECT3_HEIGHT(rectangle3_heights[298]), .RECT3_WEIGHT(rectangle3_weights[298]), .FEAT_THRES(feature_thresholds[298]), .FEAT_ABOVE(feature_aboves[298]), .FEAT_BELOW(feature_belows[298])) ac298(.scan_win(scan_win298), .scan_win_std_dev(scan_win_std_dev[298]), .feature_accum(feature_accums[298]));
  accum_calculator #(.RECT1_X(rectangle1_xs[299]), .RECT1_Y(rectangle1_ys[299]), .RECT1_WIDTH(rectangle1_widths[299]), .RECT1_HEIGHT(rectangle1_heights[299]), .RECT1_WEIGHT(rectangle1_weights[299]), .RECT2_X(rectangle2_xs[299]), .RECT2_Y(rectangle2_ys[299]), .RECT2_WIDTH(rectangle2_widths[299]), .RECT2_HEIGHT(rectangle2_heights[299]), .RECT2_WEIGHT(rectangle2_weights[299]), .RECT3_X(rectangle3_xs[299]), .RECT3_Y(rectangle3_ys[299]), .RECT3_WIDTH(rectangle3_widths[299]), .RECT3_HEIGHT(rectangle3_heights[299]), .RECT3_WEIGHT(rectangle3_weights[299]), .FEAT_THRES(feature_thresholds[299]), .FEAT_ABOVE(feature_aboves[299]), .FEAT_BELOW(feature_belows[299])) ac299(.scan_win(scan_win299), .scan_win_std_dev(scan_win_std_dev[299]), .feature_accum(feature_accums[299]));
  accum_calculator #(.RECT1_X(rectangle1_xs[300]), .RECT1_Y(rectangle1_ys[300]), .RECT1_WIDTH(rectangle1_widths[300]), .RECT1_HEIGHT(rectangle1_heights[300]), .RECT1_WEIGHT(rectangle1_weights[300]), .RECT2_X(rectangle2_xs[300]), .RECT2_Y(rectangle2_ys[300]), .RECT2_WIDTH(rectangle2_widths[300]), .RECT2_HEIGHT(rectangle2_heights[300]), .RECT2_WEIGHT(rectangle2_weights[300]), .RECT3_X(rectangle3_xs[300]), .RECT3_Y(rectangle3_ys[300]), .RECT3_WIDTH(rectangle3_widths[300]), .RECT3_HEIGHT(rectangle3_heights[300]), .RECT3_WEIGHT(rectangle3_weights[300]), .FEAT_THRES(feature_thresholds[300]), .FEAT_ABOVE(feature_aboves[300]), .FEAT_BELOW(feature_belows[300])) ac300(.scan_win(scan_win300), .scan_win_std_dev(scan_win_std_dev[300]), .feature_accum(feature_accums[300]));
  accum_calculator #(.RECT1_X(rectangle1_xs[301]), .RECT1_Y(rectangle1_ys[301]), .RECT1_WIDTH(rectangle1_widths[301]), .RECT1_HEIGHT(rectangle1_heights[301]), .RECT1_WEIGHT(rectangle1_weights[301]), .RECT2_X(rectangle2_xs[301]), .RECT2_Y(rectangle2_ys[301]), .RECT2_WIDTH(rectangle2_widths[301]), .RECT2_HEIGHT(rectangle2_heights[301]), .RECT2_WEIGHT(rectangle2_weights[301]), .RECT3_X(rectangle3_xs[301]), .RECT3_Y(rectangle3_ys[301]), .RECT3_WIDTH(rectangle3_widths[301]), .RECT3_HEIGHT(rectangle3_heights[301]), .RECT3_WEIGHT(rectangle3_weights[301]), .FEAT_THRES(feature_thresholds[301]), .FEAT_ABOVE(feature_aboves[301]), .FEAT_BELOW(feature_belows[301])) ac301(.scan_win(scan_win301), .scan_win_std_dev(scan_win_std_dev[301]), .feature_accum(feature_accums[301]));
  accum_calculator #(.RECT1_X(rectangle1_xs[302]), .RECT1_Y(rectangle1_ys[302]), .RECT1_WIDTH(rectangle1_widths[302]), .RECT1_HEIGHT(rectangle1_heights[302]), .RECT1_WEIGHT(rectangle1_weights[302]), .RECT2_X(rectangle2_xs[302]), .RECT2_Y(rectangle2_ys[302]), .RECT2_WIDTH(rectangle2_widths[302]), .RECT2_HEIGHT(rectangle2_heights[302]), .RECT2_WEIGHT(rectangle2_weights[302]), .RECT3_X(rectangle3_xs[302]), .RECT3_Y(rectangle3_ys[302]), .RECT3_WIDTH(rectangle3_widths[302]), .RECT3_HEIGHT(rectangle3_heights[302]), .RECT3_WEIGHT(rectangle3_weights[302]), .FEAT_THRES(feature_thresholds[302]), .FEAT_ABOVE(feature_aboves[302]), .FEAT_BELOW(feature_belows[302])) ac302(.scan_win(scan_win302), .scan_win_std_dev(scan_win_std_dev[302]), .feature_accum(feature_accums[302]));
  accum_calculator #(.RECT1_X(rectangle1_xs[303]), .RECT1_Y(rectangle1_ys[303]), .RECT1_WIDTH(rectangle1_widths[303]), .RECT1_HEIGHT(rectangle1_heights[303]), .RECT1_WEIGHT(rectangle1_weights[303]), .RECT2_X(rectangle2_xs[303]), .RECT2_Y(rectangle2_ys[303]), .RECT2_WIDTH(rectangle2_widths[303]), .RECT2_HEIGHT(rectangle2_heights[303]), .RECT2_WEIGHT(rectangle2_weights[303]), .RECT3_X(rectangle3_xs[303]), .RECT3_Y(rectangle3_ys[303]), .RECT3_WIDTH(rectangle3_widths[303]), .RECT3_HEIGHT(rectangle3_heights[303]), .RECT3_WEIGHT(rectangle3_weights[303]), .FEAT_THRES(feature_thresholds[303]), .FEAT_ABOVE(feature_aboves[303]), .FEAT_BELOW(feature_belows[303])) ac303(.scan_win(scan_win303), .scan_win_std_dev(scan_win_std_dev[303]), .feature_accum(feature_accums[303]));
  accum_calculator #(.RECT1_X(rectangle1_xs[304]), .RECT1_Y(rectangle1_ys[304]), .RECT1_WIDTH(rectangle1_widths[304]), .RECT1_HEIGHT(rectangle1_heights[304]), .RECT1_WEIGHT(rectangle1_weights[304]), .RECT2_X(rectangle2_xs[304]), .RECT2_Y(rectangle2_ys[304]), .RECT2_WIDTH(rectangle2_widths[304]), .RECT2_HEIGHT(rectangle2_heights[304]), .RECT2_WEIGHT(rectangle2_weights[304]), .RECT3_X(rectangle3_xs[304]), .RECT3_Y(rectangle3_ys[304]), .RECT3_WIDTH(rectangle3_widths[304]), .RECT3_HEIGHT(rectangle3_heights[304]), .RECT3_WEIGHT(rectangle3_weights[304]), .FEAT_THRES(feature_thresholds[304]), .FEAT_ABOVE(feature_aboves[304]), .FEAT_BELOW(feature_belows[304])) ac304(.scan_win(scan_win304), .scan_win_std_dev(scan_win_std_dev[304]), .feature_accum(feature_accums[304]));
  accum_calculator #(.RECT1_X(rectangle1_xs[305]), .RECT1_Y(rectangle1_ys[305]), .RECT1_WIDTH(rectangle1_widths[305]), .RECT1_HEIGHT(rectangle1_heights[305]), .RECT1_WEIGHT(rectangle1_weights[305]), .RECT2_X(rectangle2_xs[305]), .RECT2_Y(rectangle2_ys[305]), .RECT2_WIDTH(rectangle2_widths[305]), .RECT2_HEIGHT(rectangle2_heights[305]), .RECT2_WEIGHT(rectangle2_weights[305]), .RECT3_X(rectangle3_xs[305]), .RECT3_Y(rectangle3_ys[305]), .RECT3_WIDTH(rectangle3_widths[305]), .RECT3_HEIGHT(rectangle3_heights[305]), .RECT3_WEIGHT(rectangle3_weights[305]), .FEAT_THRES(feature_thresholds[305]), .FEAT_ABOVE(feature_aboves[305]), .FEAT_BELOW(feature_belows[305])) ac305(.scan_win(scan_win305), .scan_win_std_dev(scan_win_std_dev[305]), .feature_accum(feature_accums[305]));
  accum_calculator #(.RECT1_X(rectangle1_xs[306]), .RECT1_Y(rectangle1_ys[306]), .RECT1_WIDTH(rectangle1_widths[306]), .RECT1_HEIGHT(rectangle1_heights[306]), .RECT1_WEIGHT(rectangle1_weights[306]), .RECT2_X(rectangle2_xs[306]), .RECT2_Y(rectangle2_ys[306]), .RECT2_WIDTH(rectangle2_widths[306]), .RECT2_HEIGHT(rectangle2_heights[306]), .RECT2_WEIGHT(rectangle2_weights[306]), .RECT3_X(rectangle3_xs[306]), .RECT3_Y(rectangle3_ys[306]), .RECT3_WIDTH(rectangle3_widths[306]), .RECT3_HEIGHT(rectangle3_heights[306]), .RECT3_WEIGHT(rectangle3_weights[306]), .FEAT_THRES(feature_thresholds[306]), .FEAT_ABOVE(feature_aboves[306]), .FEAT_BELOW(feature_belows[306])) ac306(.scan_win(scan_win306), .scan_win_std_dev(scan_win_std_dev[306]), .feature_accum(feature_accums[306]));
  accum_calculator #(.RECT1_X(rectangle1_xs[307]), .RECT1_Y(rectangle1_ys[307]), .RECT1_WIDTH(rectangle1_widths[307]), .RECT1_HEIGHT(rectangle1_heights[307]), .RECT1_WEIGHT(rectangle1_weights[307]), .RECT2_X(rectangle2_xs[307]), .RECT2_Y(rectangle2_ys[307]), .RECT2_WIDTH(rectangle2_widths[307]), .RECT2_HEIGHT(rectangle2_heights[307]), .RECT2_WEIGHT(rectangle2_weights[307]), .RECT3_X(rectangle3_xs[307]), .RECT3_Y(rectangle3_ys[307]), .RECT3_WIDTH(rectangle3_widths[307]), .RECT3_HEIGHT(rectangle3_heights[307]), .RECT3_WEIGHT(rectangle3_weights[307]), .FEAT_THRES(feature_thresholds[307]), .FEAT_ABOVE(feature_aboves[307]), .FEAT_BELOW(feature_belows[307])) ac307(.scan_win(scan_win307), .scan_win_std_dev(scan_win_std_dev[307]), .feature_accum(feature_accums[307]));
  accum_calculator #(.RECT1_X(rectangle1_xs[308]), .RECT1_Y(rectangle1_ys[308]), .RECT1_WIDTH(rectangle1_widths[308]), .RECT1_HEIGHT(rectangle1_heights[308]), .RECT1_WEIGHT(rectangle1_weights[308]), .RECT2_X(rectangle2_xs[308]), .RECT2_Y(rectangle2_ys[308]), .RECT2_WIDTH(rectangle2_widths[308]), .RECT2_HEIGHT(rectangle2_heights[308]), .RECT2_WEIGHT(rectangle2_weights[308]), .RECT3_X(rectangle3_xs[308]), .RECT3_Y(rectangle3_ys[308]), .RECT3_WIDTH(rectangle3_widths[308]), .RECT3_HEIGHT(rectangle3_heights[308]), .RECT3_WEIGHT(rectangle3_weights[308]), .FEAT_THRES(feature_thresholds[308]), .FEAT_ABOVE(feature_aboves[308]), .FEAT_BELOW(feature_belows[308])) ac308(.scan_win(scan_win308), .scan_win_std_dev(scan_win_std_dev[308]), .feature_accum(feature_accums[308]));
  accum_calculator #(.RECT1_X(rectangle1_xs[309]), .RECT1_Y(rectangle1_ys[309]), .RECT1_WIDTH(rectangle1_widths[309]), .RECT1_HEIGHT(rectangle1_heights[309]), .RECT1_WEIGHT(rectangle1_weights[309]), .RECT2_X(rectangle2_xs[309]), .RECT2_Y(rectangle2_ys[309]), .RECT2_WIDTH(rectangle2_widths[309]), .RECT2_HEIGHT(rectangle2_heights[309]), .RECT2_WEIGHT(rectangle2_weights[309]), .RECT3_X(rectangle3_xs[309]), .RECT3_Y(rectangle3_ys[309]), .RECT3_WIDTH(rectangle3_widths[309]), .RECT3_HEIGHT(rectangle3_heights[309]), .RECT3_WEIGHT(rectangle3_weights[309]), .FEAT_THRES(feature_thresholds[309]), .FEAT_ABOVE(feature_aboves[309]), .FEAT_BELOW(feature_belows[309])) ac309(.scan_win(scan_win309), .scan_win_std_dev(scan_win_std_dev[309]), .feature_accum(feature_accums[309]));
  accum_calculator #(.RECT1_X(rectangle1_xs[310]), .RECT1_Y(rectangle1_ys[310]), .RECT1_WIDTH(rectangle1_widths[310]), .RECT1_HEIGHT(rectangle1_heights[310]), .RECT1_WEIGHT(rectangle1_weights[310]), .RECT2_X(rectangle2_xs[310]), .RECT2_Y(rectangle2_ys[310]), .RECT2_WIDTH(rectangle2_widths[310]), .RECT2_HEIGHT(rectangle2_heights[310]), .RECT2_WEIGHT(rectangle2_weights[310]), .RECT3_X(rectangle3_xs[310]), .RECT3_Y(rectangle3_ys[310]), .RECT3_WIDTH(rectangle3_widths[310]), .RECT3_HEIGHT(rectangle3_heights[310]), .RECT3_WEIGHT(rectangle3_weights[310]), .FEAT_THRES(feature_thresholds[310]), .FEAT_ABOVE(feature_aboves[310]), .FEAT_BELOW(feature_belows[310])) ac310(.scan_win(scan_win310), .scan_win_std_dev(scan_win_std_dev[310]), .feature_accum(feature_accums[310]));
  accum_calculator #(.RECT1_X(rectangle1_xs[311]), .RECT1_Y(rectangle1_ys[311]), .RECT1_WIDTH(rectangle1_widths[311]), .RECT1_HEIGHT(rectangle1_heights[311]), .RECT1_WEIGHT(rectangle1_weights[311]), .RECT2_X(rectangle2_xs[311]), .RECT2_Y(rectangle2_ys[311]), .RECT2_WIDTH(rectangle2_widths[311]), .RECT2_HEIGHT(rectangle2_heights[311]), .RECT2_WEIGHT(rectangle2_weights[311]), .RECT3_X(rectangle3_xs[311]), .RECT3_Y(rectangle3_ys[311]), .RECT3_WIDTH(rectangle3_widths[311]), .RECT3_HEIGHT(rectangle3_heights[311]), .RECT3_WEIGHT(rectangle3_weights[311]), .FEAT_THRES(feature_thresholds[311]), .FEAT_ABOVE(feature_aboves[311]), .FEAT_BELOW(feature_belows[311])) ac311(.scan_win(scan_win311), .scan_win_std_dev(scan_win_std_dev[311]), .feature_accum(feature_accums[311]));
  accum_calculator #(.RECT1_X(rectangle1_xs[312]), .RECT1_Y(rectangle1_ys[312]), .RECT1_WIDTH(rectangle1_widths[312]), .RECT1_HEIGHT(rectangle1_heights[312]), .RECT1_WEIGHT(rectangle1_weights[312]), .RECT2_X(rectangle2_xs[312]), .RECT2_Y(rectangle2_ys[312]), .RECT2_WIDTH(rectangle2_widths[312]), .RECT2_HEIGHT(rectangle2_heights[312]), .RECT2_WEIGHT(rectangle2_weights[312]), .RECT3_X(rectangle3_xs[312]), .RECT3_Y(rectangle3_ys[312]), .RECT3_WIDTH(rectangle3_widths[312]), .RECT3_HEIGHT(rectangle3_heights[312]), .RECT3_WEIGHT(rectangle3_weights[312]), .FEAT_THRES(feature_thresholds[312]), .FEAT_ABOVE(feature_aboves[312]), .FEAT_BELOW(feature_belows[312])) ac312(.scan_win(scan_win312), .scan_win_std_dev(scan_win_std_dev[312]), .feature_accum(feature_accums[312]));
  accum_calculator #(.RECT1_X(rectangle1_xs[313]), .RECT1_Y(rectangle1_ys[313]), .RECT1_WIDTH(rectangle1_widths[313]), .RECT1_HEIGHT(rectangle1_heights[313]), .RECT1_WEIGHT(rectangle1_weights[313]), .RECT2_X(rectangle2_xs[313]), .RECT2_Y(rectangle2_ys[313]), .RECT2_WIDTH(rectangle2_widths[313]), .RECT2_HEIGHT(rectangle2_heights[313]), .RECT2_WEIGHT(rectangle2_weights[313]), .RECT3_X(rectangle3_xs[313]), .RECT3_Y(rectangle3_ys[313]), .RECT3_WIDTH(rectangle3_widths[313]), .RECT3_HEIGHT(rectangle3_heights[313]), .RECT3_WEIGHT(rectangle3_weights[313]), .FEAT_THRES(feature_thresholds[313]), .FEAT_ABOVE(feature_aboves[313]), .FEAT_BELOW(feature_belows[313])) ac313(.scan_win(scan_win313), .scan_win_std_dev(scan_win_std_dev[313]), .feature_accum(feature_accums[313]));
  accum_calculator #(.RECT1_X(rectangle1_xs[314]), .RECT1_Y(rectangle1_ys[314]), .RECT1_WIDTH(rectangle1_widths[314]), .RECT1_HEIGHT(rectangle1_heights[314]), .RECT1_WEIGHT(rectangle1_weights[314]), .RECT2_X(rectangle2_xs[314]), .RECT2_Y(rectangle2_ys[314]), .RECT2_WIDTH(rectangle2_widths[314]), .RECT2_HEIGHT(rectangle2_heights[314]), .RECT2_WEIGHT(rectangle2_weights[314]), .RECT3_X(rectangle3_xs[314]), .RECT3_Y(rectangle3_ys[314]), .RECT3_WIDTH(rectangle3_widths[314]), .RECT3_HEIGHT(rectangle3_heights[314]), .RECT3_WEIGHT(rectangle3_weights[314]), .FEAT_THRES(feature_thresholds[314]), .FEAT_ABOVE(feature_aboves[314]), .FEAT_BELOW(feature_belows[314])) ac314(.scan_win(scan_win314), .scan_win_std_dev(scan_win_std_dev[314]), .feature_accum(feature_accums[314]));
  accum_calculator #(.RECT1_X(rectangle1_xs[315]), .RECT1_Y(rectangle1_ys[315]), .RECT1_WIDTH(rectangle1_widths[315]), .RECT1_HEIGHT(rectangle1_heights[315]), .RECT1_WEIGHT(rectangle1_weights[315]), .RECT2_X(rectangle2_xs[315]), .RECT2_Y(rectangle2_ys[315]), .RECT2_WIDTH(rectangle2_widths[315]), .RECT2_HEIGHT(rectangle2_heights[315]), .RECT2_WEIGHT(rectangle2_weights[315]), .RECT3_X(rectangle3_xs[315]), .RECT3_Y(rectangle3_ys[315]), .RECT3_WIDTH(rectangle3_widths[315]), .RECT3_HEIGHT(rectangle3_heights[315]), .RECT3_WEIGHT(rectangle3_weights[315]), .FEAT_THRES(feature_thresholds[315]), .FEAT_ABOVE(feature_aboves[315]), .FEAT_BELOW(feature_belows[315])) ac315(.scan_win(scan_win315), .scan_win_std_dev(scan_win_std_dev[315]), .feature_accum(feature_accums[315]));
  accum_calculator #(.RECT1_X(rectangle1_xs[316]), .RECT1_Y(rectangle1_ys[316]), .RECT1_WIDTH(rectangle1_widths[316]), .RECT1_HEIGHT(rectangle1_heights[316]), .RECT1_WEIGHT(rectangle1_weights[316]), .RECT2_X(rectangle2_xs[316]), .RECT2_Y(rectangle2_ys[316]), .RECT2_WIDTH(rectangle2_widths[316]), .RECT2_HEIGHT(rectangle2_heights[316]), .RECT2_WEIGHT(rectangle2_weights[316]), .RECT3_X(rectangle3_xs[316]), .RECT3_Y(rectangle3_ys[316]), .RECT3_WIDTH(rectangle3_widths[316]), .RECT3_HEIGHT(rectangle3_heights[316]), .RECT3_WEIGHT(rectangle3_weights[316]), .FEAT_THRES(feature_thresholds[316]), .FEAT_ABOVE(feature_aboves[316]), .FEAT_BELOW(feature_belows[316])) ac316(.scan_win(scan_win316), .scan_win_std_dev(scan_win_std_dev[316]), .feature_accum(feature_accums[316]));
  accum_calculator #(.RECT1_X(rectangle1_xs[317]), .RECT1_Y(rectangle1_ys[317]), .RECT1_WIDTH(rectangle1_widths[317]), .RECT1_HEIGHT(rectangle1_heights[317]), .RECT1_WEIGHT(rectangle1_weights[317]), .RECT2_X(rectangle2_xs[317]), .RECT2_Y(rectangle2_ys[317]), .RECT2_WIDTH(rectangle2_widths[317]), .RECT2_HEIGHT(rectangle2_heights[317]), .RECT2_WEIGHT(rectangle2_weights[317]), .RECT3_X(rectangle3_xs[317]), .RECT3_Y(rectangle3_ys[317]), .RECT3_WIDTH(rectangle3_widths[317]), .RECT3_HEIGHT(rectangle3_heights[317]), .RECT3_WEIGHT(rectangle3_weights[317]), .FEAT_THRES(feature_thresholds[317]), .FEAT_ABOVE(feature_aboves[317]), .FEAT_BELOW(feature_belows[317])) ac317(.scan_win(scan_win317), .scan_win_std_dev(scan_win_std_dev[317]), .feature_accum(feature_accums[317]));
  accum_calculator #(.RECT1_X(rectangle1_xs[318]), .RECT1_Y(rectangle1_ys[318]), .RECT1_WIDTH(rectangle1_widths[318]), .RECT1_HEIGHT(rectangle1_heights[318]), .RECT1_WEIGHT(rectangle1_weights[318]), .RECT2_X(rectangle2_xs[318]), .RECT2_Y(rectangle2_ys[318]), .RECT2_WIDTH(rectangle2_widths[318]), .RECT2_HEIGHT(rectangle2_heights[318]), .RECT2_WEIGHT(rectangle2_weights[318]), .RECT3_X(rectangle3_xs[318]), .RECT3_Y(rectangle3_ys[318]), .RECT3_WIDTH(rectangle3_widths[318]), .RECT3_HEIGHT(rectangle3_heights[318]), .RECT3_WEIGHT(rectangle3_weights[318]), .FEAT_THRES(feature_thresholds[318]), .FEAT_ABOVE(feature_aboves[318]), .FEAT_BELOW(feature_belows[318])) ac318(.scan_win(scan_win318), .scan_win_std_dev(scan_win_std_dev[318]), .feature_accum(feature_accums[318]));
  accum_calculator #(.RECT1_X(rectangle1_xs[319]), .RECT1_Y(rectangle1_ys[319]), .RECT1_WIDTH(rectangle1_widths[319]), .RECT1_HEIGHT(rectangle1_heights[319]), .RECT1_WEIGHT(rectangle1_weights[319]), .RECT2_X(rectangle2_xs[319]), .RECT2_Y(rectangle2_ys[319]), .RECT2_WIDTH(rectangle2_widths[319]), .RECT2_HEIGHT(rectangle2_heights[319]), .RECT2_WEIGHT(rectangle2_weights[319]), .RECT3_X(rectangle3_xs[319]), .RECT3_Y(rectangle3_ys[319]), .RECT3_WIDTH(rectangle3_widths[319]), .RECT3_HEIGHT(rectangle3_heights[319]), .RECT3_WEIGHT(rectangle3_weights[319]), .FEAT_THRES(feature_thresholds[319]), .FEAT_ABOVE(feature_aboves[319]), .FEAT_BELOW(feature_belows[319])) ac319(.scan_win(scan_win319), .scan_win_std_dev(scan_win_std_dev[319]), .feature_accum(feature_accums[319]));
  accum_calculator #(.RECT1_X(rectangle1_xs[320]), .RECT1_Y(rectangle1_ys[320]), .RECT1_WIDTH(rectangle1_widths[320]), .RECT1_HEIGHT(rectangle1_heights[320]), .RECT1_WEIGHT(rectangle1_weights[320]), .RECT2_X(rectangle2_xs[320]), .RECT2_Y(rectangle2_ys[320]), .RECT2_WIDTH(rectangle2_widths[320]), .RECT2_HEIGHT(rectangle2_heights[320]), .RECT2_WEIGHT(rectangle2_weights[320]), .RECT3_X(rectangle3_xs[320]), .RECT3_Y(rectangle3_ys[320]), .RECT3_WIDTH(rectangle3_widths[320]), .RECT3_HEIGHT(rectangle3_heights[320]), .RECT3_WEIGHT(rectangle3_weights[320]), .FEAT_THRES(feature_thresholds[320]), .FEAT_ABOVE(feature_aboves[320]), .FEAT_BELOW(feature_belows[320])) ac320(.scan_win(scan_win320), .scan_win_std_dev(scan_win_std_dev[320]), .feature_accum(feature_accums[320]));
  accum_calculator #(.RECT1_X(rectangle1_xs[321]), .RECT1_Y(rectangle1_ys[321]), .RECT1_WIDTH(rectangle1_widths[321]), .RECT1_HEIGHT(rectangle1_heights[321]), .RECT1_WEIGHT(rectangle1_weights[321]), .RECT2_X(rectangle2_xs[321]), .RECT2_Y(rectangle2_ys[321]), .RECT2_WIDTH(rectangle2_widths[321]), .RECT2_HEIGHT(rectangle2_heights[321]), .RECT2_WEIGHT(rectangle2_weights[321]), .RECT3_X(rectangle3_xs[321]), .RECT3_Y(rectangle3_ys[321]), .RECT3_WIDTH(rectangle3_widths[321]), .RECT3_HEIGHT(rectangle3_heights[321]), .RECT3_WEIGHT(rectangle3_weights[321]), .FEAT_THRES(feature_thresholds[321]), .FEAT_ABOVE(feature_aboves[321]), .FEAT_BELOW(feature_belows[321])) ac321(.scan_win(scan_win321), .scan_win_std_dev(scan_win_std_dev[321]), .feature_accum(feature_accums[321]));
  accum_calculator #(.RECT1_X(rectangle1_xs[322]), .RECT1_Y(rectangle1_ys[322]), .RECT1_WIDTH(rectangle1_widths[322]), .RECT1_HEIGHT(rectangle1_heights[322]), .RECT1_WEIGHT(rectangle1_weights[322]), .RECT2_X(rectangle2_xs[322]), .RECT2_Y(rectangle2_ys[322]), .RECT2_WIDTH(rectangle2_widths[322]), .RECT2_HEIGHT(rectangle2_heights[322]), .RECT2_WEIGHT(rectangle2_weights[322]), .RECT3_X(rectangle3_xs[322]), .RECT3_Y(rectangle3_ys[322]), .RECT3_WIDTH(rectangle3_widths[322]), .RECT3_HEIGHT(rectangle3_heights[322]), .RECT3_WEIGHT(rectangle3_weights[322]), .FEAT_THRES(feature_thresholds[322]), .FEAT_ABOVE(feature_aboves[322]), .FEAT_BELOW(feature_belows[322])) ac322(.scan_win(scan_win322), .scan_win_std_dev(scan_win_std_dev[322]), .feature_accum(feature_accums[322]));
  accum_calculator #(.RECT1_X(rectangle1_xs[323]), .RECT1_Y(rectangle1_ys[323]), .RECT1_WIDTH(rectangle1_widths[323]), .RECT1_HEIGHT(rectangle1_heights[323]), .RECT1_WEIGHT(rectangle1_weights[323]), .RECT2_X(rectangle2_xs[323]), .RECT2_Y(rectangle2_ys[323]), .RECT2_WIDTH(rectangle2_widths[323]), .RECT2_HEIGHT(rectangle2_heights[323]), .RECT2_WEIGHT(rectangle2_weights[323]), .RECT3_X(rectangle3_xs[323]), .RECT3_Y(rectangle3_ys[323]), .RECT3_WIDTH(rectangle3_widths[323]), .RECT3_HEIGHT(rectangle3_heights[323]), .RECT3_WEIGHT(rectangle3_weights[323]), .FEAT_THRES(feature_thresholds[323]), .FEAT_ABOVE(feature_aboves[323]), .FEAT_BELOW(feature_belows[323])) ac323(.scan_win(scan_win323), .scan_win_std_dev(scan_win_std_dev[323]), .feature_accum(feature_accums[323]));
  accum_calculator #(.RECT1_X(rectangle1_xs[324]), .RECT1_Y(rectangle1_ys[324]), .RECT1_WIDTH(rectangle1_widths[324]), .RECT1_HEIGHT(rectangle1_heights[324]), .RECT1_WEIGHT(rectangle1_weights[324]), .RECT2_X(rectangle2_xs[324]), .RECT2_Y(rectangle2_ys[324]), .RECT2_WIDTH(rectangle2_widths[324]), .RECT2_HEIGHT(rectangle2_heights[324]), .RECT2_WEIGHT(rectangle2_weights[324]), .RECT3_X(rectangle3_xs[324]), .RECT3_Y(rectangle3_ys[324]), .RECT3_WIDTH(rectangle3_widths[324]), .RECT3_HEIGHT(rectangle3_heights[324]), .RECT3_WEIGHT(rectangle3_weights[324]), .FEAT_THRES(feature_thresholds[324]), .FEAT_ABOVE(feature_aboves[324]), .FEAT_BELOW(feature_belows[324])) ac324(.scan_win(scan_win324), .scan_win_std_dev(scan_win_std_dev[324]), .feature_accum(feature_accums[324]));
  accum_calculator #(.RECT1_X(rectangle1_xs[325]), .RECT1_Y(rectangle1_ys[325]), .RECT1_WIDTH(rectangle1_widths[325]), .RECT1_HEIGHT(rectangle1_heights[325]), .RECT1_WEIGHT(rectangle1_weights[325]), .RECT2_X(rectangle2_xs[325]), .RECT2_Y(rectangle2_ys[325]), .RECT2_WIDTH(rectangle2_widths[325]), .RECT2_HEIGHT(rectangle2_heights[325]), .RECT2_WEIGHT(rectangle2_weights[325]), .RECT3_X(rectangle3_xs[325]), .RECT3_Y(rectangle3_ys[325]), .RECT3_WIDTH(rectangle3_widths[325]), .RECT3_HEIGHT(rectangle3_heights[325]), .RECT3_WEIGHT(rectangle3_weights[325]), .FEAT_THRES(feature_thresholds[325]), .FEAT_ABOVE(feature_aboves[325]), .FEAT_BELOW(feature_belows[325])) ac325(.scan_win(scan_win325), .scan_win_std_dev(scan_win_std_dev[325]), .feature_accum(feature_accums[325]));
  accum_calculator #(.RECT1_X(rectangle1_xs[326]), .RECT1_Y(rectangle1_ys[326]), .RECT1_WIDTH(rectangle1_widths[326]), .RECT1_HEIGHT(rectangle1_heights[326]), .RECT1_WEIGHT(rectangle1_weights[326]), .RECT2_X(rectangle2_xs[326]), .RECT2_Y(rectangle2_ys[326]), .RECT2_WIDTH(rectangle2_widths[326]), .RECT2_HEIGHT(rectangle2_heights[326]), .RECT2_WEIGHT(rectangle2_weights[326]), .RECT3_X(rectangle3_xs[326]), .RECT3_Y(rectangle3_ys[326]), .RECT3_WIDTH(rectangle3_widths[326]), .RECT3_HEIGHT(rectangle3_heights[326]), .RECT3_WEIGHT(rectangle3_weights[326]), .FEAT_THRES(feature_thresholds[326]), .FEAT_ABOVE(feature_aboves[326]), .FEAT_BELOW(feature_belows[326])) ac326(.scan_win(scan_win326), .scan_win_std_dev(scan_win_std_dev[326]), .feature_accum(feature_accums[326]));
  accum_calculator #(.RECT1_X(rectangle1_xs[327]), .RECT1_Y(rectangle1_ys[327]), .RECT1_WIDTH(rectangle1_widths[327]), .RECT1_HEIGHT(rectangle1_heights[327]), .RECT1_WEIGHT(rectangle1_weights[327]), .RECT2_X(rectangle2_xs[327]), .RECT2_Y(rectangle2_ys[327]), .RECT2_WIDTH(rectangle2_widths[327]), .RECT2_HEIGHT(rectangle2_heights[327]), .RECT2_WEIGHT(rectangle2_weights[327]), .RECT3_X(rectangle3_xs[327]), .RECT3_Y(rectangle3_ys[327]), .RECT3_WIDTH(rectangle3_widths[327]), .RECT3_HEIGHT(rectangle3_heights[327]), .RECT3_WEIGHT(rectangle3_weights[327]), .FEAT_THRES(feature_thresholds[327]), .FEAT_ABOVE(feature_aboves[327]), .FEAT_BELOW(feature_belows[327])) ac327(.scan_win(scan_win327), .scan_win_std_dev(scan_win_std_dev[327]), .feature_accum(feature_accums[327]));
  accum_calculator #(.RECT1_X(rectangle1_xs[328]), .RECT1_Y(rectangle1_ys[328]), .RECT1_WIDTH(rectangle1_widths[328]), .RECT1_HEIGHT(rectangle1_heights[328]), .RECT1_WEIGHT(rectangle1_weights[328]), .RECT2_X(rectangle2_xs[328]), .RECT2_Y(rectangle2_ys[328]), .RECT2_WIDTH(rectangle2_widths[328]), .RECT2_HEIGHT(rectangle2_heights[328]), .RECT2_WEIGHT(rectangle2_weights[328]), .RECT3_X(rectangle3_xs[328]), .RECT3_Y(rectangle3_ys[328]), .RECT3_WIDTH(rectangle3_widths[328]), .RECT3_HEIGHT(rectangle3_heights[328]), .RECT3_WEIGHT(rectangle3_weights[328]), .FEAT_THRES(feature_thresholds[328]), .FEAT_ABOVE(feature_aboves[328]), .FEAT_BELOW(feature_belows[328])) ac328(.scan_win(scan_win328), .scan_win_std_dev(scan_win_std_dev[328]), .feature_accum(feature_accums[328]));
  accum_calculator #(.RECT1_X(rectangle1_xs[329]), .RECT1_Y(rectangle1_ys[329]), .RECT1_WIDTH(rectangle1_widths[329]), .RECT1_HEIGHT(rectangle1_heights[329]), .RECT1_WEIGHT(rectangle1_weights[329]), .RECT2_X(rectangle2_xs[329]), .RECT2_Y(rectangle2_ys[329]), .RECT2_WIDTH(rectangle2_widths[329]), .RECT2_HEIGHT(rectangle2_heights[329]), .RECT2_WEIGHT(rectangle2_weights[329]), .RECT3_X(rectangle3_xs[329]), .RECT3_Y(rectangle3_ys[329]), .RECT3_WIDTH(rectangle3_widths[329]), .RECT3_HEIGHT(rectangle3_heights[329]), .RECT3_WEIGHT(rectangle3_weights[329]), .FEAT_THRES(feature_thresholds[329]), .FEAT_ABOVE(feature_aboves[329]), .FEAT_BELOW(feature_belows[329])) ac329(.scan_win(scan_win329), .scan_win_std_dev(scan_win_std_dev[329]), .feature_accum(feature_accums[329]));
  accum_calculator #(.RECT1_X(rectangle1_xs[330]), .RECT1_Y(rectangle1_ys[330]), .RECT1_WIDTH(rectangle1_widths[330]), .RECT1_HEIGHT(rectangle1_heights[330]), .RECT1_WEIGHT(rectangle1_weights[330]), .RECT2_X(rectangle2_xs[330]), .RECT2_Y(rectangle2_ys[330]), .RECT2_WIDTH(rectangle2_widths[330]), .RECT2_HEIGHT(rectangle2_heights[330]), .RECT2_WEIGHT(rectangle2_weights[330]), .RECT3_X(rectangle3_xs[330]), .RECT3_Y(rectangle3_ys[330]), .RECT3_WIDTH(rectangle3_widths[330]), .RECT3_HEIGHT(rectangle3_heights[330]), .RECT3_WEIGHT(rectangle3_weights[330]), .FEAT_THRES(feature_thresholds[330]), .FEAT_ABOVE(feature_aboves[330]), .FEAT_BELOW(feature_belows[330])) ac330(.scan_win(scan_win330), .scan_win_std_dev(scan_win_std_dev[330]), .feature_accum(feature_accums[330]));
  accum_calculator #(.RECT1_X(rectangle1_xs[331]), .RECT1_Y(rectangle1_ys[331]), .RECT1_WIDTH(rectangle1_widths[331]), .RECT1_HEIGHT(rectangle1_heights[331]), .RECT1_WEIGHT(rectangle1_weights[331]), .RECT2_X(rectangle2_xs[331]), .RECT2_Y(rectangle2_ys[331]), .RECT2_WIDTH(rectangle2_widths[331]), .RECT2_HEIGHT(rectangle2_heights[331]), .RECT2_WEIGHT(rectangle2_weights[331]), .RECT3_X(rectangle3_xs[331]), .RECT3_Y(rectangle3_ys[331]), .RECT3_WIDTH(rectangle3_widths[331]), .RECT3_HEIGHT(rectangle3_heights[331]), .RECT3_WEIGHT(rectangle3_weights[331]), .FEAT_THRES(feature_thresholds[331]), .FEAT_ABOVE(feature_aboves[331]), .FEAT_BELOW(feature_belows[331])) ac331(.scan_win(scan_win331), .scan_win_std_dev(scan_win_std_dev[331]), .feature_accum(feature_accums[331]));
  accum_calculator #(.RECT1_X(rectangle1_xs[332]), .RECT1_Y(rectangle1_ys[332]), .RECT1_WIDTH(rectangle1_widths[332]), .RECT1_HEIGHT(rectangle1_heights[332]), .RECT1_WEIGHT(rectangle1_weights[332]), .RECT2_X(rectangle2_xs[332]), .RECT2_Y(rectangle2_ys[332]), .RECT2_WIDTH(rectangle2_widths[332]), .RECT2_HEIGHT(rectangle2_heights[332]), .RECT2_WEIGHT(rectangle2_weights[332]), .RECT3_X(rectangle3_xs[332]), .RECT3_Y(rectangle3_ys[332]), .RECT3_WIDTH(rectangle3_widths[332]), .RECT3_HEIGHT(rectangle3_heights[332]), .RECT3_WEIGHT(rectangle3_weights[332]), .FEAT_THRES(feature_thresholds[332]), .FEAT_ABOVE(feature_aboves[332]), .FEAT_BELOW(feature_belows[332])) ac332(.scan_win(scan_win332), .scan_win_std_dev(scan_win_std_dev[332]), .feature_accum(feature_accums[332]));
  accum_calculator #(.RECT1_X(rectangle1_xs[333]), .RECT1_Y(rectangle1_ys[333]), .RECT1_WIDTH(rectangle1_widths[333]), .RECT1_HEIGHT(rectangle1_heights[333]), .RECT1_WEIGHT(rectangle1_weights[333]), .RECT2_X(rectangle2_xs[333]), .RECT2_Y(rectangle2_ys[333]), .RECT2_WIDTH(rectangle2_widths[333]), .RECT2_HEIGHT(rectangle2_heights[333]), .RECT2_WEIGHT(rectangle2_weights[333]), .RECT3_X(rectangle3_xs[333]), .RECT3_Y(rectangle3_ys[333]), .RECT3_WIDTH(rectangle3_widths[333]), .RECT3_HEIGHT(rectangle3_heights[333]), .RECT3_WEIGHT(rectangle3_weights[333]), .FEAT_THRES(feature_thresholds[333]), .FEAT_ABOVE(feature_aboves[333]), .FEAT_BELOW(feature_belows[333])) ac333(.scan_win(scan_win333), .scan_win_std_dev(scan_win_std_dev[333]), .feature_accum(feature_accums[333]));
  accum_calculator #(.RECT1_X(rectangle1_xs[334]), .RECT1_Y(rectangle1_ys[334]), .RECT1_WIDTH(rectangle1_widths[334]), .RECT1_HEIGHT(rectangle1_heights[334]), .RECT1_WEIGHT(rectangle1_weights[334]), .RECT2_X(rectangle2_xs[334]), .RECT2_Y(rectangle2_ys[334]), .RECT2_WIDTH(rectangle2_widths[334]), .RECT2_HEIGHT(rectangle2_heights[334]), .RECT2_WEIGHT(rectangle2_weights[334]), .RECT3_X(rectangle3_xs[334]), .RECT3_Y(rectangle3_ys[334]), .RECT3_WIDTH(rectangle3_widths[334]), .RECT3_HEIGHT(rectangle3_heights[334]), .RECT3_WEIGHT(rectangle3_weights[334]), .FEAT_THRES(feature_thresholds[334]), .FEAT_ABOVE(feature_aboves[334]), .FEAT_BELOW(feature_belows[334])) ac334(.scan_win(scan_win334), .scan_win_std_dev(scan_win_std_dev[334]), .feature_accum(feature_accums[334]));
  accum_calculator #(.RECT1_X(rectangle1_xs[335]), .RECT1_Y(rectangle1_ys[335]), .RECT1_WIDTH(rectangle1_widths[335]), .RECT1_HEIGHT(rectangle1_heights[335]), .RECT1_WEIGHT(rectangle1_weights[335]), .RECT2_X(rectangle2_xs[335]), .RECT2_Y(rectangle2_ys[335]), .RECT2_WIDTH(rectangle2_widths[335]), .RECT2_HEIGHT(rectangle2_heights[335]), .RECT2_WEIGHT(rectangle2_weights[335]), .RECT3_X(rectangle3_xs[335]), .RECT3_Y(rectangle3_ys[335]), .RECT3_WIDTH(rectangle3_widths[335]), .RECT3_HEIGHT(rectangle3_heights[335]), .RECT3_WEIGHT(rectangle3_weights[335]), .FEAT_THRES(feature_thresholds[335]), .FEAT_ABOVE(feature_aboves[335]), .FEAT_BELOW(feature_belows[335])) ac335(.scan_win(scan_win335), .scan_win_std_dev(scan_win_std_dev[335]), .feature_accum(feature_accums[335]));
  accum_calculator #(.RECT1_X(rectangle1_xs[336]), .RECT1_Y(rectangle1_ys[336]), .RECT1_WIDTH(rectangle1_widths[336]), .RECT1_HEIGHT(rectangle1_heights[336]), .RECT1_WEIGHT(rectangle1_weights[336]), .RECT2_X(rectangle2_xs[336]), .RECT2_Y(rectangle2_ys[336]), .RECT2_WIDTH(rectangle2_widths[336]), .RECT2_HEIGHT(rectangle2_heights[336]), .RECT2_WEIGHT(rectangle2_weights[336]), .RECT3_X(rectangle3_xs[336]), .RECT3_Y(rectangle3_ys[336]), .RECT3_WIDTH(rectangle3_widths[336]), .RECT3_HEIGHT(rectangle3_heights[336]), .RECT3_WEIGHT(rectangle3_weights[336]), .FEAT_THRES(feature_thresholds[336]), .FEAT_ABOVE(feature_aboves[336]), .FEAT_BELOW(feature_belows[336])) ac336(.scan_win(scan_win336), .scan_win_std_dev(scan_win_std_dev[336]), .feature_accum(feature_accums[336]));
  accum_calculator #(.RECT1_X(rectangle1_xs[337]), .RECT1_Y(rectangle1_ys[337]), .RECT1_WIDTH(rectangle1_widths[337]), .RECT1_HEIGHT(rectangle1_heights[337]), .RECT1_WEIGHT(rectangle1_weights[337]), .RECT2_X(rectangle2_xs[337]), .RECT2_Y(rectangle2_ys[337]), .RECT2_WIDTH(rectangle2_widths[337]), .RECT2_HEIGHT(rectangle2_heights[337]), .RECT2_WEIGHT(rectangle2_weights[337]), .RECT3_X(rectangle3_xs[337]), .RECT3_Y(rectangle3_ys[337]), .RECT3_WIDTH(rectangle3_widths[337]), .RECT3_HEIGHT(rectangle3_heights[337]), .RECT3_WEIGHT(rectangle3_weights[337]), .FEAT_THRES(feature_thresholds[337]), .FEAT_ABOVE(feature_aboves[337]), .FEAT_BELOW(feature_belows[337])) ac337(.scan_win(scan_win337), .scan_win_std_dev(scan_win_std_dev[337]), .feature_accum(feature_accums[337]));
  accum_calculator #(.RECT1_X(rectangle1_xs[338]), .RECT1_Y(rectangle1_ys[338]), .RECT1_WIDTH(rectangle1_widths[338]), .RECT1_HEIGHT(rectangle1_heights[338]), .RECT1_WEIGHT(rectangle1_weights[338]), .RECT2_X(rectangle2_xs[338]), .RECT2_Y(rectangle2_ys[338]), .RECT2_WIDTH(rectangle2_widths[338]), .RECT2_HEIGHT(rectangle2_heights[338]), .RECT2_WEIGHT(rectangle2_weights[338]), .RECT3_X(rectangle3_xs[338]), .RECT3_Y(rectangle3_ys[338]), .RECT3_WIDTH(rectangle3_widths[338]), .RECT3_HEIGHT(rectangle3_heights[338]), .RECT3_WEIGHT(rectangle3_weights[338]), .FEAT_THRES(feature_thresholds[338]), .FEAT_ABOVE(feature_aboves[338]), .FEAT_BELOW(feature_belows[338])) ac338(.scan_win(scan_win338), .scan_win_std_dev(scan_win_std_dev[338]), .feature_accum(feature_accums[338]));
  accum_calculator #(.RECT1_X(rectangle1_xs[339]), .RECT1_Y(rectangle1_ys[339]), .RECT1_WIDTH(rectangle1_widths[339]), .RECT1_HEIGHT(rectangle1_heights[339]), .RECT1_WEIGHT(rectangle1_weights[339]), .RECT2_X(rectangle2_xs[339]), .RECT2_Y(rectangle2_ys[339]), .RECT2_WIDTH(rectangle2_widths[339]), .RECT2_HEIGHT(rectangle2_heights[339]), .RECT2_WEIGHT(rectangle2_weights[339]), .RECT3_X(rectangle3_xs[339]), .RECT3_Y(rectangle3_ys[339]), .RECT3_WIDTH(rectangle3_widths[339]), .RECT3_HEIGHT(rectangle3_heights[339]), .RECT3_WEIGHT(rectangle3_weights[339]), .FEAT_THRES(feature_thresholds[339]), .FEAT_ABOVE(feature_aboves[339]), .FEAT_BELOW(feature_belows[339])) ac339(.scan_win(scan_win339), .scan_win_std_dev(scan_win_std_dev[339]), .feature_accum(feature_accums[339]));
  accum_calculator #(.RECT1_X(rectangle1_xs[340]), .RECT1_Y(rectangle1_ys[340]), .RECT1_WIDTH(rectangle1_widths[340]), .RECT1_HEIGHT(rectangle1_heights[340]), .RECT1_WEIGHT(rectangle1_weights[340]), .RECT2_X(rectangle2_xs[340]), .RECT2_Y(rectangle2_ys[340]), .RECT2_WIDTH(rectangle2_widths[340]), .RECT2_HEIGHT(rectangle2_heights[340]), .RECT2_WEIGHT(rectangle2_weights[340]), .RECT3_X(rectangle3_xs[340]), .RECT3_Y(rectangle3_ys[340]), .RECT3_WIDTH(rectangle3_widths[340]), .RECT3_HEIGHT(rectangle3_heights[340]), .RECT3_WEIGHT(rectangle3_weights[340]), .FEAT_THRES(feature_thresholds[340]), .FEAT_ABOVE(feature_aboves[340]), .FEAT_BELOW(feature_belows[340])) ac340(.scan_win(scan_win340), .scan_win_std_dev(scan_win_std_dev[340]), .feature_accum(feature_accums[340]));
  accum_calculator #(.RECT1_X(rectangle1_xs[341]), .RECT1_Y(rectangle1_ys[341]), .RECT1_WIDTH(rectangle1_widths[341]), .RECT1_HEIGHT(rectangle1_heights[341]), .RECT1_WEIGHT(rectangle1_weights[341]), .RECT2_X(rectangle2_xs[341]), .RECT2_Y(rectangle2_ys[341]), .RECT2_WIDTH(rectangle2_widths[341]), .RECT2_HEIGHT(rectangle2_heights[341]), .RECT2_WEIGHT(rectangle2_weights[341]), .RECT3_X(rectangle3_xs[341]), .RECT3_Y(rectangle3_ys[341]), .RECT3_WIDTH(rectangle3_widths[341]), .RECT3_HEIGHT(rectangle3_heights[341]), .RECT3_WEIGHT(rectangle3_weights[341]), .FEAT_THRES(feature_thresholds[341]), .FEAT_ABOVE(feature_aboves[341]), .FEAT_BELOW(feature_belows[341])) ac341(.scan_win(scan_win341), .scan_win_std_dev(scan_win_std_dev[341]), .feature_accum(feature_accums[341]));
  accum_calculator #(.RECT1_X(rectangle1_xs[342]), .RECT1_Y(rectangle1_ys[342]), .RECT1_WIDTH(rectangle1_widths[342]), .RECT1_HEIGHT(rectangle1_heights[342]), .RECT1_WEIGHT(rectangle1_weights[342]), .RECT2_X(rectangle2_xs[342]), .RECT2_Y(rectangle2_ys[342]), .RECT2_WIDTH(rectangle2_widths[342]), .RECT2_HEIGHT(rectangle2_heights[342]), .RECT2_WEIGHT(rectangle2_weights[342]), .RECT3_X(rectangle3_xs[342]), .RECT3_Y(rectangle3_ys[342]), .RECT3_WIDTH(rectangle3_widths[342]), .RECT3_HEIGHT(rectangle3_heights[342]), .RECT3_WEIGHT(rectangle3_weights[342]), .FEAT_THRES(feature_thresholds[342]), .FEAT_ABOVE(feature_aboves[342]), .FEAT_BELOW(feature_belows[342])) ac342(.scan_win(scan_win342), .scan_win_std_dev(scan_win_std_dev[342]), .feature_accum(feature_accums[342]));
  accum_calculator #(.RECT1_X(rectangle1_xs[343]), .RECT1_Y(rectangle1_ys[343]), .RECT1_WIDTH(rectangle1_widths[343]), .RECT1_HEIGHT(rectangle1_heights[343]), .RECT1_WEIGHT(rectangle1_weights[343]), .RECT2_X(rectangle2_xs[343]), .RECT2_Y(rectangle2_ys[343]), .RECT2_WIDTH(rectangle2_widths[343]), .RECT2_HEIGHT(rectangle2_heights[343]), .RECT2_WEIGHT(rectangle2_weights[343]), .RECT3_X(rectangle3_xs[343]), .RECT3_Y(rectangle3_ys[343]), .RECT3_WIDTH(rectangle3_widths[343]), .RECT3_HEIGHT(rectangle3_heights[343]), .RECT3_WEIGHT(rectangle3_weights[343]), .FEAT_THRES(feature_thresholds[343]), .FEAT_ABOVE(feature_aboves[343]), .FEAT_BELOW(feature_belows[343])) ac343(.scan_win(scan_win343), .scan_win_std_dev(scan_win_std_dev[343]), .feature_accum(feature_accums[343]));
  accum_calculator #(.RECT1_X(rectangle1_xs[344]), .RECT1_Y(rectangle1_ys[344]), .RECT1_WIDTH(rectangle1_widths[344]), .RECT1_HEIGHT(rectangle1_heights[344]), .RECT1_WEIGHT(rectangle1_weights[344]), .RECT2_X(rectangle2_xs[344]), .RECT2_Y(rectangle2_ys[344]), .RECT2_WIDTH(rectangle2_widths[344]), .RECT2_HEIGHT(rectangle2_heights[344]), .RECT2_WEIGHT(rectangle2_weights[344]), .RECT3_X(rectangle3_xs[344]), .RECT3_Y(rectangle3_ys[344]), .RECT3_WIDTH(rectangle3_widths[344]), .RECT3_HEIGHT(rectangle3_heights[344]), .RECT3_WEIGHT(rectangle3_weights[344]), .FEAT_THRES(feature_thresholds[344]), .FEAT_ABOVE(feature_aboves[344]), .FEAT_BELOW(feature_belows[344])) ac344(.scan_win(scan_win344), .scan_win_std_dev(scan_win_std_dev[344]), .feature_accum(feature_accums[344]));
  accum_calculator #(.RECT1_X(rectangle1_xs[345]), .RECT1_Y(rectangle1_ys[345]), .RECT1_WIDTH(rectangle1_widths[345]), .RECT1_HEIGHT(rectangle1_heights[345]), .RECT1_WEIGHT(rectangle1_weights[345]), .RECT2_X(rectangle2_xs[345]), .RECT2_Y(rectangle2_ys[345]), .RECT2_WIDTH(rectangle2_widths[345]), .RECT2_HEIGHT(rectangle2_heights[345]), .RECT2_WEIGHT(rectangle2_weights[345]), .RECT3_X(rectangle3_xs[345]), .RECT3_Y(rectangle3_ys[345]), .RECT3_WIDTH(rectangle3_widths[345]), .RECT3_HEIGHT(rectangle3_heights[345]), .RECT3_WEIGHT(rectangle3_weights[345]), .FEAT_THRES(feature_thresholds[345]), .FEAT_ABOVE(feature_aboves[345]), .FEAT_BELOW(feature_belows[345])) ac345(.scan_win(scan_win345), .scan_win_std_dev(scan_win_std_dev[345]), .feature_accum(feature_accums[345]));
  accum_calculator #(.RECT1_X(rectangle1_xs[346]), .RECT1_Y(rectangle1_ys[346]), .RECT1_WIDTH(rectangle1_widths[346]), .RECT1_HEIGHT(rectangle1_heights[346]), .RECT1_WEIGHT(rectangle1_weights[346]), .RECT2_X(rectangle2_xs[346]), .RECT2_Y(rectangle2_ys[346]), .RECT2_WIDTH(rectangle2_widths[346]), .RECT2_HEIGHT(rectangle2_heights[346]), .RECT2_WEIGHT(rectangle2_weights[346]), .RECT3_X(rectangle3_xs[346]), .RECT3_Y(rectangle3_ys[346]), .RECT3_WIDTH(rectangle3_widths[346]), .RECT3_HEIGHT(rectangle3_heights[346]), .RECT3_WEIGHT(rectangle3_weights[346]), .FEAT_THRES(feature_thresholds[346]), .FEAT_ABOVE(feature_aboves[346]), .FEAT_BELOW(feature_belows[346])) ac346(.scan_win(scan_win346), .scan_win_std_dev(scan_win_std_dev[346]), .feature_accum(feature_accums[346]));
  accum_calculator #(.RECT1_X(rectangle1_xs[347]), .RECT1_Y(rectangle1_ys[347]), .RECT1_WIDTH(rectangle1_widths[347]), .RECT1_HEIGHT(rectangle1_heights[347]), .RECT1_WEIGHT(rectangle1_weights[347]), .RECT2_X(rectangle2_xs[347]), .RECT2_Y(rectangle2_ys[347]), .RECT2_WIDTH(rectangle2_widths[347]), .RECT2_HEIGHT(rectangle2_heights[347]), .RECT2_WEIGHT(rectangle2_weights[347]), .RECT3_X(rectangle3_xs[347]), .RECT3_Y(rectangle3_ys[347]), .RECT3_WIDTH(rectangle3_widths[347]), .RECT3_HEIGHT(rectangle3_heights[347]), .RECT3_WEIGHT(rectangle3_weights[347]), .FEAT_THRES(feature_thresholds[347]), .FEAT_ABOVE(feature_aboves[347]), .FEAT_BELOW(feature_belows[347])) ac347(.scan_win(scan_win347), .scan_win_std_dev(scan_win_std_dev[347]), .feature_accum(feature_accums[347]));
  accum_calculator #(.RECT1_X(rectangle1_xs[348]), .RECT1_Y(rectangle1_ys[348]), .RECT1_WIDTH(rectangle1_widths[348]), .RECT1_HEIGHT(rectangle1_heights[348]), .RECT1_WEIGHT(rectangle1_weights[348]), .RECT2_X(rectangle2_xs[348]), .RECT2_Y(rectangle2_ys[348]), .RECT2_WIDTH(rectangle2_widths[348]), .RECT2_HEIGHT(rectangle2_heights[348]), .RECT2_WEIGHT(rectangle2_weights[348]), .RECT3_X(rectangle3_xs[348]), .RECT3_Y(rectangle3_ys[348]), .RECT3_WIDTH(rectangle3_widths[348]), .RECT3_HEIGHT(rectangle3_heights[348]), .RECT3_WEIGHT(rectangle3_weights[348]), .FEAT_THRES(feature_thresholds[348]), .FEAT_ABOVE(feature_aboves[348]), .FEAT_BELOW(feature_belows[348])) ac348(.scan_win(scan_win348), .scan_win_std_dev(scan_win_std_dev[348]), .feature_accum(feature_accums[348]));
  accum_calculator #(.RECT1_X(rectangle1_xs[349]), .RECT1_Y(rectangle1_ys[349]), .RECT1_WIDTH(rectangle1_widths[349]), .RECT1_HEIGHT(rectangle1_heights[349]), .RECT1_WEIGHT(rectangle1_weights[349]), .RECT2_X(rectangle2_xs[349]), .RECT2_Y(rectangle2_ys[349]), .RECT2_WIDTH(rectangle2_widths[349]), .RECT2_HEIGHT(rectangle2_heights[349]), .RECT2_WEIGHT(rectangle2_weights[349]), .RECT3_X(rectangle3_xs[349]), .RECT3_Y(rectangle3_ys[349]), .RECT3_WIDTH(rectangle3_widths[349]), .RECT3_HEIGHT(rectangle3_heights[349]), .RECT3_WEIGHT(rectangle3_weights[349]), .FEAT_THRES(feature_thresholds[349]), .FEAT_ABOVE(feature_aboves[349]), .FEAT_BELOW(feature_belows[349])) ac349(.scan_win(scan_win349), .scan_win_std_dev(scan_win_std_dev[349]), .feature_accum(feature_accums[349]));
  accum_calculator #(.RECT1_X(rectangle1_xs[350]), .RECT1_Y(rectangle1_ys[350]), .RECT1_WIDTH(rectangle1_widths[350]), .RECT1_HEIGHT(rectangle1_heights[350]), .RECT1_WEIGHT(rectangle1_weights[350]), .RECT2_X(rectangle2_xs[350]), .RECT2_Y(rectangle2_ys[350]), .RECT2_WIDTH(rectangle2_widths[350]), .RECT2_HEIGHT(rectangle2_heights[350]), .RECT2_WEIGHT(rectangle2_weights[350]), .RECT3_X(rectangle3_xs[350]), .RECT3_Y(rectangle3_ys[350]), .RECT3_WIDTH(rectangle3_widths[350]), .RECT3_HEIGHT(rectangle3_heights[350]), .RECT3_WEIGHT(rectangle3_weights[350]), .FEAT_THRES(feature_thresholds[350]), .FEAT_ABOVE(feature_aboves[350]), .FEAT_BELOW(feature_belows[350])) ac350(.scan_win(scan_win350), .scan_win_std_dev(scan_win_std_dev[350]), .feature_accum(feature_accums[350]));
  accum_calculator #(.RECT1_X(rectangle1_xs[351]), .RECT1_Y(rectangle1_ys[351]), .RECT1_WIDTH(rectangle1_widths[351]), .RECT1_HEIGHT(rectangle1_heights[351]), .RECT1_WEIGHT(rectangle1_weights[351]), .RECT2_X(rectangle2_xs[351]), .RECT2_Y(rectangle2_ys[351]), .RECT2_WIDTH(rectangle2_widths[351]), .RECT2_HEIGHT(rectangle2_heights[351]), .RECT2_WEIGHT(rectangle2_weights[351]), .RECT3_X(rectangle3_xs[351]), .RECT3_Y(rectangle3_ys[351]), .RECT3_WIDTH(rectangle3_widths[351]), .RECT3_HEIGHT(rectangle3_heights[351]), .RECT3_WEIGHT(rectangle3_weights[351]), .FEAT_THRES(feature_thresholds[351]), .FEAT_ABOVE(feature_aboves[351]), .FEAT_BELOW(feature_belows[351])) ac351(.scan_win(scan_win351), .scan_win_std_dev(scan_win_std_dev[351]), .feature_accum(feature_accums[351]));
  accum_calculator #(.RECT1_X(rectangle1_xs[352]), .RECT1_Y(rectangle1_ys[352]), .RECT1_WIDTH(rectangle1_widths[352]), .RECT1_HEIGHT(rectangle1_heights[352]), .RECT1_WEIGHT(rectangle1_weights[352]), .RECT2_X(rectangle2_xs[352]), .RECT2_Y(rectangle2_ys[352]), .RECT2_WIDTH(rectangle2_widths[352]), .RECT2_HEIGHT(rectangle2_heights[352]), .RECT2_WEIGHT(rectangle2_weights[352]), .RECT3_X(rectangle3_xs[352]), .RECT3_Y(rectangle3_ys[352]), .RECT3_WIDTH(rectangle3_widths[352]), .RECT3_HEIGHT(rectangle3_heights[352]), .RECT3_WEIGHT(rectangle3_weights[352]), .FEAT_THRES(feature_thresholds[352]), .FEAT_ABOVE(feature_aboves[352]), .FEAT_BELOW(feature_belows[352])) ac352(.scan_win(scan_win352), .scan_win_std_dev(scan_win_std_dev[352]), .feature_accum(feature_accums[352]));
  accum_calculator #(.RECT1_X(rectangle1_xs[353]), .RECT1_Y(rectangle1_ys[353]), .RECT1_WIDTH(rectangle1_widths[353]), .RECT1_HEIGHT(rectangle1_heights[353]), .RECT1_WEIGHT(rectangle1_weights[353]), .RECT2_X(rectangle2_xs[353]), .RECT2_Y(rectangle2_ys[353]), .RECT2_WIDTH(rectangle2_widths[353]), .RECT2_HEIGHT(rectangle2_heights[353]), .RECT2_WEIGHT(rectangle2_weights[353]), .RECT3_X(rectangle3_xs[353]), .RECT3_Y(rectangle3_ys[353]), .RECT3_WIDTH(rectangle3_widths[353]), .RECT3_HEIGHT(rectangle3_heights[353]), .RECT3_WEIGHT(rectangle3_weights[353]), .FEAT_THRES(feature_thresholds[353]), .FEAT_ABOVE(feature_aboves[353]), .FEAT_BELOW(feature_belows[353])) ac353(.scan_win(scan_win353), .scan_win_std_dev(scan_win_std_dev[353]), .feature_accum(feature_accums[353]));
  accum_calculator #(.RECT1_X(rectangle1_xs[354]), .RECT1_Y(rectangle1_ys[354]), .RECT1_WIDTH(rectangle1_widths[354]), .RECT1_HEIGHT(rectangle1_heights[354]), .RECT1_WEIGHT(rectangle1_weights[354]), .RECT2_X(rectangle2_xs[354]), .RECT2_Y(rectangle2_ys[354]), .RECT2_WIDTH(rectangle2_widths[354]), .RECT2_HEIGHT(rectangle2_heights[354]), .RECT2_WEIGHT(rectangle2_weights[354]), .RECT3_X(rectangle3_xs[354]), .RECT3_Y(rectangle3_ys[354]), .RECT3_WIDTH(rectangle3_widths[354]), .RECT3_HEIGHT(rectangle3_heights[354]), .RECT3_WEIGHT(rectangle3_weights[354]), .FEAT_THRES(feature_thresholds[354]), .FEAT_ABOVE(feature_aboves[354]), .FEAT_BELOW(feature_belows[354])) ac354(.scan_win(scan_win354), .scan_win_std_dev(scan_win_std_dev[354]), .feature_accum(feature_accums[354]));
  accum_calculator #(.RECT1_X(rectangle1_xs[355]), .RECT1_Y(rectangle1_ys[355]), .RECT1_WIDTH(rectangle1_widths[355]), .RECT1_HEIGHT(rectangle1_heights[355]), .RECT1_WEIGHT(rectangle1_weights[355]), .RECT2_X(rectangle2_xs[355]), .RECT2_Y(rectangle2_ys[355]), .RECT2_WIDTH(rectangle2_widths[355]), .RECT2_HEIGHT(rectangle2_heights[355]), .RECT2_WEIGHT(rectangle2_weights[355]), .RECT3_X(rectangle3_xs[355]), .RECT3_Y(rectangle3_ys[355]), .RECT3_WIDTH(rectangle3_widths[355]), .RECT3_HEIGHT(rectangle3_heights[355]), .RECT3_WEIGHT(rectangle3_weights[355]), .FEAT_THRES(feature_thresholds[355]), .FEAT_ABOVE(feature_aboves[355]), .FEAT_BELOW(feature_belows[355])) ac355(.scan_win(scan_win355), .scan_win_std_dev(scan_win_std_dev[355]), .feature_accum(feature_accums[355]));
  accum_calculator #(.RECT1_X(rectangle1_xs[356]), .RECT1_Y(rectangle1_ys[356]), .RECT1_WIDTH(rectangle1_widths[356]), .RECT1_HEIGHT(rectangle1_heights[356]), .RECT1_WEIGHT(rectangle1_weights[356]), .RECT2_X(rectangle2_xs[356]), .RECT2_Y(rectangle2_ys[356]), .RECT2_WIDTH(rectangle2_widths[356]), .RECT2_HEIGHT(rectangle2_heights[356]), .RECT2_WEIGHT(rectangle2_weights[356]), .RECT3_X(rectangle3_xs[356]), .RECT3_Y(rectangle3_ys[356]), .RECT3_WIDTH(rectangle3_widths[356]), .RECT3_HEIGHT(rectangle3_heights[356]), .RECT3_WEIGHT(rectangle3_weights[356]), .FEAT_THRES(feature_thresholds[356]), .FEAT_ABOVE(feature_aboves[356]), .FEAT_BELOW(feature_belows[356])) ac356(.scan_win(scan_win356), .scan_win_std_dev(scan_win_std_dev[356]), .feature_accum(feature_accums[356]));
  accum_calculator #(.RECT1_X(rectangle1_xs[357]), .RECT1_Y(rectangle1_ys[357]), .RECT1_WIDTH(rectangle1_widths[357]), .RECT1_HEIGHT(rectangle1_heights[357]), .RECT1_WEIGHT(rectangle1_weights[357]), .RECT2_X(rectangle2_xs[357]), .RECT2_Y(rectangle2_ys[357]), .RECT2_WIDTH(rectangle2_widths[357]), .RECT2_HEIGHT(rectangle2_heights[357]), .RECT2_WEIGHT(rectangle2_weights[357]), .RECT3_X(rectangle3_xs[357]), .RECT3_Y(rectangle3_ys[357]), .RECT3_WIDTH(rectangle3_widths[357]), .RECT3_HEIGHT(rectangle3_heights[357]), .RECT3_WEIGHT(rectangle3_weights[357]), .FEAT_THRES(feature_thresholds[357]), .FEAT_ABOVE(feature_aboves[357]), .FEAT_BELOW(feature_belows[357])) ac357(.scan_win(scan_win357), .scan_win_std_dev(scan_win_std_dev[357]), .feature_accum(feature_accums[357]));
  accum_calculator #(.RECT1_X(rectangle1_xs[358]), .RECT1_Y(rectangle1_ys[358]), .RECT1_WIDTH(rectangle1_widths[358]), .RECT1_HEIGHT(rectangle1_heights[358]), .RECT1_WEIGHT(rectangle1_weights[358]), .RECT2_X(rectangle2_xs[358]), .RECT2_Y(rectangle2_ys[358]), .RECT2_WIDTH(rectangle2_widths[358]), .RECT2_HEIGHT(rectangle2_heights[358]), .RECT2_WEIGHT(rectangle2_weights[358]), .RECT3_X(rectangle3_xs[358]), .RECT3_Y(rectangle3_ys[358]), .RECT3_WIDTH(rectangle3_widths[358]), .RECT3_HEIGHT(rectangle3_heights[358]), .RECT3_WEIGHT(rectangle3_weights[358]), .FEAT_THRES(feature_thresholds[358]), .FEAT_ABOVE(feature_aboves[358]), .FEAT_BELOW(feature_belows[358])) ac358(.scan_win(scan_win358), .scan_win_std_dev(scan_win_std_dev[358]), .feature_accum(feature_accums[358]));
  accum_calculator #(.RECT1_X(rectangle1_xs[359]), .RECT1_Y(rectangle1_ys[359]), .RECT1_WIDTH(rectangle1_widths[359]), .RECT1_HEIGHT(rectangle1_heights[359]), .RECT1_WEIGHT(rectangle1_weights[359]), .RECT2_X(rectangle2_xs[359]), .RECT2_Y(rectangle2_ys[359]), .RECT2_WIDTH(rectangle2_widths[359]), .RECT2_HEIGHT(rectangle2_heights[359]), .RECT2_WEIGHT(rectangle2_weights[359]), .RECT3_X(rectangle3_xs[359]), .RECT3_Y(rectangle3_ys[359]), .RECT3_WIDTH(rectangle3_widths[359]), .RECT3_HEIGHT(rectangle3_heights[359]), .RECT3_WEIGHT(rectangle3_weights[359]), .FEAT_THRES(feature_thresholds[359]), .FEAT_ABOVE(feature_aboves[359]), .FEAT_BELOW(feature_belows[359])) ac359(.scan_win(scan_win359), .scan_win_std_dev(scan_win_std_dev[359]), .feature_accum(feature_accums[359]));
  accum_calculator #(.RECT1_X(rectangle1_xs[360]), .RECT1_Y(rectangle1_ys[360]), .RECT1_WIDTH(rectangle1_widths[360]), .RECT1_HEIGHT(rectangle1_heights[360]), .RECT1_WEIGHT(rectangle1_weights[360]), .RECT2_X(rectangle2_xs[360]), .RECT2_Y(rectangle2_ys[360]), .RECT2_WIDTH(rectangle2_widths[360]), .RECT2_HEIGHT(rectangle2_heights[360]), .RECT2_WEIGHT(rectangle2_weights[360]), .RECT3_X(rectangle3_xs[360]), .RECT3_Y(rectangle3_ys[360]), .RECT3_WIDTH(rectangle3_widths[360]), .RECT3_HEIGHT(rectangle3_heights[360]), .RECT3_WEIGHT(rectangle3_weights[360]), .FEAT_THRES(feature_thresholds[360]), .FEAT_ABOVE(feature_aboves[360]), .FEAT_BELOW(feature_belows[360])) ac360(.scan_win(scan_win360), .scan_win_std_dev(scan_win_std_dev[360]), .feature_accum(feature_accums[360]));
  accum_calculator #(.RECT1_X(rectangle1_xs[361]), .RECT1_Y(rectangle1_ys[361]), .RECT1_WIDTH(rectangle1_widths[361]), .RECT1_HEIGHT(rectangle1_heights[361]), .RECT1_WEIGHT(rectangle1_weights[361]), .RECT2_X(rectangle2_xs[361]), .RECT2_Y(rectangle2_ys[361]), .RECT2_WIDTH(rectangle2_widths[361]), .RECT2_HEIGHT(rectangle2_heights[361]), .RECT2_WEIGHT(rectangle2_weights[361]), .RECT3_X(rectangle3_xs[361]), .RECT3_Y(rectangle3_ys[361]), .RECT3_WIDTH(rectangle3_widths[361]), .RECT3_HEIGHT(rectangle3_heights[361]), .RECT3_WEIGHT(rectangle3_weights[361]), .FEAT_THRES(feature_thresholds[361]), .FEAT_ABOVE(feature_aboves[361]), .FEAT_BELOW(feature_belows[361])) ac361(.scan_win(scan_win361), .scan_win_std_dev(scan_win_std_dev[361]), .feature_accum(feature_accums[361]));
  accum_calculator #(.RECT1_X(rectangle1_xs[362]), .RECT1_Y(rectangle1_ys[362]), .RECT1_WIDTH(rectangle1_widths[362]), .RECT1_HEIGHT(rectangle1_heights[362]), .RECT1_WEIGHT(rectangle1_weights[362]), .RECT2_X(rectangle2_xs[362]), .RECT2_Y(rectangle2_ys[362]), .RECT2_WIDTH(rectangle2_widths[362]), .RECT2_HEIGHT(rectangle2_heights[362]), .RECT2_WEIGHT(rectangle2_weights[362]), .RECT3_X(rectangle3_xs[362]), .RECT3_Y(rectangle3_ys[362]), .RECT3_WIDTH(rectangle3_widths[362]), .RECT3_HEIGHT(rectangle3_heights[362]), .RECT3_WEIGHT(rectangle3_weights[362]), .FEAT_THRES(feature_thresholds[362]), .FEAT_ABOVE(feature_aboves[362]), .FEAT_BELOW(feature_belows[362])) ac362(.scan_win(scan_win362), .scan_win_std_dev(scan_win_std_dev[362]), .feature_accum(feature_accums[362]));
  accum_calculator #(.RECT1_X(rectangle1_xs[363]), .RECT1_Y(rectangle1_ys[363]), .RECT1_WIDTH(rectangle1_widths[363]), .RECT1_HEIGHT(rectangle1_heights[363]), .RECT1_WEIGHT(rectangle1_weights[363]), .RECT2_X(rectangle2_xs[363]), .RECT2_Y(rectangle2_ys[363]), .RECT2_WIDTH(rectangle2_widths[363]), .RECT2_HEIGHT(rectangle2_heights[363]), .RECT2_WEIGHT(rectangle2_weights[363]), .RECT3_X(rectangle3_xs[363]), .RECT3_Y(rectangle3_ys[363]), .RECT3_WIDTH(rectangle3_widths[363]), .RECT3_HEIGHT(rectangle3_heights[363]), .RECT3_WEIGHT(rectangle3_weights[363]), .FEAT_THRES(feature_thresholds[363]), .FEAT_ABOVE(feature_aboves[363]), .FEAT_BELOW(feature_belows[363])) ac363(.scan_win(scan_win363), .scan_win_std_dev(scan_win_std_dev[363]), .feature_accum(feature_accums[363]));
  accum_calculator #(.RECT1_X(rectangle1_xs[364]), .RECT1_Y(rectangle1_ys[364]), .RECT1_WIDTH(rectangle1_widths[364]), .RECT1_HEIGHT(rectangle1_heights[364]), .RECT1_WEIGHT(rectangle1_weights[364]), .RECT2_X(rectangle2_xs[364]), .RECT2_Y(rectangle2_ys[364]), .RECT2_WIDTH(rectangle2_widths[364]), .RECT2_HEIGHT(rectangle2_heights[364]), .RECT2_WEIGHT(rectangle2_weights[364]), .RECT3_X(rectangle3_xs[364]), .RECT3_Y(rectangle3_ys[364]), .RECT3_WIDTH(rectangle3_widths[364]), .RECT3_HEIGHT(rectangle3_heights[364]), .RECT3_WEIGHT(rectangle3_weights[364]), .FEAT_THRES(feature_thresholds[364]), .FEAT_ABOVE(feature_aboves[364]), .FEAT_BELOW(feature_belows[364])) ac364(.scan_win(scan_win364), .scan_win_std_dev(scan_win_std_dev[364]), .feature_accum(feature_accums[364]));
  accum_calculator #(.RECT1_X(rectangle1_xs[365]), .RECT1_Y(rectangle1_ys[365]), .RECT1_WIDTH(rectangle1_widths[365]), .RECT1_HEIGHT(rectangle1_heights[365]), .RECT1_WEIGHT(rectangle1_weights[365]), .RECT2_X(rectangle2_xs[365]), .RECT2_Y(rectangle2_ys[365]), .RECT2_WIDTH(rectangle2_widths[365]), .RECT2_HEIGHT(rectangle2_heights[365]), .RECT2_WEIGHT(rectangle2_weights[365]), .RECT3_X(rectangle3_xs[365]), .RECT3_Y(rectangle3_ys[365]), .RECT3_WIDTH(rectangle3_widths[365]), .RECT3_HEIGHT(rectangle3_heights[365]), .RECT3_WEIGHT(rectangle3_weights[365]), .FEAT_THRES(feature_thresholds[365]), .FEAT_ABOVE(feature_aboves[365]), .FEAT_BELOW(feature_belows[365])) ac365(.scan_win(scan_win365), .scan_win_std_dev(scan_win_std_dev[365]), .feature_accum(feature_accums[365]));
  accum_calculator #(.RECT1_X(rectangle1_xs[366]), .RECT1_Y(rectangle1_ys[366]), .RECT1_WIDTH(rectangle1_widths[366]), .RECT1_HEIGHT(rectangle1_heights[366]), .RECT1_WEIGHT(rectangle1_weights[366]), .RECT2_X(rectangle2_xs[366]), .RECT2_Y(rectangle2_ys[366]), .RECT2_WIDTH(rectangle2_widths[366]), .RECT2_HEIGHT(rectangle2_heights[366]), .RECT2_WEIGHT(rectangle2_weights[366]), .RECT3_X(rectangle3_xs[366]), .RECT3_Y(rectangle3_ys[366]), .RECT3_WIDTH(rectangle3_widths[366]), .RECT3_HEIGHT(rectangle3_heights[366]), .RECT3_WEIGHT(rectangle3_weights[366]), .FEAT_THRES(feature_thresholds[366]), .FEAT_ABOVE(feature_aboves[366]), .FEAT_BELOW(feature_belows[366])) ac366(.scan_win(scan_win366), .scan_win_std_dev(scan_win_std_dev[366]), .feature_accum(feature_accums[366]));
  accum_calculator #(.RECT1_X(rectangle1_xs[367]), .RECT1_Y(rectangle1_ys[367]), .RECT1_WIDTH(rectangle1_widths[367]), .RECT1_HEIGHT(rectangle1_heights[367]), .RECT1_WEIGHT(rectangle1_weights[367]), .RECT2_X(rectangle2_xs[367]), .RECT2_Y(rectangle2_ys[367]), .RECT2_WIDTH(rectangle2_widths[367]), .RECT2_HEIGHT(rectangle2_heights[367]), .RECT2_WEIGHT(rectangle2_weights[367]), .RECT3_X(rectangle3_xs[367]), .RECT3_Y(rectangle3_ys[367]), .RECT3_WIDTH(rectangle3_widths[367]), .RECT3_HEIGHT(rectangle3_heights[367]), .RECT3_WEIGHT(rectangle3_weights[367]), .FEAT_THRES(feature_thresholds[367]), .FEAT_ABOVE(feature_aboves[367]), .FEAT_BELOW(feature_belows[367])) ac367(.scan_win(scan_win367), .scan_win_std_dev(scan_win_std_dev[367]), .feature_accum(feature_accums[367]));
  accum_calculator #(.RECT1_X(rectangle1_xs[368]), .RECT1_Y(rectangle1_ys[368]), .RECT1_WIDTH(rectangle1_widths[368]), .RECT1_HEIGHT(rectangle1_heights[368]), .RECT1_WEIGHT(rectangle1_weights[368]), .RECT2_X(rectangle2_xs[368]), .RECT2_Y(rectangle2_ys[368]), .RECT2_WIDTH(rectangle2_widths[368]), .RECT2_HEIGHT(rectangle2_heights[368]), .RECT2_WEIGHT(rectangle2_weights[368]), .RECT3_X(rectangle3_xs[368]), .RECT3_Y(rectangle3_ys[368]), .RECT3_WIDTH(rectangle3_widths[368]), .RECT3_HEIGHT(rectangle3_heights[368]), .RECT3_WEIGHT(rectangle3_weights[368]), .FEAT_THRES(feature_thresholds[368]), .FEAT_ABOVE(feature_aboves[368]), .FEAT_BELOW(feature_belows[368])) ac368(.scan_win(scan_win368), .scan_win_std_dev(scan_win_std_dev[368]), .feature_accum(feature_accums[368]));
  accum_calculator #(.RECT1_X(rectangle1_xs[369]), .RECT1_Y(rectangle1_ys[369]), .RECT1_WIDTH(rectangle1_widths[369]), .RECT1_HEIGHT(rectangle1_heights[369]), .RECT1_WEIGHT(rectangle1_weights[369]), .RECT2_X(rectangle2_xs[369]), .RECT2_Y(rectangle2_ys[369]), .RECT2_WIDTH(rectangle2_widths[369]), .RECT2_HEIGHT(rectangle2_heights[369]), .RECT2_WEIGHT(rectangle2_weights[369]), .RECT3_X(rectangle3_xs[369]), .RECT3_Y(rectangle3_ys[369]), .RECT3_WIDTH(rectangle3_widths[369]), .RECT3_HEIGHT(rectangle3_heights[369]), .RECT3_WEIGHT(rectangle3_weights[369]), .FEAT_THRES(feature_thresholds[369]), .FEAT_ABOVE(feature_aboves[369]), .FEAT_BELOW(feature_belows[369])) ac369(.scan_win(scan_win369), .scan_win_std_dev(scan_win_std_dev[369]), .feature_accum(feature_accums[369]));
  accum_calculator #(.RECT1_X(rectangle1_xs[370]), .RECT1_Y(rectangle1_ys[370]), .RECT1_WIDTH(rectangle1_widths[370]), .RECT1_HEIGHT(rectangle1_heights[370]), .RECT1_WEIGHT(rectangle1_weights[370]), .RECT2_X(rectangle2_xs[370]), .RECT2_Y(rectangle2_ys[370]), .RECT2_WIDTH(rectangle2_widths[370]), .RECT2_HEIGHT(rectangle2_heights[370]), .RECT2_WEIGHT(rectangle2_weights[370]), .RECT3_X(rectangle3_xs[370]), .RECT3_Y(rectangle3_ys[370]), .RECT3_WIDTH(rectangle3_widths[370]), .RECT3_HEIGHT(rectangle3_heights[370]), .RECT3_WEIGHT(rectangle3_weights[370]), .FEAT_THRES(feature_thresholds[370]), .FEAT_ABOVE(feature_aboves[370]), .FEAT_BELOW(feature_belows[370])) ac370(.scan_win(scan_win370), .scan_win_std_dev(scan_win_std_dev[370]), .feature_accum(feature_accums[370]));
  accum_calculator #(.RECT1_X(rectangle1_xs[371]), .RECT1_Y(rectangle1_ys[371]), .RECT1_WIDTH(rectangle1_widths[371]), .RECT1_HEIGHT(rectangle1_heights[371]), .RECT1_WEIGHT(rectangle1_weights[371]), .RECT2_X(rectangle2_xs[371]), .RECT2_Y(rectangle2_ys[371]), .RECT2_WIDTH(rectangle2_widths[371]), .RECT2_HEIGHT(rectangle2_heights[371]), .RECT2_WEIGHT(rectangle2_weights[371]), .RECT3_X(rectangle3_xs[371]), .RECT3_Y(rectangle3_ys[371]), .RECT3_WIDTH(rectangle3_widths[371]), .RECT3_HEIGHT(rectangle3_heights[371]), .RECT3_WEIGHT(rectangle3_weights[371]), .FEAT_THRES(feature_thresholds[371]), .FEAT_ABOVE(feature_aboves[371]), .FEAT_BELOW(feature_belows[371])) ac371(.scan_win(scan_win371), .scan_win_std_dev(scan_win_std_dev[371]), .feature_accum(feature_accums[371]));
  accum_calculator #(.RECT1_X(rectangle1_xs[372]), .RECT1_Y(rectangle1_ys[372]), .RECT1_WIDTH(rectangle1_widths[372]), .RECT1_HEIGHT(rectangle1_heights[372]), .RECT1_WEIGHT(rectangle1_weights[372]), .RECT2_X(rectangle2_xs[372]), .RECT2_Y(rectangle2_ys[372]), .RECT2_WIDTH(rectangle2_widths[372]), .RECT2_HEIGHT(rectangle2_heights[372]), .RECT2_WEIGHT(rectangle2_weights[372]), .RECT3_X(rectangle3_xs[372]), .RECT3_Y(rectangle3_ys[372]), .RECT3_WIDTH(rectangle3_widths[372]), .RECT3_HEIGHT(rectangle3_heights[372]), .RECT3_WEIGHT(rectangle3_weights[372]), .FEAT_THRES(feature_thresholds[372]), .FEAT_ABOVE(feature_aboves[372]), .FEAT_BELOW(feature_belows[372])) ac372(.scan_win(scan_win372), .scan_win_std_dev(scan_win_std_dev[372]), .feature_accum(feature_accums[372]));
  accum_calculator #(.RECT1_X(rectangle1_xs[373]), .RECT1_Y(rectangle1_ys[373]), .RECT1_WIDTH(rectangle1_widths[373]), .RECT1_HEIGHT(rectangle1_heights[373]), .RECT1_WEIGHT(rectangle1_weights[373]), .RECT2_X(rectangle2_xs[373]), .RECT2_Y(rectangle2_ys[373]), .RECT2_WIDTH(rectangle2_widths[373]), .RECT2_HEIGHT(rectangle2_heights[373]), .RECT2_WEIGHT(rectangle2_weights[373]), .RECT3_X(rectangle3_xs[373]), .RECT3_Y(rectangle3_ys[373]), .RECT3_WIDTH(rectangle3_widths[373]), .RECT3_HEIGHT(rectangle3_heights[373]), .RECT3_WEIGHT(rectangle3_weights[373]), .FEAT_THRES(feature_thresholds[373]), .FEAT_ABOVE(feature_aboves[373]), .FEAT_BELOW(feature_belows[373])) ac373(.scan_win(scan_win373), .scan_win_std_dev(scan_win_std_dev[373]), .feature_accum(feature_accums[373]));
  accum_calculator #(.RECT1_X(rectangle1_xs[374]), .RECT1_Y(rectangle1_ys[374]), .RECT1_WIDTH(rectangle1_widths[374]), .RECT1_HEIGHT(rectangle1_heights[374]), .RECT1_WEIGHT(rectangle1_weights[374]), .RECT2_X(rectangle2_xs[374]), .RECT2_Y(rectangle2_ys[374]), .RECT2_WIDTH(rectangle2_widths[374]), .RECT2_HEIGHT(rectangle2_heights[374]), .RECT2_WEIGHT(rectangle2_weights[374]), .RECT3_X(rectangle3_xs[374]), .RECT3_Y(rectangle3_ys[374]), .RECT3_WIDTH(rectangle3_widths[374]), .RECT3_HEIGHT(rectangle3_heights[374]), .RECT3_WEIGHT(rectangle3_weights[374]), .FEAT_THRES(feature_thresholds[374]), .FEAT_ABOVE(feature_aboves[374]), .FEAT_BELOW(feature_belows[374])) ac374(.scan_win(scan_win374), .scan_win_std_dev(scan_win_std_dev[374]), .feature_accum(feature_accums[374]));
  accum_calculator #(.RECT1_X(rectangle1_xs[375]), .RECT1_Y(rectangle1_ys[375]), .RECT1_WIDTH(rectangle1_widths[375]), .RECT1_HEIGHT(rectangle1_heights[375]), .RECT1_WEIGHT(rectangle1_weights[375]), .RECT2_X(rectangle2_xs[375]), .RECT2_Y(rectangle2_ys[375]), .RECT2_WIDTH(rectangle2_widths[375]), .RECT2_HEIGHT(rectangle2_heights[375]), .RECT2_WEIGHT(rectangle2_weights[375]), .RECT3_X(rectangle3_xs[375]), .RECT3_Y(rectangle3_ys[375]), .RECT3_WIDTH(rectangle3_widths[375]), .RECT3_HEIGHT(rectangle3_heights[375]), .RECT3_WEIGHT(rectangle3_weights[375]), .FEAT_THRES(feature_thresholds[375]), .FEAT_ABOVE(feature_aboves[375]), .FEAT_BELOW(feature_belows[375])) ac375(.scan_win(scan_win375), .scan_win_std_dev(scan_win_std_dev[375]), .feature_accum(feature_accums[375]));
  accum_calculator #(.RECT1_X(rectangle1_xs[376]), .RECT1_Y(rectangle1_ys[376]), .RECT1_WIDTH(rectangle1_widths[376]), .RECT1_HEIGHT(rectangle1_heights[376]), .RECT1_WEIGHT(rectangle1_weights[376]), .RECT2_X(rectangle2_xs[376]), .RECT2_Y(rectangle2_ys[376]), .RECT2_WIDTH(rectangle2_widths[376]), .RECT2_HEIGHT(rectangle2_heights[376]), .RECT2_WEIGHT(rectangle2_weights[376]), .RECT3_X(rectangle3_xs[376]), .RECT3_Y(rectangle3_ys[376]), .RECT3_WIDTH(rectangle3_widths[376]), .RECT3_HEIGHT(rectangle3_heights[376]), .RECT3_WEIGHT(rectangle3_weights[376]), .FEAT_THRES(feature_thresholds[376]), .FEAT_ABOVE(feature_aboves[376]), .FEAT_BELOW(feature_belows[376])) ac376(.scan_win(scan_win376), .scan_win_std_dev(scan_win_std_dev[376]), .feature_accum(feature_accums[376]));
  accum_calculator #(.RECT1_X(rectangle1_xs[377]), .RECT1_Y(rectangle1_ys[377]), .RECT1_WIDTH(rectangle1_widths[377]), .RECT1_HEIGHT(rectangle1_heights[377]), .RECT1_WEIGHT(rectangle1_weights[377]), .RECT2_X(rectangle2_xs[377]), .RECT2_Y(rectangle2_ys[377]), .RECT2_WIDTH(rectangle2_widths[377]), .RECT2_HEIGHT(rectangle2_heights[377]), .RECT2_WEIGHT(rectangle2_weights[377]), .RECT3_X(rectangle3_xs[377]), .RECT3_Y(rectangle3_ys[377]), .RECT3_WIDTH(rectangle3_widths[377]), .RECT3_HEIGHT(rectangle3_heights[377]), .RECT3_WEIGHT(rectangle3_weights[377]), .FEAT_THRES(feature_thresholds[377]), .FEAT_ABOVE(feature_aboves[377]), .FEAT_BELOW(feature_belows[377])) ac377(.scan_win(scan_win377), .scan_win_std_dev(scan_win_std_dev[377]), .feature_accum(feature_accums[377]));
  accum_calculator #(.RECT1_X(rectangle1_xs[378]), .RECT1_Y(rectangle1_ys[378]), .RECT1_WIDTH(rectangle1_widths[378]), .RECT1_HEIGHT(rectangle1_heights[378]), .RECT1_WEIGHT(rectangle1_weights[378]), .RECT2_X(rectangle2_xs[378]), .RECT2_Y(rectangle2_ys[378]), .RECT2_WIDTH(rectangle2_widths[378]), .RECT2_HEIGHT(rectangle2_heights[378]), .RECT2_WEIGHT(rectangle2_weights[378]), .RECT3_X(rectangle3_xs[378]), .RECT3_Y(rectangle3_ys[378]), .RECT3_WIDTH(rectangle3_widths[378]), .RECT3_HEIGHT(rectangle3_heights[378]), .RECT3_WEIGHT(rectangle3_weights[378]), .FEAT_THRES(feature_thresholds[378]), .FEAT_ABOVE(feature_aboves[378]), .FEAT_BELOW(feature_belows[378])) ac378(.scan_win(scan_win378), .scan_win_std_dev(scan_win_std_dev[378]), .feature_accum(feature_accums[378]));
  accum_calculator #(.RECT1_X(rectangle1_xs[379]), .RECT1_Y(rectangle1_ys[379]), .RECT1_WIDTH(rectangle1_widths[379]), .RECT1_HEIGHT(rectangle1_heights[379]), .RECT1_WEIGHT(rectangle1_weights[379]), .RECT2_X(rectangle2_xs[379]), .RECT2_Y(rectangle2_ys[379]), .RECT2_WIDTH(rectangle2_widths[379]), .RECT2_HEIGHT(rectangle2_heights[379]), .RECT2_WEIGHT(rectangle2_weights[379]), .RECT3_X(rectangle3_xs[379]), .RECT3_Y(rectangle3_ys[379]), .RECT3_WIDTH(rectangle3_widths[379]), .RECT3_HEIGHT(rectangle3_heights[379]), .RECT3_WEIGHT(rectangle3_weights[379]), .FEAT_THRES(feature_thresholds[379]), .FEAT_ABOVE(feature_aboves[379]), .FEAT_BELOW(feature_belows[379])) ac379(.scan_win(scan_win379), .scan_win_std_dev(scan_win_std_dev[379]), .feature_accum(feature_accums[379]));
  accum_calculator #(.RECT1_X(rectangle1_xs[380]), .RECT1_Y(rectangle1_ys[380]), .RECT1_WIDTH(rectangle1_widths[380]), .RECT1_HEIGHT(rectangle1_heights[380]), .RECT1_WEIGHT(rectangle1_weights[380]), .RECT2_X(rectangle2_xs[380]), .RECT2_Y(rectangle2_ys[380]), .RECT2_WIDTH(rectangle2_widths[380]), .RECT2_HEIGHT(rectangle2_heights[380]), .RECT2_WEIGHT(rectangle2_weights[380]), .RECT3_X(rectangle3_xs[380]), .RECT3_Y(rectangle3_ys[380]), .RECT3_WIDTH(rectangle3_widths[380]), .RECT3_HEIGHT(rectangle3_heights[380]), .RECT3_WEIGHT(rectangle3_weights[380]), .FEAT_THRES(feature_thresholds[380]), .FEAT_ABOVE(feature_aboves[380]), .FEAT_BELOW(feature_belows[380])) ac380(.scan_win(scan_win380), .scan_win_std_dev(scan_win_std_dev[380]), .feature_accum(feature_accums[380]));
  accum_calculator #(.RECT1_X(rectangle1_xs[381]), .RECT1_Y(rectangle1_ys[381]), .RECT1_WIDTH(rectangle1_widths[381]), .RECT1_HEIGHT(rectangle1_heights[381]), .RECT1_WEIGHT(rectangle1_weights[381]), .RECT2_X(rectangle2_xs[381]), .RECT2_Y(rectangle2_ys[381]), .RECT2_WIDTH(rectangle2_widths[381]), .RECT2_HEIGHT(rectangle2_heights[381]), .RECT2_WEIGHT(rectangle2_weights[381]), .RECT3_X(rectangle3_xs[381]), .RECT3_Y(rectangle3_ys[381]), .RECT3_WIDTH(rectangle3_widths[381]), .RECT3_HEIGHT(rectangle3_heights[381]), .RECT3_WEIGHT(rectangle3_weights[381]), .FEAT_THRES(feature_thresholds[381]), .FEAT_ABOVE(feature_aboves[381]), .FEAT_BELOW(feature_belows[381])) ac381(.scan_win(scan_win381), .scan_win_std_dev(scan_win_std_dev[381]), .feature_accum(feature_accums[381]));
  accum_calculator #(.RECT1_X(rectangle1_xs[382]), .RECT1_Y(rectangle1_ys[382]), .RECT1_WIDTH(rectangle1_widths[382]), .RECT1_HEIGHT(rectangle1_heights[382]), .RECT1_WEIGHT(rectangle1_weights[382]), .RECT2_X(rectangle2_xs[382]), .RECT2_Y(rectangle2_ys[382]), .RECT2_WIDTH(rectangle2_widths[382]), .RECT2_HEIGHT(rectangle2_heights[382]), .RECT2_WEIGHT(rectangle2_weights[382]), .RECT3_X(rectangle3_xs[382]), .RECT3_Y(rectangle3_ys[382]), .RECT3_WIDTH(rectangle3_widths[382]), .RECT3_HEIGHT(rectangle3_heights[382]), .RECT3_WEIGHT(rectangle3_weights[382]), .FEAT_THRES(feature_thresholds[382]), .FEAT_ABOVE(feature_aboves[382]), .FEAT_BELOW(feature_belows[382])) ac382(.scan_win(scan_win382), .scan_win_std_dev(scan_win_std_dev[382]), .feature_accum(feature_accums[382]));
  accum_calculator #(.RECT1_X(rectangle1_xs[383]), .RECT1_Y(rectangle1_ys[383]), .RECT1_WIDTH(rectangle1_widths[383]), .RECT1_HEIGHT(rectangle1_heights[383]), .RECT1_WEIGHT(rectangle1_weights[383]), .RECT2_X(rectangle2_xs[383]), .RECT2_Y(rectangle2_ys[383]), .RECT2_WIDTH(rectangle2_widths[383]), .RECT2_HEIGHT(rectangle2_heights[383]), .RECT2_WEIGHT(rectangle2_weights[383]), .RECT3_X(rectangle3_xs[383]), .RECT3_Y(rectangle3_ys[383]), .RECT3_WIDTH(rectangle3_widths[383]), .RECT3_HEIGHT(rectangle3_heights[383]), .RECT3_WEIGHT(rectangle3_weights[383]), .FEAT_THRES(feature_thresholds[383]), .FEAT_ABOVE(feature_aboves[383]), .FEAT_BELOW(feature_belows[383])) ac383(.scan_win(scan_win383), .scan_win_std_dev(scan_win_std_dev[383]), .feature_accum(feature_accums[383]));
  accum_calculator #(.RECT1_X(rectangle1_xs[384]), .RECT1_Y(rectangle1_ys[384]), .RECT1_WIDTH(rectangle1_widths[384]), .RECT1_HEIGHT(rectangle1_heights[384]), .RECT1_WEIGHT(rectangle1_weights[384]), .RECT2_X(rectangle2_xs[384]), .RECT2_Y(rectangle2_ys[384]), .RECT2_WIDTH(rectangle2_widths[384]), .RECT2_HEIGHT(rectangle2_heights[384]), .RECT2_WEIGHT(rectangle2_weights[384]), .RECT3_X(rectangle3_xs[384]), .RECT3_Y(rectangle3_ys[384]), .RECT3_WIDTH(rectangle3_widths[384]), .RECT3_HEIGHT(rectangle3_heights[384]), .RECT3_WEIGHT(rectangle3_weights[384]), .FEAT_THRES(feature_thresholds[384]), .FEAT_ABOVE(feature_aboves[384]), .FEAT_BELOW(feature_belows[384])) ac384(.scan_win(scan_win384), .scan_win_std_dev(scan_win_std_dev[384]), .feature_accum(feature_accums[384]));
  accum_calculator #(.RECT1_X(rectangle1_xs[385]), .RECT1_Y(rectangle1_ys[385]), .RECT1_WIDTH(rectangle1_widths[385]), .RECT1_HEIGHT(rectangle1_heights[385]), .RECT1_WEIGHT(rectangle1_weights[385]), .RECT2_X(rectangle2_xs[385]), .RECT2_Y(rectangle2_ys[385]), .RECT2_WIDTH(rectangle2_widths[385]), .RECT2_HEIGHT(rectangle2_heights[385]), .RECT2_WEIGHT(rectangle2_weights[385]), .RECT3_X(rectangle3_xs[385]), .RECT3_Y(rectangle3_ys[385]), .RECT3_WIDTH(rectangle3_widths[385]), .RECT3_HEIGHT(rectangle3_heights[385]), .RECT3_WEIGHT(rectangle3_weights[385]), .FEAT_THRES(feature_thresholds[385]), .FEAT_ABOVE(feature_aboves[385]), .FEAT_BELOW(feature_belows[385])) ac385(.scan_win(scan_win385), .scan_win_std_dev(scan_win_std_dev[385]), .feature_accum(feature_accums[385]));
  accum_calculator #(.RECT1_X(rectangle1_xs[386]), .RECT1_Y(rectangle1_ys[386]), .RECT1_WIDTH(rectangle1_widths[386]), .RECT1_HEIGHT(rectangle1_heights[386]), .RECT1_WEIGHT(rectangle1_weights[386]), .RECT2_X(rectangle2_xs[386]), .RECT2_Y(rectangle2_ys[386]), .RECT2_WIDTH(rectangle2_widths[386]), .RECT2_HEIGHT(rectangle2_heights[386]), .RECT2_WEIGHT(rectangle2_weights[386]), .RECT3_X(rectangle3_xs[386]), .RECT3_Y(rectangle3_ys[386]), .RECT3_WIDTH(rectangle3_widths[386]), .RECT3_HEIGHT(rectangle3_heights[386]), .RECT3_WEIGHT(rectangle3_weights[386]), .FEAT_THRES(feature_thresholds[386]), .FEAT_ABOVE(feature_aboves[386]), .FEAT_BELOW(feature_belows[386])) ac386(.scan_win(scan_win386), .scan_win_std_dev(scan_win_std_dev[386]), .feature_accum(feature_accums[386]));
  accum_calculator #(.RECT1_X(rectangle1_xs[387]), .RECT1_Y(rectangle1_ys[387]), .RECT1_WIDTH(rectangle1_widths[387]), .RECT1_HEIGHT(rectangle1_heights[387]), .RECT1_WEIGHT(rectangle1_weights[387]), .RECT2_X(rectangle2_xs[387]), .RECT2_Y(rectangle2_ys[387]), .RECT2_WIDTH(rectangle2_widths[387]), .RECT2_HEIGHT(rectangle2_heights[387]), .RECT2_WEIGHT(rectangle2_weights[387]), .RECT3_X(rectangle3_xs[387]), .RECT3_Y(rectangle3_ys[387]), .RECT3_WIDTH(rectangle3_widths[387]), .RECT3_HEIGHT(rectangle3_heights[387]), .RECT3_WEIGHT(rectangle3_weights[387]), .FEAT_THRES(feature_thresholds[387]), .FEAT_ABOVE(feature_aboves[387]), .FEAT_BELOW(feature_belows[387])) ac387(.scan_win(scan_win387), .scan_win_std_dev(scan_win_std_dev[387]), .feature_accum(feature_accums[387]));
  accum_calculator #(.RECT1_X(rectangle1_xs[388]), .RECT1_Y(rectangle1_ys[388]), .RECT1_WIDTH(rectangle1_widths[388]), .RECT1_HEIGHT(rectangle1_heights[388]), .RECT1_WEIGHT(rectangle1_weights[388]), .RECT2_X(rectangle2_xs[388]), .RECT2_Y(rectangle2_ys[388]), .RECT2_WIDTH(rectangle2_widths[388]), .RECT2_HEIGHT(rectangle2_heights[388]), .RECT2_WEIGHT(rectangle2_weights[388]), .RECT3_X(rectangle3_xs[388]), .RECT3_Y(rectangle3_ys[388]), .RECT3_WIDTH(rectangle3_widths[388]), .RECT3_HEIGHT(rectangle3_heights[388]), .RECT3_WEIGHT(rectangle3_weights[388]), .FEAT_THRES(feature_thresholds[388]), .FEAT_ABOVE(feature_aboves[388]), .FEAT_BELOW(feature_belows[388])) ac388(.scan_win(scan_win388), .scan_win_std_dev(scan_win_std_dev[388]), .feature_accum(feature_accums[388]));
  accum_calculator #(.RECT1_X(rectangle1_xs[389]), .RECT1_Y(rectangle1_ys[389]), .RECT1_WIDTH(rectangle1_widths[389]), .RECT1_HEIGHT(rectangle1_heights[389]), .RECT1_WEIGHT(rectangle1_weights[389]), .RECT2_X(rectangle2_xs[389]), .RECT2_Y(rectangle2_ys[389]), .RECT2_WIDTH(rectangle2_widths[389]), .RECT2_HEIGHT(rectangle2_heights[389]), .RECT2_WEIGHT(rectangle2_weights[389]), .RECT3_X(rectangle3_xs[389]), .RECT3_Y(rectangle3_ys[389]), .RECT3_WIDTH(rectangle3_widths[389]), .RECT3_HEIGHT(rectangle3_heights[389]), .RECT3_WEIGHT(rectangle3_weights[389]), .FEAT_THRES(feature_thresholds[389]), .FEAT_ABOVE(feature_aboves[389]), .FEAT_BELOW(feature_belows[389])) ac389(.scan_win(scan_win389), .scan_win_std_dev(scan_win_std_dev[389]), .feature_accum(feature_accums[389]));
  accum_calculator #(.RECT1_X(rectangle1_xs[390]), .RECT1_Y(rectangle1_ys[390]), .RECT1_WIDTH(rectangle1_widths[390]), .RECT1_HEIGHT(rectangle1_heights[390]), .RECT1_WEIGHT(rectangle1_weights[390]), .RECT2_X(rectangle2_xs[390]), .RECT2_Y(rectangle2_ys[390]), .RECT2_WIDTH(rectangle2_widths[390]), .RECT2_HEIGHT(rectangle2_heights[390]), .RECT2_WEIGHT(rectangle2_weights[390]), .RECT3_X(rectangle3_xs[390]), .RECT3_Y(rectangle3_ys[390]), .RECT3_WIDTH(rectangle3_widths[390]), .RECT3_HEIGHT(rectangle3_heights[390]), .RECT3_WEIGHT(rectangle3_weights[390]), .FEAT_THRES(feature_thresholds[390]), .FEAT_ABOVE(feature_aboves[390]), .FEAT_BELOW(feature_belows[390])) ac390(.scan_win(scan_win390), .scan_win_std_dev(scan_win_std_dev[390]), .feature_accum(feature_accums[390]));
  accum_calculator #(.RECT1_X(rectangle1_xs[391]), .RECT1_Y(rectangle1_ys[391]), .RECT1_WIDTH(rectangle1_widths[391]), .RECT1_HEIGHT(rectangle1_heights[391]), .RECT1_WEIGHT(rectangle1_weights[391]), .RECT2_X(rectangle2_xs[391]), .RECT2_Y(rectangle2_ys[391]), .RECT2_WIDTH(rectangle2_widths[391]), .RECT2_HEIGHT(rectangle2_heights[391]), .RECT2_WEIGHT(rectangle2_weights[391]), .RECT3_X(rectangle3_xs[391]), .RECT3_Y(rectangle3_ys[391]), .RECT3_WIDTH(rectangle3_widths[391]), .RECT3_HEIGHT(rectangle3_heights[391]), .RECT3_WEIGHT(rectangle3_weights[391]), .FEAT_THRES(feature_thresholds[391]), .FEAT_ABOVE(feature_aboves[391]), .FEAT_BELOW(feature_belows[391])) ac391(.scan_win(scan_win391), .scan_win_std_dev(scan_win_std_dev[391]), .feature_accum(feature_accums[391]));
  accum_calculator #(.RECT1_X(rectangle1_xs[392]), .RECT1_Y(rectangle1_ys[392]), .RECT1_WIDTH(rectangle1_widths[392]), .RECT1_HEIGHT(rectangle1_heights[392]), .RECT1_WEIGHT(rectangle1_weights[392]), .RECT2_X(rectangle2_xs[392]), .RECT2_Y(rectangle2_ys[392]), .RECT2_WIDTH(rectangle2_widths[392]), .RECT2_HEIGHT(rectangle2_heights[392]), .RECT2_WEIGHT(rectangle2_weights[392]), .RECT3_X(rectangle3_xs[392]), .RECT3_Y(rectangle3_ys[392]), .RECT3_WIDTH(rectangle3_widths[392]), .RECT3_HEIGHT(rectangle3_heights[392]), .RECT3_WEIGHT(rectangle3_weights[392]), .FEAT_THRES(feature_thresholds[392]), .FEAT_ABOVE(feature_aboves[392]), .FEAT_BELOW(feature_belows[392])) ac392(.scan_win(scan_win392), .scan_win_std_dev(scan_win_std_dev[392]), .feature_accum(feature_accums[392]));
  accum_calculator #(.RECT1_X(rectangle1_xs[393]), .RECT1_Y(rectangle1_ys[393]), .RECT1_WIDTH(rectangle1_widths[393]), .RECT1_HEIGHT(rectangle1_heights[393]), .RECT1_WEIGHT(rectangle1_weights[393]), .RECT2_X(rectangle2_xs[393]), .RECT2_Y(rectangle2_ys[393]), .RECT2_WIDTH(rectangle2_widths[393]), .RECT2_HEIGHT(rectangle2_heights[393]), .RECT2_WEIGHT(rectangle2_weights[393]), .RECT3_X(rectangle3_xs[393]), .RECT3_Y(rectangle3_ys[393]), .RECT3_WIDTH(rectangle3_widths[393]), .RECT3_HEIGHT(rectangle3_heights[393]), .RECT3_WEIGHT(rectangle3_weights[393]), .FEAT_THRES(feature_thresholds[393]), .FEAT_ABOVE(feature_aboves[393]), .FEAT_BELOW(feature_belows[393])) ac393(.scan_win(scan_win393), .scan_win_std_dev(scan_win_std_dev[393]), .feature_accum(feature_accums[393]));
  accum_calculator #(.RECT1_X(rectangle1_xs[394]), .RECT1_Y(rectangle1_ys[394]), .RECT1_WIDTH(rectangle1_widths[394]), .RECT1_HEIGHT(rectangle1_heights[394]), .RECT1_WEIGHT(rectangle1_weights[394]), .RECT2_X(rectangle2_xs[394]), .RECT2_Y(rectangle2_ys[394]), .RECT2_WIDTH(rectangle2_widths[394]), .RECT2_HEIGHT(rectangle2_heights[394]), .RECT2_WEIGHT(rectangle2_weights[394]), .RECT3_X(rectangle3_xs[394]), .RECT3_Y(rectangle3_ys[394]), .RECT3_WIDTH(rectangle3_widths[394]), .RECT3_HEIGHT(rectangle3_heights[394]), .RECT3_WEIGHT(rectangle3_weights[394]), .FEAT_THRES(feature_thresholds[394]), .FEAT_ABOVE(feature_aboves[394]), .FEAT_BELOW(feature_belows[394])) ac394(.scan_win(scan_win394), .scan_win_std_dev(scan_win_std_dev[394]), .feature_accum(feature_accums[394]));
  accum_calculator #(.RECT1_X(rectangle1_xs[395]), .RECT1_Y(rectangle1_ys[395]), .RECT1_WIDTH(rectangle1_widths[395]), .RECT1_HEIGHT(rectangle1_heights[395]), .RECT1_WEIGHT(rectangle1_weights[395]), .RECT2_X(rectangle2_xs[395]), .RECT2_Y(rectangle2_ys[395]), .RECT2_WIDTH(rectangle2_widths[395]), .RECT2_HEIGHT(rectangle2_heights[395]), .RECT2_WEIGHT(rectangle2_weights[395]), .RECT3_X(rectangle3_xs[395]), .RECT3_Y(rectangle3_ys[395]), .RECT3_WIDTH(rectangle3_widths[395]), .RECT3_HEIGHT(rectangle3_heights[395]), .RECT3_WEIGHT(rectangle3_weights[395]), .FEAT_THRES(feature_thresholds[395]), .FEAT_ABOVE(feature_aboves[395]), .FEAT_BELOW(feature_belows[395])) ac395(.scan_win(scan_win395), .scan_win_std_dev(scan_win_std_dev[395]), .feature_accum(feature_accums[395]));
  accum_calculator #(.RECT1_X(rectangle1_xs[396]), .RECT1_Y(rectangle1_ys[396]), .RECT1_WIDTH(rectangle1_widths[396]), .RECT1_HEIGHT(rectangle1_heights[396]), .RECT1_WEIGHT(rectangle1_weights[396]), .RECT2_X(rectangle2_xs[396]), .RECT2_Y(rectangle2_ys[396]), .RECT2_WIDTH(rectangle2_widths[396]), .RECT2_HEIGHT(rectangle2_heights[396]), .RECT2_WEIGHT(rectangle2_weights[396]), .RECT3_X(rectangle3_xs[396]), .RECT3_Y(rectangle3_ys[396]), .RECT3_WIDTH(rectangle3_widths[396]), .RECT3_HEIGHT(rectangle3_heights[396]), .RECT3_WEIGHT(rectangle3_weights[396]), .FEAT_THRES(feature_thresholds[396]), .FEAT_ABOVE(feature_aboves[396]), .FEAT_BELOW(feature_belows[396])) ac396(.scan_win(scan_win396), .scan_win_std_dev(scan_win_std_dev[396]), .feature_accum(feature_accums[396]));
  accum_calculator #(.RECT1_X(rectangle1_xs[397]), .RECT1_Y(rectangle1_ys[397]), .RECT1_WIDTH(rectangle1_widths[397]), .RECT1_HEIGHT(rectangle1_heights[397]), .RECT1_WEIGHT(rectangle1_weights[397]), .RECT2_X(rectangle2_xs[397]), .RECT2_Y(rectangle2_ys[397]), .RECT2_WIDTH(rectangle2_widths[397]), .RECT2_HEIGHT(rectangle2_heights[397]), .RECT2_WEIGHT(rectangle2_weights[397]), .RECT3_X(rectangle3_xs[397]), .RECT3_Y(rectangle3_ys[397]), .RECT3_WIDTH(rectangle3_widths[397]), .RECT3_HEIGHT(rectangle3_heights[397]), .RECT3_WEIGHT(rectangle3_weights[397]), .FEAT_THRES(feature_thresholds[397]), .FEAT_ABOVE(feature_aboves[397]), .FEAT_BELOW(feature_belows[397])) ac397(.scan_win(scan_win397), .scan_win_std_dev(scan_win_std_dev[397]), .feature_accum(feature_accums[397]));
  accum_calculator #(.RECT1_X(rectangle1_xs[398]), .RECT1_Y(rectangle1_ys[398]), .RECT1_WIDTH(rectangle1_widths[398]), .RECT1_HEIGHT(rectangle1_heights[398]), .RECT1_WEIGHT(rectangle1_weights[398]), .RECT2_X(rectangle2_xs[398]), .RECT2_Y(rectangle2_ys[398]), .RECT2_WIDTH(rectangle2_widths[398]), .RECT2_HEIGHT(rectangle2_heights[398]), .RECT2_WEIGHT(rectangle2_weights[398]), .RECT3_X(rectangle3_xs[398]), .RECT3_Y(rectangle3_ys[398]), .RECT3_WIDTH(rectangle3_widths[398]), .RECT3_HEIGHT(rectangle3_heights[398]), .RECT3_WEIGHT(rectangle3_weights[398]), .FEAT_THRES(feature_thresholds[398]), .FEAT_ABOVE(feature_aboves[398]), .FEAT_BELOW(feature_belows[398])) ac398(.scan_win(scan_win398), .scan_win_std_dev(scan_win_std_dev[398]), .feature_accum(feature_accums[398]));
  accum_calculator #(.RECT1_X(rectangle1_xs[399]), .RECT1_Y(rectangle1_ys[399]), .RECT1_WIDTH(rectangle1_widths[399]), .RECT1_HEIGHT(rectangle1_heights[399]), .RECT1_WEIGHT(rectangle1_weights[399]), .RECT2_X(rectangle2_xs[399]), .RECT2_Y(rectangle2_ys[399]), .RECT2_WIDTH(rectangle2_widths[399]), .RECT2_HEIGHT(rectangle2_heights[399]), .RECT2_WEIGHT(rectangle2_weights[399]), .RECT3_X(rectangle3_xs[399]), .RECT3_Y(rectangle3_ys[399]), .RECT3_WIDTH(rectangle3_widths[399]), .RECT3_HEIGHT(rectangle3_heights[399]), .RECT3_WEIGHT(rectangle3_weights[399]), .FEAT_THRES(feature_thresholds[399]), .FEAT_ABOVE(feature_aboves[399]), .FEAT_BELOW(feature_belows[399])) ac399(.scan_win(scan_win399), .scan_win_std_dev(scan_win_std_dev[399]), .feature_accum(feature_accums[399]));
  accum_calculator #(.RECT1_X(rectangle1_xs[400]), .RECT1_Y(rectangle1_ys[400]), .RECT1_WIDTH(rectangle1_widths[400]), .RECT1_HEIGHT(rectangle1_heights[400]), .RECT1_WEIGHT(rectangle1_weights[400]), .RECT2_X(rectangle2_xs[400]), .RECT2_Y(rectangle2_ys[400]), .RECT2_WIDTH(rectangle2_widths[400]), .RECT2_HEIGHT(rectangle2_heights[400]), .RECT2_WEIGHT(rectangle2_weights[400]), .RECT3_X(rectangle3_xs[400]), .RECT3_Y(rectangle3_ys[400]), .RECT3_WIDTH(rectangle3_widths[400]), .RECT3_HEIGHT(rectangle3_heights[400]), .RECT3_WEIGHT(rectangle3_weights[400]), .FEAT_THRES(feature_thresholds[400]), .FEAT_ABOVE(feature_aboves[400]), .FEAT_BELOW(feature_belows[400])) ac400(.scan_win(scan_win400), .scan_win_std_dev(scan_win_std_dev[400]), .feature_accum(feature_accums[400]));
  accum_calculator #(.RECT1_X(rectangle1_xs[401]), .RECT1_Y(rectangle1_ys[401]), .RECT1_WIDTH(rectangle1_widths[401]), .RECT1_HEIGHT(rectangle1_heights[401]), .RECT1_WEIGHT(rectangle1_weights[401]), .RECT2_X(rectangle2_xs[401]), .RECT2_Y(rectangle2_ys[401]), .RECT2_WIDTH(rectangle2_widths[401]), .RECT2_HEIGHT(rectangle2_heights[401]), .RECT2_WEIGHT(rectangle2_weights[401]), .RECT3_X(rectangle3_xs[401]), .RECT3_Y(rectangle3_ys[401]), .RECT3_WIDTH(rectangle3_widths[401]), .RECT3_HEIGHT(rectangle3_heights[401]), .RECT3_WEIGHT(rectangle3_weights[401]), .FEAT_THRES(feature_thresholds[401]), .FEAT_ABOVE(feature_aboves[401]), .FEAT_BELOW(feature_belows[401])) ac401(.scan_win(scan_win401), .scan_win_std_dev(scan_win_std_dev[401]), .feature_accum(feature_accums[401]));
  accum_calculator #(.RECT1_X(rectangle1_xs[402]), .RECT1_Y(rectangle1_ys[402]), .RECT1_WIDTH(rectangle1_widths[402]), .RECT1_HEIGHT(rectangle1_heights[402]), .RECT1_WEIGHT(rectangle1_weights[402]), .RECT2_X(rectangle2_xs[402]), .RECT2_Y(rectangle2_ys[402]), .RECT2_WIDTH(rectangle2_widths[402]), .RECT2_HEIGHT(rectangle2_heights[402]), .RECT2_WEIGHT(rectangle2_weights[402]), .RECT3_X(rectangle3_xs[402]), .RECT3_Y(rectangle3_ys[402]), .RECT3_WIDTH(rectangle3_widths[402]), .RECT3_HEIGHT(rectangle3_heights[402]), .RECT3_WEIGHT(rectangle3_weights[402]), .FEAT_THRES(feature_thresholds[402]), .FEAT_ABOVE(feature_aboves[402]), .FEAT_BELOW(feature_belows[402])) ac402(.scan_win(scan_win402), .scan_win_std_dev(scan_win_std_dev[402]), .feature_accum(feature_accums[402]));
  accum_calculator #(.RECT1_X(rectangle1_xs[403]), .RECT1_Y(rectangle1_ys[403]), .RECT1_WIDTH(rectangle1_widths[403]), .RECT1_HEIGHT(rectangle1_heights[403]), .RECT1_WEIGHT(rectangle1_weights[403]), .RECT2_X(rectangle2_xs[403]), .RECT2_Y(rectangle2_ys[403]), .RECT2_WIDTH(rectangle2_widths[403]), .RECT2_HEIGHT(rectangle2_heights[403]), .RECT2_WEIGHT(rectangle2_weights[403]), .RECT3_X(rectangle3_xs[403]), .RECT3_Y(rectangle3_ys[403]), .RECT3_WIDTH(rectangle3_widths[403]), .RECT3_HEIGHT(rectangle3_heights[403]), .RECT3_WEIGHT(rectangle3_weights[403]), .FEAT_THRES(feature_thresholds[403]), .FEAT_ABOVE(feature_aboves[403]), .FEAT_BELOW(feature_belows[403])) ac403(.scan_win(scan_win403), .scan_win_std_dev(scan_win_std_dev[403]), .feature_accum(feature_accums[403]));
  accum_calculator #(.RECT1_X(rectangle1_xs[404]), .RECT1_Y(rectangle1_ys[404]), .RECT1_WIDTH(rectangle1_widths[404]), .RECT1_HEIGHT(rectangle1_heights[404]), .RECT1_WEIGHT(rectangle1_weights[404]), .RECT2_X(rectangle2_xs[404]), .RECT2_Y(rectangle2_ys[404]), .RECT2_WIDTH(rectangle2_widths[404]), .RECT2_HEIGHT(rectangle2_heights[404]), .RECT2_WEIGHT(rectangle2_weights[404]), .RECT3_X(rectangle3_xs[404]), .RECT3_Y(rectangle3_ys[404]), .RECT3_WIDTH(rectangle3_widths[404]), .RECT3_HEIGHT(rectangle3_heights[404]), .RECT3_WEIGHT(rectangle3_weights[404]), .FEAT_THRES(feature_thresholds[404]), .FEAT_ABOVE(feature_aboves[404]), .FEAT_BELOW(feature_belows[404])) ac404(.scan_win(scan_win404), .scan_win_std_dev(scan_win_std_dev[404]), .feature_accum(feature_accums[404]));
  accum_calculator #(.RECT1_X(rectangle1_xs[405]), .RECT1_Y(rectangle1_ys[405]), .RECT1_WIDTH(rectangle1_widths[405]), .RECT1_HEIGHT(rectangle1_heights[405]), .RECT1_WEIGHT(rectangle1_weights[405]), .RECT2_X(rectangle2_xs[405]), .RECT2_Y(rectangle2_ys[405]), .RECT2_WIDTH(rectangle2_widths[405]), .RECT2_HEIGHT(rectangle2_heights[405]), .RECT2_WEIGHT(rectangle2_weights[405]), .RECT3_X(rectangle3_xs[405]), .RECT3_Y(rectangle3_ys[405]), .RECT3_WIDTH(rectangle3_widths[405]), .RECT3_HEIGHT(rectangle3_heights[405]), .RECT3_WEIGHT(rectangle3_weights[405]), .FEAT_THRES(feature_thresholds[405]), .FEAT_ABOVE(feature_aboves[405]), .FEAT_BELOW(feature_belows[405])) ac405(.scan_win(scan_win405), .scan_win_std_dev(scan_win_std_dev[405]), .feature_accum(feature_accums[405]));
  accum_calculator #(.RECT1_X(rectangle1_xs[406]), .RECT1_Y(rectangle1_ys[406]), .RECT1_WIDTH(rectangle1_widths[406]), .RECT1_HEIGHT(rectangle1_heights[406]), .RECT1_WEIGHT(rectangle1_weights[406]), .RECT2_X(rectangle2_xs[406]), .RECT2_Y(rectangle2_ys[406]), .RECT2_WIDTH(rectangle2_widths[406]), .RECT2_HEIGHT(rectangle2_heights[406]), .RECT2_WEIGHT(rectangle2_weights[406]), .RECT3_X(rectangle3_xs[406]), .RECT3_Y(rectangle3_ys[406]), .RECT3_WIDTH(rectangle3_widths[406]), .RECT3_HEIGHT(rectangle3_heights[406]), .RECT3_WEIGHT(rectangle3_weights[406]), .FEAT_THRES(feature_thresholds[406]), .FEAT_ABOVE(feature_aboves[406]), .FEAT_BELOW(feature_belows[406])) ac406(.scan_win(scan_win406), .scan_win_std_dev(scan_win_std_dev[406]), .feature_accum(feature_accums[406]));
  accum_calculator #(.RECT1_X(rectangle1_xs[407]), .RECT1_Y(rectangle1_ys[407]), .RECT1_WIDTH(rectangle1_widths[407]), .RECT1_HEIGHT(rectangle1_heights[407]), .RECT1_WEIGHT(rectangle1_weights[407]), .RECT2_X(rectangle2_xs[407]), .RECT2_Y(rectangle2_ys[407]), .RECT2_WIDTH(rectangle2_widths[407]), .RECT2_HEIGHT(rectangle2_heights[407]), .RECT2_WEIGHT(rectangle2_weights[407]), .RECT3_X(rectangle3_xs[407]), .RECT3_Y(rectangle3_ys[407]), .RECT3_WIDTH(rectangle3_widths[407]), .RECT3_HEIGHT(rectangle3_heights[407]), .RECT3_WEIGHT(rectangle3_weights[407]), .FEAT_THRES(feature_thresholds[407]), .FEAT_ABOVE(feature_aboves[407]), .FEAT_BELOW(feature_belows[407])) ac407(.scan_win(scan_win407), .scan_win_std_dev(scan_win_std_dev[407]), .feature_accum(feature_accums[407]));
  accum_calculator #(.RECT1_X(rectangle1_xs[408]), .RECT1_Y(rectangle1_ys[408]), .RECT1_WIDTH(rectangle1_widths[408]), .RECT1_HEIGHT(rectangle1_heights[408]), .RECT1_WEIGHT(rectangle1_weights[408]), .RECT2_X(rectangle2_xs[408]), .RECT2_Y(rectangle2_ys[408]), .RECT2_WIDTH(rectangle2_widths[408]), .RECT2_HEIGHT(rectangle2_heights[408]), .RECT2_WEIGHT(rectangle2_weights[408]), .RECT3_X(rectangle3_xs[408]), .RECT3_Y(rectangle3_ys[408]), .RECT3_WIDTH(rectangle3_widths[408]), .RECT3_HEIGHT(rectangle3_heights[408]), .RECT3_WEIGHT(rectangle3_weights[408]), .FEAT_THRES(feature_thresholds[408]), .FEAT_ABOVE(feature_aboves[408]), .FEAT_BELOW(feature_belows[408])) ac408(.scan_win(scan_win408), .scan_win_std_dev(scan_win_std_dev[408]), .feature_accum(feature_accums[408]));
  accum_calculator #(.RECT1_X(rectangle1_xs[409]), .RECT1_Y(rectangle1_ys[409]), .RECT1_WIDTH(rectangle1_widths[409]), .RECT1_HEIGHT(rectangle1_heights[409]), .RECT1_WEIGHT(rectangle1_weights[409]), .RECT2_X(rectangle2_xs[409]), .RECT2_Y(rectangle2_ys[409]), .RECT2_WIDTH(rectangle2_widths[409]), .RECT2_HEIGHT(rectangle2_heights[409]), .RECT2_WEIGHT(rectangle2_weights[409]), .RECT3_X(rectangle3_xs[409]), .RECT3_Y(rectangle3_ys[409]), .RECT3_WIDTH(rectangle3_widths[409]), .RECT3_HEIGHT(rectangle3_heights[409]), .RECT3_WEIGHT(rectangle3_weights[409]), .FEAT_THRES(feature_thresholds[409]), .FEAT_ABOVE(feature_aboves[409]), .FEAT_BELOW(feature_belows[409])) ac409(.scan_win(scan_win409), .scan_win_std_dev(scan_win_std_dev[409]), .feature_accum(feature_accums[409]));
  accum_calculator #(.RECT1_X(rectangle1_xs[410]), .RECT1_Y(rectangle1_ys[410]), .RECT1_WIDTH(rectangle1_widths[410]), .RECT1_HEIGHT(rectangle1_heights[410]), .RECT1_WEIGHT(rectangle1_weights[410]), .RECT2_X(rectangle2_xs[410]), .RECT2_Y(rectangle2_ys[410]), .RECT2_WIDTH(rectangle2_widths[410]), .RECT2_HEIGHT(rectangle2_heights[410]), .RECT2_WEIGHT(rectangle2_weights[410]), .RECT3_X(rectangle3_xs[410]), .RECT3_Y(rectangle3_ys[410]), .RECT3_WIDTH(rectangle3_widths[410]), .RECT3_HEIGHT(rectangle3_heights[410]), .RECT3_WEIGHT(rectangle3_weights[410]), .FEAT_THRES(feature_thresholds[410]), .FEAT_ABOVE(feature_aboves[410]), .FEAT_BELOW(feature_belows[410])) ac410(.scan_win(scan_win410), .scan_win_std_dev(scan_win_std_dev[410]), .feature_accum(feature_accums[410]));
  accum_calculator #(.RECT1_X(rectangle1_xs[411]), .RECT1_Y(rectangle1_ys[411]), .RECT1_WIDTH(rectangle1_widths[411]), .RECT1_HEIGHT(rectangle1_heights[411]), .RECT1_WEIGHT(rectangle1_weights[411]), .RECT2_X(rectangle2_xs[411]), .RECT2_Y(rectangle2_ys[411]), .RECT2_WIDTH(rectangle2_widths[411]), .RECT2_HEIGHT(rectangle2_heights[411]), .RECT2_WEIGHT(rectangle2_weights[411]), .RECT3_X(rectangle3_xs[411]), .RECT3_Y(rectangle3_ys[411]), .RECT3_WIDTH(rectangle3_widths[411]), .RECT3_HEIGHT(rectangle3_heights[411]), .RECT3_WEIGHT(rectangle3_weights[411]), .FEAT_THRES(feature_thresholds[411]), .FEAT_ABOVE(feature_aboves[411]), .FEAT_BELOW(feature_belows[411])) ac411(.scan_win(scan_win411), .scan_win_std_dev(scan_win_std_dev[411]), .feature_accum(feature_accums[411]));
  accum_calculator #(.RECT1_X(rectangle1_xs[412]), .RECT1_Y(rectangle1_ys[412]), .RECT1_WIDTH(rectangle1_widths[412]), .RECT1_HEIGHT(rectangle1_heights[412]), .RECT1_WEIGHT(rectangle1_weights[412]), .RECT2_X(rectangle2_xs[412]), .RECT2_Y(rectangle2_ys[412]), .RECT2_WIDTH(rectangle2_widths[412]), .RECT2_HEIGHT(rectangle2_heights[412]), .RECT2_WEIGHT(rectangle2_weights[412]), .RECT3_X(rectangle3_xs[412]), .RECT3_Y(rectangle3_ys[412]), .RECT3_WIDTH(rectangle3_widths[412]), .RECT3_HEIGHT(rectangle3_heights[412]), .RECT3_WEIGHT(rectangle3_weights[412]), .FEAT_THRES(feature_thresholds[412]), .FEAT_ABOVE(feature_aboves[412]), .FEAT_BELOW(feature_belows[412])) ac412(.scan_win(scan_win412), .scan_win_std_dev(scan_win_std_dev[412]), .feature_accum(feature_accums[412]));
  accum_calculator #(.RECT1_X(rectangle1_xs[413]), .RECT1_Y(rectangle1_ys[413]), .RECT1_WIDTH(rectangle1_widths[413]), .RECT1_HEIGHT(rectangle1_heights[413]), .RECT1_WEIGHT(rectangle1_weights[413]), .RECT2_X(rectangle2_xs[413]), .RECT2_Y(rectangle2_ys[413]), .RECT2_WIDTH(rectangle2_widths[413]), .RECT2_HEIGHT(rectangle2_heights[413]), .RECT2_WEIGHT(rectangle2_weights[413]), .RECT3_X(rectangle3_xs[413]), .RECT3_Y(rectangle3_ys[413]), .RECT3_WIDTH(rectangle3_widths[413]), .RECT3_HEIGHT(rectangle3_heights[413]), .RECT3_WEIGHT(rectangle3_weights[413]), .FEAT_THRES(feature_thresholds[413]), .FEAT_ABOVE(feature_aboves[413]), .FEAT_BELOW(feature_belows[413])) ac413(.scan_win(scan_win413), .scan_win_std_dev(scan_win_std_dev[413]), .feature_accum(feature_accums[413]));
  accum_calculator #(.RECT1_X(rectangle1_xs[414]), .RECT1_Y(rectangle1_ys[414]), .RECT1_WIDTH(rectangle1_widths[414]), .RECT1_HEIGHT(rectangle1_heights[414]), .RECT1_WEIGHT(rectangle1_weights[414]), .RECT2_X(rectangle2_xs[414]), .RECT2_Y(rectangle2_ys[414]), .RECT2_WIDTH(rectangle2_widths[414]), .RECT2_HEIGHT(rectangle2_heights[414]), .RECT2_WEIGHT(rectangle2_weights[414]), .RECT3_X(rectangle3_xs[414]), .RECT3_Y(rectangle3_ys[414]), .RECT3_WIDTH(rectangle3_widths[414]), .RECT3_HEIGHT(rectangle3_heights[414]), .RECT3_WEIGHT(rectangle3_weights[414]), .FEAT_THRES(feature_thresholds[414]), .FEAT_ABOVE(feature_aboves[414]), .FEAT_BELOW(feature_belows[414])) ac414(.scan_win(scan_win414), .scan_win_std_dev(scan_win_std_dev[414]), .feature_accum(feature_accums[414]));
  accum_calculator #(.RECT1_X(rectangle1_xs[415]), .RECT1_Y(rectangle1_ys[415]), .RECT1_WIDTH(rectangle1_widths[415]), .RECT1_HEIGHT(rectangle1_heights[415]), .RECT1_WEIGHT(rectangle1_weights[415]), .RECT2_X(rectangle2_xs[415]), .RECT2_Y(rectangle2_ys[415]), .RECT2_WIDTH(rectangle2_widths[415]), .RECT2_HEIGHT(rectangle2_heights[415]), .RECT2_WEIGHT(rectangle2_weights[415]), .RECT3_X(rectangle3_xs[415]), .RECT3_Y(rectangle3_ys[415]), .RECT3_WIDTH(rectangle3_widths[415]), .RECT3_HEIGHT(rectangle3_heights[415]), .RECT3_WEIGHT(rectangle3_weights[415]), .FEAT_THRES(feature_thresholds[415]), .FEAT_ABOVE(feature_aboves[415]), .FEAT_BELOW(feature_belows[415])) ac415(.scan_win(scan_win415), .scan_win_std_dev(scan_win_std_dev[415]), .feature_accum(feature_accums[415]));
  accum_calculator #(.RECT1_X(rectangle1_xs[416]), .RECT1_Y(rectangle1_ys[416]), .RECT1_WIDTH(rectangle1_widths[416]), .RECT1_HEIGHT(rectangle1_heights[416]), .RECT1_WEIGHT(rectangle1_weights[416]), .RECT2_X(rectangle2_xs[416]), .RECT2_Y(rectangle2_ys[416]), .RECT2_WIDTH(rectangle2_widths[416]), .RECT2_HEIGHT(rectangle2_heights[416]), .RECT2_WEIGHT(rectangle2_weights[416]), .RECT3_X(rectangle3_xs[416]), .RECT3_Y(rectangle3_ys[416]), .RECT3_WIDTH(rectangle3_widths[416]), .RECT3_HEIGHT(rectangle3_heights[416]), .RECT3_WEIGHT(rectangle3_weights[416]), .FEAT_THRES(feature_thresholds[416]), .FEAT_ABOVE(feature_aboves[416]), .FEAT_BELOW(feature_belows[416])) ac416(.scan_win(scan_win416), .scan_win_std_dev(scan_win_std_dev[416]), .feature_accum(feature_accums[416]));
  accum_calculator #(.RECT1_X(rectangle1_xs[417]), .RECT1_Y(rectangle1_ys[417]), .RECT1_WIDTH(rectangle1_widths[417]), .RECT1_HEIGHT(rectangle1_heights[417]), .RECT1_WEIGHT(rectangle1_weights[417]), .RECT2_X(rectangle2_xs[417]), .RECT2_Y(rectangle2_ys[417]), .RECT2_WIDTH(rectangle2_widths[417]), .RECT2_HEIGHT(rectangle2_heights[417]), .RECT2_WEIGHT(rectangle2_weights[417]), .RECT3_X(rectangle3_xs[417]), .RECT3_Y(rectangle3_ys[417]), .RECT3_WIDTH(rectangle3_widths[417]), .RECT3_HEIGHT(rectangle3_heights[417]), .RECT3_WEIGHT(rectangle3_weights[417]), .FEAT_THRES(feature_thresholds[417]), .FEAT_ABOVE(feature_aboves[417]), .FEAT_BELOW(feature_belows[417])) ac417(.scan_win(scan_win417), .scan_win_std_dev(scan_win_std_dev[417]), .feature_accum(feature_accums[417]));
  accum_calculator #(.RECT1_X(rectangle1_xs[418]), .RECT1_Y(rectangle1_ys[418]), .RECT1_WIDTH(rectangle1_widths[418]), .RECT1_HEIGHT(rectangle1_heights[418]), .RECT1_WEIGHT(rectangle1_weights[418]), .RECT2_X(rectangle2_xs[418]), .RECT2_Y(rectangle2_ys[418]), .RECT2_WIDTH(rectangle2_widths[418]), .RECT2_HEIGHT(rectangle2_heights[418]), .RECT2_WEIGHT(rectangle2_weights[418]), .RECT3_X(rectangle3_xs[418]), .RECT3_Y(rectangle3_ys[418]), .RECT3_WIDTH(rectangle3_widths[418]), .RECT3_HEIGHT(rectangle3_heights[418]), .RECT3_WEIGHT(rectangle3_weights[418]), .FEAT_THRES(feature_thresholds[418]), .FEAT_ABOVE(feature_aboves[418]), .FEAT_BELOW(feature_belows[418])) ac418(.scan_win(scan_win418), .scan_win_std_dev(scan_win_std_dev[418]), .feature_accum(feature_accums[418]));
  accum_calculator #(.RECT1_X(rectangle1_xs[419]), .RECT1_Y(rectangle1_ys[419]), .RECT1_WIDTH(rectangle1_widths[419]), .RECT1_HEIGHT(rectangle1_heights[419]), .RECT1_WEIGHT(rectangle1_weights[419]), .RECT2_X(rectangle2_xs[419]), .RECT2_Y(rectangle2_ys[419]), .RECT2_WIDTH(rectangle2_widths[419]), .RECT2_HEIGHT(rectangle2_heights[419]), .RECT2_WEIGHT(rectangle2_weights[419]), .RECT3_X(rectangle3_xs[419]), .RECT3_Y(rectangle3_ys[419]), .RECT3_WIDTH(rectangle3_widths[419]), .RECT3_HEIGHT(rectangle3_heights[419]), .RECT3_WEIGHT(rectangle3_weights[419]), .FEAT_THRES(feature_thresholds[419]), .FEAT_ABOVE(feature_aboves[419]), .FEAT_BELOW(feature_belows[419])) ac419(.scan_win(scan_win419), .scan_win_std_dev(scan_win_std_dev[419]), .feature_accum(feature_accums[419]));
  accum_calculator #(.RECT1_X(rectangle1_xs[420]), .RECT1_Y(rectangle1_ys[420]), .RECT1_WIDTH(rectangle1_widths[420]), .RECT1_HEIGHT(rectangle1_heights[420]), .RECT1_WEIGHT(rectangle1_weights[420]), .RECT2_X(rectangle2_xs[420]), .RECT2_Y(rectangle2_ys[420]), .RECT2_WIDTH(rectangle2_widths[420]), .RECT2_HEIGHT(rectangle2_heights[420]), .RECT2_WEIGHT(rectangle2_weights[420]), .RECT3_X(rectangle3_xs[420]), .RECT3_Y(rectangle3_ys[420]), .RECT3_WIDTH(rectangle3_widths[420]), .RECT3_HEIGHT(rectangle3_heights[420]), .RECT3_WEIGHT(rectangle3_weights[420]), .FEAT_THRES(feature_thresholds[420]), .FEAT_ABOVE(feature_aboves[420]), .FEAT_BELOW(feature_belows[420])) ac420(.scan_win(scan_win420), .scan_win_std_dev(scan_win_std_dev[420]), .feature_accum(feature_accums[420]));
  accum_calculator #(.RECT1_X(rectangle1_xs[421]), .RECT1_Y(rectangle1_ys[421]), .RECT1_WIDTH(rectangle1_widths[421]), .RECT1_HEIGHT(rectangle1_heights[421]), .RECT1_WEIGHT(rectangle1_weights[421]), .RECT2_X(rectangle2_xs[421]), .RECT2_Y(rectangle2_ys[421]), .RECT2_WIDTH(rectangle2_widths[421]), .RECT2_HEIGHT(rectangle2_heights[421]), .RECT2_WEIGHT(rectangle2_weights[421]), .RECT3_X(rectangle3_xs[421]), .RECT3_Y(rectangle3_ys[421]), .RECT3_WIDTH(rectangle3_widths[421]), .RECT3_HEIGHT(rectangle3_heights[421]), .RECT3_WEIGHT(rectangle3_weights[421]), .FEAT_THRES(feature_thresholds[421]), .FEAT_ABOVE(feature_aboves[421]), .FEAT_BELOW(feature_belows[421])) ac421(.scan_win(scan_win421), .scan_win_std_dev(scan_win_std_dev[421]), .feature_accum(feature_accums[421]));
  accum_calculator #(.RECT1_X(rectangle1_xs[422]), .RECT1_Y(rectangle1_ys[422]), .RECT1_WIDTH(rectangle1_widths[422]), .RECT1_HEIGHT(rectangle1_heights[422]), .RECT1_WEIGHT(rectangle1_weights[422]), .RECT2_X(rectangle2_xs[422]), .RECT2_Y(rectangle2_ys[422]), .RECT2_WIDTH(rectangle2_widths[422]), .RECT2_HEIGHT(rectangle2_heights[422]), .RECT2_WEIGHT(rectangle2_weights[422]), .RECT3_X(rectangle3_xs[422]), .RECT3_Y(rectangle3_ys[422]), .RECT3_WIDTH(rectangle3_widths[422]), .RECT3_HEIGHT(rectangle3_heights[422]), .RECT3_WEIGHT(rectangle3_weights[422]), .FEAT_THRES(feature_thresholds[422]), .FEAT_ABOVE(feature_aboves[422]), .FEAT_BELOW(feature_belows[422])) ac422(.scan_win(scan_win422), .scan_win_std_dev(scan_win_std_dev[422]), .feature_accum(feature_accums[422]));
  accum_calculator #(.RECT1_X(rectangle1_xs[423]), .RECT1_Y(rectangle1_ys[423]), .RECT1_WIDTH(rectangle1_widths[423]), .RECT1_HEIGHT(rectangle1_heights[423]), .RECT1_WEIGHT(rectangle1_weights[423]), .RECT2_X(rectangle2_xs[423]), .RECT2_Y(rectangle2_ys[423]), .RECT2_WIDTH(rectangle2_widths[423]), .RECT2_HEIGHT(rectangle2_heights[423]), .RECT2_WEIGHT(rectangle2_weights[423]), .RECT3_X(rectangle3_xs[423]), .RECT3_Y(rectangle3_ys[423]), .RECT3_WIDTH(rectangle3_widths[423]), .RECT3_HEIGHT(rectangle3_heights[423]), .RECT3_WEIGHT(rectangle3_weights[423]), .FEAT_THRES(feature_thresholds[423]), .FEAT_ABOVE(feature_aboves[423]), .FEAT_BELOW(feature_belows[423])) ac423(.scan_win(scan_win423), .scan_win_std_dev(scan_win_std_dev[423]), .feature_accum(feature_accums[423]));
  accum_calculator #(.RECT1_X(rectangle1_xs[424]), .RECT1_Y(rectangle1_ys[424]), .RECT1_WIDTH(rectangle1_widths[424]), .RECT1_HEIGHT(rectangle1_heights[424]), .RECT1_WEIGHT(rectangle1_weights[424]), .RECT2_X(rectangle2_xs[424]), .RECT2_Y(rectangle2_ys[424]), .RECT2_WIDTH(rectangle2_widths[424]), .RECT2_HEIGHT(rectangle2_heights[424]), .RECT2_WEIGHT(rectangle2_weights[424]), .RECT3_X(rectangle3_xs[424]), .RECT3_Y(rectangle3_ys[424]), .RECT3_WIDTH(rectangle3_widths[424]), .RECT3_HEIGHT(rectangle3_heights[424]), .RECT3_WEIGHT(rectangle3_weights[424]), .FEAT_THRES(feature_thresholds[424]), .FEAT_ABOVE(feature_aboves[424]), .FEAT_BELOW(feature_belows[424])) ac424(.scan_win(scan_win424), .scan_win_std_dev(scan_win_std_dev[424]), .feature_accum(feature_accums[424]));
  accum_calculator #(.RECT1_X(rectangle1_xs[425]), .RECT1_Y(rectangle1_ys[425]), .RECT1_WIDTH(rectangle1_widths[425]), .RECT1_HEIGHT(rectangle1_heights[425]), .RECT1_WEIGHT(rectangle1_weights[425]), .RECT2_X(rectangle2_xs[425]), .RECT2_Y(rectangle2_ys[425]), .RECT2_WIDTH(rectangle2_widths[425]), .RECT2_HEIGHT(rectangle2_heights[425]), .RECT2_WEIGHT(rectangle2_weights[425]), .RECT3_X(rectangle3_xs[425]), .RECT3_Y(rectangle3_ys[425]), .RECT3_WIDTH(rectangle3_widths[425]), .RECT3_HEIGHT(rectangle3_heights[425]), .RECT3_WEIGHT(rectangle3_weights[425]), .FEAT_THRES(feature_thresholds[425]), .FEAT_ABOVE(feature_aboves[425]), .FEAT_BELOW(feature_belows[425])) ac425(.scan_win(scan_win425), .scan_win_std_dev(scan_win_std_dev[425]), .feature_accum(feature_accums[425]));
  accum_calculator #(.RECT1_X(rectangle1_xs[426]), .RECT1_Y(rectangle1_ys[426]), .RECT1_WIDTH(rectangle1_widths[426]), .RECT1_HEIGHT(rectangle1_heights[426]), .RECT1_WEIGHT(rectangle1_weights[426]), .RECT2_X(rectangle2_xs[426]), .RECT2_Y(rectangle2_ys[426]), .RECT2_WIDTH(rectangle2_widths[426]), .RECT2_HEIGHT(rectangle2_heights[426]), .RECT2_WEIGHT(rectangle2_weights[426]), .RECT3_X(rectangle3_xs[426]), .RECT3_Y(rectangle3_ys[426]), .RECT3_WIDTH(rectangle3_widths[426]), .RECT3_HEIGHT(rectangle3_heights[426]), .RECT3_WEIGHT(rectangle3_weights[426]), .FEAT_THRES(feature_thresholds[426]), .FEAT_ABOVE(feature_aboves[426]), .FEAT_BELOW(feature_belows[426])) ac426(.scan_win(scan_win426), .scan_win_std_dev(scan_win_std_dev[426]), .feature_accum(feature_accums[426]));
  accum_calculator #(.RECT1_X(rectangle1_xs[427]), .RECT1_Y(rectangle1_ys[427]), .RECT1_WIDTH(rectangle1_widths[427]), .RECT1_HEIGHT(rectangle1_heights[427]), .RECT1_WEIGHT(rectangle1_weights[427]), .RECT2_X(rectangle2_xs[427]), .RECT2_Y(rectangle2_ys[427]), .RECT2_WIDTH(rectangle2_widths[427]), .RECT2_HEIGHT(rectangle2_heights[427]), .RECT2_WEIGHT(rectangle2_weights[427]), .RECT3_X(rectangle3_xs[427]), .RECT3_Y(rectangle3_ys[427]), .RECT3_WIDTH(rectangle3_widths[427]), .RECT3_HEIGHT(rectangle3_heights[427]), .RECT3_WEIGHT(rectangle3_weights[427]), .FEAT_THRES(feature_thresholds[427]), .FEAT_ABOVE(feature_aboves[427]), .FEAT_BELOW(feature_belows[427])) ac427(.scan_win(scan_win427), .scan_win_std_dev(scan_win_std_dev[427]), .feature_accum(feature_accums[427]));
  accum_calculator #(.RECT1_X(rectangle1_xs[428]), .RECT1_Y(rectangle1_ys[428]), .RECT1_WIDTH(rectangle1_widths[428]), .RECT1_HEIGHT(rectangle1_heights[428]), .RECT1_WEIGHT(rectangle1_weights[428]), .RECT2_X(rectangle2_xs[428]), .RECT2_Y(rectangle2_ys[428]), .RECT2_WIDTH(rectangle2_widths[428]), .RECT2_HEIGHT(rectangle2_heights[428]), .RECT2_WEIGHT(rectangle2_weights[428]), .RECT3_X(rectangle3_xs[428]), .RECT3_Y(rectangle3_ys[428]), .RECT3_WIDTH(rectangle3_widths[428]), .RECT3_HEIGHT(rectangle3_heights[428]), .RECT3_WEIGHT(rectangle3_weights[428]), .FEAT_THRES(feature_thresholds[428]), .FEAT_ABOVE(feature_aboves[428]), .FEAT_BELOW(feature_belows[428])) ac428(.scan_win(scan_win428), .scan_win_std_dev(scan_win_std_dev[428]), .feature_accum(feature_accums[428]));
  accum_calculator #(.RECT1_X(rectangle1_xs[429]), .RECT1_Y(rectangle1_ys[429]), .RECT1_WIDTH(rectangle1_widths[429]), .RECT1_HEIGHT(rectangle1_heights[429]), .RECT1_WEIGHT(rectangle1_weights[429]), .RECT2_X(rectangle2_xs[429]), .RECT2_Y(rectangle2_ys[429]), .RECT2_WIDTH(rectangle2_widths[429]), .RECT2_HEIGHT(rectangle2_heights[429]), .RECT2_WEIGHT(rectangle2_weights[429]), .RECT3_X(rectangle3_xs[429]), .RECT3_Y(rectangle3_ys[429]), .RECT3_WIDTH(rectangle3_widths[429]), .RECT3_HEIGHT(rectangle3_heights[429]), .RECT3_WEIGHT(rectangle3_weights[429]), .FEAT_THRES(feature_thresholds[429]), .FEAT_ABOVE(feature_aboves[429]), .FEAT_BELOW(feature_belows[429])) ac429(.scan_win(scan_win429), .scan_win_std_dev(scan_win_std_dev[429]), .feature_accum(feature_accums[429]));
  accum_calculator #(.RECT1_X(rectangle1_xs[430]), .RECT1_Y(rectangle1_ys[430]), .RECT1_WIDTH(rectangle1_widths[430]), .RECT1_HEIGHT(rectangle1_heights[430]), .RECT1_WEIGHT(rectangle1_weights[430]), .RECT2_X(rectangle2_xs[430]), .RECT2_Y(rectangle2_ys[430]), .RECT2_WIDTH(rectangle2_widths[430]), .RECT2_HEIGHT(rectangle2_heights[430]), .RECT2_WEIGHT(rectangle2_weights[430]), .RECT3_X(rectangle3_xs[430]), .RECT3_Y(rectangle3_ys[430]), .RECT3_WIDTH(rectangle3_widths[430]), .RECT3_HEIGHT(rectangle3_heights[430]), .RECT3_WEIGHT(rectangle3_weights[430]), .FEAT_THRES(feature_thresholds[430]), .FEAT_ABOVE(feature_aboves[430]), .FEAT_BELOW(feature_belows[430])) ac430(.scan_win(scan_win430), .scan_win_std_dev(scan_win_std_dev[430]), .feature_accum(feature_accums[430]));
  accum_calculator #(.RECT1_X(rectangle1_xs[431]), .RECT1_Y(rectangle1_ys[431]), .RECT1_WIDTH(rectangle1_widths[431]), .RECT1_HEIGHT(rectangle1_heights[431]), .RECT1_WEIGHT(rectangle1_weights[431]), .RECT2_X(rectangle2_xs[431]), .RECT2_Y(rectangle2_ys[431]), .RECT2_WIDTH(rectangle2_widths[431]), .RECT2_HEIGHT(rectangle2_heights[431]), .RECT2_WEIGHT(rectangle2_weights[431]), .RECT3_X(rectangle3_xs[431]), .RECT3_Y(rectangle3_ys[431]), .RECT3_WIDTH(rectangle3_widths[431]), .RECT3_HEIGHT(rectangle3_heights[431]), .RECT3_WEIGHT(rectangle3_weights[431]), .FEAT_THRES(feature_thresholds[431]), .FEAT_ABOVE(feature_aboves[431]), .FEAT_BELOW(feature_belows[431])) ac431(.scan_win(scan_win431), .scan_win_std_dev(scan_win_std_dev[431]), .feature_accum(feature_accums[431]));
  accum_calculator #(.RECT1_X(rectangle1_xs[432]), .RECT1_Y(rectangle1_ys[432]), .RECT1_WIDTH(rectangle1_widths[432]), .RECT1_HEIGHT(rectangle1_heights[432]), .RECT1_WEIGHT(rectangle1_weights[432]), .RECT2_X(rectangle2_xs[432]), .RECT2_Y(rectangle2_ys[432]), .RECT2_WIDTH(rectangle2_widths[432]), .RECT2_HEIGHT(rectangle2_heights[432]), .RECT2_WEIGHT(rectangle2_weights[432]), .RECT3_X(rectangle3_xs[432]), .RECT3_Y(rectangle3_ys[432]), .RECT3_WIDTH(rectangle3_widths[432]), .RECT3_HEIGHT(rectangle3_heights[432]), .RECT3_WEIGHT(rectangle3_weights[432]), .FEAT_THRES(feature_thresholds[432]), .FEAT_ABOVE(feature_aboves[432]), .FEAT_BELOW(feature_belows[432])) ac432(.scan_win(scan_win432), .scan_win_std_dev(scan_win_std_dev[432]), .feature_accum(feature_accums[432]));
  accum_calculator #(.RECT1_X(rectangle1_xs[433]), .RECT1_Y(rectangle1_ys[433]), .RECT1_WIDTH(rectangle1_widths[433]), .RECT1_HEIGHT(rectangle1_heights[433]), .RECT1_WEIGHT(rectangle1_weights[433]), .RECT2_X(rectangle2_xs[433]), .RECT2_Y(rectangle2_ys[433]), .RECT2_WIDTH(rectangle2_widths[433]), .RECT2_HEIGHT(rectangle2_heights[433]), .RECT2_WEIGHT(rectangle2_weights[433]), .RECT3_X(rectangle3_xs[433]), .RECT3_Y(rectangle3_ys[433]), .RECT3_WIDTH(rectangle3_widths[433]), .RECT3_HEIGHT(rectangle3_heights[433]), .RECT3_WEIGHT(rectangle3_weights[433]), .FEAT_THRES(feature_thresholds[433]), .FEAT_ABOVE(feature_aboves[433]), .FEAT_BELOW(feature_belows[433])) ac433(.scan_win(scan_win433), .scan_win_std_dev(scan_win_std_dev[433]), .feature_accum(feature_accums[433]));
  accum_calculator #(.RECT1_X(rectangle1_xs[434]), .RECT1_Y(rectangle1_ys[434]), .RECT1_WIDTH(rectangle1_widths[434]), .RECT1_HEIGHT(rectangle1_heights[434]), .RECT1_WEIGHT(rectangle1_weights[434]), .RECT2_X(rectangle2_xs[434]), .RECT2_Y(rectangle2_ys[434]), .RECT2_WIDTH(rectangle2_widths[434]), .RECT2_HEIGHT(rectangle2_heights[434]), .RECT2_WEIGHT(rectangle2_weights[434]), .RECT3_X(rectangle3_xs[434]), .RECT3_Y(rectangle3_ys[434]), .RECT3_WIDTH(rectangle3_widths[434]), .RECT3_HEIGHT(rectangle3_heights[434]), .RECT3_WEIGHT(rectangle3_weights[434]), .FEAT_THRES(feature_thresholds[434]), .FEAT_ABOVE(feature_aboves[434]), .FEAT_BELOW(feature_belows[434])) ac434(.scan_win(scan_win434), .scan_win_std_dev(scan_win_std_dev[434]), .feature_accum(feature_accums[434]));
  accum_calculator #(.RECT1_X(rectangle1_xs[435]), .RECT1_Y(rectangle1_ys[435]), .RECT1_WIDTH(rectangle1_widths[435]), .RECT1_HEIGHT(rectangle1_heights[435]), .RECT1_WEIGHT(rectangle1_weights[435]), .RECT2_X(rectangle2_xs[435]), .RECT2_Y(rectangle2_ys[435]), .RECT2_WIDTH(rectangle2_widths[435]), .RECT2_HEIGHT(rectangle2_heights[435]), .RECT2_WEIGHT(rectangle2_weights[435]), .RECT3_X(rectangle3_xs[435]), .RECT3_Y(rectangle3_ys[435]), .RECT3_WIDTH(rectangle3_widths[435]), .RECT3_HEIGHT(rectangle3_heights[435]), .RECT3_WEIGHT(rectangle3_weights[435]), .FEAT_THRES(feature_thresholds[435]), .FEAT_ABOVE(feature_aboves[435]), .FEAT_BELOW(feature_belows[435])) ac435(.scan_win(scan_win435), .scan_win_std_dev(scan_win_std_dev[435]), .feature_accum(feature_accums[435]));
  accum_calculator #(.RECT1_X(rectangle1_xs[436]), .RECT1_Y(rectangle1_ys[436]), .RECT1_WIDTH(rectangle1_widths[436]), .RECT1_HEIGHT(rectangle1_heights[436]), .RECT1_WEIGHT(rectangle1_weights[436]), .RECT2_X(rectangle2_xs[436]), .RECT2_Y(rectangle2_ys[436]), .RECT2_WIDTH(rectangle2_widths[436]), .RECT2_HEIGHT(rectangle2_heights[436]), .RECT2_WEIGHT(rectangle2_weights[436]), .RECT3_X(rectangle3_xs[436]), .RECT3_Y(rectangle3_ys[436]), .RECT3_WIDTH(rectangle3_widths[436]), .RECT3_HEIGHT(rectangle3_heights[436]), .RECT3_WEIGHT(rectangle3_weights[436]), .FEAT_THRES(feature_thresholds[436]), .FEAT_ABOVE(feature_aboves[436]), .FEAT_BELOW(feature_belows[436])) ac436(.scan_win(scan_win436), .scan_win_std_dev(scan_win_std_dev[436]), .feature_accum(feature_accums[436]));
  accum_calculator #(.RECT1_X(rectangle1_xs[437]), .RECT1_Y(rectangle1_ys[437]), .RECT1_WIDTH(rectangle1_widths[437]), .RECT1_HEIGHT(rectangle1_heights[437]), .RECT1_WEIGHT(rectangle1_weights[437]), .RECT2_X(rectangle2_xs[437]), .RECT2_Y(rectangle2_ys[437]), .RECT2_WIDTH(rectangle2_widths[437]), .RECT2_HEIGHT(rectangle2_heights[437]), .RECT2_WEIGHT(rectangle2_weights[437]), .RECT3_X(rectangle3_xs[437]), .RECT3_Y(rectangle3_ys[437]), .RECT3_WIDTH(rectangle3_widths[437]), .RECT3_HEIGHT(rectangle3_heights[437]), .RECT3_WEIGHT(rectangle3_weights[437]), .FEAT_THRES(feature_thresholds[437]), .FEAT_ABOVE(feature_aboves[437]), .FEAT_BELOW(feature_belows[437])) ac437(.scan_win(scan_win437), .scan_win_std_dev(scan_win_std_dev[437]), .feature_accum(feature_accums[437]));
  accum_calculator #(.RECT1_X(rectangle1_xs[438]), .RECT1_Y(rectangle1_ys[438]), .RECT1_WIDTH(rectangle1_widths[438]), .RECT1_HEIGHT(rectangle1_heights[438]), .RECT1_WEIGHT(rectangle1_weights[438]), .RECT2_X(rectangle2_xs[438]), .RECT2_Y(rectangle2_ys[438]), .RECT2_WIDTH(rectangle2_widths[438]), .RECT2_HEIGHT(rectangle2_heights[438]), .RECT2_WEIGHT(rectangle2_weights[438]), .RECT3_X(rectangle3_xs[438]), .RECT3_Y(rectangle3_ys[438]), .RECT3_WIDTH(rectangle3_widths[438]), .RECT3_HEIGHT(rectangle3_heights[438]), .RECT3_WEIGHT(rectangle3_weights[438]), .FEAT_THRES(feature_thresholds[438]), .FEAT_ABOVE(feature_aboves[438]), .FEAT_BELOW(feature_belows[438])) ac438(.scan_win(scan_win438), .scan_win_std_dev(scan_win_std_dev[438]), .feature_accum(feature_accums[438]));
  accum_calculator #(.RECT1_X(rectangle1_xs[439]), .RECT1_Y(rectangle1_ys[439]), .RECT1_WIDTH(rectangle1_widths[439]), .RECT1_HEIGHT(rectangle1_heights[439]), .RECT1_WEIGHT(rectangle1_weights[439]), .RECT2_X(rectangle2_xs[439]), .RECT2_Y(rectangle2_ys[439]), .RECT2_WIDTH(rectangle2_widths[439]), .RECT2_HEIGHT(rectangle2_heights[439]), .RECT2_WEIGHT(rectangle2_weights[439]), .RECT3_X(rectangle3_xs[439]), .RECT3_Y(rectangle3_ys[439]), .RECT3_WIDTH(rectangle3_widths[439]), .RECT3_HEIGHT(rectangle3_heights[439]), .RECT3_WEIGHT(rectangle3_weights[439]), .FEAT_THRES(feature_thresholds[439]), .FEAT_ABOVE(feature_aboves[439]), .FEAT_BELOW(feature_belows[439])) ac439(.scan_win(scan_win439), .scan_win_std_dev(scan_win_std_dev[439]), .feature_accum(feature_accums[439]));
  accum_calculator #(.RECT1_X(rectangle1_xs[440]), .RECT1_Y(rectangle1_ys[440]), .RECT1_WIDTH(rectangle1_widths[440]), .RECT1_HEIGHT(rectangle1_heights[440]), .RECT1_WEIGHT(rectangle1_weights[440]), .RECT2_X(rectangle2_xs[440]), .RECT2_Y(rectangle2_ys[440]), .RECT2_WIDTH(rectangle2_widths[440]), .RECT2_HEIGHT(rectangle2_heights[440]), .RECT2_WEIGHT(rectangle2_weights[440]), .RECT3_X(rectangle3_xs[440]), .RECT3_Y(rectangle3_ys[440]), .RECT3_WIDTH(rectangle3_widths[440]), .RECT3_HEIGHT(rectangle3_heights[440]), .RECT3_WEIGHT(rectangle3_weights[440]), .FEAT_THRES(feature_thresholds[440]), .FEAT_ABOVE(feature_aboves[440]), .FEAT_BELOW(feature_belows[440])) ac440(.scan_win(scan_win440), .scan_win_std_dev(scan_win_std_dev[440]), .feature_accum(feature_accums[440]));
  accum_calculator #(.RECT1_X(rectangle1_xs[441]), .RECT1_Y(rectangle1_ys[441]), .RECT1_WIDTH(rectangle1_widths[441]), .RECT1_HEIGHT(rectangle1_heights[441]), .RECT1_WEIGHT(rectangle1_weights[441]), .RECT2_X(rectangle2_xs[441]), .RECT2_Y(rectangle2_ys[441]), .RECT2_WIDTH(rectangle2_widths[441]), .RECT2_HEIGHT(rectangle2_heights[441]), .RECT2_WEIGHT(rectangle2_weights[441]), .RECT3_X(rectangle3_xs[441]), .RECT3_Y(rectangle3_ys[441]), .RECT3_WIDTH(rectangle3_widths[441]), .RECT3_HEIGHT(rectangle3_heights[441]), .RECT3_WEIGHT(rectangle3_weights[441]), .FEAT_THRES(feature_thresholds[441]), .FEAT_ABOVE(feature_aboves[441]), .FEAT_BELOW(feature_belows[441])) ac441(.scan_win(scan_win441), .scan_win_std_dev(scan_win_std_dev[441]), .feature_accum(feature_accums[441]));
  accum_calculator #(.RECT1_X(rectangle1_xs[442]), .RECT1_Y(rectangle1_ys[442]), .RECT1_WIDTH(rectangle1_widths[442]), .RECT1_HEIGHT(rectangle1_heights[442]), .RECT1_WEIGHT(rectangle1_weights[442]), .RECT2_X(rectangle2_xs[442]), .RECT2_Y(rectangle2_ys[442]), .RECT2_WIDTH(rectangle2_widths[442]), .RECT2_HEIGHT(rectangle2_heights[442]), .RECT2_WEIGHT(rectangle2_weights[442]), .RECT3_X(rectangle3_xs[442]), .RECT3_Y(rectangle3_ys[442]), .RECT3_WIDTH(rectangle3_widths[442]), .RECT3_HEIGHT(rectangle3_heights[442]), .RECT3_WEIGHT(rectangle3_weights[442]), .FEAT_THRES(feature_thresholds[442]), .FEAT_ABOVE(feature_aboves[442]), .FEAT_BELOW(feature_belows[442])) ac442(.scan_win(scan_win442), .scan_win_std_dev(scan_win_std_dev[442]), .feature_accum(feature_accums[442]));
  accum_calculator #(.RECT1_X(rectangle1_xs[443]), .RECT1_Y(rectangle1_ys[443]), .RECT1_WIDTH(rectangle1_widths[443]), .RECT1_HEIGHT(rectangle1_heights[443]), .RECT1_WEIGHT(rectangle1_weights[443]), .RECT2_X(rectangle2_xs[443]), .RECT2_Y(rectangle2_ys[443]), .RECT2_WIDTH(rectangle2_widths[443]), .RECT2_HEIGHT(rectangle2_heights[443]), .RECT2_WEIGHT(rectangle2_weights[443]), .RECT3_X(rectangle3_xs[443]), .RECT3_Y(rectangle3_ys[443]), .RECT3_WIDTH(rectangle3_widths[443]), .RECT3_HEIGHT(rectangle3_heights[443]), .RECT3_WEIGHT(rectangle3_weights[443]), .FEAT_THRES(feature_thresholds[443]), .FEAT_ABOVE(feature_aboves[443]), .FEAT_BELOW(feature_belows[443])) ac443(.scan_win(scan_win443), .scan_win_std_dev(scan_win_std_dev[443]), .feature_accum(feature_accums[443]));
  accum_calculator #(.RECT1_X(rectangle1_xs[444]), .RECT1_Y(rectangle1_ys[444]), .RECT1_WIDTH(rectangle1_widths[444]), .RECT1_HEIGHT(rectangle1_heights[444]), .RECT1_WEIGHT(rectangle1_weights[444]), .RECT2_X(rectangle2_xs[444]), .RECT2_Y(rectangle2_ys[444]), .RECT2_WIDTH(rectangle2_widths[444]), .RECT2_HEIGHT(rectangle2_heights[444]), .RECT2_WEIGHT(rectangle2_weights[444]), .RECT3_X(rectangle3_xs[444]), .RECT3_Y(rectangle3_ys[444]), .RECT3_WIDTH(rectangle3_widths[444]), .RECT3_HEIGHT(rectangle3_heights[444]), .RECT3_WEIGHT(rectangle3_weights[444]), .FEAT_THRES(feature_thresholds[444]), .FEAT_ABOVE(feature_aboves[444]), .FEAT_BELOW(feature_belows[444])) ac444(.scan_win(scan_win444), .scan_win_std_dev(scan_win_std_dev[444]), .feature_accum(feature_accums[444]));
  accum_calculator #(.RECT1_X(rectangle1_xs[445]), .RECT1_Y(rectangle1_ys[445]), .RECT1_WIDTH(rectangle1_widths[445]), .RECT1_HEIGHT(rectangle1_heights[445]), .RECT1_WEIGHT(rectangle1_weights[445]), .RECT2_X(rectangle2_xs[445]), .RECT2_Y(rectangle2_ys[445]), .RECT2_WIDTH(rectangle2_widths[445]), .RECT2_HEIGHT(rectangle2_heights[445]), .RECT2_WEIGHT(rectangle2_weights[445]), .RECT3_X(rectangle3_xs[445]), .RECT3_Y(rectangle3_ys[445]), .RECT3_WIDTH(rectangle3_widths[445]), .RECT3_HEIGHT(rectangle3_heights[445]), .RECT3_WEIGHT(rectangle3_weights[445]), .FEAT_THRES(feature_thresholds[445]), .FEAT_ABOVE(feature_aboves[445]), .FEAT_BELOW(feature_belows[445])) ac445(.scan_win(scan_win445), .scan_win_std_dev(scan_win_std_dev[445]), .feature_accum(feature_accums[445]));
  accum_calculator #(.RECT1_X(rectangle1_xs[446]), .RECT1_Y(rectangle1_ys[446]), .RECT1_WIDTH(rectangle1_widths[446]), .RECT1_HEIGHT(rectangle1_heights[446]), .RECT1_WEIGHT(rectangle1_weights[446]), .RECT2_X(rectangle2_xs[446]), .RECT2_Y(rectangle2_ys[446]), .RECT2_WIDTH(rectangle2_widths[446]), .RECT2_HEIGHT(rectangle2_heights[446]), .RECT2_WEIGHT(rectangle2_weights[446]), .RECT3_X(rectangle3_xs[446]), .RECT3_Y(rectangle3_ys[446]), .RECT3_WIDTH(rectangle3_widths[446]), .RECT3_HEIGHT(rectangle3_heights[446]), .RECT3_WEIGHT(rectangle3_weights[446]), .FEAT_THRES(feature_thresholds[446]), .FEAT_ABOVE(feature_aboves[446]), .FEAT_BELOW(feature_belows[446])) ac446(.scan_win(scan_win446), .scan_win_std_dev(scan_win_std_dev[446]), .feature_accum(feature_accums[446]));
  accum_calculator #(.RECT1_X(rectangle1_xs[447]), .RECT1_Y(rectangle1_ys[447]), .RECT1_WIDTH(rectangle1_widths[447]), .RECT1_HEIGHT(rectangle1_heights[447]), .RECT1_WEIGHT(rectangle1_weights[447]), .RECT2_X(rectangle2_xs[447]), .RECT2_Y(rectangle2_ys[447]), .RECT2_WIDTH(rectangle2_widths[447]), .RECT2_HEIGHT(rectangle2_heights[447]), .RECT2_WEIGHT(rectangle2_weights[447]), .RECT3_X(rectangle3_xs[447]), .RECT3_Y(rectangle3_ys[447]), .RECT3_WIDTH(rectangle3_widths[447]), .RECT3_HEIGHT(rectangle3_heights[447]), .RECT3_WEIGHT(rectangle3_weights[447]), .FEAT_THRES(feature_thresholds[447]), .FEAT_ABOVE(feature_aboves[447]), .FEAT_BELOW(feature_belows[447])) ac447(.scan_win(scan_win447), .scan_win_std_dev(scan_win_std_dev[447]), .feature_accum(feature_accums[447]));
  accum_calculator #(.RECT1_X(rectangle1_xs[448]), .RECT1_Y(rectangle1_ys[448]), .RECT1_WIDTH(rectangle1_widths[448]), .RECT1_HEIGHT(rectangle1_heights[448]), .RECT1_WEIGHT(rectangle1_weights[448]), .RECT2_X(rectangle2_xs[448]), .RECT2_Y(rectangle2_ys[448]), .RECT2_WIDTH(rectangle2_widths[448]), .RECT2_HEIGHT(rectangle2_heights[448]), .RECT2_WEIGHT(rectangle2_weights[448]), .RECT3_X(rectangle3_xs[448]), .RECT3_Y(rectangle3_ys[448]), .RECT3_WIDTH(rectangle3_widths[448]), .RECT3_HEIGHT(rectangle3_heights[448]), .RECT3_WEIGHT(rectangle3_weights[448]), .FEAT_THRES(feature_thresholds[448]), .FEAT_ABOVE(feature_aboves[448]), .FEAT_BELOW(feature_belows[448])) ac448(.scan_win(scan_win448), .scan_win_std_dev(scan_win_std_dev[448]), .feature_accum(feature_accums[448]));
  accum_calculator #(.RECT1_X(rectangle1_xs[449]), .RECT1_Y(rectangle1_ys[449]), .RECT1_WIDTH(rectangle1_widths[449]), .RECT1_HEIGHT(rectangle1_heights[449]), .RECT1_WEIGHT(rectangle1_weights[449]), .RECT2_X(rectangle2_xs[449]), .RECT2_Y(rectangle2_ys[449]), .RECT2_WIDTH(rectangle2_widths[449]), .RECT2_HEIGHT(rectangle2_heights[449]), .RECT2_WEIGHT(rectangle2_weights[449]), .RECT3_X(rectangle3_xs[449]), .RECT3_Y(rectangle3_ys[449]), .RECT3_WIDTH(rectangle3_widths[449]), .RECT3_HEIGHT(rectangle3_heights[449]), .RECT3_WEIGHT(rectangle3_weights[449]), .FEAT_THRES(feature_thresholds[449]), .FEAT_ABOVE(feature_aboves[449]), .FEAT_BELOW(feature_belows[449])) ac449(.scan_win(scan_win449), .scan_win_std_dev(scan_win_std_dev[449]), .feature_accum(feature_accums[449]));
  accum_calculator #(.RECT1_X(rectangle1_xs[450]), .RECT1_Y(rectangle1_ys[450]), .RECT1_WIDTH(rectangle1_widths[450]), .RECT1_HEIGHT(rectangle1_heights[450]), .RECT1_WEIGHT(rectangle1_weights[450]), .RECT2_X(rectangle2_xs[450]), .RECT2_Y(rectangle2_ys[450]), .RECT2_WIDTH(rectangle2_widths[450]), .RECT2_HEIGHT(rectangle2_heights[450]), .RECT2_WEIGHT(rectangle2_weights[450]), .RECT3_X(rectangle3_xs[450]), .RECT3_Y(rectangle3_ys[450]), .RECT3_WIDTH(rectangle3_widths[450]), .RECT3_HEIGHT(rectangle3_heights[450]), .RECT3_WEIGHT(rectangle3_weights[450]), .FEAT_THRES(feature_thresholds[450]), .FEAT_ABOVE(feature_aboves[450]), .FEAT_BELOW(feature_belows[450])) ac450(.scan_win(scan_win450), .scan_win_std_dev(scan_win_std_dev[450]), .feature_accum(feature_accums[450]));
  accum_calculator #(.RECT1_X(rectangle1_xs[451]), .RECT1_Y(rectangle1_ys[451]), .RECT1_WIDTH(rectangle1_widths[451]), .RECT1_HEIGHT(rectangle1_heights[451]), .RECT1_WEIGHT(rectangle1_weights[451]), .RECT2_X(rectangle2_xs[451]), .RECT2_Y(rectangle2_ys[451]), .RECT2_WIDTH(rectangle2_widths[451]), .RECT2_HEIGHT(rectangle2_heights[451]), .RECT2_WEIGHT(rectangle2_weights[451]), .RECT3_X(rectangle3_xs[451]), .RECT3_Y(rectangle3_ys[451]), .RECT3_WIDTH(rectangle3_widths[451]), .RECT3_HEIGHT(rectangle3_heights[451]), .RECT3_WEIGHT(rectangle3_weights[451]), .FEAT_THRES(feature_thresholds[451]), .FEAT_ABOVE(feature_aboves[451]), .FEAT_BELOW(feature_belows[451])) ac451(.scan_win(scan_win451), .scan_win_std_dev(scan_win_std_dev[451]), .feature_accum(feature_accums[451]));
  accum_calculator #(.RECT1_X(rectangle1_xs[452]), .RECT1_Y(rectangle1_ys[452]), .RECT1_WIDTH(rectangle1_widths[452]), .RECT1_HEIGHT(rectangle1_heights[452]), .RECT1_WEIGHT(rectangle1_weights[452]), .RECT2_X(rectangle2_xs[452]), .RECT2_Y(rectangle2_ys[452]), .RECT2_WIDTH(rectangle2_widths[452]), .RECT2_HEIGHT(rectangle2_heights[452]), .RECT2_WEIGHT(rectangle2_weights[452]), .RECT3_X(rectangle3_xs[452]), .RECT3_Y(rectangle3_ys[452]), .RECT3_WIDTH(rectangle3_widths[452]), .RECT3_HEIGHT(rectangle3_heights[452]), .RECT3_WEIGHT(rectangle3_weights[452]), .FEAT_THRES(feature_thresholds[452]), .FEAT_ABOVE(feature_aboves[452]), .FEAT_BELOW(feature_belows[452])) ac452(.scan_win(scan_win452), .scan_win_std_dev(scan_win_std_dev[452]), .feature_accum(feature_accums[452]));
  accum_calculator #(.RECT1_X(rectangle1_xs[453]), .RECT1_Y(rectangle1_ys[453]), .RECT1_WIDTH(rectangle1_widths[453]), .RECT1_HEIGHT(rectangle1_heights[453]), .RECT1_WEIGHT(rectangle1_weights[453]), .RECT2_X(rectangle2_xs[453]), .RECT2_Y(rectangle2_ys[453]), .RECT2_WIDTH(rectangle2_widths[453]), .RECT2_HEIGHT(rectangle2_heights[453]), .RECT2_WEIGHT(rectangle2_weights[453]), .RECT3_X(rectangle3_xs[453]), .RECT3_Y(rectangle3_ys[453]), .RECT3_WIDTH(rectangle3_widths[453]), .RECT3_HEIGHT(rectangle3_heights[453]), .RECT3_WEIGHT(rectangle3_weights[453]), .FEAT_THRES(feature_thresholds[453]), .FEAT_ABOVE(feature_aboves[453]), .FEAT_BELOW(feature_belows[453])) ac453(.scan_win(scan_win453), .scan_win_std_dev(scan_win_std_dev[453]), .feature_accum(feature_accums[453]));
  accum_calculator #(.RECT1_X(rectangle1_xs[454]), .RECT1_Y(rectangle1_ys[454]), .RECT1_WIDTH(rectangle1_widths[454]), .RECT1_HEIGHT(rectangle1_heights[454]), .RECT1_WEIGHT(rectangle1_weights[454]), .RECT2_X(rectangle2_xs[454]), .RECT2_Y(rectangle2_ys[454]), .RECT2_WIDTH(rectangle2_widths[454]), .RECT2_HEIGHT(rectangle2_heights[454]), .RECT2_WEIGHT(rectangle2_weights[454]), .RECT3_X(rectangle3_xs[454]), .RECT3_Y(rectangle3_ys[454]), .RECT3_WIDTH(rectangle3_widths[454]), .RECT3_HEIGHT(rectangle3_heights[454]), .RECT3_WEIGHT(rectangle3_weights[454]), .FEAT_THRES(feature_thresholds[454]), .FEAT_ABOVE(feature_aboves[454]), .FEAT_BELOW(feature_belows[454])) ac454(.scan_win(scan_win454), .scan_win_std_dev(scan_win_std_dev[454]), .feature_accum(feature_accums[454]));
  accum_calculator #(.RECT1_X(rectangle1_xs[455]), .RECT1_Y(rectangle1_ys[455]), .RECT1_WIDTH(rectangle1_widths[455]), .RECT1_HEIGHT(rectangle1_heights[455]), .RECT1_WEIGHT(rectangle1_weights[455]), .RECT2_X(rectangle2_xs[455]), .RECT2_Y(rectangle2_ys[455]), .RECT2_WIDTH(rectangle2_widths[455]), .RECT2_HEIGHT(rectangle2_heights[455]), .RECT2_WEIGHT(rectangle2_weights[455]), .RECT3_X(rectangle3_xs[455]), .RECT3_Y(rectangle3_ys[455]), .RECT3_WIDTH(rectangle3_widths[455]), .RECT3_HEIGHT(rectangle3_heights[455]), .RECT3_WEIGHT(rectangle3_weights[455]), .FEAT_THRES(feature_thresholds[455]), .FEAT_ABOVE(feature_aboves[455]), .FEAT_BELOW(feature_belows[455])) ac455(.scan_win(scan_win455), .scan_win_std_dev(scan_win_std_dev[455]), .feature_accum(feature_accums[455]));
  accum_calculator #(.RECT1_X(rectangle1_xs[456]), .RECT1_Y(rectangle1_ys[456]), .RECT1_WIDTH(rectangle1_widths[456]), .RECT1_HEIGHT(rectangle1_heights[456]), .RECT1_WEIGHT(rectangle1_weights[456]), .RECT2_X(rectangle2_xs[456]), .RECT2_Y(rectangle2_ys[456]), .RECT2_WIDTH(rectangle2_widths[456]), .RECT2_HEIGHT(rectangle2_heights[456]), .RECT2_WEIGHT(rectangle2_weights[456]), .RECT3_X(rectangle3_xs[456]), .RECT3_Y(rectangle3_ys[456]), .RECT3_WIDTH(rectangle3_widths[456]), .RECT3_HEIGHT(rectangle3_heights[456]), .RECT3_WEIGHT(rectangle3_weights[456]), .FEAT_THRES(feature_thresholds[456]), .FEAT_ABOVE(feature_aboves[456]), .FEAT_BELOW(feature_belows[456])) ac456(.scan_win(scan_win456), .scan_win_std_dev(scan_win_std_dev[456]), .feature_accum(feature_accums[456]));
  accum_calculator #(.RECT1_X(rectangle1_xs[457]), .RECT1_Y(rectangle1_ys[457]), .RECT1_WIDTH(rectangle1_widths[457]), .RECT1_HEIGHT(rectangle1_heights[457]), .RECT1_WEIGHT(rectangle1_weights[457]), .RECT2_X(rectangle2_xs[457]), .RECT2_Y(rectangle2_ys[457]), .RECT2_WIDTH(rectangle2_widths[457]), .RECT2_HEIGHT(rectangle2_heights[457]), .RECT2_WEIGHT(rectangle2_weights[457]), .RECT3_X(rectangle3_xs[457]), .RECT3_Y(rectangle3_ys[457]), .RECT3_WIDTH(rectangle3_widths[457]), .RECT3_HEIGHT(rectangle3_heights[457]), .RECT3_WEIGHT(rectangle3_weights[457]), .FEAT_THRES(feature_thresholds[457]), .FEAT_ABOVE(feature_aboves[457]), .FEAT_BELOW(feature_belows[457])) ac457(.scan_win(scan_win457), .scan_win_std_dev(scan_win_std_dev[457]), .feature_accum(feature_accums[457]));
  accum_calculator #(.RECT1_X(rectangle1_xs[458]), .RECT1_Y(rectangle1_ys[458]), .RECT1_WIDTH(rectangle1_widths[458]), .RECT1_HEIGHT(rectangle1_heights[458]), .RECT1_WEIGHT(rectangle1_weights[458]), .RECT2_X(rectangle2_xs[458]), .RECT2_Y(rectangle2_ys[458]), .RECT2_WIDTH(rectangle2_widths[458]), .RECT2_HEIGHT(rectangle2_heights[458]), .RECT2_WEIGHT(rectangle2_weights[458]), .RECT3_X(rectangle3_xs[458]), .RECT3_Y(rectangle3_ys[458]), .RECT3_WIDTH(rectangle3_widths[458]), .RECT3_HEIGHT(rectangle3_heights[458]), .RECT3_WEIGHT(rectangle3_weights[458]), .FEAT_THRES(feature_thresholds[458]), .FEAT_ABOVE(feature_aboves[458]), .FEAT_BELOW(feature_belows[458])) ac458(.scan_win(scan_win458), .scan_win_std_dev(scan_win_std_dev[458]), .feature_accum(feature_accums[458]));
  accum_calculator #(.RECT1_X(rectangle1_xs[459]), .RECT1_Y(rectangle1_ys[459]), .RECT1_WIDTH(rectangle1_widths[459]), .RECT1_HEIGHT(rectangle1_heights[459]), .RECT1_WEIGHT(rectangle1_weights[459]), .RECT2_X(rectangle2_xs[459]), .RECT2_Y(rectangle2_ys[459]), .RECT2_WIDTH(rectangle2_widths[459]), .RECT2_HEIGHT(rectangle2_heights[459]), .RECT2_WEIGHT(rectangle2_weights[459]), .RECT3_X(rectangle3_xs[459]), .RECT3_Y(rectangle3_ys[459]), .RECT3_WIDTH(rectangle3_widths[459]), .RECT3_HEIGHT(rectangle3_heights[459]), .RECT3_WEIGHT(rectangle3_weights[459]), .FEAT_THRES(feature_thresholds[459]), .FEAT_ABOVE(feature_aboves[459]), .FEAT_BELOW(feature_belows[459])) ac459(.scan_win(scan_win459), .scan_win_std_dev(scan_win_std_dev[459]), .feature_accum(feature_accums[459]));
  accum_calculator #(.RECT1_X(rectangle1_xs[460]), .RECT1_Y(rectangle1_ys[460]), .RECT1_WIDTH(rectangle1_widths[460]), .RECT1_HEIGHT(rectangle1_heights[460]), .RECT1_WEIGHT(rectangle1_weights[460]), .RECT2_X(rectangle2_xs[460]), .RECT2_Y(rectangle2_ys[460]), .RECT2_WIDTH(rectangle2_widths[460]), .RECT2_HEIGHT(rectangle2_heights[460]), .RECT2_WEIGHT(rectangle2_weights[460]), .RECT3_X(rectangle3_xs[460]), .RECT3_Y(rectangle3_ys[460]), .RECT3_WIDTH(rectangle3_widths[460]), .RECT3_HEIGHT(rectangle3_heights[460]), .RECT3_WEIGHT(rectangle3_weights[460]), .FEAT_THRES(feature_thresholds[460]), .FEAT_ABOVE(feature_aboves[460]), .FEAT_BELOW(feature_belows[460])) ac460(.scan_win(scan_win460), .scan_win_std_dev(scan_win_std_dev[460]), .feature_accum(feature_accums[460]));
  accum_calculator #(.RECT1_X(rectangle1_xs[461]), .RECT1_Y(rectangle1_ys[461]), .RECT1_WIDTH(rectangle1_widths[461]), .RECT1_HEIGHT(rectangle1_heights[461]), .RECT1_WEIGHT(rectangle1_weights[461]), .RECT2_X(rectangle2_xs[461]), .RECT2_Y(rectangle2_ys[461]), .RECT2_WIDTH(rectangle2_widths[461]), .RECT2_HEIGHT(rectangle2_heights[461]), .RECT2_WEIGHT(rectangle2_weights[461]), .RECT3_X(rectangle3_xs[461]), .RECT3_Y(rectangle3_ys[461]), .RECT3_WIDTH(rectangle3_widths[461]), .RECT3_HEIGHT(rectangle3_heights[461]), .RECT3_WEIGHT(rectangle3_weights[461]), .FEAT_THRES(feature_thresholds[461]), .FEAT_ABOVE(feature_aboves[461]), .FEAT_BELOW(feature_belows[461])) ac461(.scan_win(scan_win461), .scan_win_std_dev(scan_win_std_dev[461]), .feature_accum(feature_accums[461]));
  accum_calculator #(.RECT1_X(rectangle1_xs[462]), .RECT1_Y(rectangle1_ys[462]), .RECT1_WIDTH(rectangle1_widths[462]), .RECT1_HEIGHT(rectangle1_heights[462]), .RECT1_WEIGHT(rectangle1_weights[462]), .RECT2_X(rectangle2_xs[462]), .RECT2_Y(rectangle2_ys[462]), .RECT2_WIDTH(rectangle2_widths[462]), .RECT2_HEIGHT(rectangle2_heights[462]), .RECT2_WEIGHT(rectangle2_weights[462]), .RECT3_X(rectangle3_xs[462]), .RECT3_Y(rectangle3_ys[462]), .RECT3_WIDTH(rectangle3_widths[462]), .RECT3_HEIGHT(rectangle3_heights[462]), .RECT3_WEIGHT(rectangle3_weights[462]), .FEAT_THRES(feature_thresholds[462]), .FEAT_ABOVE(feature_aboves[462]), .FEAT_BELOW(feature_belows[462])) ac462(.scan_win(scan_win462), .scan_win_std_dev(scan_win_std_dev[462]), .feature_accum(feature_accums[462]));
  accum_calculator #(.RECT1_X(rectangle1_xs[463]), .RECT1_Y(rectangle1_ys[463]), .RECT1_WIDTH(rectangle1_widths[463]), .RECT1_HEIGHT(rectangle1_heights[463]), .RECT1_WEIGHT(rectangle1_weights[463]), .RECT2_X(rectangle2_xs[463]), .RECT2_Y(rectangle2_ys[463]), .RECT2_WIDTH(rectangle2_widths[463]), .RECT2_HEIGHT(rectangle2_heights[463]), .RECT2_WEIGHT(rectangle2_weights[463]), .RECT3_X(rectangle3_xs[463]), .RECT3_Y(rectangle3_ys[463]), .RECT3_WIDTH(rectangle3_widths[463]), .RECT3_HEIGHT(rectangle3_heights[463]), .RECT3_WEIGHT(rectangle3_weights[463]), .FEAT_THRES(feature_thresholds[463]), .FEAT_ABOVE(feature_aboves[463]), .FEAT_BELOW(feature_belows[463])) ac463(.scan_win(scan_win463), .scan_win_std_dev(scan_win_std_dev[463]), .feature_accum(feature_accums[463]));
  accum_calculator #(.RECT1_X(rectangle1_xs[464]), .RECT1_Y(rectangle1_ys[464]), .RECT1_WIDTH(rectangle1_widths[464]), .RECT1_HEIGHT(rectangle1_heights[464]), .RECT1_WEIGHT(rectangle1_weights[464]), .RECT2_X(rectangle2_xs[464]), .RECT2_Y(rectangle2_ys[464]), .RECT2_WIDTH(rectangle2_widths[464]), .RECT2_HEIGHT(rectangle2_heights[464]), .RECT2_WEIGHT(rectangle2_weights[464]), .RECT3_X(rectangle3_xs[464]), .RECT3_Y(rectangle3_ys[464]), .RECT3_WIDTH(rectangle3_widths[464]), .RECT3_HEIGHT(rectangle3_heights[464]), .RECT3_WEIGHT(rectangle3_weights[464]), .FEAT_THRES(feature_thresholds[464]), .FEAT_ABOVE(feature_aboves[464]), .FEAT_BELOW(feature_belows[464])) ac464(.scan_win(scan_win464), .scan_win_std_dev(scan_win_std_dev[464]), .feature_accum(feature_accums[464]));
  accum_calculator #(.RECT1_X(rectangle1_xs[465]), .RECT1_Y(rectangle1_ys[465]), .RECT1_WIDTH(rectangle1_widths[465]), .RECT1_HEIGHT(rectangle1_heights[465]), .RECT1_WEIGHT(rectangle1_weights[465]), .RECT2_X(rectangle2_xs[465]), .RECT2_Y(rectangle2_ys[465]), .RECT2_WIDTH(rectangle2_widths[465]), .RECT2_HEIGHT(rectangle2_heights[465]), .RECT2_WEIGHT(rectangle2_weights[465]), .RECT3_X(rectangle3_xs[465]), .RECT3_Y(rectangle3_ys[465]), .RECT3_WIDTH(rectangle3_widths[465]), .RECT3_HEIGHT(rectangle3_heights[465]), .RECT3_WEIGHT(rectangle3_weights[465]), .FEAT_THRES(feature_thresholds[465]), .FEAT_ABOVE(feature_aboves[465]), .FEAT_BELOW(feature_belows[465])) ac465(.scan_win(scan_win465), .scan_win_std_dev(scan_win_std_dev[465]), .feature_accum(feature_accums[465]));
  accum_calculator #(.RECT1_X(rectangle1_xs[466]), .RECT1_Y(rectangle1_ys[466]), .RECT1_WIDTH(rectangle1_widths[466]), .RECT1_HEIGHT(rectangle1_heights[466]), .RECT1_WEIGHT(rectangle1_weights[466]), .RECT2_X(rectangle2_xs[466]), .RECT2_Y(rectangle2_ys[466]), .RECT2_WIDTH(rectangle2_widths[466]), .RECT2_HEIGHT(rectangle2_heights[466]), .RECT2_WEIGHT(rectangle2_weights[466]), .RECT3_X(rectangle3_xs[466]), .RECT3_Y(rectangle3_ys[466]), .RECT3_WIDTH(rectangle3_widths[466]), .RECT3_HEIGHT(rectangle3_heights[466]), .RECT3_WEIGHT(rectangle3_weights[466]), .FEAT_THRES(feature_thresholds[466]), .FEAT_ABOVE(feature_aboves[466]), .FEAT_BELOW(feature_belows[466])) ac466(.scan_win(scan_win466), .scan_win_std_dev(scan_win_std_dev[466]), .feature_accum(feature_accums[466]));
  accum_calculator #(.RECT1_X(rectangle1_xs[467]), .RECT1_Y(rectangle1_ys[467]), .RECT1_WIDTH(rectangle1_widths[467]), .RECT1_HEIGHT(rectangle1_heights[467]), .RECT1_WEIGHT(rectangle1_weights[467]), .RECT2_X(rectangle2_xs[467]), .RECT2_Y(rectangle2_ys[467]), .RECT2_WIDTH(rectangle2_widths[467]), .RECT2_HEIGHT(rectangle2_heights[467]), .RECT2_WEIGHT(rectangle2_weights[467]), .RECT3_X(rectangle3_xs[467]), .RECT3_Y(rectangle3_ys[467]), .RECT3_WIDTH(rectangle3_widths[467]), .RECT3_HEIGHT(rectangle3_heights[467]), .RECT3_WEIGHT(rectangle3_weights[467]), .FEAT_THRES(feature_thresholds[467]), .FEAT_ABOVE(feature_aboves[467]), .FEAT_BELOW(feature_belows[467])) ac467(.scan_win(scan_win467), .scan_win_std_dev(scan_win_std_dev[467]), .feature_accum(feature_accums[467]));
  accum_calculator #(.RECT1_X(rectangle1_xs[468]), .RECT1_Y(rectangle1_ys[468]), .RECT1_WIDTH(rectangle1_widths[468]), .RECT1_HEIGHT(rectangle1_heights[468]), .RECT1_WEIGHT(rectangle1_weights[468]), .RECT2_X(rectangle2_xs[468]), .RECT2_Y(rectangle2_ys[468]), .RECT2_WIDTH(rectangle2_widths[468]), .RECT2_HEIGHT(rectangle2_heights[468]), .RECT2_WEIGHT(rectangle2_weights[468]), .RECT3_X(rectangle3_xs[468]), .RECT3_Y(rectangle3_ys[468]), .RECT3_WIDTH(rectangle3_widths[468]), .RECT3_HEIGHT(rectangle3_heights[468]), .RECT3_WEIGHT(rectangle3_weights[468]), .FEAT_THRES(feature_thresholds[468]), .FEAT_ABOVE(feature_aboves[468]), .FEAT_BELOW(feature_belows[468])) ac468(.scan_win(scan_win468), .scan_win_std_dev(scan_win_std_dev[468]), .feature_accum(feature_accums[468]));
  accum_calculator #(.RECT1_X(rectangle1_xs[469]), .RECT1_Y(rectangle1_ys[469]), .RECT1_WIDTH(rectangle1_widths[469]), .RECT1_HEIGHT(rectangle1_heights[469]), .RECT1_WEIGHT(rectangle1_weights[469]), .RECT2_X(rectangle2_xs[469]), .RECT2_Y(rectangle2_ys[469]), .RECT2_WIDTH(rectangle2_widths[469]), .RECT2_HEIGHT(rectangle2_heights[469]), .RECT2_WEIGHT(rectangle2_weights[469]), .RECT3_X(rectangle3_xs[469]), .RECT3_Y(rectangle3_ys[469]), .RECT3_WIDTH(rectangle3_widths[469]), .RECT3_HEIGHT(rectangle3_heights[469]), .RECT3_WEIGHT(rectangle3_weights[469]), .FEAT_THRES(feature_thresholds[469]), .FEAT_ABOVE(feature_aboves[469]), .FEAT_BELOW(feature_belows[469])) ac469(.scan_win(scan_win469), .scan_win_std_dev(scan_win_std_dev[469]), .feature_accum(feature_accums[469]));
  accum_calculator #(.RECT1_X(rectangle1_xs[470]), .RECT1_Y(rectangle1_ys[470]), .RECT1_WIDTH(rectangle1_widths[470]), .RECT1_HEIGHT(rectangle1_heights[470]), .RECT1_WEIGHT(rectangle1_weights[470]), .RECT2_X(rectangle2_xs[470]), .RECT2_Y(rectangle2_ys[470]), .RECT2_WIDTH(rectangle2_widths[470]), .RECT2_HEIGHT(rectangle2_heights[470]), .RECT2_WEIGHT(rectangle2_weights[470]), .RECT3_X(rectangle3_xs[470]), .RECT3_Y(rectangle3_ys[470]), .RECT3_WIDTH(rectangle3_widths[470]), .RECT3_HEIGHT(rectangle3_heights[470]), .RECT3_WEIGHT(rectangle3_weights[470]), .FEAT_THRES(feature_thresholds[470]), .FEAT_ABOVE(feature_aboves[470]), .FEAT_BELOW(feature_belows[470])) ac470(.scan_win(scan_win470), .scan_win_std_dev(scan_win_std_dev[470]), .feature_accum(feature_accums[470]));
  accum_calculator #(.RECT1_X(rectangle1_xs[471]), .RECT1_Y(rectangle1_ys[471]), .RECT1_WIDTH(rectangle1_widths[471]), .RECT1_HEIGHT(rectangle1_heights[471]), .RECT1_WEIGHT(rectangle1_weights[471]), .RECT2_X(rectangle2_xs[471]), .RECT2_Y(rectangle2_ys[471]), .RECT2_WIDTH(rectangle2_widths[471]), .RECT2_HEIGHT(rectangle2_heights[471]), .RECT2_WEIGHT(rectangle2_weights[471]), .RECT3_X(rectangle3_xs[471]), .RECT3_Y(rectangle3_ys[471]), .RECT3_WIDTH(rectangle3_widths[471]), .RECT3_HEIGHT(rectangle3_heights[471]), .RECT3_WEIGHT(rectangle3_weights[471]), .FEAT_THRES(feature_thresholds[471]), .FEAT_ABOVE(feature_aboves[471]), .FEAT_BELOW(feature_belows[471])) ac471(.scan_win(scan_win471), .scan_win_std_dev(scan_win_std_dev[471]), .feature_accum(feature_accums[471]));
  accum_calculator #(.RECT1_X(rectangle1_xs[472]), .RECT1_Y(rectangle1_ys[472]), .RECT1_WIDTH(rectangle1_widths[472]), .RECT1_HEIGHT(rectangle1_heights[472]), .RECT1_WEIGHT(rectangle1_weights[472]), .RECT2_X(rectangle2_xs[472]), .RECT2_Y(rectangle2_ys[472]), .RECT2_WIDTH(rectangle2_widths[472]), .RECT2_HEIGHT(rectangle2_heights[472]), .RECT2_WEIGHT(rectangle2_weights[472]), .RECT3_X(rectangle3_xs[472]), .RECT3_Y(rectangle3_ys[472]), .RECT3_WIDTH(rectangle3_widths[472]), .RECT3_HEIGHT(rectangle3_heights[472]), .RECT3_WEIGHT(rectangle3_weights[472]), .FEAT_THRES(feature_thresholds[472]), .FEAT_ABOVE(feature_aboves[472]), .FEAT_BELOW(feature_belows[472])) ac472(.scan_win(scan_win472), .scan_win_std_dev(scan_win_std_dev[472]), .feature_accum(feature_accums[472]));
  accum_calculator #(.RECT1_X(rectangle1_xs[473]), .RECT1_Y(rectangle1_ys[473]), .RECT1_WIDTH(rectangle1_widths[473]), .RECT1_HEIGHT(rectangle1_heights[473]), .RECT1_WEIGHT(rectangle1_weights[473]), .RECT2_X(rectangle2_xs[473]), .RECT2_Y(rectangle2_ys[473]), .RECT2_WIDTH(rectangle2_widths[473]), .RECT2_HEIGHT(rectangle2_heights[473]), .RECT2_WEIGHT(rectangle2_weights[473]), .RECT3_X(rectangle3_xs[473]), .RECT3_Y(rectangle3_ys[473]), .RECT3_WIDTH(rectangle3_widths[473]), .RECT3_HEIGHT(rectangle3_heights[473]), .RECT3_WEIGHT(rectangle3_weights[473]), .FEAT_THRES(feature_thresholds[473]), .FEAT_ABOVE(feature_aboves[473]), .FEAT_BELOW(feature_belows[473])) ac473(.scan_win(scan_win473), .scan_win_std_dev(scan_win_std_dev[473]), .feature_accum(feature_accums[473]));
  accum_calculator #(.RECT1_X(rectangle1_xs[474]), .RECT1_Y(rectangle1_ys[474]), .RECT1_WIDTH(rectangle1_widths[474]), .RECT1_HEIGHT(rectangle1_heights[474]), .RECT1_WEIGHT(rectangle1_weights[474]), .RECT2_X(rectangle2_xs[474]), .RECT2_Y(rectangle2_ys[474]), .RECT2_WIDTH(rectangle2_widths[474]), .RECT2_HEIGHT(rectangle2_heights[474]), .RECT2_WEIGHT(rectangle2_weights[474]), .RECT3_X(rectangle3_xs[474]), .RECT3_Y(rectangle3_ys[474]), .RECT3_WIDTH(rectangle3_widths[474]), .RECT3_HEIGHT(rectangle3_heights[474]), .RECT3_WEIGHT(rectangle3_weights[474]), .FEAT_THRES(feature_thresholds[474]), .FEAT_ABOVE(feature_aboves[474]), .FEAT_BELOW(feature_belows[474])) ac474(.scan_win(scan_win474), .scan_win_std_dev(scan_win_std_dev[474]), .feature_accum(feature_accums[474]));
  accum_calculator #(.RECT1_X(rectangle1_xs[475]), .RECT1_Y(rectangle1_ys[475]), .RECT1_WIDTH(rectangle1_widths[475]), .RECT1_HEIGHT(rectangle1_heights[475]), .RECT1_WEIGHT(rectangle1_weights[475]), .RECT2_X(rectangle2_xs[475]), .RECT2_Y(rectangle2_ys[475]), .RECT2_WIDTH(rectangle2_widths[475]), .RECT2_HEIGHT(rectangle2_heights[475]), .RECT2_WEIGHT(rectangle2_weights[475]), .RECT3_X(rectangle3_xs[475]), .RECT3_Y(rectangle3_ys[475]), .RECT3_WIDTH(rectangle3_widths[475]), .RECT3_HEIGHT(rectangle3_heights[475]), .RECT3_WEIGHT(rectangle3_weights[475]), .FEAT_THRES(feature_thresholds[475]), .FEAT_ABOVE(feature_aboves[475]), .FEAT_BELOW(feature_belows[475])) ac475(.scan_win(scan_win475), .scan_win_std_dev(scan_win_std_dev[475]), .feature_accum(feature_accums[475]));
  accum_calculator #(.RECT1_X(rectangle1_xs[476]), .RECT1_Y(rectangle1_ys[476]), .RECT1_WIDTH(rectangle1_widths[476]), .RECT1_HEIGHT(rectangle1_heights[476]), .RECT1_WEIGHT(rectangle1_weights[476]), .RECT2_X(rectangle2_xs[476]), .RECT2_Y(rectangle2_ys[476]), .RECT2_WIDTH(rectangle2_widths[476]), .RECT2_HEIGHT(rectangle2_heights[476]), .RECT2_WEIGHT(rectangle2_weights[476]), .RECT3_X(rectangle3_xs[476]), .RECT3_Y(rectangle3_ys[476]), .RECT3_WIDTH(rectangle3_widths[476]), .RECT3_HEIGHT(rectangle3_heights[476]), .RECT3_WEIGHT(rectangle3_weights[476]), .FEAT_THRES(feature_thresholds[476]), .FEAT_ABOVE(feature_aboves[476]), .FEAT_BELOW(feature_belows[476])) ac476(.scan_win(scan_win476), .scan_win_std_dev(scan_win_std_dev[476]), .feature_accum(feature_accums[476]));
  accum_calculator #(.RECT1_X(rectangle1_xs[477]), .RECT1_Y(rectangle1_ys[477]), .RECT1_WIDTH(rectangle1_widths[477]), .RECT1_HEIGHT(rectangle1_heights[477]), .RECT1_WEIGHT(rectangle1_weights[477]), .RECT2_X(rectangle2_xs[477]), .RECT2_Y(rectangle2_ys[477]), .RECT2_WIDTH(rectangle2_widths[477]), .RECT2_HEIGHT(rectangle2_heights[477]), .RECT2_WEIGHT(rectangle2_weights[477]), .RECT3_X(rectangle3_xs[477]), .RECT3_Y(rectangle3_ys[477]), .RECT3_WIDTH(rectangle3_widths[477]), .RECT3_HEIGHT(rectangle3_heights[477]), .RECT3_WEIGHT(rectangle3_weights[477]), .FEAT_THRES(feature_thresholds[477]), .FEAT_ABOVE(feature_aboves[477]), .FEAT_BELOW(feature_belows[477])) ac477(.scan_win(scan_win477), .scan_win_std_dev(scan_win_std_dev[477]), .feature_accum(feature_accums[477]));
  accum_calculator #(.RECT1_X(rectangle1_xs[478]), .RECT1_Y(rectangle1_ys[478]), .RECT1_WIDTH(rectangle1_widths[478]), .RECT1_HEIGHT(rectangle1_heights[478]), .RECT1_WEIGHT(rectangle1_weights[478]), .RECT2_X(rectangle2_xs[478]), .RECT2_Y(rectangle2_ys[478]), .RECT2_WIDTH(rectangle2_widths[478]), .RECT2_HEIGHT(rectangle2_heights[478]), .RECT2_WEIGHT(rectangle2_weights[478]), .RECT3_X(rectangle3_xs[478]), .RECT3_Y(rectangle3_ys[478]), .RECT3_WIDTH(rectangle3_widths[478]), .RECT3_HEIGHT(rectangle3_heights[478]), .RECT3_WEIGHT(rectangle3_weights[478]), .FEAT_THRES(feature_thresholds[478]), .FEAT_ABOVE(feature_aboves[478]), .FEAT_BELOW(feature_belows[478])) ac478(.scan_win(scan_win478), .scan_win_std_dev(scan_win_std_dev[478]), .feature_accum(feature_accums[478]));
  accum_calculator #(.RECT1_X(rectangle1_xs[479]), .RECT1_Y(rectangle1_ys[479]), .RECT1_WIDTH(rectangle1_widths[479]), .RECT1_HEIGHT(rectangle1_heights[479]), .RECT1_WEIGHT(rectangle1_weights[479]), .RECT2_X(rectangle2_xs[479]), .RECT2_Y(rectangle2_ys[479]), .RECT2_WIDTH(rectangle2_widths[479]), .RECT2_HEIGHT(rectangle2_heights[479]), .RECT2_WEIGHT(rectangle2_weights[479]), .RECT3_X(rectangle3_xs[479]), .RECT3_Y(rectangle3_ys[479]), .RECT3_WIDTH(rectangle3_widths[479]), .RECT3_HEIGHT(rectangle3_heights[479]), .RECT3_WEIGHT(rectangle3_weights[479]), .FEAT_THRES(feature_thresholds[479]), .FEAT_ABOVE(feature_aboves[479]), .FEAT_BELOW(feature_belows[479])) ac479(.scan_win(scan_win479), .scan_win_std_dev(scan_win_std_dev[479]), .feature_accum(feature_accums[479]));
  accum_calculator #(.RECT1_X(rectangle1_xs[480]), .RECT1_Y(rectangle1_ys[480]), .RECT1_WIDTH(rectangle1_widths[480]), .RECT1_HEIGHT(rectangle1_heights[480]), .RECT1_WEIGHT(rectangle1_weights[480]), .RECT2_X(rectangle2_xs[480]), .RECT2_Y(rectangle2_ys[480]), .RECT2_WIDTH(rectangle2_widths[480]), .RECT2_HEIGHT(rectangle2_heights[480]), .RECT2_WEIGHT(rectangle2_weights[480]), .RECT3_X(rectangle3_xs[480]), .RECT3_Y(rectangle3_ys[480]), .RECT3_WIDTH(rectangle3_widths[480]), .RECT3_HEIGHT(rectangle3_heights[480]), .RECT3_WEIGHT(rectangle3_weights[480]), .FEAT_THRES(feature_thresholds[480]), .FEAT_ABOVE(feature_aboves[480]), .FEAT_BELOW(feature_belows[480])) ac480(.scan_win(scan_win480), .scan_win_std_dev(scan_win_std_dev[480]), .feature_accum(feature_accums[480]));
  accum_calculator #(.RECT1_X(rectangle1_xs[481]), .RECT1_Y(rectangle1_ys[481]), .RECT1_WIDTH(rectangle1_widths[481]), .RECT1_HEIGHT(rectangle1_heights[481]), .RECT1_WEIGHT(rectangle1_weights[481]), .RECT2_X(rectangle2_xs[481]), .RECT2_Y(rectangle2_ys[481]), .RECT2_WIDTH(rectangle2_widths[481]), .RECT2_HEIGHT(rectangle2_heights[481]), .RECT2_WEIGHT(rectangle2_weights[481]), .RECT3_X(rectangle3_xs[481]), .RECT3_Y(rectangle3_ys[481]), .RECT3_WIDTH(rectangle3_widths[481]), .RECT3_HEIGHT(rectangle3_heights[481]), .RECT3_WEIGHT(rectangle3_weights[481]), .FEAT_THRES(feature_thresholds[481]), .FEAT_ABOVE(feature_aboves[481]), .FEAT_BELOW(feature_belows[481])) ac481(.scan_win(scan_win481), .scan_win_std_dev(scan_win_std_dev[481]), .feature_accum(feature_accums[481]));
  accum_calculator #(.RECT1_X(rectangle1_xs[482]), .RECT1_Y(rectangle1_ys[482]), .RECT1_WIDTH(rectangle1_widths[482]), .RECT1_HEIGHT(rectangle1_heights[482]), .RECT1_WEIGHT(rectangle1_weights[482]), .RECT2_X(rectangle2_xs[482]), .RECT2_Y(rectangle2_ys[482]), .RECT2_WIDTH(rectangle2_widths[482]), .RECT2_HEIGHT(rectangle2_heights[482]), .RECT2_WEIGHT(rectangle2_weights[482]), .RECT3_X(rectangle3_xs[482]), .RECT3_Y(rectangle3_ys[482]), .RECT3_WIDTH(rectangle3_widths[482]), .RECT3_HEIGHT(rectangle3_heights[482]), .RECT3_WEIGHT(rectangle3_weights[482]), .FEAT_THRES(feature_thresholds[482]), .FEAT_ABOVE(feature_aboves[482]), .FEAT_BELOW(feature_belows[482])) ac482(.scan_win(scan_win482), .scan_win_std_dev(scan_win_std_dev[482]), .feature_accum(feature_accums[482]));
  accum_calculator #(.RECT1_X(rectangle1_xs[483]), .RECT1_Y(rectangle1_ys[483]), .RECT1_WIDTH(rectangle1_widths[483]), .RECT1_HEIGHT(rectangle1_heights[483]), .RECT1_WEIGHT(rectangle1_weights[483]), .RECT2_X(rectangle2_xs[483]), .RECT2_Y(rectangle2_ys[483]), .RECT2_WIDTH(rectangle2_widths[483]), .RECT2_HEIGHT(rectangle2_heights[483]), .RECT2_WEIGHT(rectangle2_weights[483]), .RECT3_X(rectangle3_xs[483]), .RECT3_Y(rectangle3_ys[483]), .RECT3_WIDTH(rectangle3_widths[483]), .RECT3_HEIGHT(rectangle3_heights[483]), .RECT3_WEIGHT(rectangle3_weights[483]), .FEAT_THRES(feature_thresholds[483]), .FEAT_ABOVE(feature_aboves[483]), .FEAT_BELOW(feature_belows[483])) ac483(.scan_win(scan_win483), .scan_win_std_dev(scan_win_std_dev[483]), .feature_accum(feature_accums[483]));
  accum_calculator #(.RECT1_X(rectangle1_xs[484]), .RECT1_Y(rectangle1_ys[484]), .RECT1_WIDTH(rectangle1_widths[484]), .RECT1_HEIGHT(rectangle1_heights[484]), .RECT1_WEIGHT(rectangle1_weights[484]), .RECT2_X(rectangle2_xs[484]), .RECT2_Y(rectangle2_ys[484]), .RECT2_WIDTH(rectangle2_widths[484]), .RECT2_HEIGHT(rectangle2_heights[484]), .RECT2_WEIGHT(rectangle2_weights[484]), .RECT3_X(rectangle3_xs[484]), .RECT3_Y(rectangle3_ys[484]), .RECT3_WIDTH(rectangle3_widths[484]), .RECT3_HEIGHT(rectangle3_heights[484]), .RECT3_WEIGHT(rectangle3_weights[484]), .FEAT_THRES(feature_thresholds[484]), .FEAT_ABOVE(feature_aboves[484]), .FEAT_BELOW(feature_belows[484])) ac484(.scan_win(scan_win484), .scan_win_std_dev(scan_win_std_dev[484]), .feature_accum(feature_accums[484]));
  accum_calculator #(.RECT1_X(rectangle1_xs[485]), .RECT1_Y(rectangle1_ys[485]), .RECT1_WIDTH(rectangle1_widths[485]), .RECT1_HEIGHT(rectangle1_heights[485]), .RECT1_WEIGHT(rectangle1_weights[485]), .RECT2_X(rectangle2_xs[485]), .RECT2_Y(rectangle2_ys[485]), .RECT2_WIDTH(rectangle2_widths[485]), .RECT2_HEIGHT(rectangle2_heights[485]), .RECT2_WEIGHT(rectangle2_weights[485]), .RECT3_X(rectangle3_xs[485]), .RECT3_Y(rectangle3_ys[485]), .RECT3_WIDTH(rectangle3_widths[485]), .RECT3_HEIGHT(rectangle3_heights[485]), .RECT3_WEIGHT(rectangle3_weights[485]), .FEAT_THRES(feature_thresholds[485]), .FEAT_ABOVE(feature_aboves[485]), .FEAT_BELOW(feature_belows[485])) ac485(.scan_win(scan_win485), .scan_win_std_dev(scan_win_std_dev[485]), .feature_accum(feature_accums[485]));
  accum_calculator #(.RECT1_X(rectangle1_xs[486]), .RECT1_Y(rectangle1_ys[486]), .RECT1_WIDTH(rectangle1_widths[486]), .RECT1_HEIGHT(rectangle1_heights[486]), .RECT1_WEIGHT(rectangle1_weights[486]), .RECT2_X(rectangle2_xs[486]), .RECT2_Y(rectangle2_ys[486]), .RECT2_WIDTH(rectangle2_widths[486]), .RECT2_HEIGHT(rectangle2_heights[486]), .RECT2_WEIGHT(rectangle2_weights[486]), .RECT3_X(rectangle3_xs[486]), .RECT3_Y(rectangle3_ys[486]), .RECT3_WIDTH(rectangle3_widths[486]), .RECT3_HEIGHT(rectangle3_heights[486]), .RECT3_WEIGHT(rectangle3_weights[486]), .FEAT_THRES(feature_thresholds[486]), .FEAT_ABOVE(feature_aboves[486]), .FEAT_BELOW(feature_belows[486])) ac486(.scan_win(scan_win486), .scan_win_std_dev(scan_win_std_dev[486]), .feature_accum(feature_accums[486]));
  accum_calculator #(.RECT1_X(rectangle1_xs[487]), .RECT1_Y(rectangle1_ys[487]), .RECT1_WIDTH(rectangle1_widths[487]), .RECT1_HEIGHT(rectangle1_heights[487]), .RECT1_WEIGHT(rectangle1_weights[487]), .RECT2_X(rectangle2_xs[487]), .RECT2_Y(rectangle2_ys[487]), .RECT2_WIDTH(rectangle2_widths[487]), .RECT2_HEIGHT(rectangle2_heights[487]), .RECT2_WEIGHT(rectangle2_weights[487]), .RECT3_X(rectangle3_xs[487]), .RECT3_Y(rectangle3_ys[487]), .RECT3_WIDTH(rectangle3_widths[487]), .RECT3_HEIGHT(rectangle3_heights[487]), .RECT3_WEIGHT(rectangle3_weights[487]), .FEAT_THRES(feature_thresholds[487]), .FEAT_ABOVE(feature_aboves[487]), .FEAT_BELOW(feature_belows[487])) ac487(.scan_win(scan_win487), .scan_win_std_dev(scan_win_std_dev[487]), .feature_accum(feature_accums[487]));
  accum_calculator #(.RECT1_X(rectangle1_xs[488]), .RECT1_Y(rectangle1_ys[488]), .RECT1_WIDTH(rectangle1_widths[488]), .RECT1_HEIGHT(rectangle1_heights[488]), .RECT1_WEIGHT(rectangle1_weights[488]), .RECT2_X(rectangle2_xs[488]), .RECT2_Y(rectangle2_ys[488]), .RECT2_WIDTH(rectangle2_widths[488]), .RECT2_HEIGHT(rectangle2_heights[488]), .RECT2_WEIGHT(rectangle2_weights[488]), .RECT3_X(rectangle3_xs[488]), .RECT3_Y(rectangle3_ys[488]), .RECT3_WIDTH(rectangle3_widths[488]), .RECT3_HEIGHT(rectangle3_heights[488]), .RECT3_WEIGHT(rectangle3_weights[488]), .FEAT_THRES(feature_thresholds[488]), .FEAT_ABOVE(feature_aboves[488]), .FEAT_BELOW(feature_belows[488])) ac488(.scan_win(scan_win488), .scan_win_std_dev(scan_win_std_dev[488]), .feature_accum(feature_accums[488]));
  accum_calculator #(.RECT1_X(rectangle1_xs[489]), .RECT1_Y(rectangle1_ys[489]), .RECT1_WIDTH(rectangle1_widths[489]), .RECT1_HEIGHT(rectangle1_heights[489]), .RECT1_WEIGHT(rectangle1_weights[489]), .RECT2_X(rectangle2_xs[489]), .RECT2_Y(rectangle2_ys[489]), .RECT2_WIDTH(rectangle2_widths[489]), .RECT2_HEIGHT(rectangle2_heights[489]), .RECT2_WEIGHT(rectangle2_weights[489]), .RECT3_X(rectangle3_xs[489]), .RECT3_Y(rectangle3_ys[489]), .RECT3_WIDTH(rectangle3_widths[489]), .RECT3_HEIGHT(rectangle3_heights[489]), .RECT3_WEIGHT(rectangle3_weights[489]), .FEAT_THRES(feature_thresholds[489]), .FEAT_ABOVE(feature_aboves[489]), .FEAT_BELOW(feature_belows[489])) ac489(.scan_win(scan_win489), .scan_win_std_dev(scan_win_std_dev[489]), .feature_accum(feature_accums[489]));
  accum_calculator #(.RECT1_X(rectangle1_xs[490]), .RECT1_Y(rectangle1_ys[490]), .RECT1_WIDTH(rectangle1_widths[490]), .RECT1_HEIGHT(rectangle1_heights[490]), .RECT1_WEIGHT(rectangle1_weights[490]), .RECT2_X(rectangle2_xs[490]), .RECT2_Y(rectangle2_ys[490]), .RECT2_WIDTH(rectangle2_widths[490]), .RECT2_HEIGHT(rectangle2_heights[490]), .RECT2_WEIGHT(rectangle2_weights[490]), .RECT3_X(rectangle3_xs[490]), .RECT3_Y(rectangle3_ys[490]), .RECT3_WIDTH(rectangle3_widths[490]), .RECT3_HEIGHT(rectangle3_heights[490]), .RECT3_WEIGHT(rectangle3_weights[490]), .FEAT_THRES(feature_thresholds[490]), .FEAT_ABOVE(feature_aboves[490]), .FEAT_BELOW(feature_belows[490])) ac490(.scan_win(scan_win490), .scan_win_std_dev(scan_win_std_dev[490]), .feature_accum(feature_accums[490]));
  accum_calculator #(.RECT1_X(rectangle1_xs[491]), .RECT1_Y(rectangle1_ys[491]), .RECT1_WIDTH(rectangle1_widths[491]), .RECT1_HEIGHT(rectangle1_heights[491]), .RECT1_WEIGHT(rectangle1_weights[491]), .RECT2_X(rectangle2_xs[491]), .RECT2_Y(rectangle2_ys[491]), .RECT2_WIDTH(rectangle2_widths[491]), .RECT2_HEIGHT(rectangle2_heights[491]), .RECT2_WEIGHT(rectangle2_weights[491]), .RECT3_X(rectangle3_xs[491]), .RECT3_Y(rectangle3_ys[491]), .RECT3_WIDTH(rectangle3_widths[491]), .RECT3_HEIGHT(rectangle3_heights[491]), .RECT3_WEIGHT(rectangle3_weights[491]), .FEAT_THRES(feature_thresholds[491]), .FEAT_ABOVE(feature_aboves[491]), .FEAT_BELOW(feature_belows[491])) ac491(.scan_win(scan_win491), .scan_win_std_dev(scan_win_std_dev[491]), .feature_accum(feature_accums[491]));
  accum_calculator #(.RECT1_X(rectangle1_xs[492]), .RECT1_Y(rectangle1_ys[492]), .RECT1_WIDTH(rectangle1_widths[492]), .RECT1_HEIGHT(rectangle1_heights[492]), .RECT1_WEIGHT(rectangle1_weights[492]), .RECT2_X(rectangle2_xs[492]), .RECT2_Y(rectangle2_ys[492]), .RECT2_WIDTH(rectangle2_widths[492]), .RECT2_HEIGHT(rectangle2_heights[492]), .RECT2_WEIGHT(rectangle2_weights[492]), .RECT3_X(rectangle3_xs[492]), .RECT3_Y(rectangle3_ys[492]), .RECT3_WIDTH(rectangle3_widths[492]), .RECT3_HEIGHT(rectangle3_heights[492]), .RECT3_WEIGHT(rectangle3_weights[492]), .FEAT_THRES(feature_thresholds[492]), .FEAT_ABOVE(feature_aboves[492]), .FEAT_BELOW(feature_belows[492])) ac492(.scan_win(scan_win492), .scan_win_std_dev(scan_win_std_dev[492]), .feature_accum(feature_accums[492]));
  accum_calculator #(.RECT1_X(rectangle1_xs[493]), .RECT1_Y(rectangle1_ys[493]), .RECT1_WIDTH(rectangle1_widths[493]), .RECT1_HEIGHT(rectangle1_heights[493]), .RECT1_WEIGHT(rectangle1_weights[493]), .RECT2_X(rectangle2_xs[493]), .RECT2_Y(rectangle2_ys[493]), .RECT2_WIDTH(rectangle2_widths[493]), .RECT2_HEIGHT(rectangle2_heights[493]), .RECT2_WEIGHT(rectangle2_weights[493]), .RECT3_X(rectangle3_xs[493]), .RECT3_Y(rectangle3_ys[493]), .RECT3_WIDTH(rectangle3_widths[493]), .RECT3_HEIGHT(rectangle3_heights[493]), .RECT3_WEIGHT(rectangle3_weights[493]), .FEAT_THRES(feature_thresholds[493]), .FEAT_ABOVE(feature_aboves[493]), .FEAT_BELOW(feature_belows[493])) ac493(.scan_win(scan_win493), .scan_win_std_dev(scan_win_std_dev[493]), .feature_accum(feature_accums[493]));
  accum_calculator #(.RECT1_X(rectangle1_xs[494]), .RECT1_Y(rectangle1_ys[494]), .RECT1_WIDTH(rectangle1_widths[494]), .RECT1_HEIGHT(rectangle1_heights[494]), .RECT1_WEIGHT(rectangle1_weights[494]), .RECT2_X(rectangle2_xs[494]), .RECT2_Y(rectangle2_ys[494]), .RECT2_WIDTH(rectangle2_widths[494]), .RECT2_HEIGHT(rectangle2_heights[494]), .RECT2_WEIGHT(rectangle2_weights[494]), .RECT3_X(rectangle3_xs[494]), .RECT3_Y(rectangle3_ys[494]), .RECT3_WIDTH(rectangle3_widths[494]), .RECT3_HEIGHT(rectangle3_heights[494]), .RECT3_WEIGHT(rectangle3_weights[494]), .FEAT_THRES(feature_thresholds[494]), .FEAT_ABOVE(feature_aboves[494]), .FEAT_BELOW(feature_belows[494])) ac494(.scan_win(scan_win494), .scan_win_std_dev(scan_win_std_dev[494]), .feature_accum(feature_accums[494]));
  accum_calculator #(.RECT1_X(rectangle1_xs[495]), .RECT1_Y(rectangle1_ys[495]), .RECT1_WIDTH(rectangle1_widths[495]), .RECT1_HEIGHT(rectangle1_heights[495]), .RECT1_WEIGHT(rectangle1_weights[495]), .RECT2_X(rectangle2_xs[495]), .RECT2_Y(rectangle2_ys[495]), .RECT2_WIDTH(rectangle2_widths[495]), .RECT2_HEIGHT(rectangle2_heights[495]), .RECT2_WEIGHT(rectangle2_weights[495]), .RECT3_X(rectangle3_xs[495]), .RECT3_Y(rectangle3_ys[495]), .RECT3_WIDTH(rectangle3_widths[495]), .RECT3_HEIGHT(rectangle3_heights[495]), .RECT3_WEIGHT(rectangle3_weights[495]), .FEAT_THRES(feature_thresholds[495]), .FEAT_ABOVE(feature_aboves[495]), .FEAT_BELOW(feature_belows[495])) ac495(.scan_win(scan_win495), .scan_win_std_dev(scan_win_std_dev[495]), .feature_accum(feature_accums[495]));
  accum_calculator #(.RECT1_X(rectangle1_xs[496]), .RECT1_Y(rectangle1_ys[496]), .RECT1_WIDTH(rectangle1_widths[496]), .RECT1_HEIGHT(rectangle1_heights[496]), .RECT1_WEIGHT(rectangle1_weights[496]), .RECT2_X(rectangle2_xs[496]), .RECT2_Y(rectangle2_ys[496]), .RECT2_WIDTH(rectangle2_widths[496]), .RECT2_HEIGHT(rectangle2_heights[496]), .RECT2_WEIGHT(rectangle2_weights[496]), .RECT3_X(rectangle3_xs[496]), .RECT3_Y(rectangle3_ys[496]), .RECT3_WIDTH(rectangle3_widths[496]), .RECT3_HEIGHT(rectangle3_heights[496]), .RECT3_WEIGHT(rectangle3_weights[496]), .FEAT_THRES(feature_thresholds[496]), .FEAT_ABOVE(feature_aboves[496]), .FEAT_BELOW(feature_belows[496])) ac496(.scan_win(scan_win496), .scan_win_std_dev(scan_win_std_dev[496]), .feature_accum(feature_accums[496]));
  accum_calculator #(.RECT1_X(rectangle1_xs[497]), .RECT1_Y(rectangle1_ys[497]), .RECT1_WIDTH(rectangle1_widths[497]), .RECT1_HEIGHT(rectangle1_heights[497]), .RECT1_WEIGHT(rectangle1_weights[497]), .RECT2_X(rectangle2_xs[497]), .RECT2_Y(rectangle2_ys[497]), .RECT2_WIDTH(rectangle2_widths[497]), .RECT2_HEIGHT(rectangle2_heights[497]), .RECT2_WEIGHT(rectangle2_weights[497]), .RECT3_X(rectangle3_xs[497]), .RECT3_Y(rectangle3_ys[497]), .RECT3_WIDTH(rectangle3_widths[497]), .RECT3_HEIGHT(rectangle3_heights[497]), .RECT3_WEIGHT(rectangle3_weights[497]), .FEAT_THRES(feature_thresholds[497]), .FEAT_ABOVE(feature_aboves[497]), .FEAT_BELOW(feature_belows[497])) ac497(.scan_win(scan_win497), .scan_win_std_dev(scan_win_std_dev[497]), .feature_accum(feature_accums[497]));
  accum_calculator #(.RECT1_X(rectangle1_xs[498]), .RECT1_Y(rectangle1_ys[498]), .RECT1_WIDTH(rectangle1_widths[498]), .RECT1_HEIGHT(rectangle1_heights[498]), .RECT1_WEIGHT(rectangle1_weights[498]), .RECT2_X(rectangle2_xs[498]), .RECT2_Y(rectangle2_ys[498]), .RECT2_WIDTH(rectangle2_widths[498]), .RECT2_HEIGHT(rectangle2_heights[498]), .RECT2_WEIGHT(rectangle2_weights[498]), .RECT3_X(rectangle3_xs[498]), .RECT3_Y(rectangle3_ys[498]), .RECT3_WIDTH(rectangle3_widths[498]), .RECT3_HEIGHT(rectangle3_heights[498]), .RECT3_WEIGHT(rectangle3_weights[498]), .FEAT_THRES(feature_thresholds[498]), .FEAT_ABOVE(feature_aboves[498]), .FEAT_BELOW(feature_belows[498])) ac498(.scan_win(scan_win498), .scan_win_std_dev(scan_win_std_dev[498]), .feature_accum(feature_accums[498]));
  accum_calculator #(.RECT1_X(rectangle1_xs[499]), .RECT1_Y(rectangle1_ys[499]), .RECT1_WIDTH(rectangle1_widths[499]), .RECT1_HEIGHT(rectangle1_heights[499]), .RECT1_WEIGHT(rectangle1_weights[499]), .RECT2_X(rectangle2_xs[499]), .RECT2_Y(rectangle2_ys[499]), .RECT2_WIDTH(rectangle2_widths[499]), .RECT2_HEIGHT(rectangle2_heights[499]), .RECT2_WEIGHT(rectangle2_weights[499]), .RECT3_X(rectangle3_xs[499]), .RECT3_Y(rectangle3_ys[499]), .RECT3_WIDTH(rectangle3_widths[499]), .RECT3_HEIGHT(rectangle3_heights[499]), .RECT3_WEIGHT(rectangle3_weights[499]), .FEAT_THRES(feature_thresholds[499]), .FEAT_ABOVE(feature_aboves[499]), .FEAT_BELOW(feature_belows[499])) ac499(.scan_win(scan_win499), .scan_win_std_dev(scan_win_std_dev[499]), .feature_accum(feature_accums[499]));
  accum_calculator #(.RECT1_X(rectangle1_xs[500]), .RECT1_Y(rectangle1_ys[500]), .RECT1_WIDTH(rectangle1_widths[500]), .RECT1_HEIGHT(rectangle1_heights[500]), .RECT1_WEIGHT(rectangle1_weights[500]), .RECT2_X(rectangle2_xs[500]), .RECT2_Y(rectangle2_ys[500]), .RECT2_WIDTH(rectangle2_widths[500]), .RECT2_HEIGHT(rectangle2_heights[500]), .RECT2_WEIGHT(rectangle2_weights[500]), .RECT3_X(rectangle3_xs[500]), .RECT3_Y(rectangle3_ys[500]), .RECT3_WIDTH(rectangle3_widths[500]), .RECT3_HEIGHT(rectangle3_heights[500]), .RECT3_WEIGHT(rectangle3_weights[500]), .FEAT_THRES(feature_thresholds[500]), .FEAT_ABOVE(feature_aboves[500]), .FEAT_BELOW(feature_belows[500])) ac500(.scan_win(scan_win500), .scan_win_std_dev(scan_win_std_dev[500]), .feature_accum(feature_accums[500]));
  accum_calculator #(.RECT1_X(rectangle1_xs[501]), .RECT1_Y(rectangle1_ys[501]), .RECT1_WIDTH(rectangle1_widths[501]), .RECT1_HEIGHT(rectangle1_heights[501]), .RECT1_WEIGHT(rectangle1_weights[501]), .RECT2_X(rectangle2_xs[501]), .RECT2_Y(rectangle2_ys[501]), .RECT2_WIDTH(rectangle2_widths[501]), .RECT2_HEIGHT(rectangle2_heights[501]), .RECT2_WEIGHT(rectangle2_weights[501]), .RECT3_X(rectangle3_xs[501]), .RECT3_Y(rectangle3_ys[501]), .RECT3_WIDTH(rectangle3_widths[501]), .RECT3_HEIGHT(rectangle3_heights[501]), .RECT3_WEIGHT(rectangle3_weights[501]), .FEAT_THRES(feature_thresholds[501]), .FEAT_ABOVE(feature_aboves[501]), .FEAT_BELOW(feature_belows[501])) ac501(.scan_win(scan_win501), .scan_win_std_dev(scan_win_std_dev[501]), .feature_accum(feature_accums[501]));
  accum_calculator #(.RECT1_X(rectangle1_xs[502]), .RECT1_Y(rectangle1_ys[502]), .RECT1_WIDTH(rectangle1_widths[502]), .RECT1_HEIGHT(rectangle1_heights[502]), .RECT1_WEIGHT(rectangle1_weights[502]), .RECT2_X(rectangle2_xs[502]), .RECT2_Y(rectangle2_ys[502]), .RECT2_WIDTH(rectangle2_widths[502]), .RECT2_HEIGHT(rectangle2_heights[502]), .RECT2_WEIGHT(rectangle2_weights[502]), .RECT3_X(rectangle3_xs[502]), .RECT3_Y(rectangle3_ys[502]), .RECT3_WIDTH(rectangle3_widths[502]), .RECT3_HEIGHT(rectangle3_heights[502]), .RECT3_WEIGHT(rectangle3_weights[502]), .FEAT_THRES(feature_thresholds[502]), .FEAT_ABOVE(feature_aboves[502]), .FEAT_BELOW(feature_belows[502])) ac502(.scan_win(scan_win502), .scan_win_std_dev(scan_win_std_dev[502]), .feature_accum(feature_accums[502]));
  accum_calculator #(.RECT1_X(rectangle1_xs[503]), .RECT1_Y(rectangle1_ys[503]), .RECT1_WIDTH(rectangle1_widths[503]), .RECT1_HEIGHT(rectangle1_heights[503]), .RECT1_WEIGHT(rectangle1_weights[503]), .RECT2_X(rectangle2_xs[503]), .RECT2_Y(rectangle2_ys[503]), .RECT2_WIDTH(rectangle2_widths[503]), .RECT2_HEIGHT(rectangle2_heights[503]), .RECT2_WEIGHT(rectangle2_weights[503]), .RECT3_X(rectangle3_xs[503]), .RECT3_Y(rectangle3_ys[503]), .RECT3_WIDTH(rectangle3_widths[503]), .RECT3_HEIGHT(rectangle3_heights[503]), .RECT3_WEIGHT(rectangle3_weights[503]), .FEAT_THRES(feature_thresholds[503]), .FEAT_ABOVE(feature_aboves[503]), .FEAT_BELOW(feature_belows[503])) ac503(.scan_win(scan_win503), .scan_win_std_dev(scan_win_std_dev[503]), .feature_accum(feature_accums[503]));
  accum_calculator #(.RECT1_X(rectangle1_xs[504]), .RECT1_Y(rectangle1_ys[504]), .RECT1_WIDTH(rectangle1_widths[504]), .RECT1_HEIGHT(rectangle1_heights[504]), .RECT1_WEIGHT(rectangle1_weights[504]), .RECT2_X(rectangle2_xs[504]), .RECT2_Y(rectangle2_ys[504]), .RECT2_WIDTH(rectangle2_widths[504]), .RECT2_HEIGHT(rectangle2_heights[504]), .RECT2_WEIGHT(rectangle2_weights[504]), .RECT3_X(rectangle3_xs[504]), .RECT3_Y(rectangle3_ys[504]), .RECT3_WIDTH(rectangle3_widths[504]), .RECT3_HEIGHT(rectangle3_heights[504]), .RECT3_WEIGHT(rectangle3_weights[504]), .FEAT_THRES(feature_thresholds[504]), .FEAT_ABOVE(feature_aboves[504]), .FEAT_BELOW(feature_belows[504])) ac504(.scan_win(scan_win504), .scan_win_std_dev(scan_win_std_dev[504]), .feature_accum(feature_accums[504]));
  accum_calculator #(.RECT1_X(rectangle1_xs[505]), .RECT1_Y(rectangle1_ys[505]), .RECT1_WIDTH(rectangle1_widths[505]), .RECT1_HEIGHT(rectangle1_heights[505]), .RECT1_WEIGHT(rectangle1_weights[505]), .RECT2_X(rectangle2_xs[505]), .RECT2_Y(rectangle2_ys[505]), .RECT2_WIDTH(rectangle2_widths[505]), .RECT2_HEIGHT(rectangle2_heights[505]), .RECT2_WEIGHT(rectangle2_weights[505]), .RECT3_X(rectangle3_xs[505]), .RECT3_Y(rectangle3_ys[505]), .RECT3_WIDTH(rectangle3_widths[505]), .RECT3_HEIGHT(rectangle3_heights[505]), .RECT3_WEIGHT(rectangle3_weights[505]), .FEAT_THRES(feature_thresholds[505]), .FEAT_ABOVE(feature_aboves[505]), .FEAT_BELOW(feature_belows[505])) ac505(.scan_win(scan_win505), .scan_win_std_dev(scan_win_std_dev[505]), .feature_accum(feature_accums[505]));
  accum_calculator #(.RECT1_X(rectangle1_xs[506]), .RECT1_Y(rectangle1_ys[506]), .RECT1_WIDTH(rectangle1_widths[506]), .RECT1_HEIGHT(rectangle1_heights[506]), .RECT1_WEIGHT(rectangle1_weights[506]), .RECT2_X(rectangle2_xs[506]), .RECT2_Y(rectangle2_ys[506]), .RECT2_WIDTH(rectangle2_widths[506]), .RECT2_HEIGHT(rectangle2_heights[506]), .RECT2_WEIGHT(rectangle2_weights[506]), .RECT3_X(rectangle3_xs[506]), .RECT3_Y(rectangle3_ys[506]), .RECT3_WIDTH(rectangle3_widths[506]), .RECT3_HEIGHT(rectangle3_heights[506]), .RECT3_WEIGHT(rectangle3_weights[506]), .FEAT_THRES(feature_thresholds[506]), .FEAT_ABOVE(feature_aboves[506]), .FEAT_BELOW(feature_belows[506])) ac506(.scan_win(scan_win506), .scan_win_std_dev(scan_win_std_dev[506]), .feature_accum(feature_accums[506]));
  accum_calculator #(.RECT1_X(rectangle1_xs[507]), .RECT1_Y(rectangle1_ys[507]), .RECT1_WIDTH(rectangle1_widths[507]), .RECT1_HEIGHT(rectangle1_heights[507]), .RECT1_WEIGHT(rectangle1_weights[507]), .RECT2_X(rectangle2_xs[507]), .RECT2_Y(rectangle2_ys[507]), .RECT2_WIDTH(rectangle2_widths[507]), .RECT2_HEIGHT(rectangle2_heights[507]), .RECT2_WEIGHT(rectangle2_weights[507]), .RECT3_X(rectangle3_xs[507]), .RECT3_Y(rectangle3_ys[507]), .RECT3_WIDTH(rectangle3_widths[507]), .RECT3_HEIGHT(rectangle3_heights[507]), .RECT3_WEIGHT(rectangle3_weights[507]), .FEAT_THRES(feature_thresholds[507]), .FEAT_ABOVE(feature_aboves[507]), .FEAT_BELOW(feature_belows[507])) ac507(.scan_win(scan_win507), .scan_win_std_dev(scan_win_std_dev[507]), .feature_accum(feature_accums[507]));
  accum_calculator #(.RECT1_X(rectangle1_xs[508]), .RECT1_Y(rectangle1_ys[508]), .RECT1_WIDTH(rectangle1_widths[508]), .RECT1_HEIGHT(rectangle1_heights[508]), .RECT1_WEIGHT(rectangle1_weights[508]), .RECT2_X(rectangle2_xs[508]), .RECT2_Y(rectangle2_ys[508]), .RECT2_WIDTH(rectangle2_widths[508]), .RECT2_HEIGHT(rectangle2_heights[508]), .RECT2_WEIGHT(rectangle2_weights[508]), .RECT3_X(rectangle3_xs[508]), .RECT3_Y(rectangle3_ys[508]), .RECT3_WIDTH(rectangle3_widths[508]), .RECT3_HEIGHT(rectangle3_heights[508]), .RECT3_WEIGHT(rectangle3_weights[508]), .FEAT_THRES(feature_thresholds[508]), .FEAT_ABOVE(feature_aboves[508]), .FEAT_BELOW(feature_belows[508])) ac508(.scan_win(scan_win508), .scan_win_std_dev(scan_win_std_dev[508]), .feature_accum(feature_accums[508]));
  accum_calculator #(.RECT1_X(rectangle1_xs[509]), .RECT1_Y(rectangle1_ys[509]), .RECT1_WIDTH(rectangle1_widths[509]), .RECT1_HEIGHT(rectangle1_heights[509]), .RECT1_WEIGHT(rectangle1_weights[509]), .RECT2_X(rectangle2_xs[509]), .RECT2_Y(rectangle2_ys[509]), .RECT2_WIDTH(rectangle2_widths[509]), .RECT2_HEIGHT(rectangle2_heights[509]), .RECT2_WEIGHT(rectangle2_weights[509]), .RECT3_X(rectangle3_xs[509]), .RECT3_Y(rectangle3_ys[509]), .RECT3_WIDTH(rectangle3_widths[509]), .RECT3_HEIGHT(rectangle3_heights[509]), .RECT3_WEIGHT(rectangle3_weights[509]), .FEAT_THRES(feature_thresholds[509]), .FEAT_ABOVE(feature_aboves[509]), .FEAT_BELOW(feature_belows[509])) ac509(.scan_win(scan_win509), .scan_win_std_dev(scan_win_std_dev[509]), .feature_accum(feature_accums[509]));
  accum_calculator #(.RECT1_X(rectangle1_xs[510]), .RECT1_Y(rectangle1_ys[510]), .RECT1_WIDTH(rectangle1_widths[510]), .RECT1_HEIGHT(rectangle1_heights[510]), .RECT1_WEIGHT(rectangle1_weights[510]), .RECT2_X(rectangle2_xs[510]), .RECT2_Y(rectangle2_ys[510]), .RECT2_WIDTH(rectangle2_widths[510]), .RECT2_HEIGHT(rectangle2_heights[510]), .RECT2_WEIGHT(rectangle2_weights[510]), .RECT3_X(rectangle3_xs[510]), .RECT3_Y(rectangle3_ys[510]), .RECT3_WIDTH(rectangle3_widths[510]), .RECT3_HEIGHT(rectangle3_heights[510]), .RECT3_WEIGHT(rectangle3_weights[510]), .FEAT_THRES(feature_thresholds[510]), .FEAT_ABOVE(feature_aboves[510]), .FEAT_BELOW(feature_belows[510])) ac510(.scan_win(scan_win510), .scan_win_std_dev(scan_win_std_dev[510]), .feature_accum(feature_accums[510]));
  accum_calculator #(.RECT1_X(rectangle1_xs[511]), .RECT1_Y(rectangle1_ys[511]), .RECT1_WIDTH(rectangle1_widths[511]), .RECT1_HEIGHT(rectangle1_heights[511]), .RECT1_WEIGHT(rectangle1_weights[511]), .RECT2_X(rectangle2_xs[511]), .RECT2_Y(rectangle2_ys[511]), .RECT2_WIDTH(rectangle2_widths[511]), .RECT2_HEIGHT(rectangle2_heights[511]), .RECT2_WEIGHT(rectangle2_weights[511]), .RECT3_X(rectangle3_xs[511]), .RECT3_Y(rectangle3_ys[511]), .RECT3_WIDTH(rectangle3_widths[511]), .RECT3_HEIGHT(rectangle3_heights[511]), .RECT3_WEIGHT(rectangle3_weights[511]), .FEAT_THRES(feature_thresholds[511]), .FEAT_ABOVE(feature_aboves[511]), .FEAT_BELOW(feature_belows[511])) ac511(.scan_win(scan_win511), .scan_win_std_dev(scan_win_std_dev[511]), .feature_accum(feature_accums[511]));
  accum_calculator #(.RECT1_X(rectangle1_xs[512]), .RECT1_Y(rectangle1_ys[512]), .RECT1_WIDTH(rectangle1_widths[512]), .RECT1_HEIGHT(rectangle1_heights[512]), .RECT1_WEIGHT(rectangle1_weights[512]), .RECT2_X(rectangle2_xs[512]), .RECT2_Y(rectangle2_ys[512]), .RECT2_WIDTH(rectangle2_widths[512]), .RECT2_HEIGHT(rectangle2_heights[512]), .RECT2_WEIGHT(rectangle2_weights[512]), .RECT3_X(rectangle3_xs[512]), .RECT3_Y(rectangle3_ys[512]), .RECT3_WIDTH(rectangle3_widths[512]), .RECT3_HEIGHT(rectangle3_heights[512]), .RECT3_WEIGHT(rectangle3_weights[512]), .FEAT_THRES(feature_thresholds[512]), .FEAT_ABOVE(feature_aboves[512]), .FEAT_BELOW(feature_belows[512])) ac512(.scan_win(scan_win512), .scan_win_std_dev(scan_win_std_dev[512]), .feature_accum(feature_accums[512]));
  accum_calculator #(.RECT1_X(rectangle1_xs[513]), .RECT1_Y(rectangle1_ys[513]), .RECT1_WIDTH(rectangle1_widths[513]), .RECT1_HEIGHT(rectangle1_heights[513]), .RECT1_WEIGHT(rectangle1_weights[513]), .RECT2_X(rectangle2_xs[513]), .RECT2_Y(rectangle2_ys[513]), .RECT2_WIDTH(rectangle2_widths[513]), .RECT2_HEIGHT(rectangle2_heights[513]), .RECT2_WEIGHT(rectangle2_weights[513]), .RECT3_X(rectangle3_xs[513]), .RECT3_Y(rectangle3_ys[513]), .RECT3_WIDTH(rectangle3_widths[513]), .RECT3_HEIGHT(rectangle3_heights[513]), .RECT3_WEIGHT(rectangle3_weights[513]), .FEAT_THRES(feature_thresholds[513]), .FEAT_ABOVE(feature_aboves[513]), .FEAT_BELOW(feature_belows[513])) ac513(.scan_win(scan_win513), .scan_win_std_dev(scan_win_std_dev[513]), .feature_accum(feature_accums[513]));
  accum_calculator #(.RECT1_X(rectangle1_xs[514]), .RECT1_Y(rectangle1_ys[514]), .RECT1_WIDTH(rectangle1_widths[514]), .RECT1_HEIGHT(rectangle1_heights[514]), .RECT1_WEIGHT(rectangle1_weights[514]), .RECT2_X(rectangle2_xs[514]), .RECT2_Y(rectangle2_ys[514]), .RECT2_WIDTH(rectangle2_widths[514]), .RECT2_HEIGHT(rectangle2_heights[514]), .RECT2_WEIGHT(rectangle2_weights[514]), .RECT3_X(rectangle3_xs[514]), .RECT3_Y(rectangle3_ys[514]), .RECT3_WIDTH(rectangle3_widths[514]), .RECT3_HEIGHT(rectangle3_heights[514]), .RECT3_WEIGHT(rectangle3_weights[514]), .FEAT_THRES(feature_thresholds[514]), .FEAT_ABOVE(feature_aboves[514]), .FEAT_BELOW(feature_belows[514])) ac514(.scan_win(scan_win514), .scan_win_std_dev(scan_win_std_dev[514]), .feature_accum(feature_accums[514]));
  accum_calculator #(.RECT1_X(rectangle1_xs[515]), .RECT1_Y(rectangle1_ys[515]), .RECT1_WIDTH(rectangle1_widths[515]), .RECT1_HEIGHT(rectangle1_heights[515]), .RECT1_WEIGHT(rectangle1_weights[515]), .RECT2_X(rectangle2_xs[515]), .RECT2_Y(rectangle2_ys[515]), .RECT2_WIDTH(rectangle2_widths[515]), .RECT2_HEIGHT(rectangle2_heights[515]), .RECT2_WEIGHT(rectangle2_weights[515]), .RECT3_X(rectangle3_xs[515]), .RECT3_Y(rectangle3_ys[515]), .RECT3_WIDTH(rectangle3_widths[515]), .RECT3_HEIGHT(rectangle3_heights[515]), .RECT3_WEIGHT(rectangle3_weights[515]), .FEAT_THRES(feature_thresholds[515]), .FEAT_ABOVE(feature_aboves[515]), .FEAT_BELOW(feature_belows[515])) ac515(.scan_win(scan_win515), .scan_win_std_dev(scan_win_std_dev[515]), .feature_accum(feature_accums[515]));
  accum_calculator #(.RECT1_X(rectangle1_xs[516]), .RECT1_Y(rectangle1_ys[516]), .RECT1_WIDTH(rectangle1_widths[516]), .RECT1_HEIGHT(rectangle1_heights[516]), .RECT1_WEIGHT(rectangle1_weights[516]), .RECT2_X(rectangle2_xs[516]), .RECT2_Y(rectangle2_ys[516]), .RECT2_WIDTH(rectangle2_widths[516]), .RECT2_HEIGHT(rectangle2_heights[516]), .RECT2_WEIGHT(rectangle2_weights[516]), .RECT3_X(rectangle3_xs[516]), .RECT3_Y(rectangle3_ys[516]), .RECT3_WIDTH(rectangle3_widths[516]), .RECT3_HEIGHT(rectangle3_heights[516]), .RECT3_WEIGHT(rectangle3_weights[516]), .FEAT_THRES(feature_thresholds[516]), .FEAT_ABOVE(feature_aboves[516]), .FEAT_BELOW(feature_belows[516])) ac516(.scan_win(scan_win516), .scan_win_std_dev(scan_win_std_dev[516]), .feature_accum(feature_accums[516]));
  accum_calculator #(.RECT1_X(rectangle1_xs[517]), .RECT1_Y(rectangle1_ys[517]), .RECT1_WIDTH(rectangle1_widths[517]), .RECT1_HEIGHT(rectangle1_heights[517]), .RECT1_WEIGHT(rectangle1_weights[517]), .RECT2_X(rectangle2_xs[517]), .RECT2_Y(rectangle2_ys[517]), .RECT2_WIDTH(rectangle2_widths[517]), .RECT2_HEIGHT(rectangle2_heights[517]), .RECT2_WEIGHT(rectangle2_weights[517]), .RECT3_X(rectangle3_xs[517]), .RECT3_Y(rectangle3_ys[517]), .RECT3_WIDTH(rectangle3_widths[517]), .RECT3_HEIGHT(rectangle3_heights[517]), .RECT3_WEIGHT(rectangle3_weights[517]), .FEAT_THRES(feature_thresholds[517]), .FEAT_ABOVE(feature_aboves[517]), .FEAT_BELOW(feature_belows[517])) ac517(.scan_win(scan_win517), .scan_win_std_dev(scan_win_std_dev[517]), .feature_accum(feature_accums[517]));
  accum_calculator #(.RECT1_X(rectangle1_xs[518]), .RECT1_Y(rectangle1_ys[518]), .RECT1_WIDTH(rectangle1_widths[518]), .RECT1_HEIGHT(rectangle1_heights[518]), .RECT1_WEIGHT(rectangle1_weights[518]), .RECT2_X(rectangle2_xs[518]), .RECT2_Y(rectangle2_ys[518]), .RECT2_WIDTH(rectangle2_widths[518]), .RECT2_HEIGHT(rectangle2_heights[518]), .RECT2_WEIGHT(rectangle2_weights[518]), .RECT3_X(rectangle3_xs[518]), .RECT3_Y(rectangle3_ys[518]), .RECT3_WIDTH(rectangle3_widths[518]), .RECT3_HEIGHT(rectangle3_heights[518]), .RECT3_WEIGHT(rectangle3_weights[518]), .FEAT_THRES(feature_thresholds[518]), .FEAT_ABOVE(feature_aboves[518]), .FEAT_BELOW(feature_belows[518])) ac518(.scan_win(scan_win518), .scan_win_std_dev(scan_win_std_dev[518]), .feature_accum(feature_accums[518]));
  accum_calculator #(.RECT1_X(rectangle1_xs[519]), .RECT1_Y(rectangle1_ys[519]), .RECT1_WIDTH(rectangle1_widths[519]), .RECT1_HEIGHT(rectangle1_heights[519]), .RECT1_WEIGHT(rectangle1_weights[519]), .RECT2_X(rectangle2_xs[519]), .RECT2_Y(rectangle2_ys[519]), .RECT2_WIDTH(rectangle2_widths[519]), .RECT2_HEIGHT(rectangle2_heights[519]), .RECT2_WEIGHT(rectangle2_weights[519]), .RECT3_X(rectangle3_xs[519]), .RECT3_Y(rectangle3_ys[519]), .RECT3_WIDTH(rectangle3_widths[519]), .RECT3_HEIGHT(rectangle3_heights[519]), .RECT3_WEIGHT(rectangle3_weights[519]), .FEAT_THRES(feature_thresholds[519]), .FEAT_ABOVE(feature_aboves[519]), .FEAT_BELOW(feature_belows[519])) ac519(.scan_win(scan_win519), .scan_win_std_dev(scan_win_std_dev[519]), .feature_accum(feature_accums[519]));
  accum_calculator #(.RECT1_X(rectangle1_xs[520]), .RECT1_Y(rectangle1_ys[520]), .RECT1_WIDTH(rectangle1_widths[520]), .RECT1_HEIGHT(rectangle1_heights[520]), .RECT1_WEIGHT(rectangle1_weights[520]), .RECT2_X(rectangle2_xs[520]), .RECT2_Y(rectangle2_ys[520]), .RECT2_WIDTH(rectangle2_widths[520]), .RECT2_HEIGHT(rectangle2_heights[520]), .RECT2_WEIGHT(rectangle2_weights[520]), .RECT3_X(rectangle3_xs[520]), .RECT3_Y(rectangle3_ys[520]), .RECT3_WIDTH(rectangle3_widths[520]), .RECT3_HEIGHT(rectangle3_heights[520]), .RECT3_WEIGHT(rectangle3_weights[520]), .FEAT_THRES(feature_thresholds[520]), .FEAT_ABOVE(feature_aboves[520]), .FEAT_BELOW(feature_belows[520])) ac520(.scan_win(scan_win520), .scan_win_std_dev(scan_win_std_dev[520]), .feature_accum(feature_accums[520]));
  accum_calculator #(.RECT1_X(rectangle1_xs[521]), .RECT1_Y(rectangle1_ys[521]), .RECT1_WIDTH(rectangle1_widths[521]), .RECT1_HEIGHT(rectangle1_heights[521]), .RECT1_WEIGHT(rectangle1_weights[521]), .RECT2_X(rectangle2_xs[521]), .RECT2_Y(rectangle2_ys[521]), .RECT2_WIDTH(rectangle2_widths[521]), .RECT2_HEIGHT(rectangle2_heights[521]), .RECT2_WEIGHT(rectangle2_weights[521]), .RECT3_X(rectangle3_xs[521]), .RECT3_Y(rectangle3_ys[521]), .RECT3_WIDTH(rectangle3_widths[521]), .RECT3_HEIGHT(rectangle3_heights[521]), .RECT3_WEIGHT(rectangle3_weights[521]), .FEAT_THRES(feature_thresholds[521]), .FEAT_ABOVE(feature_aboves[521]), .FEAT_BELOW(feature_belows[521])) ac521(.scan_win(scan_win521), .scan_win_std_dev(scan_win_std_dev[521]), .feature_accum(feature_accums[521]));
  accum_calculator #(.RECT1_X(rectangle1_xs[522]), .RECT1_Y(rectangle1_ys[522]), .RECT1_WIDTH(rectangle1_widths[522]), .RECT1_HEIGHT(rectangle1_heights[522]), .RECT1_WEIGHT(rectangle1_weights[522]), .RECT2_X(rectangle2_xs[522]), .RECT2_Y(rectangle2_ys[522]), .RECT2_WIDTH(rectangle2_widths[522]), .RECT2_HEIGHT(rectangle2_heights[522]), .RECT2_WEIGHT(rectangle2_weights[522]), .RECT3_X(rectangle3_xs[522]), .RECT3_Y(rectangle3_ys[522]), .RECT3_WIDTH(rectangle3_widths[522]), .RECT3_HEIGHT(rectangle3_heights[522]), .RECT3_WEIGHT(rectangle3_weights[522]), .FEAT_THRES(feature_thresholds[522]), .FEAT_ABOVE(feature_aboves[522]), .FEAT_BELOW(feature_belows[522])) ac522(.scan_win(scan_win522), .scan_win_std_dev(scan_win_std_dev[522]), .feature_accum(feature_accums[522]));
  accum_calculator #(.RECT1_X(rectangle1_xs[523]), .RECT1_Y(rectangle1_ys[523]), .RECT1_WIDTH(rectangle1_widths[523]), .RECT1_HEIGHT(rectangle1_heights[523]), .RECT1_WEIGHT(rectangle1_weights[523]), .RECT2_X(rectangle2_xs[523]), .RECT2_Y(rectangle2_ys[523]), .RECT2_WIDTH(rectangle2_widths[523]), .RECT2_HEIGHT(rectangle2_heights[523]), .RECT2_WEIGHT(rectangle2_weights[523]), .RECT3_X(rectangle3_xs[523]), .RECT3_Y(rectangle3_ys[523]), .RECT3_WIDTH(rectangle3_widths[523]), .RECT3_HEIGHT(rectangle3_heights[523]), .RECT3_WEIGHT(rectangle3_weights[523]), .FEAT_THRES(feature_thresholds[523]), .FEAT_ABOVE(feature_aboves[523]), .FEAT_BELOW(feature_belows[523])) ac523(.scan_win(scan_win523), .scan_win_std_dev(scan_win_std_dev[523]), .feature_accum(feature_accums[523]));
  accum_calculator #(.RECT1_X(rectangle1_xs[524]), .RECT1_Y(rectangle1_ys[524]), .RECT1_WIDTH(rectangle1_widths[524]), .RECT1_HEIGHT(rectangle1_heights[524]), .RECT1_WEIGHT(rectangle1_weights[524]), .RECT2_X(rectangle2_xs[524]), .RECT2_Y(rectangle2_ys[524]), .RECT2_WIDTH(rectangle2_widths[524]), .RECT2_HEIGHT(rectangle2_heights[524]), .RECT2_WEIGHT(rectangle2_weights[524]), .RECT3_X(rectangle3_xs[524]), .RECT3_Y(rectangle3_ys[524]), .RECT3_WIDTH(rectangle3_widths[524]), .RECT3_HEIGHT(rectangle3_heights[524]), .RECT3_WEIGHT(rectangle3_weights[524]), .FEAT_THRES(feature_thresholds[524]), .FEAT_ABOVE(feature_aboves[524]), .FEAT_BELOW(feature_belows[524])) ac524(.scan_win(scan_win524), .scan_win_std_dev(scan_win_std_dev[524]), .feature_accum(feature_accums[524]));
  accum_calculator #(.RECT1_X(rectangle1_xs[525]), .RECT1_Y(rectangle1_ys[525]), .RECT1_WIDTH(rectangle1_widths[525]), .RECT1_HEIGHT(rectangle1_heights[525]), .RECT1_WEIGHT(rectangle1_weights[525]), .RECT2_X(rectangle2_xs[525]), .RECT2_Y(rectangle2_ys[525]), .RECT2_WIDTH(rectangle2_widths[525]), .RECT2_HEIGHT(rectangle2_heights[525]), .RECT2_WEIGHT(rectangle2_weights[525]), .RECT3_X(rectangle3_xs[525]), .RECT3_Y(rectangle3_ys[525]), .RECT3_WIDTH(rectangle3_widths[525]), .RECT3_HEIGHT(rectangle3_heights[525]), .RECT3_WEIGHT(rectangle3_weights[525]), .FEAT_THRES(feature_thresholds[525]), .FEAT_ABOVE(feature_aboves[525]), .FEAT_BELOW(feature_belows[525])) ac525(.scan_win(scan_win525), .scan_win_std_dev(scan_win_std_dev[525]), .feature_accum(feature_accums[525]));
  accum_calculator #(.RECT1_X(rectangle1_xs[526]), .RECT1_Y(rectangle1_ys[526]), .RECT1_WIDTH(rectangle1_widths[526]), .RECT1_HEIGHT(rectangle1_heights[526]), .RECT1_WEIGHT(rectangle1_weights[526]), .RECT2_X(rectangle2_xs[526]), .RECT2_Y(rectangle2_ys[526]), .RECT2_WIDTH(rectangle2_widths[526]), .RECT2_HEIGHT(rectangle2_heights[526]), .RECT2_WEIGHT(rectangle2_weights[526]), .RECT3_X(rectangle3_xs[526]), .RECT3_Y(rectangle3_ys[526]), .RECT3_WIDTH(rectangle3_widths[526]), .RECT3_HEIGHT(rectangle3_heights[526]), .RECT3_WEIGHT(rectangle3_weights[526]), .FEAT_THRES(feature_thresholds[526]), .FEAT_ABOVE(feature_aboves[526]), .FEAT_BELOW(feature_belows[526])) ac526(.scan_win(scan_win526), .scan_win_std_dev(scan_win_std_dev[526]), .feature_accum(feature_accums[526]));
  accum_calculator #(.RECT1_X(rectangle1_xs[527]), .RECT1_Y(rectangle1_ys[527]), .RECT1_WIDTH(rectangle1_widths[527]), .RECT1_HEIGHT(rectangle1_heights[527]), .RECT1_WEIGHT(rectangle1_weights[527]), .RECT2_X(rectangle2_xs[527]), .RECT2_Y(rectangle2_ys[527]), .RECT2_WIDTH(rectangle2_widths[527]), .RECT2_HEIGHT(rectangle2_heights[527]), .RECT2_WEIGHT(rectangle2_weights[527]), .RECT3_X(rectangle3_xs[527]), .RECT3_Y(rectangle3_ys[527]), .RECT3_WIDTH(rectangle3_widths[527]), .RECT3_HEIGHT(rectangle3_heights[527]), .RECT3_WEIGHT(rectangle3_weights[527]), .FEAT_THRES(feature_thresholds[527]), .FEAT_ABOVE(feature_aboves[527]), .FEAT_BELOW(feature_belows[527])) ac527(.scan_win(scan_win527), .scan_win_std_dev(scan_win_std_dev[527]), .feature_accum(feature_accums[527]));
  accum_calculator #(.RECT1_X(rectangle1_xs[528]), .RECT1_Y(rectangle1_ys[528]), .RECT1_WIDTH(rectangle1_widths[528]), .RECT1_HEIGHT(rectangle1_heights[528]), .RECT1_WEIGHT(rectangle1_weights[528]), .RECT2_X(rectangle2_xs[528]), .RECT2_Y(rectangle2_ys[528]), .RECT2_WIDTH(rectangle2_widths[528]), .RECT2_HEIGHT(rectangle2_heights[528]), .RECT2_WEIGHT(rectangle2_weights[528]), .RECT3_X(rectangle3_xs[528]), .RECT3_Y(rectangle3_ys[528]), .RECT3_WIDTH(rectangle3_widths[528]), .RECT3_HEIGHT(rectangle3_heights[528]), .RECT3_WEIGHT(rectangle3_weights[528]), .FEAT_THRES(feature_thresholds[528]), .FEAT_ABOVE(feature_aboves[528]), .FEAT_BELOW(feature_belows[528])) ac528(.scan_win(scan_win528), .scan_win_std_dev(scan_win_std_dev[528]), .feature_accum(feature_accums[528]));
  accum_calculator #(.RECT1_X(rectangle1_xs[529]), .RECT1_Y(rectangle1_ys[529]), .RECT1_WIDTH(rectangle1_widths[529]), .RECT1_HEIGHT(rectangle1_heights[529]), .RECT1_WEIGHT(rectangle1_weights[529]), .RECT2_X(rectangle2_xs[529]), .RECT2_Y(rectangle2_ys[529]), .RECT2_WIDTH(rectangle2_widths[529]), .RECT2_HEIGHT(rectangle2_heights[529]), .RECT2_WEIGHT(rectangle2_weights[529]), .RECT3_X(rectangle3_xs[529]), .RECT3_Y(rectangle3_ys[529]), .RECT3_WIDTH(rectangle3_widths[529]), .RECT3_HEIGHT(rectangle3_heights[529]), .RECT3_WEIGHT(rectangle3_weights[529]), .FEAT_THRES(feature_thresholds[529]), .FEAT_ABOVE(feature_aboves[529]), .FEAT_BELOW(feature_belows[529])) ac529(.scan_win(scan_win529), .scan_win_std_dev(scan_win_std_dev[529]), .feature_accum(feature_accums[529]));
  accum_calculator #(.RECT1_X(rectangle1_xs[530]), .RECT1_Y(rectangle1_ys[530]), .RECT1_WIDTH(rectangle1_widths[530]), .RECT1_HEIGHT(rectangle1_heights[530]), .RECT1_WEIGHT(rectangle1_weights[530]), .RECT2_X(rectangle2_xs[530]), .RECT2_Y(rectangle2_ys[530]), .RECT2_WIDTH(rectangle2_widths[530]), .RECT2_HEIGHT(rectangle2_heights[530]), .RECT2_WEIGHT(rectangle2_weights[530]), .RECT3_X(rectangle3_xs[530]), .RECT3_Y(rectangle3_ys[530]), .RECT3_WIDTH(rectangle3_widths[530]), .RECT3_HEIGHT(rectangle3_heights[530]), .RECT3_WEIGHT(rectangle3_weights[530]), .FEAT_THRES(feature_thresholds[530]), .FEAT_ABOVE(feature_aboves[530]), .FEAT_BELOW(feature_belows[530])) ac530(.scan_win(scan_win530), .scan_win_std_dev(scan_win_std_dev[530]), .feature_accum(feature_accums[530]));
  accum_calculator #(.RECT1_X(rectangle1_xs[531]), .RECT1_Y(rectangle1_ys[531]), .RECT1_WIDTH(rectangle1_widths[531]), .RECT1_HEIGHT(rectangle1_heights[531]), .RECT1_WEIGHT(rectangle1_weights[531]), .RECT2_X(rectangle2_xs[531]), .RECT2_Y(rectangle2_ys[531]), .RECT2_WIDTH(rectangle2_widths[531]), .RECT2_HEIGHT(rectangle2_heights[531]), .RECT2_WEIGHT(rectangle2_weights[531]), .RECT3_X(rectangle3_xs[531]), .RECT3_Y(rectangle3_ys[531]), .RECT3_WIDTH(rectangle3_widths[531]), .RECT3_HEIGHT(rectangle3_heights[531]), .RECT3_WEIGHT(rectangle3_weights[531]), .FEAT_THRES(feature_thresholds[531]), .FEAT_ABOVE(feature_aboves[531]), .FEAT_BELOW(feature_belows[531])) ac531(.scan_win(scan_win531), .scan_win_std_dev(scan_win_std_dev[531]), .feature_accum(feature_accums[531]));
  accum_calculator #(.RECT1_X(rectangle1_xs[532]), .RECT1_Y(rectangle1_ys[532]), .RECT1_WIDTH(rectangle1_widths[532]), .RECT1_HEIGHT(rectangle1_heights[532]), .RECT1_WEIGHT(rectangle1_weights[532]), .RECT2_X(rectangle2_xs[532]), .RECT2_Y(rectangle2_ys[532]), .RECT2_WIDTH(rectangle2_widths[532]), .RECT2_HEIGHT(rectangle2_heights[532]), .RECT2_WEIGHT(rectangle2_weights[532]), .RECT3_X(rectangle3_xs[532]), .RECT3_Y(rectangle3_ys[532]), .RECT3_WIDTH(rectangle3_widths[532]), .RECT3_HEIGHT(rectangle3_heights[532]), .RECT3_WEIGHT(rectangle3_weights[532]), .FEAT_THRES(feature_thresholds[532]), .FEAT_ABOVE(feature_aboves[532]), .FEAT_BELOW(feature_belows[532])) ac532(.scan_win(scan_win532), .scan_win_std_dev(scan_win_std_dev[532]), .feature_accum(feature_accums[532]));
  accum_calculator #(.RECT1_X(rectangle1_xs[533]), .RECT1_Y(rectangle1_ys[533]), .RECT1_WIDTH(rectangle1_widths[533]), .RECT1_HEIGHT(rectangle1_heights[533]), .RECT1_WEIGHT(rectangle1_weights[533]), .RECT2_X(rectangle2_xs[533]), .RECT2_Y(rectangle2_ys[533]), .RECT2_WIDTH(rectangle2_widths[533]), .RECT2_HEIGHT(rectangle2_heights[533]), .RECT2_WEIGHT(rectangle2_weights[533]), .RECT3_X(rectangle3_xs[533]), .RECT3_Y(rectangle3_ys[533]), .RECT3_WIDTH(rectangle3_widths[533]), .RECT3_HEIGHT(rectangle3_heights[533]), .RECT3_WEIGHT(rectangle3_weights[533]), .FEAT_THRES(feature_thresholds[533]), .FEAT_ABOVE(feature_aboves[533]), .FEAT_BELOW(feature_belows[533])) ac533(.scan_win(scan_win533), .scan_win_std_dev(scan_win_std_dev[533]), .feature_accum(feature_accums[533]));
  accum_calculator #(.RECT1_X(rectangle1_xs[534]), .RECT1_Y(rectangle1_ys[534]), .RECT1_WIDTH(rectangle1_widths[534]), .RECT1_HEIGHT(rectangle1_heights[534]), .RECT1_WEIGHT(rectangle1_weights[534]), .RECT2_X(rectangle2_xs[534]), .RECT2_Y(rectangle2_ys[534]), .RECT2_WIDTH(rectangle2_widths[534]), .RECT2_HEIGHT(rectangle2_heights[534]), .RECT2_WEIGHT(rectangle2_weights[534]), .RECT3_X(rectangle3_xs[534]), .RECT3_Y(rectangle3_ys[534]), .RECT3_WIDTH(rectangle3_widths[534]), .RECT3_HEIGHT(rectangle3_heights[534]), .RECT3_WEIGHT(rectangle3_weights[534]), .FEAT_THRES(feature_thresholds[534]), .FEAT_ABOVE(feature_aboves[534]), .FEAT_BELOW(feature_belows[534])) ac534(.scan_win(scan_win534), .scan_win_std_dev(scan_win_std_dev[534]), .feature_accum(feature_accums[534]));
  accum_calculator #(.RECT1_X(rectangle1_xs[535]), .RECT1_Y(rectangle1_ys[535]), .RECT1_WIDTH(rectangle1_widths[535]), .RECT1_HEIGHT(rectangle1_heights[535]), .RECT1_WEIGHT(rectangle1_weights[535]), .RECT2_X(rectangle2_xs[535]), .RECT2_Y(rectangle2_ys[535]), .RECT2_WIDTH(rectangle2_widths[535]), .RECT2_HEIGHT(rectangle2_heights[535]), .RECT2_WEIGHT(rectangle2_weights[535]), .RECT3_X(rectangle3_xs[535]), .RECT3_Y(rectangle3_ys[535]), .RECT3_WIDTH(rectangle3_widths[535]), .RECT3_HEIGHT(rectangle3_heights[535]), .RECT3_WEIGHT(rectangle3_weights[535]), .FEAT_THRES(feature_thresholds[535]), .FEAT_ABOVE(feature_aboves[535]), .FEAT_BELOW(feature_belows[535])) ac535(.scan_win(scan_win535), .scan_win_std_dev(scan_win_std_dev[535]), .feature_accum(feature_accums[535]));
  accum_calculator #(.RECT1_X(rectangle1_xs[536]), .RECT1_Y(rectangle1_ys[536]), .RECT1_WIDTH(rectangle1_widths[536]), .RECT1_HEIGHT(rectangle1_heights[536]), .RECT1_WEIGHT(rectangle1_weights[536]), .RECT2_X(rectangle2_xs[536]), .RECT2_Y(rectangle2_ys[536]), .RECT2_WIDTH(rectangle2_widths[536]), .RECT2_HEIGHT(rectangle2_heights[536]), .RECT2_WEIGHT(rectangle2_weights[536]), .RECT3_X(rectangle3_xs[536]), .RECT3_Y(rectangle3_ys[536]), .RECT3_WIDTH(rectangle3_widths[536]), .RECT3_HEIGHT(rectangle3_heights[536]), .RECT3_WEIGHT(rectangle3_weights[536]), .FEAT_THRES(feature_thresholds[536]), .FEAT_ABOVE(feature_aboves[536]), .FEAT_BELOW(feature_belows[536])) ac536(.scan_win(scan_win536), .scan_win_std_dev(scan_win_std_dev[536]), .feature_accum(feature_accums[536]));
  accum_calculator #(.RECT1_X(rectangle1_xs[537]), .RECT1_Y(rectangle1_ys[537]), .RECT1_WIDTH(rectangle1_widths[537]), .RECT1_HEIGHT(rectangle1_heights[537]), .RECT1_WEIGHT(rectangle1_weights[537]), .RECT2_X(rectangle2_xs[537]), .RECT2_Y(rectangle2_ys[537]), .RECT2_WIDTH(rectangle2_widths[537]), .RECT2_HEIGHT(rectangle2_heights[537]), .RECT2_WEIGHT(rectangle2_weights[537]), .RECT3_X(rectangle3_xs[537]), .RECT3_Y(rectangle3_ys[537]), .RECT3_WIDTH(rectangle3_widths[537]), .RECT3_HEIGHT(rectangle3_heights[537]), .RECT3_WEIGHT(rectangle3_weights[537]), .FEAT_THRES(feature_thresholds[537]), .FEAT_ABOVE(feature_aboves[537]), .FEAT_BELOW(feature_belows[537])) ac537(.scan_win(scan_win537), .scan_win_std_dev(scan_win_std_dev[537]), .feature_accum(feature_accums[537]));
  accum_calculator #(.RECT1_X(rectangle1_xs[538]), .RECT1_Y(rectangle1_ys[538]), .RECT1_WIDTH(rectangle1_widths[538]), .RECT1_HEIGHT(rectangle1_heights[538]), .RECT1_WEIGHT(rectangle1_weights[538]), .RECT2_X(rectangle2_xs[538]), .RECT2_Y(rectangle2_ys[538]), .RECT2_WIDTH(rectangle2_widths[538]), .RECT2_HEIGHT(rectangle2_heights[538]), .RECT2_WEIGHT(rectangle2_weights[538]), .RECT3_X(rectangle3_xs[538]), .RECT3_Y(rectangle3_ys[538]), .RECT3_WIDTH(rectangle3_widths[538]), .RECT3_HEIGHT(rectangle3_heights[538]), .RECT3_WEIGHT(rectangle3_weights[538]), .FEAT_THRES(feature_thresholds[538]), .FEAT_ABOVE(feature_aboves[538]), .FEAT_BELOW(feature_belows[538])) ac538(.scan_win(scan_win538), .scan_win_std_dev(scan_win_std_dev[538]), .feature_accum(feature_accums[538]));
  accum_calculator #(.RECT1_X(rectangle1_xs[539]), .RECT1_Y(rectangle1_ys[539]), .RECT1_WIDTH(rectangle1_widths[539]), .RECT1_HEIGHT(rectangle1_heights[539]), .RECT1_WEIGHT(rectangle1_weights[539]), .RECT2_X(rectangle2_xs[539]), .RECT2_Y(rectangle2_ys[539]), .RECT2_WIDTH(rectangle2_widths[539]), .RECT2_HEIGHT(rectangle2_heights[539]), .RECT2_WEIGHT(rectangle2_weights[539]), .RECT3_X(rectangle3_xs[539]), .RECT3_Y(rectangle3_ys[539]), .RECT3_WIDTH(rectangle3_widths[539]), .RECT3_HEIGHT(rectangle3_heights[539]), .RECT3_WEIGHT(rectangle3_weights[539]), .FEAT_THRES(feature_thresholds[539]), .FEAT_ABOVE(feature_aboves[539]), .FEAT_BELOW(feature_belows[539])) ac539(.scan_win(scan_win539), .scan_win_std_dev(scan_win_std_dev[539]), .feature_accum(feature_accums[539]));
  accum_calculator #(.RECT1_X(rectangle1_xs[540]), .RECT1_Y(rectangle1_ys[540]), .RECT1_WIDTH(rectangle1_widths[540]), .RECT1_HEIGHT(rectangle1_heights[540]), .RECT1_WEIGHT(rectangle1_weights[540]), .RECT2_X(rectangle2_xs[540]), .RECT2_Y(rectangle2_ys[540]), .RECT2_WIDTH(rectangle2_widths[540]), .RECT2_HEIGHT(rectangle2_heights[540]), .RECT2_WEIGHT(rectangle2_weights[540]), .RECT3_X(rectangle3_xs[540]), .RECT3_Y(rectangle3_ys[540]), .RECT3_WIDTH(rectangle3_widths[540]), .RECT3_HEIGHT(rectangle3_heights[540]), .RECT3_WEIGHT(rectangle3_weights[540]), .FEAT_THRES(feature_thresholds[540]), .FEAT_ABOVE(feature_aboves[540]), .FEAT_BELOW(feature_belows[540])) ac540(.scan_win(scan_win540), .scan_win_std_dev(scan_win_std_dev[540]), .feature_accum(feature_accums[540]));
  accum_calculator #(.RECT1_X(rectangle1_xs[541]), .RECT1_Y(rectangle1_ys[541]), .RECT1_WIDTH(rectangle1_widths[541]), .RECT1_HEIGHT(rectangle1_heights[541]), .RECT1_WEIGHT(rectangle1_weights[541]), .RECT2_X(rectangle2_xs[541]), .RECT2_Y(rectangle2_ys[541]), .RECT2_WIDTH(rectangle2_widths[541]), .RECT2_HEIGHT(rectangle2_heights[541]), .RECT2_WEIGHT(rectangle2_weights[541]), .RECT3_X(rectangle3_xs[541]), .RECT3_Y(rectangle3_ys[541]), .RECT3_WIDTH(rectangle3_widths[541]), .RECT3_HEIGHT(rectangle3_heights[541]), .RECT3_WEIGHT(rectangle3_weights[541]), .FEAT_THRES(feature_thresholds[541]), .FEAT_ABOVE(feature_aboves[541]), .FEAT_BELOW(feature_belows[541])) ac541(.scan_win(scan_win541), .scan_win_std_dev(scan_win_std_dev[541]), .feature_accum(feature_accums[541]));
  accum_calculator #(.RECT1_X(rectangle1_xs[542]), .RECT1_Y(rectangle1_ys[542]), .RECT1_WIDTH(rectangle1_widths[542]), .RECT1_HEIGHT(rectangle1_heights[542]), .RECT1_WEIGHT(rectangle1_weights[542]), .RECT2_X(rectangle2_xs[542]), .RECT2_Y(rectangle2_ys[542]), .RECT2_WIDTH(rectangle2_widths[542]), .RECT2_HEIGHT(rectangle2_heights[542]), .RECT2_WEIGHT(rectangle2_weights[542]), .RECT3_X(rectangle3_xs[542]), .RECT3_Y(rectangle3_ys[542]), .RECT3_WIDTH(rectangle3_widths[542]), .RECT3_HEIGHT(rectangle3_heights[542]), .RECT3_WEIGHT(rectangle3_weights[542]), .FEAT_THRES(feature_thresholds[542]), .FEAT_ABOVE(feature_aboves[542]), .FEAT_BELOW(feature_belows[542])) ac542(.scan_win(scan_win542), .scan_win_std_dev(scan_win_std_dev[542]), .feature_accum(feature_accums[542]));
  accum_calculator #(.RECT1_X(rectangle1_xs[543]), .RECT1_Y(rectangle1_ys[543]), .RECT1_WIDTH(rectangle1_widths[543]), .RECT1_HEIGHT(rectangle1_heights[543]), .RECT1_WEIGHT(rectangle1_weights[543]), .RECT2_X(rectangle2_xs[543]), .RECT2_Y(rectangle2_ys[543]), .RECT2_WIDTH(rectangle2_widths[543]), .RECT2_HEIGHT(rectangle2_heights[543]), .RECT2_WEIGHT(rectangle2_weights[543]), .RECT3_X(rectangle3_xs[543]), .RECT3_Y(rectangle3_ys[543]), .RECT3_WIDTH(rectangle3_widths[543]), .RECT3_HEIGHT(rectangle3_heights[543]), .RECT3_WEIGHT(rectangle3_weights[543]), .FEAT_THRES(feature_thresholds[543]), .FEAT_ABOVE(feature_aboves[543]), .FEAT_BELOW(feature_belows[543])) ac543(.scan_win(scan_win543), .scan_win_std_dev(scan_win_std_dev[543]), .feature_accum(feature_accums[543]));
  accum_calculator #(.RECT1_X(rectangle1_xs[544]), .RECT1_Y(rectangle1_ys[544]), .RECT1_WIDTH(rectangle1_widths[544]), .RECT1_HEIGHT(rectangle1_heights[544]), .RECT1_WEIGHT(rectangle1_weights[544]), .RECT2_X(rectangle2_xs[544]), .RECT2_Y(rectangle2_ys[544]), .RECT2_WIDTH(rectangle2_widths[544]), .RECT2_HEIGHT(rectangle2_heights[544]), .RECT2_WEIGHT(rectangle2_weights[544]), .RECT3_X(rectangle3_xs[544]), .RECT3_Y(rectangle3_ys[544]), .RECT3_WIDTH(rectangle3_widths[544]), .RECT3_HEIGHT(rectangle3_heights[544]), .RECT3_WEIGHT(rectangle3_weights[544]), .FEAT_THRES(feature_thresholds[544]), .FEAT_ABOVE(feature_aboves[544]), .FEAT_BELOW(feature_belows[544])) ac544(.scan_win(scan_win544), .scan_win_std_dev(scan_win_std_dev[544]), .feature_accum(feature_accums[544]));
  accum_calculator #(.RECT1_X(rectangle1_xs[545]), .RECT1_Y(rectangle1_ys[545]), .RECT1_WIDTH(rectangle1_widths[545]), .RECT1_HEIGHT(rectangle1_heights[545]), .RECT1_WEIGHT(rectangle1_weights[545]), .RECT2_X(rectangle2_xs[545]), .RECT2_Y(rectangle2_ys[545]), .RECT2_WIDTH(rectangle2_widths[545]), .RECT2_HEIGHT(rectangle2_heights[545]), .RECT2_WEIGHT(rectangle2_weights[545]), .RECT3_X(rectangle3_xs[545]), .RECT3_Y(rectangle3_ys[545]), .RECT3_WIDTH(rectangle3_widths[545]), .RECT3_HEIGHT(rectangle3_heights[545]), .RECT3_WEIGHT(rectangle3_weights[545]), .FEAT_THRES(feature_thresholds[545]), .FEAT_ABOVE(feature_aboves[545]), .FEAT_BELOW(feature_belows[545])) ac545(.scan_win(scan_win545), .scan_win_std_dev(scan_win_std_dev[545]), .feature_accum(feature_accums[545]));
  accum_calculator #(.RECT1_X(rectangle1_xs[546]), .RECT1_Y(rectangle1_ys[546]), .RECT1_WIDTH(rectangle1_widths[546]), .RECT1_HEIGHT(rectangle1_heights[546]), .RECT1_WEIGHT(rectangle1_weights[546]), .RECT2_X(rectangle2_xs[546]), .RECT2_Y(rectangle2_ys[546]), .RECT2_WIDTH(rectangle2_widths[546]), .RECT2_HEIGHT(rectangle2_heights[546]), .RECT2_WEIGHT(rectangle2_weights[546]), .RECT3_X(rectangle3_xs[546]), .RECT3_Y(rectangle3_ys[546]), .RECT3_WIDTH(rectangle3_widths[546]), .RECT3_HEIGHT(rectangle3_heights[546]), .RECT3_WEIGHT(rectangle3_weights[546]), .FEAT_THRES(feature_thresholds[546]), .FEAT_ABOVE(feature_aboves[546]), .FEAT_BELOW(feature_belows[546])) ac546(.scan_win(scan_win546), .scan_win_std_dev(scan_win_std_dev[546]), .feature_accum(feature_accums[546]));
  accum_calculator #(.RECT1_X(rectangle1_xs[547]), .RECT1_Y(rectangle1_ys[547]), .RECT1_WIDTH(rectangle1_widths[547]), .RECT1_HEIGHT(rectangle1_heights[547]), .RECT1_WEIGHT(rectangle1_weights[547]), .RECT2_X(rectangle2_xs[547]), .RECT2_Y(rectangle2_ys[547]), .RECT2_WIDTH(rectangle2_widths[547]), .RECT2_HEIGHT(rectangle2_heights[547]), .RECT2_WEIGHT(rectangle2_weights[547]), .RECT3_X(rectangle3_xs[547]), .RECT3_Y(rectangle3_ys[547]), .RECT3_WIDTH(rectangle3_widths[547]), .RECT3_HEIGHT(rectangle3_heights[547]), .RECT3_WEIGHT(rectangle3_weights[547]), .FEAT_THRES(feature_thresholds[547]), .FEAT_ABOVE(feature_aboves[547]), .FEAT_BELOW(feature_belows[547])) ac547(.scan_win(scan_win547), .scan_win_std_dev(scan_win_std_dev[547]), .feature_accum(feature_accums[547]));
  accum_calculator #(.RECT1_X(rectangle1_xs[548]), .RECT1_Y(rectangle1_ys[548]), .RECT1_WIDTH(rectangle1_widths[548]), .RECT1_HEIGHT(rectangle1_heights[548]), .RECT1_WEIGHT(rectangle1_weights[548]), .RECT2_X(rectangle2_xs[548]), .RECT2_Y(rectangle2_ys[548]), .RECT2_WIDTH(rectangle2_widths[548]), .RECT2_HEIGHT(rectangle2_heights[548]), .RECT2_WEIGHT(rectangle2_weights[548]), .RECT3_X(rectangle3_xs[548]), .RECT3_Y(rectangle3_ys[548]), .RECT3_WIDTH(rectangle3_widths[548]), .RECT3_HEIGHT(rectangle3_heights[548]), .RECT3_WEIGHT(rectangle3_weights[548]), .FEAT_THRES(feature_thresholds[548]), .FEAT_ABOVE(feature_aboves[548]), .FEAT_BELOW(feature_belows[548])) ac548(.scan_win(scan_win548), .scan_win_std_dev(scan_win_std_dev[548]), .feature_accum(feature_accums[548]));
  accum_calculator #(.RECT1_X(rectangle1_xs[549]), .RECT1_Y(rectangle1_ys[549]), .RECT1_WIDTH(rectangle1_widths[549]), .RECT1_HEIGHT(rectangle1_heights[549]), .RECT1_WEIGHT(rectangle1_weights[549]), .RECT2_X(rectangle2_xs[549]), .RECT2_Y(rectangle2_ys[549]), .RECT2_WIDTH(rectangle2_widths[549]), .RECT2_HEIGHT(rectangle2_heights[549]), .RECT2_WEIGHT(rectangle2_weights[549]), .RECT3_X(rectangle3_xs[549]), .RECT3_Y(rectangle3_ys[549]), .RECT3_WIDTH(rectangle3_widths[549]), .RECT3_HEIGHT(rectangle3_heights[549]), .RECT3_WEIGHT(rectangle3_weights[549]), .FEAT_THRES(feature_thresholds[549]), .FEAT_ABOVE(feature_aboves[549]), .FEAT_BELOW(feature_belows[549])) ac549(.scan_win(scan_win549), .scan_win_std_dev(scan_win_std_dev[549]), .feature_accum(feature_accums[549]));
  accum_calculator #(.RECT1_X(rectangle1_xs[550]), .RECT1_Y(rectangle1_ys[550]), .RECT1_WIDTH(rectangle1_widths[550]), .RECT1_HEIGHT(rectangle1_heights[550]), .RECT1_WEIGHT(rectangle1_weights[550]), .RECT2_X(rectangle2_xs[550]), .RECT2_Y(rectangle2_ys[550]), .RECT2_WIDTH(rectangle2_widths[550]), .RECT2_HEIGHT(rectangle2_heights[550]), .RECT2_WEIGHT(rectangle2_weights[550]), .RECT3_X(rectangle3_xs[550]), .RECT3_Y(rectangle3_ys[550]), .RECT3_WIDTH(rectangle3_widths[550]), .RECT3_HEIGHT(rectangle3_heights[550]), .RECT3_WEIGHT(rectangle3_weights[550]), .FEAT_THRES(feature_thresholds[550]), .FEAT_ABOVE(feature_aboves[550]), .FEAT_BELOW(feature_belows[550])) ac550(.scan_win(scan_win550), .scan_win_std_dev(scan_win_std_dev[550]), .feature_accum(feature_accums[550]));
  accum_calculator #(.RECT1_X(rectangle1_xs[551]), .RECT1_Y(rectangle1_ys[551]), .RECT1_WIDTH(rectangle1_widths[551]), .RECT1_HEIGHT(rectangle1_heights[551]), .RECT1_WEIGHT(rectangle1_weights[551]), .RECT2_X(rectangle2_xs[551]), .RECT2_Y(rectangle2_ys[551]), .RECT2_WIDTH(rectangle2_widths[551]), .RECT2_HEIGHT(rectangle2_heights[551]), .RECT2_WEIGHT(rectangle2_weights[551]), .RECT3_X(rectangle3_xs[551]), .RECT3_Y(rectangle3_ys[551]), .RECT3_WIDTH(rectangle3_widths[551]), .RECT3_HEIGHT(rectangle3_heights[551]), .RECT3_WEIGHT(rectangle3_weights[551]), .FEAT_THRES(feature_thresholds[551]), .FEAT_ABOVE(feature_aboves[551]), .FEAT_BELOW(feature_belows[551])) ac551(.scan_win(scan_win551), .scan_win_std_dev(scan_win_std_dev[551]), .feature_accum(feature_accums[551]));
  accum_calculator #(.RECT1_X(rectangle1_xs[552]), .RECT1_Y(rectangle1_ys[552]), .RECT1_WIDTH(rectangle1_widths[552]), .RECT1_HEIGHT(rectangle1_heights[552]), .RECT1_WEIGHT(rectangle1_weights[552]), .RECT2_X(rectangle2_xs[552]), .RECT2_Y(rectangle2_ys[552]), .RECT2_WIDTH(rectangle2_widths[552]), .RECT2_HEIGHT(rectangle2_heights[552]), .RECT2_WEIGHT(rectangle2_weights[552]), .RECT3_X(rectangle3_xs[552]), .RECT3_Y(rectangle3_ys[552]), .RECT3_WIDTH(rectangle3_widths[552]), .RECT3_HEIGHT(rectangle3_heights[552]), .RECT3_WEIGHT(rectangle3_weights[552]), .FEAT_THRES(feature_thresholds[552]), .FEAT_ABOVE(feature_aboves[552]), .FEAT_BELOW(feature_belows[552])) ac552(.scan_win(scan_win552), .scan_win_std_dev(scan_win_std_dev[552]), .feature_accum(feature_accums[552]));
  accum_calculator #(.RECT1_X(rectangle1_xs[553]), .RECT1_Y(rectangle1_ys[553]), .RECT1_WIDTH(rectangle1_widths[553]), .RECT1_HEIGHT(rectangle1_heights[553]), .RECT1_WEIGHT(rectangle1_weights[553]), .RECT2_X(rectangle2_xs[553]), .RECT2_Y(rectangle2_ys[553]), .RECT2_WIDTH(rectangle2_widths[553]), .RECT2_HEIGHT(rectangle2_heights[553]), .RECT2_WEIGHT(rectangle2_weights[553]), .RECT3_X(rectangle3_xs[553]), .RECT3_Y(rectangle3_ys[553]), .RECT3_WIDTH(rectangle3_widths[553]), .RECT3_HEIGHT(rectangle3_heights[553]), .RECT3_WEIGHT(rectangle3_weights[553]), .FEAT_THRES(feature_thresholds[553]), .FEAT_ABOVE(feature_aboves[553]), .FEAT_BELOW(feature_belows[553])) ac553(.scan_win(scan_win553), .scan_win_std_dev(scan_win_std_dev[553]), .feature_accum(feature_accums[553]));
  accum_calculator #(.RECT1_X(rectangle1_xs[554]), .RECT1_Y(rectangle1_ys[554]), .RECT1_WIDTH(rectangle1_widths[554]), .RECT1_HEIGHT(rectangle1_heights[554]), .RECT1_WEIGHT(rectangle1_weights[554]), .RECT2_X(rectangle2_xs[554]), .RECT2_Y(rectangle2_ys[554]), .RECT2_WIDTH(rectangle2_widths[554]), .RECT2_HEIGHT(rectangle2_heights[554]), .RECT2_WEIGHT(rectangle2_weights[554]), .RECT3_X(rectangle3_xs[554]), .RECT3_Y(rectangle3_ys[554]), .RECT3_WIDTH(rectangle3_widths[554]), .RECT3_HEIGHT(rectangle3_heights[554]), .RECT3_WEIGHT(rectangle3_weights[554]), .FEAT_THRES(feature_thresholds[554]), .FEAT_ABOVE(feature_aboves[554]), .FEAT_BELOW(feature_belows[554])) ac554(.scan_win(scan_win554), .scan_win_std_dev(scan_win_std_dev[554]), .feature_accum(feature_accums[554]));
  accum_calculator #(.RECT1_X(rectangle1_xs[555]), .RECT1_Y(rectangle1_ys[555]), .RECT1_WIDTH(rectangle1_widths[555]), .RECT1_HEIGHT(rectangle1_heights[555]), .RECT1_WEIGHT(rectangle1_weights[555]), .RECT2_X(rectangle2_xs[555]), .RECT2_Y(rectangle2_ys[555]), .RECT2_WIDTH(rectangle2_widths[555]), .RECT2_HEIGHT(rectangle2_heights[555]), .RECT2_WEIGHT(rectangle2_weights[555]), .RECT3_X(rectangle3_xs[555]), .RECT3_Y(rectangle3_ys[555]), .RECT3_WIDTH(rectangle3_widths[555]), .RECT3_HEIGHT(rectangle3_heights[555]), .RECT3_WEIGHT(rectangle3_weights[555]), .FEAT_THRES(feature_thresholds[555]), .FEAT_ABOVE(feature_aboves[555]), .FEAT_BELOW(feature_belows[555])) ac555(.scan_win(scan_win555), .scan_win_std_dev(scan_win_std_dev[555]), .feature_accum(feature_accums[555]));
  accum_calculator #(.RECT1_X(rectangle1_xs[556]), .RECT1_Y(rectangle1_ys[556]), .RECT1_WIDTH(rectangle1_widths[556]), .RECT1_HEIGHT(rectangle1_heights[556]), .RECT1_WEIGHT(rectangle1_weights[556]), .RECT2_X(rectangle2_xs[556]), .RECT2_Y(rectangle2_ys[556]), .RECT2_WIDTH(rectangle2_widths[556]), .RECT2_HEIGHT(rectangle2_heights[556]), .RECT2_WEIGHT(rectangle2_weights[556]), .RECT3_X(rectangle3_xs[556]), .RECT3_Y(rectangle3_ys[556]), .RECT3_WIDTH(rectangle3_widths[556]), .RECT3_HEIGHT(rectangle3_heights[556]), .RECT3_WEIGHT(rectangle3_weights[556]), .FEAT_THRES(feature_thresholds[556]), .FEAT_ABOVE(feature_aboves[556]), .FEAT_BELOW(feature_belows[556])) ac556(.scan_win(scan_win556), .scan_win_std_dev(scan_win_std_dev[556]), .feature_accum(feature_accums[556]));
  accum_calculator #(.RECT1_X(rectangle1_xs[557]), .RECT1_Y(rectangle1_ys[557]), .RECT1_WIDTH(rectangle1_widths[557]), .RECT1_HEIGHT(rectangle1_heights[557]), .RECT1_WEIGHT(rectangle1_weights[557]), .RECT2_X(rectangle2_xs[557]), .RECT2_Y(rectangle2_ys[557]), .RECT2_WIDTH(rectangle2_widths[557]), .RECT2_HEIGHT(rectangle2_heights[557]), .RECT2_WEIGHT(rectangle2_weights[557]), .RECT3_X(rectangle3_xs[557]), .RECT3_Y(rectangle3_ys[557]), .RECT3_WIDTH(rectangle3_widths[557]), .RECT3_HEIGHT(rectangle3_heights[557]), .RECT3_WEIGHT(rectangle3_weights[557]), .FEAT_THRES(feature_thresholds[557]), .FEAT_ABOVE(feature_aboves[557]), .FEAT_BELOW(feature_belows[557])) ac557(.scan_win(scan_win557), .scan_win_std_dev(scan_win_std_dev[557]), .feature_accum(feature_accums[557]));
  accum_calculator #(.RECT1_X(rectangle1_xs[558]), .RECT1_Y(rectangle1_ys[558]), .RECT1_WIDTH(rectangle1_widths[558]), .RECT1_HEIGHT(rectangle1_heights[558]), .RECT1_WEIGHT(rectangle1_weights[558]), .RECT2_X(rectangle2_xs[558]), .RECT2_Y(rectangle2_ys[558]), .RECT2_WIDTH(rectangle2_widths[558]), .RECT2_HEIGHT(rectangle2_heights[558]), .RECT2_WEIGHT(rectangle2_weights[558]), .RECT3_X(rectangle3_xs[558]), .RECT3_Y(rectangle3_ys[558]), .RECT3_WIDTH(rectangle3_widths[558]), .RECT3_HEIGHT(rectangle3_heights[558]), .RECT3_WEIGHT(rectangle3_weights[558]), .FEAT_THRES(feature_thresholds[558]), .FEAT_ABOVE(feature_aboves[558]), .FEAT_BELOW(feature_belows[558])) ac558(.scan_win(scan_win558), .scan_win_std_dev(scan_win_std_dev[558]), .feature_accum(feature_accums[558]));
  accum_calculator #(.RECT1_X(rectangle1_xs[559]), .RECT1_Y(rectangle1_ys[559]), .RECT1_WIDTH(rectangle1_widths[559]), .RECT1_HEIGHT(rectangle1_heights[559]), .RECT1_WEIGHT(rectangle1_weights[559]), .RECT2_X(rectangle2_xs[559]), .RECT2_Y(rectangle2_ys[559]), .RECT2_WIDTH(rectangle2_widths[559]), .RECT2_HEIGHT(rectangle2_heights[559]), .RECT2_WEIGHT(rectangle2_weights[559]), .RECT3_X(rectangle3_xs[559]), .RECT3_Y(rectangle3_ys[559]), .RECT3_WIDTH(rectangle3_widths[559]), .RECT3_HEIGHT(rectangle3_heights[559]), .RECT3_WEIGHT(rectangle3_weights[559]), .FEAT_THRES(feature_thresholds[559]), .FEAT_ABOVE(feature_aboves[559]), .FEAT_BELOW(feature_belows[559])) ac559(.scan_win(scan_win559), .scan_win_std_dev(scan_win_std_dev[559]), .feature_accum(feature_accums[559]));
  accum_calculator #(.RECT1_X(rectangle1_xs[560]), .RECT1_Y(rectangle1_ys[560]), .RECT1_WIDTH(rectangle1_widths[560]), .RECT1_HEIGHT(rectangle1_heights[560]), .RECT1_WEIGHT(rectangle1_weights[560]), .RECT2_X(rectangle2_xs[560]), .RECT2_Y(rectangle2_ys[560]), .RECT2_WIDTH(rectangle2_widths[560]), .RECT2_HEIGHT(rectangle2_heights[560]), .RECT2_WEIGHT(rectangle2_weights[560]), .RECT3_X(rectangle3_xs[560]), .RECT3_Y(rectangle3_ys[560]), .RECT3_WIDTH(rectangle3_widths[560]), .RECT3_HEIGHT(rectangle3_heights[560]), .RECT3_WEIGHT(rectangle3_weights[560]), .FEAT_THRES(feature_thresholds[560]), .FEAT_ABOVE(feature_aboves[560]), .FEAT_BELOW(feature_belows[560])) ac560(.scan_win(scan_win560), .scan_win_std_dev(scan_win_std_dev[560]), .feature_accum(feature_accums[560]));
  accum_calculator #(.RECT1_X(rectangle1_xs[561]), .RECT1_Y(rectangle1_ys[561]), .RECT1_WIDTH(rectangle1_widths[561]), .RECT1_HEIGHT(rectangle1_heights[561]), .RECT1_WEIGHT(rectangle1_weights[561]), .RECT2_X(rectangle2_xs[561]), .RECT2_Y(rectangle2_ys[561]), .RECT2_WIDTH(rectangle2_widths[561]), .RECT2_HEIGHT(rectangle2_heights[561]), .RECT2_WEIGHT(rectangle2_weights[561]), .RECT3_X(rectangle3_xs[561]), .RECT3_Y(rectangle3_ys[561]), .RECT3_WIDTH(rectangle3_widths[561]), .RECT3_HEIGHT(rectangle3_heights[561]), .RECT3_WEIGHT(rectangle3_weights[561]), .FEAT_THRES(feature_thresholds[561]), .FEAT_ABOVE(feature_aboves[561]), .FEAT_BELOW(feature_belows[561])) ac561(.scan_win(scan_win561), .scan_win_std_dev(scan_win_std_dev[561]), .feature_accum(feature_accums[561]));
  accum_calculator #(.RECT1_X(rectangle1_xs[562]), .RECT1_Y(rectangle1_ys[562]), .RECT1_WIDTH(rectangle1_widths[562]), .RECT1_HEIGHT(rectangle1_heights[562]), .RECT1_WEIGHT(rectangle1_weights[562]), .RECT2_X(rectangle2_xs[562]), .RECT2_Y(rectangle2_ys[562]), .RECT2_WIDTH(rectangle2_widths[562]), .RECT2_HEIGHT(rectangle2_heights[562]), .RECT2_WEIGHT(rectangle2_weights[562]), .RECT3_X(rectangle3_xs[562]), .RECT3_Y(rectangle3_ys[562]), .RECT3_WIDTH(rectangle3_widths[562]), .RECT3_HEIGHT(rectangle3_heights[562]), .RECT3_WEIGHT(rectangle3_weights[562]), .FEAT_THRES(feature_thresholds[562]), .FEAT_ABOVE(feature_aboves[562]), .FEAT_BELOW(feature_belows[562])) ac562(.scan_win(scan_win562), .scan_win_std_dev(scan_win_std_dev[562]), .feature_accum(feature_accums[562]));
  accum_calculator #(.RECT1_X(rectangle1_xs[563]), .RECT1_Y(rectangle1_ys[563]), .RECT1_WIDTH(rectangle1_widths[563]), .RECT1_HEIGHT(rectangle1_heights[563]), .RECT1_WEIGHT(rectangle1_weights[563]), .RECT2_X(rectangle2_xs[563]), .RECT2_Y(rectangle2_ys[563]), .RECT2_WIDTH(rectangle2_widths[563]), .RECT2_HEIGHT(rectangle2_heights[563]), .RECT2_WEIGHT(rectangle2_weights[563]), .RECT3_X(rectangle3_xs[563]), .RECT3_Y(rectangle3_ys[563]), .RECT3_WIDTH(rectangle3_widths[563]), .RECT3_HEIGHT(rectangle3_heights[563]), .RECT3_WEIGHT(rectangle3_weights[563]), .FEAT_THRES(feature_thresholds[563]), .FEAT_ABOVE(feature_aboves[563]), .FEAT_BELOW(feature_belows[563])) ac563(.scan_win(scan_win563), .scan_win_std_dev(scan_win_std_dev[563]), .feature_accum(feature_accums[563]));
  accum_calculator #(.RECT1_X(rectangle1_xs[564]), .RECT1_Y(rectangle1_ys[564]), .RECT1_WIDTH(rectangle1_widths[564]), .RECT1_HEIGHT(rectangle1_heights[564]), .RECT1_WEIGHT(rectangle1_weights[564]), .RECT2_X(rectangle2_xs[564]), .RECT2_Y(rectangle2_ys[564]), .RECT2_WIDTH(rectangle2_widths[564]), .RECT2_HEIGHT(rectangle2_heights[564]), .RECT2_WEIGHT(rectangle2_weights[564]), .RECT3_X(rectangle3_xs[564]), .RECT3_Y(rectangle3_ys[564]), .RECT3_WIDTH(rectangle3_widths[564]), .RECT3_HEIGHT(rectangle3_heights[564]), .RECT3_WEIGHT(rectangle3_weights[564]), .FEAT_THRES(feature_thresholds[564]), .FEAT_ABOVE(feature_aboves[564]), .FEAT_BELOW(feature_belows[564])) ac564(.scan_win(scan_win564), .scan_win_std_dev(scan_win_std_dev[564]), .feature_accum(feature_accums[564]));
  accum_calculator #(.RECT1_X(rectangle1_xs[565]), .RECT1_Y(rectangle1_ys[565]), .RECT1_WIDTH(rectangle1_widths[565]), .RECT1_HEIGHT(rectangle1_heights[565]), .RECT1_WEIGHT(rectangle1_weights[565]), .RECT2_X(rectangle2_xs[565]), .RECT2_Y(rectangle2_ys[565]), .RECT2_WIDTH(rectangle2_widths[565]), .RECT2_HEIGHT(rectangle2_heights[565]), .RECT2_WEIGHT(rectangle2_weights[565]), .RECT3_X(rectangle3_xs[565]), .RECT3_Y(rectangle3_ys[565]), .RECT3_WIDTH(rectangle3_widths[565]), .RECT3_HEIGHT(rectangle3_heights[565]), .RECT3_WEIGHT(rectangle3_weights[565]), .FEAT_THRES(feature_thresholds[565]), .FEAT_ABOVE(feature_aboves[565]), .FEAT_BELOW(feature_belows[565])) ac565(.scan_win(scan_win565), .scan_win_std_dev(scan_win_std_dev[565]), .feature_accum(feature_accums[565]));
  accum_calculator #(.RECT1_X(rectangle1_xs[566]), .RECT1_Y(rectangle1_ys[566]), .RECT1_WIDTH(rectangle1_widths[566]), .RECT1_HEIGHT(rectangle1_heights[566]), .RECT1_WEIGHT(rectangle1_weights[566]), .RECT2_X(rectangle2_xs[566]), .RECT2_Y(rectangle2_ys[566]), .RECT2_WIDTH(rectangle2_widths[566]), .RECT2_HEIGHT(rectangle2_heights[566]), .RECT2_WEIGHT(rectangle2_weights[566]), .RECT3_X(rectangle3_xs[566]), .RECT3_Y(rectangle3_ys[566]), .RECT3_WIDTH(rectangle3_widths[566]), .RECT3_HEIGHT(rectangle3_heights[566]), .RECT3_WEIGHT(rectangle3_weights[566]), .FEAT_THRES(feature_thresholds[566]), .FEAT_ABOVE(feature_aboves[566]), .FEAT_BELOW(feature_belows[566])) ac566(.scan_win(scan_win566), .scan_win_std_dev(scan_win_std_dev[566]), .feature_accum(feature_accums[566]));
  accum_calculator #(.RECT1_X(rectangle1_xs[567]), .RECT1_Y(rectangle1_ys[567]), .RECT1_WIDTH(rectangle1_widths[567]), .RECT1_HEIGHT(rectangle1_heights[567]), .RECT1_WEIGHT(rectangle1_weights[567]), .RECT2_X(rectangle2_xs[567]), .RECT2_Y(rectangle2_ys[567]), .RECT2_WIDTH(rectangle2_widths[567]), .RECT2_HEIGHT(rectangle2_heights[567]), .RECT2_WEIGHT(rectangle2_weights[567]), .RECT3_X(rectangle3_xs[567]), .RECT3_Y(rectangle3_ys[567]), .RECT3_WIDTH(rectangle3_widths[567]), .RECT3_HEIGHT(rectangle3_heights[567]), .RECT3_WEIGHT(rectangle3_weights[567]), .FEAT_THRES(feature_thresholds[567]), .FEAT_ABOVE(feature_aboves[567]), .FEAT_BELOW(feature_belows[567])) ac567(.scan_win(scan_win567), .scan_win_std_dev(scan_win_std_dev[567]), .feature_accum(feature_accums[567]));
  accum_calculator #(.RECT1_X(rectangle1_xs[568]), .RECT1_Y(rectangle1_ys[568]), .RECT1_WIDTH(rectangle1_widths[568]), .RECT1_HEIGHT(rectangle1_heights[568]), .RECT1_WEIGHT(rectangle1_weights[568]), .RECT2_X(rectangle2_xs[568]), .RECT2_Y(rectangle2_ys[568]), .RECT2_WIDTH(rectangle2_widths[568]), .RECT2_HEIGHT(rectangle2_heights[568]), .RECT2_WEIGHT(rectangle2_weights[568]), .RECT3_X(rectangle3_xs[568]), .RECT3_Y(rectangle3_ys[568]), .RECT3_WIDTH(rectangle3_widths[568]), .RECT3_HEIGHT(rectangle3_heights[568]), .RECT3_WEIGHT(rectangle3_weights[568]), .FEAT_THRES(feature_thresholds[568]), .FEAT_ABOVE(feature_aboves[568]), .FEAT_BELOW(feature_belows[568])) ac568(.scan_win(scan_win568), .scan_win_std_dev(scan_win_std_dev[568]), .feature_accum(feature_accums[568]));
  accum_calculator #(.RECT1_X(rectangle1_xs[569]), .RECT1_Y(rectangle1_ys[569]), .RECT1_WIDTH(rectangle1_widths[569]), .RECT1_HEIGHT(rectangle1_heights[569]), .RECT1_WEIGHT(rectangle1_weights[569]), .RECT2_X(rectangle2_xs[569]), .RECT2_Y(rectangle2_ys[569]), .RECT2_WIDTH(rectangle2_widths[569]), .RECT2_HEIGHT(rectangle2_heights[569]), .RECT2_WEIGHT(rectangle2_weights[569]), .RECT3_X(rectangle3_xs[569]), .RECT3_Y(rectangle3_ys[569]), .RECT3_WIDTH(rectangle3_widths[569]), .RECT3_HEIGHT(rectangle3_heights[569]), .RECT3_WEIGHT(rectangle3_weights[569]), .FEAT_THRES(feature_thresholds[569]), .FEAT_ABOVE(feature_aboves[569]), .FEAT_BELOW(feature_belows[569])) ac569(.scan_win(scan_win569), .scan_win_std_dev(scan_win_std_dev[569]), .feature_accum(feature_accums[569]));
  accum_calculator #(.RECT1_X(rectangle1_xs[570]), .RECT1_Y(rectangle1_ys[570]), .RECT1_WIDTH(rectangle1_widths[570]), .RECT1_HEIGHT(rectangle1_heights[570]), .RECT1_WEIGHT(rectangle1_weights[570]), .RECT2_X(rectangle2_xs[570]), .RECT2_Y(rectangle2_ys[570]), .RECT2_WIDTH(rectangle2_widths[570]), .RECT2_HEIGHT(rectangle2_heights[570]), .RECT2_WEIGHT(rectangle2_weights[570]), .RECT3_X(rectangle3_xs[570]), .RECT3_Y(rectangle3_ys[570]), .RECT3_WIDTH(rectangle3_widths[570]), .RECT3_HEIGHT(rectangle3_heights[570]), .RECT3_WEIGHT(rectangle3_weights[570]), .FEAT_THRES(feature_thresholds[570]), .FEAT_ABOVE(feature_aboves[570]), .FEAT_BELOW(feature_belows[570])) ac570(.scan_win(scan_win570), .scan_win_std_dev(scan_win_std_dev[570]), .feature_accum(feature_accums[570]));
  accum_calculator #(.RECT1_X(rectangle1_xs[571]), .RECT1_Y(rectangle1_ys[571]), .RECT1_WIDTH(rectangle1_widths[571]), .RECT1_HEIGHT(rectangle1_heights[571]), .RECT1_WEIGHT(rectangle1_weights[571]), .RECT2_X(rectangle2_xs[571]), .RECT2_Y(rectangle2_ys[571]), .RECT2_WIDTH(rectangle2_widths[571]), .RECT2_HEIGHT(rectangle2_heights[571]), .RECT2_WEIGHT(rectangle2_weights[571]), .RECT3_X(rectangle3_xs[571]), .RECT3_Y(rectangle3_ys[571]), .RECT3_WIDTH(rectangle3_widths[571]), .RECT3_HEIGHT(rectangle3_heights[571]), .RECT3_WEIGHT(rectangle3_weights[571]), .FEAT_THRES(feature_thresholds[571]), .FEAT_ABOVE(feature_aboves[571]), .FEAT_BELOW(feature_belows[571])) ac571(.scan_win(scan_win571), .scan_win_std_dev(scan_win_std_dev[571]), .feature_accum(feature_accums[571]));
  accum_calculator #(.RECT1_X(rectangle1_xs[572]), .RECT1_Y(rectangle1_ys[572]), .RECT1_WIDTH(rectangle1_widths[572]), .RECT1_HEIGHT(rectangle1_heights[572]), .RECT1_WEIGHT(rectangle1_weights[572]), .RECT2_X(rectangle2_xs[572]), .RECT2_Y(rectangle2_ys[572]), .RECT2_WIDTH(rectangle2_widths[572]), .RECT2_HEIGHT(rectangle2_heights[572]), .RECT2_WEIGHT(rectangle2_weights[572]), .RECT3_X(rectangle3_xs[572]), .RECT3_Y(rectangle3_ys[572]), .RECT3_WIDTH(rectangle3_widths[572]), .RECT3_HEIGHT(rectangle3_heights[572]), .RECT3_WEIGHT(rectangle3_weights[572]), .FEAT_THRES(feature_thresholds[572]), .FEAT_ABOVE(feature_aboves[572]), .FEAT_BELOW(feature_belows[572])) ac572(.scan_win(scan_win572), .scan_win_std_dev(scan_win_std_dev[572]), .feature_accum(feature_accums[572]));
  accum_calculator #(.RECT1_X(rectangle1_xs[573]), .RECT1_Y(rectangle1_ys[573]), .RECT1_WIDTH(rectangle1_widths[573]), .RECT1_HEIGHT(rectangle1_heights[573]), .RECT1_WEIGHT(rectangle1_weights[573]), .RECT2_X(rectangle2_xs[573]), .RECT2_Y(rectangle2_ys[573]), .RECT2_WIDTH(rectangle2_widths[573]), .RECT2_HEIGHT(rectangle2_heights[573]), .RECT2_WEIGHT(rectangle2_weights[573]), .RECT3_X(rectangle3_xs[573]), .RECT3_Y(rectangle3_ys[573]), .RECT3_WIDTH(rectangle3_widths[573]), .RECT3_HEIGHT(rectangle3_heights[573]), .RECT3_WEIGHT(rectangle3_weights[573]), .FEAT_THRES(feature_thresholds[573]), .FEAT_ABOVE(feature_aboves[573]), .FEAT_BELOW(feature_belows[573])) ac573(.scan_win(scan_win573), .scan_win_std_dev(scan_win_std_dev[573]), .feature_accum(feature_accums[573]));
  accum_calculator #(.RECT1_X(rectangle1_xs[574]), .RECT1_Y(rectangle1_ys[574]), .RECT1_WIDTH(rectangle1_widths[574]), .RECT1_HEIGHT(rectangle1_heights[574]), .RECT1_WEIGHT(rectangle1_weights[574]), .RECT2_X(rectangle2_xs[574]), .RECT2_Y(rectangle2_ys[574]), .RECT2_WIDTH(rectangle2_widths[574]), .RECT2_HEIGHT(rectangle2_heights[574]), .RECT2_WEIGHT(rectangle2_weights[574]), .RECT3_X(rectangle3_xs[574]), .RECT3_Y(rectangle3_ys[574]), .RECT3_WIDTH(rectangle3_widths[574]), .RECT3_HEIGHT(rectangle3_heights[574]), .RECT3_WEIGHT(rectangle3_weights[574]), .FEAT_THRES(feature_thresholds[574]), .FEAT_ABOVE(feature_aboves[574]), .FEAT_BELOW(feature_belows[574])) ac574(.scan_win(scan_win574), .scan_win_std_dev(scan_win_std_dev[574]), .feature_accum(feature_accums[574]));
  accum_calculator #(.RECT1_X(rectangle1_xs[575]), .RECT1_Y(rectangle1_ys[575]), .RECT1_WIDTH(rectangle1_widths[575]), .RECT1_HEIGHT(rectangle1_heights[575]), .RECT1_WEIGHT(rectangle1_weights[575]), .RECT2_X(rectangle2_xs[575]), .RECT2_Y(rectangle2_ys[575]), .RECT2_WIDTH(rectangle2_widths[575]), .RECT2_HEIGHT(rectangle2_heights[575]), .RECT2_WEIGHT(rectangle2_weights[575]), .RECT3_X(rectangle3_xs[575]), .RECT3_Y(rectangle3_ys[575]), .RECT3_WIDTH(rectangle3_widths[575]), .RECT3_HEIGHT(rectangle3_heights[575]), .RECT3_WEIGHT(rectangle3_weights[575]), .FEAT_THRES(feature_thresholds[575]), .FEAT_ABOVE(feature_aboves[575]), .FEAT_BELOW(feature_belows[575])) ac575(.scan_win(scan_win575), .scan_win_std_dev(scan_win_std_dev[575]), .feature_accum(feature_accums[575]));
  accum_calculator #(.RECT1_X(rectangle1_xs[576]), .RECT1_Y(rectangle1_ys[576]), .RECT1_WIDTH(rectangle1_widths[576]), .RECT1_HEIGHT(rectangle1_heights[576]), .RECT1_WEIGHT(rectangle1_weights[576]), .RECT2_X(rectangle2_xs[576]), .RECT2_Y(rectangle2_ys[576]), .RECT2_WIDTH(rectangle2_widths[576]), .RECT2_HEIGHT(rectangle2_heights[576]), .RECT2_WEIGHT(rectangle2_weights[576]), .RECT3_X(rectangle3_xs[576]), .RECT3_Y(rectangle3_ys[576]), .RECT3_WIDTH(rectangle3_widths[576]), .RECT3_HEIGHT(rectangle3_heights[576]), .RECT3_WEIGHT(rectangle3_weights[576]), .FEAT_THRES(feature_thresholds[576]), .FEAT_ABOVE(feature_aboves[576]), .FEAT_BELOW(feature_belows[576])) ac576(.scan_win(scan_win576), .scan_win_std_dev(scan_win_std_dev[576]), .feature_accum(feature_accums[576]));
  accum_calculator #(.RECT1_X(rectangle1_xs[577]), .RECT1_Y(rectangle1_ys[577]), .RECT1_WIDTH(rectangle1_widths[577]), .RECT1_HEIGHT(rectangle1_heights[577]), .RECT1_WEIGHT(rectangle1_weights[577]), .RECT2_X(rectangle2_xs[577]), .RECT2_Y(rectangle2_ys[577]), .RECT2_WIDTH(rectangle2_widths[577]), .RECT2_HEIGHT(rectangle2_heights[577]), .RECT2_WEIGHT(rectangle2_weights[577]), .RECT3_X(rectangle3_xs[577]), .RECT3_Y(rectangle3_ys[577]), .RECT3_WIDTH(rectangle3_widths[577]), .RECT3_HEIGHT(rectangle3_heights[577]), .RECT3_WEIGHT(rectangle3_weights[577]), .FEAT_THRES(feature_thresholds[577]), .FEAT_ABOVE(feature_aboves[577]), .FEAT_BELOW(feature_belows[577])) ac577(.scan_win(scan_win577), .scan_win_std_dev(scan_win_std_dev[577]), .feature_accum(feature_accums[577]));
  accum_calculator #(.RECT1_X(rectangle1_xs[578]), .RECT1_Y(rectangle1_ys[578]), .RECT1_WIDTH(rectangle1_widths[578]), .RECT1_HEIGHT(rectangle1_heights[578]), .RECT1_WEIGHT(rectangle1_weights[578]), .RECT2_X(rectangle2_xs[578]), .RECT2_Y(rectangle2_ys[578]), .RECT2_WIDTH(rectangle2_widths[578]), .RECT2_HEIGHT(rectangle2_heights[578]), .RECT2_WEIGHT(rectangle2_weights[578]), .RECT3_X(rectangle3_xs[578]), .RECT3_Y(rectangle3_ys[578]), .RECT3_WIDTH(rectangle3_widths[578]), .RECT3_HEIGHT(rectangle3_heights[578]), .RECT3_WEIGHT(rectangle3_weights[578]), .FEAT_THRES(feature_thresholds[578]), .FEAT_ABOVE(feature_aboves[578]), .FEAT_BELOW(feature_belows[578])) ac578(.scan_win(scan_win578), .scan_win_std_dev(scan_win_std_dev[578]), .feature_accum(feature_accums[578]));
  accum_calculator #(.RECT1_X(rectangle1_xs[579]), .RECT1_Y(rectangle1_ys[579]), .RECT1_WIDTH(rectangle1_widths[579]), .RECT1_HEIGHT(rectangle1_heights[579]), .RECT1_WEIGHT(rectangle1_weights[579]), .RECT2_X(rectangle2_xs[579]), .RECT2_Y(rectangle2_ys[579]), .RECT2_WIDTH(rectangle2_widths[579]), .RECT2_HEIGHT(rectangle2_heights[579]), .RECT2_WEIGHT(rectangle2_weights[579]), .RECT3_X(rectangle3_xs[579]), .RECT3_Y(rectangle3_ys[579]), .RECT3_WIDTH(rectangle3_widths[579]), .RECT3_HEIGHT(rectangle3_heights[579]), .RECT3_WEIGHT(rectangle3_weights[579]), .FEAT_THRES(feature_thresholds[579]), .FEAT_ABOVE(feature_aboves[579]), .FEAT_BELOW(feature_belows[579])) ac579(.scan_win(scan_win579), .scan_win_std_dev(scan_win_std_dev[579]), .feature_accum(feature_accums[579]));
  accum_calculator #(.RECT1_X(rectangle1_xs[580]), .RECT1_Y(rectangle1_ys[580]), .RECT1_WIDTH(rectangle1_widths[580]), .RECT1_HEIGHT(rectangle1_heights[580]), .RECT1_WEIGHT(rectangle1_weights[580]), .RECT2_X(rectangle2_xs[580]), .RECT2_Y(rectangle2_ys[580]), .RECT2_WIDTH(rectangle2_widths[580]), .RECT2_HEIGHT(rectangle2_heights[580]), .RECT2_WEIGHT(rectangle2_weights[580]), .RECT3_X(rectangle3_xs[580]), .RECT3_Y(rectangle3_ys[580]), .RECT3_WIDTH(rectangle3_widths[580]), .RECT3_HEIGHT(rectangle3_heights[580]), .RECT3_WEIGHT(rectangle3_weights[580]), .FEAT_THRES(feature_thresholds[580]), .FEAT_ABOVE(feature_aboves[580]), .FEAT_BELOW(feature_belows[580])) ac580(.scan_win(scan_win580), .scan_win_std_dev(scan_win_std_dev[580]), .feature_accum(feature_accums[580]));
  accum_calculator #(.RECT1_X(rectangle1_xs[581]), .RECT1_Y(rectangle1_ys[581]), .RECT1_WIDTH(rectangle1_widths[581]), .RECT1_HEIGHT(rectangle1_heights[581]), .RECT1_WEIGHT(rectangle1_weights[581]), .RECT2_X(rectangle2_xs[581]), .RECT2_Y(rectangle2_ys[581]), .RECT2_WIDTH(rectangle2_widths[581]), .RECT2_HEIGHT(rectangle2_heights[581]), .RECT2_WEIGHT(rectangle2_weights[581]), .RECT3_X(rectangle3_xs[581]), .RECT3_Y(rectangle3_ys[581]), .RECT3_WIDTH(rectangle3_widths[581]), .RECT3_HEIGHT(rectangle3_heights[581]), .RECT3_WEIGHT(rectangle3_weights[581]), .FEAT_THRES(feature_thresholds[581]), .FEAT_ABOVE(feature_aboves[581]), .FEAT_BELOW(feature_belows[581])) ac581(.scan_win(scan_win581), .scan_win_std_dev(scan_win_std_dev[581]), .feature_accum(feature_accums[581]));
  accum_calculator #(.RECT1_X(rectangle1_xs[582]), .RECT1_Y(rectangle1_ys[582]), .RECT1_WIDTH(rectangle1_widths[582]), .RECT1_HEIGHT(rectangle1_heights[582]), .RECT1_WEIGHT(rectangle1_weights[582]), .RECT2_X(rectangle2_xs[582]), .RECT2_Y(rectangle2_ys[582]), .RECT2_WIDTH(rectangle2_widths[582]), .RECT2_HEIGHT(rectangle2_heights[582]), .RECT2_WEIGHT(rectangle2_weights[582]), .RECT3_X(rectangle3_xs[582]), .RECT3_Y(rectangle3_ys[582]), .RECT3_WIDTH(rectangle3_widths[582]), .RECT3_HEIGHT(rectangle3_heights[582]), .RECT3_WEIGHT(rectangle3_weights[582]), .FEAT_THRES(feature_thresholds[582]), .FEAT_ABOVE(feature_aboves[582]), .FEAT_BELOW(feature_belows[582])) ac582(.scan_win(scan_win582), .scan_win_std_dev(scan_win_std_dev[582]), .feature_accum(feature_accums[582]));
  accum_calculator #(.RECT1_X(rectangle1_xs[583]), .RECT1_Y(rectangle1_ys[583]), .RECT1_WIDTH(rectangle1_widths[583]), .RECT1_HEIGHT(rectangle1_heights[583]), .RECT1_WEIGHT(rectangle1_weights[583]), .RECT2_X(rectangle2_xs[583]), .RECT2_Y(rectangle2_ys[583]), .RECT2_WIDTH(rectangle2_widths[583]), .RECT2_HEIGHT(rectangle2_heights[583]), .RECT2_WEIGHT(rectangle2_weights[583]), .RECT3_X(rectangle3_xs[583]), .RECT3_Y(rectangle3_ys[583]), .RECT3_WIDTH(rectangle3_widths[583]), .RECT3_HEIGHT(rectangle3_heights[583]), .RECT3_WEIGHT(rectangle3_weights[583]), .FEAT_THRES(feature_thresholds[583]), .FEAT_ABOVE(feature_aboves[583]), .FEAT_BELOW(feature_belows[583])) ac583(.scan_win(scan_win583), .scan_win_std_dev(scan_win_std_dev[583]), .feature_accum(feature_accums[583]));
  accum_calculator #(.RECT1_X(rectangle1_xs[584]), .RECT1_Y(rectangle1_ys[584]), .RECT1_WIDTH(rectangle1_widths[584]), .RECT1_HEIGHT(rectangle1_heights[584]), .RECT1_WEIGHT(rectangle1_weights[584]), .RECT2_X(rectangle2_xs[584]), .RECT2_Y(rectangle2_ys[584]), .RECT2_WIDTH(rectangle2_widths[584]), .RECT2_HEIGHT(rectangle2_heights[584]), .RECT2_WEIGHT(rectangle2_weights[584]), .RECT3_X(rectangle3_xs[584]), .RECT3_Y(rectangle3_ys[584]), .RECT3_WIDTH(rectangle3_widths[584]), .RECT3_HEIGHT(rectangle3_heights[584]), .RECT3_WEIGHT(rectangle3_weights[584]), .FEAT_THRES(feature_thresholds[584]), .FEAT_ABOVE(feature_aboves[584]), .FEAT_BELOW(feature_belows[584])) ac584(.scan_win(scan_win584), .scan_win_std_dev(scan_win_std_dev[584]), .feature_accum(feature_accums[584]));
  accum_calculator #(.RECT1_X(rectangle1_xs[585]), .RECT1_Y(rectangle1_ys[585]), .RECT1_WIDTH(rectangle1_widths[585]), .RECT1_HEIGHT(rectangle1_heights[585]), .RECT1_WEIGHT(rectangle1_weights[585]), .RECT2_X(rectangle2_xs[585]), .RECT2_Y(rectangle2_ys[585]), .RECT2_WIDTH(rectangle2_widths[585]), .RECT2_HEIGHT(rectangle2_heights[585]), .RECT2_WEIGHT(rectangle2_weights[585]), .RECT3_X(rectangle3_xs[585]), .RECT3_Y(rectangle3_ys[585]), .RECT3_WIDTH(rectangle3_widths[585]), .RECT3_HEIGHT(rectangle3_heights[585]), .RECT3_WEIGHT(rectangle3_weights[585]), .FEAT_THRES(feature_thresholds[585]), .FEAT_ABOVE(feature_aboves[585]), .FEAT_BELOW(feature_belows[585])) ac585(.scan_win(scan_win585), .scan_win_std_dev(scan_win_std_dev[585]), .feature_accum(feature_accums[585]));
  accum_calculator #(.RECT1_X(rectangle1_xs[586]), .RECT1_Y(rectangle1_ys[586]), .RECT1_WIDTH(rectangle1_widths[586]), .RECT1_HEIGHT(rectangle1_heights[586]), .RECT1_WEIGHT(rectangle1_weights[586]), .RECT2_X(rectangle2_xs[586]), .RECT2_Y(rectangle2_ys[586]), .RECT2_WIDTH(rectangle2_widths[586]), .RECT2_HEIGHT(rectangle2_heights[586]), .RECT2_WEIGHT(rectangle2_weights[586]), .RECT3_X(rectangle3_xs[586]), .RECT3_Y(rectangle3_ys[586]), .RECT3_WIDTH(rectangle3_widths[586]), .RECT3_HEIGHT(rectangle3_heights[586]), .RECT3_WEIGHT(rectangle3_weights[586]), .FEAT_THRES(feature_thresholds[586]), .FEAT_ABOVE(feature_aboves[586]), .FEAT_BELOW(feature_belows[586])) ac586(.scan_win(scan_win586), .scan_win_std_dev(scan_win_std_dev[586]), .feature_accum(feature_accums[586]));
  accum_calculator #(.RECT1_X(rectangle1_xs[587]), .RECT1_Y(rectangle1_ys[587]), .RECT1_WIDTH(rectangle1_widths[587]), .RECT1_HEIGHT(rectangle1_heights[587]), .RECT1_WEIGHT(rectangle1_weights[587]), .RECT2_X(rectangle2_xs[587]), .RECT2_Y(rectangle2_ys[587]), .RECT2_WIDTH(rectangle2_widths[587]), .RECT2_HEIGHT(rectangle2_heights[587]), .RECT2_WEIGHT(rectangle2_weights[587]), .RECT3_X(rectangle3_xs[587]), .RECT3_Y(rectangle3_ys[587]), .RECT3_WIDTH(rectangle3_widths[587]), .RECT3_HEIGHT(rectangle3_heights[587]), .RECT3_WEIGHT(rectangle3_weights[587]), .FEAT_THRES(feature_thresholds[587]), .FEAT_ABOVE(feature_aboves[587]), .FEAT_BELOW(feature_belows[587])) ac587(.scan_win(scan_win587), .scan_win_std_dev(scan_win_std_dev[587]), .feature_accum(feature_accums[587]));
  accum_calculator #(.RECT1_X(rectangle1_xs[588]), .RECT1_Y(rectangle1_ys[588]), .RECT1_WIDTH(rectangle1_widths[588]), .RECT1_HEIGHT(rectangle1_heights[588]), .RECT1_WEIGHT(rectangle1_weights[588]), .RECT2_X(rectangle2_xs[588]), .RECT2_Y(rectangle2_ys[588]), .RECT2_WIDTH(rectangle2_widths[588]), .RECT2_HEIGHT(rectangle2_heights[588]), .RECT2_WEIGHT(rectangle2_weights[588]), .RECT3_X(rectangle3_xs[588]), .RECT3_Y(rectangle3_ys[588]), .RECT3_WIDTH(rectangle3_widths[588]), .RECT3_HEIGHT(rectangle3_heights[588]), .RECT3_WEIGHT(rectangle3_weights[588]), .FEAT_THRES(feature_thresholds[588]), .FEAT_ABOVE(feature_aboves[588]), .FEAT_BELOW(feature_belows[588])) ac588(.scan_win(scan_win588), .scan_win_std_dev(scan_win_std_dev[588]), .feature_accum(feature_accums[588]));
  accum_calculator #(.RECT1_X(rectangle1_xs[589]), .RECT1_Y(rectangle1_ys[589]), .RECT1_WIDTH(rectangle1_widths[589]), .RECT1_HEIGHT(rectangle1_heights[589]), .RECT1_WEIGHT(rectangle1_weights[589]), .RECT2_X(rectangle2_xs[589]), .RECT2_Y(rectangle2_ys[589]), .RECT2_WIDTH(rectangle2_widths[589]), .RECT2_HEIGHT(rectangle2_heights[589]), .RECT2_WEIGHT(rectangle2_weights[589]), .RECT3_X(rectangle3_xs[589]), .RECT3_Y(rectangle3_ys[589]), .RECT3_WIDTH(rectangle3_widths[589]), .RECT3_HEIGHT(rectangle3_heights[589]), .RECT3_WEIGHT(rectangle3_weights[589]), .FEAT_THRES(feature_thresholds[589]), .FEAT_ABOVE(feature_aboves[589]), .FEAT_BELOW(feature_belows[589])) ac589(.scan_win(scan_win589), .scan_win_std_dev(scan_win_std_dev[589]), .feature_accum(feature_accums[589]));
  accum_calculator #(.RECT1_X(rectangle1_xs[590]), .RECT1_Y(rectangle1_ys[590]), .RECT1_WIDTH(rectangle1_widths[590]), .RECT1_HEIGHT(rectangle1_heights[590]), .RECT1_WEIGHT(rectangle1_weights[590]), .RECT2_X(rectangle2_xs[590]), .RECT2_Y(rectangle2_ys[590]), .RECT2_WIDTH(rectangle2_widths[590]), .RECT2_HEIGHT(rectangle2_heights[590]), .RECT2_WEIGHT(rectangle2_weights[590]), .RECT3_X(rectangle3_xs[590]), .RECT3_Y(rectangle3_ys[590]), .RECT3_WIDTH(rectangle3_widths[590]), .RECT3_HEIGHT(rectangle3_heights[590]), .RECT3_WEIGHT(rectangle3_weights[590]), .FEAT_THRES(feature_thresholds[590]), .FEAT_ABOVE(feature_aboves[590]), .FEAT_BELOW(feature_belows[590])) ac590(.scan_win(scan_win590), .scan_win_std_dev(scan_win_std_dev[590]), .feature_accum(feature_accums[590]));
  accum_calculator #(.RECT1_X(rectangle1_xs[591]), .RECT1_Y(rectangle1_ys[591]), .RECT1_WIDTH(rectangle1_widths[591]), .RECT1_HEIGHT(rectangle1_heights[591]), .RECT1_WEIGHT(rectangle1_weights[591]), .RECT2_X(rectangle2_xs[591]), .RECT2_Y(rectangle2_ys[591]), .RECT2_WIDTH(rectangle2_widths[591]), .RECT2_HEIGHT(rectangle2_heights[591]), .RECT2_WEIGHT(rectangle2_weights[591]), .RECT3_X(rectangle3_xs[591]), .RECT3_Y(rectangle3_ys[591]), .RECT3_WIDTH(rectangle3_widths[591]), .RECT3_HEIGHT(rectangle3_heights[591]), .RECT3_WEIGHT(rectangle3_weights[591]), .FEAT_THRES(feature_thresholds[591]), .FEAT_ABOVE(feature_aboves[591]), .FEAT_BELOW(feature_belows[591])) ac591(.scan_win(scan_win591), .scan_win_std_dev(scan_win_std_dev[591]), .feature_accum(feature_accums[591]));
  accum_calculator #(.RECT1_X(rectangle1_xs[592]), .RECT1_Y(rectangle1_ys[592]), .RECT1_WIDTH(rectangle1_widths[592]), .RECT1_HEIGHT(rectangle1_heights[592]), .RECT1_WEIGHT(rectangle1_weights[592]), .RECT2_X(rectangle2_xs[592]), .RECT2_Y(rectangle2_ys[592]), .RECT2_WIDTH(rectangle2_widths[592]), .RECT2_HEIGHT(rectangle2_heights[592]), .RECT2_WEIGHT(rectangle2_weights[592]), .RECT3_X(rectangle3_xs[592]), .RECT3_Y(rectangle3_ys[592]), .RECT3_WIDTH(rectangle3_widths[592]), .RECT3_HEIGHT(rectangle3_heights[592]), .RECT3_WEIGHT(rectangle3_weights[592]), .FEAT_THRES(feature_thresholds[592]), .FEAT_ABOVE(feature_aboves[592]), .FEAT_BELOW(feature_belows[592])) ac592(.scan_win(scan_win592), .scan_win_std_dev(scan_win_std_dev[592]), .feature_accum(feature_accums[592]));
  accum_calculator #(.RECT1_X(rectangle1_xs[593]), .RECT1_Y(rectangle1_ys[593]), .RECT1_WIDTH(rectangle1_widths[593]), .RECT1_HEIGHT(rectangle1_heights[593]), .RECT1_WEIGHT(rectangle1_weights[593]), .RECT2_X(rectangle2_xs[593]), .RECT2_Y(rectangle2_ys[593]), .RECT2_WIDTH(rectangle2_widths[593]), .RECT2_HEIGHT(rectangle2_heights[593]), .RECT2_WEIGHT(rectangle2_weights[593]), .RECT3_X(rectangle3_xs[593]), .RECT3_Y(rectangle3_ys[593]), .RECT3_WIDTH(rectangle3_widths[593]), .RECT3_HEIGHT(rectangle3_heights[593]), .RECT3_WEIGHT(rectangle3_weights[593]), .FEAT_THRES(feature_thresholds[593]), .FEAT_ABOVE(feature_aboves[593]), .FEAT_BELOW(feature_belows[593])) ac593(.scan_win(scan_win593), .scan_win_std_dev(scan_win_std_dev[593]), .feature_accum(feature_accums[593]));
  accum_calculator #(.RECT1_X(rectangle1_xs[594]), .RECT1_Y(rectangle1_ys[594]), .RECT1_WIDTH(rectangle1_widths[594]), .RECT1_HEIGHT(rectangle1_heights[594]), .RECT1_WEIGHT(rectangle1_weights[594]), .RECT2_X(rectangle2_xs[594]), .RECT2_Y(rectangle2_ys[594]), .RECT2_WIDTH(rectangle2_widths[594]), .RECT2_HEIGHT(rectangle2_heights[594]), .RECT2_WEIGHT(rectangle2_weights[594]), .RECT3_X(rectangle3_xs[594]), .RECT3_Y(rectangle3_ys[594]), .RECT3_WIDTH(rectangle3_widths[594]), .RECT3_HEIGHT(rectangle3_heights[594]), .RECT3_WEIGHT(rectangle3_weights[594]), .FEAT_THRES(feature_thresholds[594]), .FEAT_ABOVE(feature_aboves[594]), .FEAT_BELOW(feature_belows[594])) ac594(.scan_win(scan_win594), .scan_win_std_dev(scan_win_std_dev[594]), .feature_accum(feature_accums[594]));
  accum_calculator #(.RECT1_X(rectangle1_xs[595]), .RECT1_Y(rectangle1_ys[595]), .RECT1_WIDTH(rectangle1_widths[595]), .RECT1_HEIGHT(rectangle1_heights[595]), .RECT1_WEIGHT(rectangle1_weights[595]), .RECT2_X(rectangle2_xs[595]), .RECT2_Y(rectangle2_ys[595]), .RECT2_WIDTH(rectangle2_widths[595]), .RECT2_HEIGHT(rectangle2_heights[595]), .RECT2_WEIGHT(rectangle2_weights[595]), .RECT3_X(rectangle3_xs[595]), .RECT3_Y(rectangle3_ys[595]), .RECT3_WIDTH(rectangle3_widths[595]), .RECT3_HEIGHT(rectangle3_heights[595]), .RECT3_WEIGHT(rectangle3_weights[595]), .FEAT_THRES(feature_thresholds[595]), .FEAT_ABOVE(feature_aboves[595]), .FEAT_BELOW(feature_belows[595])) ac595(.scan_win(scan_win595), .scan_win_std_dev(scan_win_std_dev[595]), .feature_accum(feature_accums[595]));
  accum_calculator #(.RECT1_X(rectangle1_xs[596]), .RECT1_Y(rectangle1_ys[596]), .RECT1_WIDTH(rectangle1_widths[596]), .RECT1_HEIGHT(rectangle1_heights[596]), .RECT1_WEIGHT(rectangle1_weights[596]), .RECT2_X(rectangle2_xs[596]), .RECT2_Y(rectangle2_ys[596]), .RECT2_WIDTH(rectangle2_widths[596]), .RECT2_HEIGHT(rectangle2_heights[596]), .RECT2_WEIGHT(rectangle2_weights[596]), .RECT3_X(rectangle3_xs[596]), .RECT3_Y(rectangle3_ys[596]), .RECT3_WIDTH(rectangle3_widths[596]), .RECT3_HEIGHT(rectangle3_heights[596]), .RECT3_WEIGHT(rectangle3_weights[596]), .FEAT_THRES(feature_thresholds[596]), .FEAT_ABOVE(feature_aboves[596]), .FEAT_BELOW(feature_belows[596])) ac596(.scan_win(scan_win596), .scan_win_std_dev(scan_win_std_dev[596]), .feature_accum(feature_accums[596]));
  accum_calculator #(.RECT1_X(rectangle1_xs[597]), .RECT1_Y(rectangle1_ys[597]), .RECT1_WIDTH(rectangle1_widths[597]), .RECT1_HEIGHT(rectangle1_heights[597]), .RECT1_WEIGHT(rectangle1_weights[597]), .RECT2_X(rectangle2_xs[597]), .RECT2_Y(rectangle2_ys[597]), .RECT2_WIDTH(rectangle2_widths[597]), .RECT2_HEIGHT(rectangle2_heights[597]), .RECT2_WEIGHT(rectangle2_weights[597]), .RECT3_X(rectangle3_xs[597]), .RECT3_Y(rectangle3_ys[597]), .RECT3_WIDTH(rectangle3_widths[597]), .RECT3_HEIGHT(rectangle3_heights[597]), .RECT3_WEIGHT(rectangle3_weights[597]), .FEAT_THRES(feature_thresholds[597]), .FEAT_ABOVE(feature_aboves[597]), .FEAT_BELOW(feature_belows[597])) ac597(.scan_win(scan_win597), .scan_win_std_dev(scan_win_std_dev[597]), .feature_accum(feature_accums[597]));
  accum_calculator #(.RECT1_X(rectangle1_xs[598]), .RECT1_Y(rectangle1_ys[598]), .RECT1_WIDTH(rectangle1_widths[598]), .RECT1_HEIGHT(rectangle1_heights[598]), .RECT1_WEIGHT(rectangle1_weights[598]), .RECT2_X(rectangle2_xs[598]), .RECT2_Y(rectangle2_ys[598]), .RECT2_WIDTH(rectangle2_widths[598]), .RECT2_HEIGHT(rectangle2_heights[598]), .RECT2_WEIGHT(rectangle2_weights[598]), .RECT3_X(rectangle3_xs[598]), .RECT3_Y(rectangle3_ys[598]), .RECT3_WIDTH(rectangle3_widths[598]), .RECT3_HEIGHT(rectangle3_heights[598]), .RECT3_WEIGHT(rectangle3_weights[598]), .FEAT_THRES(feature_thresholds[598]), .FEAT_ABOVE(feature_aboves[598]), .FEAT_BELOW(feature_belows[598])) ac598(.scan_win(scan_win598), .scan_win_std_dev(scan_win_std_dev[598]), .feature_accum(feature_accums[598]));
  accum_calculator #(.RECT1_X(rectangle1_xs[599]), .RECT1_Y(rectangle1_ys[599]), .RECT1_WIDTH(rectangle1_widths[599]), .RECT1_HEIGHT(rectangle1_heights[599]), .RECT1_WEIGHT(rectangle1_weights[599]), .RECT2_X(rectangle2_xs[599]), .RECT2_Y(rectangle2_ys[599]), .RECT2_WIDTH(rectangle2_widths[599]), .RECT2_HEIGHT(rectangle2_heights[599]), .RECT2_WEIGHT(rectangle2_weights[599]), .RECT3_X(rectangle3_xs[599]), .RECT3_Y(rectangle3_ys[599]), .RECT3_WIDTH(rectangle3_widths[599]), .RECT3_HEIGHT(rectangle3_heights[599]), .RECT3_WEIGHT(rectangle3_weights[599]), .FEAT_THRES(feature_thresholds[599]), .FEAT_ABOVE(feature_aboves[599]), .FEAT_BELOW(feature_belows[599])) ac599(.scan_win(scan_win599), .scan_win_std_dev(scan_win_std_dev[599]), .feature_accum(feature_accums[599]));
  accum_calculator #(.RECT1_X(rectangle1_xs[600]), .RECT1_Y(rectangle1_ys[600]), .RECT1_WIDTH(rectangle1_widths[600]), .RECT1_HEIGHT(rectangle1_heights[600]), .RECT1_WEIGHT(rectangle1_weights[600]), .RECT2_X(rectangle2_xs[600]), .RECT2_Y(rectangle2_ys[600]), .RECT2_WIDTH(rectangle2_widths[600]), .RECT2_HEIGHT(rectangle2_heights[600]), .RECT2_WEIGHT(rectangle2_weights[600]), .RECT3_X(rectangle3_xs[600]), .RECT3_Y(rectangle3_ys[600]), .RECT3_WIDTH(rectangle3_widths[600]), .RECT3_HEIGHT(rectangle3_heights[600]), .RECT3_WEIGHT(rectangle3_weights[600]), .FEAT_THRES(feature_thresholds[600]), .FEAT_ABOVE(feature_aboves[600]), .FEAT_BELOW(feature_belows[600])) ac600(.scan_win(scan_win600), .scan_win_std_dev(scan_win_std_dev[600]), .feature_accum(feature_accums[600]));
  accum_calculator #(.RECT1_X(rectangle1_xs[601]), .RECT1_Y(rectangle1_ys[601]), .RECT1_WIDTH(rectangle1_widths[601]), .RECT1_HEIGHT(rectangle1_heights[601]), .RECT1_WEIGHT(rectangle1_weights[601]), .RECT2_X(rectangle2_xs[601]), .RECT2_Y(rectangle2_ys[601]), .RECT2_WIDTH(rectangle2_widths[601]), .RECT2_HEIGHT(rectangle2_heights[601]), .RECT2_WEIGHT(rectangle2_weights[601]), .RECT3_X(rectangle3_xs[601]), .RECT3_Y(rectangle3_ys[601]), .RECT3_WIDTH(rectangle3_widths[601]), .RECT3_HEIGHT(rectangle3_heights[601]), .RECT3_WEIGHT(rectangle3_weights[601]), .FEAT_THRES(feature_thresholds[601]), .FEAT_ABOVE(feature_aboves[601]), .FEAT_BELOW(feature_belows[601])) ac601(.scan_win(scan_win601), .scan_win_std_dev(scan_win_std_dev[601]), .feature_accum(feature_accums[601]));
  accum_calculator #(.RECT1_X(rectangle1_xs[602]), .RECT1_Y(rectangle1_ys[602]), .RECT1_WIDTH(rectangle1_widths[602]), .RECT1_HEIGHT(rectangle1_heights[602]), .RECT1_WEIGHT(rectangle1_weights[602]), .RECT2_X(rectangle2_xs[602]), .RECT2_Y(rectangle2_ys[602]), .RECT2_WIDTH(rectangle2_widths[602]), .RECT2_HEIGHT(rectangle2_heights[602]), .RECT2_WEIGHT(rectangle2_weights[602]), .RECT3_X(rectangle3_xs[602]), .RECT3_Y(rectangle3_ys[602]), .RECT3_WIDTH(rectangle3_widths[602]), .RECT3_HEIGHT(rectangle3_heights[602]), .RECT3_WEIGHT(rectangle3_weights[602]), .FEAT_THRES(feature_thresholds[602]), .FEAT_ABOVE(feature_aboves[602]), .FEAT_BELOW(feature_belows[602])) ac602(.scan_win(scan_win602), .scan_win_std_dev(scan_win_std_dev[602]), .feature_accum(feature_accums[602]));
  accum_calculator #(.RECT1_X(rectangle1_xs[603]), .RECT1_Y(rectangle1_ys[603]), .RECT1_WIDTH(rectangle1_widths[603]), .RECT1_HEIGHT(rectangle1_heights[603]), .RECT1_WEIGHT(rectangle1_weights[603]), .RECT2_X(rectangle2_xs[603]), .RECT2_Y(rectangle2_ys[603]), .RECT2_WIDTH(rectangle2_widths[603]), .RECT2_HEIGHT(rectangle2_heights[603]), .RECT2_WEIGHT(rectangle2_weights[603]), .RECT3_X(rectangle3_xs[603]), .RECT3_Y(rectangle3_ys[603]), .RECT3_WIDTH(rectangle3_widths[603]), .RECT3_HEIGHT(rectangle3_heights[603]), .RECT3_WEIGHT(rectangle3_weights[603]), .FEAT_THRES(feature_thresholds[603]), .FEAT_ABOVE(feature_aboves[603]), .FEAT_BELOW(feature_belows[603])) ac603(.scan_win(scan_win603), .scan_win_std_dev(scan_win_std_dev[603]), .feature_accum(feature_accums[603]));
  accum_calculator #(.RECT1_X(rectangle1_xs[604]), .RECT1_Y(rectangle1_ys[604]), .RECT1_WIDTH(rectangle1_widths[604]), .RECT1_HEIGHT(rectangle1_heights[604]), .RECT1_WEIGHT(rectangle1_weights[604]), .RECT2_X(rectangle2_xs[604]), .RECT2_Y(rectangle2_ys[604]), .RECT2_WIDTH(rectangle2_widths[604]), .RECT2_HEIGHT(rectangle2_heights[604]), .RECT2_WEIGHT(rectangle2_weights[604]), .RECT3_X(rectangle3_xs[604]), .RECT3_Y(rectangle3_ys[604]), .RECT3_WIDTH(rectangle3_widths[604]), .RECT3_HEIGHT(rectangle3_heights[604]), .RECT3_WEIGHT(rectangle3_weights[604]), .FEAT_THRES(feature_thresholds[604]), .FEAT_ABOVE(feature_aboves[604]), .FEAT_BELOW(feature_belows[604])) ac604(.scan_win(scan_win604), .scan_win_std_dev(scan_win_std_dev[604]), .feature_accum(feature_accums[604]));
  accum_calculator #(.RECT1_X(rectangle1_xs[605]), .RECT1_Y(rectangle1_ys[605]), .RECT1_WIDTH(rectangle1_widths[605]), .RECT1_HEIGHT(rectangle1_heights[605]), .RECT1_WEIGHT(rectangle1_weights[605]), .RECT2_X(rectangle2_xs[605]), .RECT2_Y(rectangle2_ys[605]), .RECT2_WIDTH(rectangle2_widths[605]), .RECT2_HEIGHT(rectangle2_heights[605]), .RECT2_WEIGHT(rectangle2_weights[605]), .RECT3_X(rectangle3_xs[605]), .RECT3_Y(rectangle3_ys[605]), .RECT3_WIDTH(rectangle3_widths[605]), .RECT3_HEIGHT(rectangle3_heights[605]), .RECT3_WEIGHT(rectangle3_weights[605]), .FEAT_THRES(feature_thresholds[605]), .FEAT_ABOVE(feature_aboves[605]), .FEAT_BELOW(feature_belows[605])) ac605(.scan_win(scan_win605), .scan_win_std_dev(scan_win_std_dev[605]), .feature_accum(feature_accums[605]));
  accum_calculator #(.RECT1_X(rectangle1_xs[606]), .RECT1_Y(rectangle1_ys[606]), .RECT1_WIDTH(rectangle1_widths[606]), .RECT1_HEIGHT(rectangle1_heights[606]), .RECT1_WEIGHT(rectangle1_weights[606]), .RECT2_X(rectangle2_xs[606]), .RECT2_Y(rectangle2_ys[606]), .RECT2_WIDTH(rectangle2_widths[606]), .RECT2_HEIGHT(rectangle2_heights[606]), .RECT2_WEIGHT(rectangle2_weights[606]), .RECT3_X(rectangle3_xs[606]), .RECT3_Y(rectangle3_ys[606]), .RECT3_WIDTH(rectangle3_widths[606]), .RECT3_HEIGHT(rectangle3_heights[606]), .RECT3_WEIGHT(rectangle3_weights[606]), .FEAT_THRES(feature_thresholds[606]), .FEAT_ABOVE(feature_aboves[606]), .FEAT_BELOW(feature_belows[606])) ac606(.scan_win(scan_win606), .scan_win_std_dev(scan_win_std_dev[606]), .feature_accum(feature_accums[606]));
  accum_calculator #(.RECT1_X(rectangle1_xs[607]), .RECT1_Y(rectangle1_ys[607]), .RECT1_WIDTH(rectangle1_widths[607]), .RECT1_HEIGHT(rectangle1_heights[607]), .RECT1_WEIGHT(rectangle1_weights[607]), .RECT2_X(rectangle2_xs[607]), .RECT2_Y(rectangle2_ys[607]), .RECT2_WIDTH(rectangle2_widths[607]), .RECT2_HEIGHT(rectangle2_heights[607]), .RECT2_WEIGHT(rectangle2_weights[607]), .RECT3_X(rectangle3_xs[607]), .RECT3_Y(rectangle3_ys[607]), .RECT3_WIDTH(rectangle3_widths[607]), .RECT3_HEIGHT(rectangle3_heights[607]), .RECT3_WEIGHT(rectangle3_weights[607]), .FEAT_THRES(feature_thresholds[607]), .FEAT_ABOVE(feature_aboves[607]), .FEAT_BELOW(feature_belows[607])) ac607(.scan_win(scan_win607), .scan_win_std_dev(scan_win_std_dev[607]), .feature_accum(feature_accums[607]));
  accum_calculator #(.RECT1_X(rectangle1_xs[608]), .RECT1_Y(rectangle1_ys[608]), .RECT1_WIDTH(rectangle1_widths[608]), .RECT1_HEIGHT(rectangle1_heights[608]), .RECT1_WEIGHT(rectangle1_weights[608]), .RECT2_X(rectangle2_xs[608]), .RECT2_Y(rectangle2_ys[608]), .RECT2_WIDTH(rectangle2_widths[608]), .RECT2_HEIGHT(rectangle2_heights[608]), .RECT2_WEIGHT(rectangle2_weights[608]), .RECT3_X(rectangle3_xs[608]), .RECT3_Y(rectangle3_ys[608]), .RECT3_WIDTH(rectangle3_widths[608]), .RECT3_HEIGHT(rectangle3_heights[608]), .RECT3_WEIGHT(rectangle3_weights[608]), .FEAT_THRES(feature_thresholds[608]), .FEAT_ABOVE(feature_aboves[608]), .FEAT_BELOW(feature_belows[608])) ac608(.scan_win(scan_win608), .scan_win_std_dev(scan_win_std_dev[608]), .feature_accum(feature_accums[608]));
  accum_calculator #(.RECT1_X(rectangle1_xs[609]), .RECT1_Y(rectangle1_ys[609]), .RECT1_WIDTH(rectangle1_widths[609]), .RECT1_HEIGHT(rectangle1_heights[609]), .RECT1_WEIGHT(rectangle1_weights[609]), .RECT2_X(rectangle2_xs[609]), .RECT2_Y(rectangle2_ys[609]), .RECT2_WIDTH(rectangle2_widths[609]), .RECT2_HEIGHT(rectangle2_heights[609]), .RECT2_WEIGHT(rectangle2_weights[609]), .RECT3_X(rectangle3_xs[609]), .RECT3_Y(rectangle3_ys[609]), .RECT3_WIDTH(rectangle3_widths[609]), .RECT3_HEIGHT(rectangle3_heights[609]), .RECT3_WEIGHT(rectangle3_weights[609]), .FEAT_THRES(feature_thresholds[609]), .FEAT_ABOVE(feature_aboves[609]), .FEAT_BELOW(feature_belows[609])) ac609(.scan_win(scan_win609), .scan_win_std_dev(scan_win_std_dev[609]), .feature_accum(feature_accums[609]));
  accum_calculator #(.RECT1_X(rectangle1_xs[610]), .RECT1_Y(rectangle1_ys[610]), .RECT1_WIDTH(rectangle1_widths[610]), .RECT1_HEIGHT(rectangle1_heights[610]), .RECT1_WEIGHT(rectangle1_weights[610]), .RECT2_X(rectangle2_xs[610]), .RECT2_Y(rectangle2_ys[610]), .RECT2_WIDTH(rectangle2_widths[610]), .RECT2_HEIGHT(rectangle2_heights[610]), .RECT2_WEIGHT(rectangle2_weights[610]), .RECT3_X(rectangle3_xs[610]), .RECT3_Y(rectangle3_ys[610]), .RECT3_WIDTH(rectangle3_widths[610]), .RECT3_HEIGHT(rectangle3_heights[610]), .RECT3_WEIGHT(rectangle3_weights[610]), .FEAT_THRES(feature_thresholds[610]), .FEAT_ABOVE(feature_aboves[610]), .FEAT_BELOW(feature_belows[610])) ac610(.scan_win(scan_win610), .scan_win_std_dev(scan_win_std_dev[610]), .feature_accum(feature_accums[610]));
  accum_calculator #(.RECT1_X(rectangle1_xs[611]), .RECT1_Y(rectangle1_ys[611]), .RECT1_WIDTH(rectangle1_widths[611]), .RECT1_HEIGHT(rectangle1_heights[611]), .RECT1_WEIGHT(rectangle1_weights[611]), .RECT2_X(rectangle2_xs[611]), .RECT2_Y(rectangle2_ys[611]), .RECT2_WIDTH(rectangle2_widths[611]), .RECT2_HEIGHT(rectangle2_heights[611]), .RECT2_WEIGHT(rectangle2_weights[611]), .RECT3_X(rectangle3_xs[611]), .RECT3_Y(rectangle3_ys[611]), .RECT3_WIDTH(rectangle3_widths[611]), .RECT3_HEIGHT(rectangle3_heights[611]), .RECT3_WEIGHT(rectangle3_weights[611]), .FEAT_THRES(feature_thresholds[611]), .FEAT_ABOVE(feature_aboves[611]), .FEAT_BELOW(feature_belows[611])) ac611(.scan_win(scan_win611), .scan_win_std_dev(scan_win_std_dev[611]), .feature_accum(feature_accums[611]));
  accum_calculator #(.RECT1_X(rectangle1_xs[612]), .RECT1_Y(rectangle1_ys[612]), .RECT1_WIDTH(rectangle1_widths[612]), .RECT1_HEIGHT(rectangle1_heights[612]), .RECT1_WEIGHT(rectangle1_weights[612]), .RECT2_X(rectangle2_xs[612]), .RECT2_Y(rectangle2_ys[612]), .RECT2_WIDTH(rectangle2_widths[612]), .RECT2_HEIGHT(rectangle2_heights[612]), .RECT2_WEIGHT(rectangle2_weights[612]), .RECT3_X(rectangle3_xs[612]), .RECT3_Y(rectangle3_ys[612]), .RECT3_WIDTH(rectangle3_widths[612]), .RECT3_HEIGHT(rectangle3_heights[612]), .RECT3_WEIGHT(rectangle3_weights[612]), .FEAT_THRES(feature_thresholds[612]), .FEAT_ABOVE(feature_aboves[612]), .FEAT_BELOW(feature_belows[612])) ac612(.scan_win(scan_win612), .scan_win_std_dev(scan_win_std_dev[612]), .feature_accum(feature_accums[612]));
  accum_calculator #(.RECT1_X(rectangle1_xs[613]), .RECT1_Y(rectangle1_ys[613]), .RECT1_WIDTH(rectangle1_widths[613]), .RECT1_HEIGHT(rectangle1_heights[613]), .RECT1_WEIGHT(rectangle1_weights[613]), .RECT2_X(rectangle2_xs[613]), .RECT2_Y(rectangle2_ys[613]), .RECT2_WIDTH(rectangle2_widths[613]), .RECT2_HEIGHT(rectangle2_heights[613]), .RECT2_WEIGHT(rectangle2_weights[613]), .RECT3_X(rectangle3_xs[613]), .RECT3_Y(rectangle3_ys[613]), .RECT3_WIDTH(rectangle3_widths[613]), .RECT3_HEIGHT(rectangle3_heights[613]), .RECT3_WEIGHT(rectangle3_weights[613]), .FEAT_THRES(feature_thresholds[613]), .FEAT_ABOVE(feature_aboves[613]), .FEAT_BELOW(feature_belows[613])) ac613(.scan_win(scan_win613), .scan_win_std_dev(scan_win_std_dev[613]), .feature_accum(feature_accums[613]));
  accum_calculator #(.RECT1_X(rectangle1_xs[614]), .RECT1_Y(rectangle1_ys[614]), .RECT1_WIDTH(rectangle1_widths[614]), .RECT1_HEIGHT(rectangle1_heights[614]), .RECT1_WEIGHT(rectangle1_weights[614]), .RECT2_X(rectangle2_xs[614]), .RECT2_Y(rectangle2_ys[614]), .RECT2_WIDTH(rectangle2_widths[614]), .RECT2_HEIGHT(rectangle2_heights[614]), .RECT2_WEIGHT(rectangle2_weights[614]), .RECT3_X(rectangle3_xs[614]), .RECT3_Y(rectangle3_ys[614]), .RECT3_WIDTH(rectangle3_widths[614]), .RECT3_HEIGHT(rectangle3_heights[614]), .RECT3_WEIGHT(rectangle3_weights[614]), .FEAT_THRES(feature_thresholds[614]), .FEAT_ABOVE(feature_aboves[614]), .FEAT_BELOW(feature_belows[614])) ac614(.scan_win(scan_win614), .scan_win_std_dev(scan_win_std_dev[614]), .feature_accum(feature_accums[614]));
  accum_calculator #(.RECT1_X(rectangle1_xs[615]), .RECT1_Y(rectangle1_ys[615]), .RECT1_WIDTH(rectangle1_widths[615]), .RECT1_HEIGHT(rectangle1_heights[615]), .RECT1_WEIGHT(rectangle1_weights[615]), .RECT2_X(rectangle2_xs[615]), .RECT2_Y(rectangle2_ys[615]), .RECT2_WIDTH(rectangle2_widths[615]), .RECT2_HEIGHT(rectangle2_heights[615]), .RECT2_WEIGHT(rectangle2_weights[615]), .RECT3_X(rectangle3_xs[615]), .RECT3_Y(rectangle3_ys[615]), .RECT3_WIDTH(rectangle3_widths[615]), .RECT3_HEIGHT(rectangle3_heights[615]), .RECT3_WEIGHT(rectangle3_weights[615]), .FEAT_THRES(feature_thresholds[615]), .FEAT_ABOVE(feature_aboves[615]), .FEAT_BELOW(feature_belows[615])) ac615(.scan_win(scan_win615), .scan_win_std_dev(scan_win_std_dev[615]), .feature_accum(feature_accums[615]));
  accum_calculator #(.RECT1_X(rectangle1_xs[616]), .RECT1_Y(rectangle1_ys[616]), .RECT1_WIDTH(rectangle1_widths[616]), .RECT1_HEIGHT(rectangle1_heights[616]), .RECT1_WEIGHT(rectangle1_weights[616]), .RECT2_X(rectangle2_xs[616]), .RECT2_Y(rectangle2_ys[616]), .RECT2_WIDTH(rectangle2_widths[616]), .RECT2_HEIGHT(rectangle2_heights[616]), .RECT2_WEIGHT(rectangle2_weights[616]), .RECT3_X(rectangle3_xs[616]), .RECT3_Y(rectangle3_ys[616]), .RECT3_WIDTH(rectangle3_widths[616]), .RECT3_HEIGHT(rectangle3_heights[616]), .RECT3_WEIGHT(rectangle3_weights[616]), .FEAT_THRES(feature_thresholds[616]), .FEAT_ABOVE(feature_aboves[616]), .FEAT_BELOW(feature_belows[616])) ac616(.scan_win(scan_win616), .scan_win_std_dev(scan_win_std_dev[616]), .feature_accum(feature_accums[616]));
  accum_calculator #(.RECT1_X(rectangle1_xs[617]), .RECT1_Y(rectangle1_ys[617]), .RECT1_WIDTH(rectangle1_widths[617]), .RECT1_HEIGHT(rectangle1_heights[617]), .RECT1_WEIGHT(rectangle1_weights[617]), .RECT2_X(rectangle2_xs[617]), .RECT2_Y(rectangle2_ys[617]), .RECT2_WIDTH(rectangle2_widths[617]), .RECT2_HEIGHT(rectangle2_heights[617]), .RECT2_WEIGHT(rectangle2_weights[617]), .RECT3_X(rectangle3_xs[617]), .RECT3_Y(rectangle3_ys[617]), .RECT3_WIDTH(rectangle3_widths[617]), .RECT3_HEIGHT(rectangle3_heights[617]), .RECT3_WEIGHT(rectangle3_weights[617]), .FEAT_THRES(feature_thresholds[617]), .FEAT_ABOVE(feature_aboves[617]), .FEAT_BELOW(feature_belows[617])) ac617(.scan_win(scan_win617), .scan_win_std_dev(scan_win_std_dev[617]), .feature_accum(feature_accums[617]));
  accum_calculator #(.RECT1_X(rectangle1_xs[618]), .RECT1_Y(rectangle1_ys[618]), .RECT1_WIDTH(rectangle1_widths[618]), .RECT1_HEIGHT(rectangle1_heights[618]), .RECT1_WEIGHT(rectangle1_weights[618]), .RECT2_X(rectangle2_xs[618]), .RECT2_Y(rectangle2_ys[618]), .RECT2_WIDTH(rectangle2_widths[618]), .RECT2_HEIGHT(rectangle2_heights[618]), .RECT2_WEIGHT(rectangle2_weights[618]), .RECT3_X(rectangle3_xs[618]), .RECT3_Y(rectangle3_ys[618]), .RECT3_WIDTH(rectangle3_widths[618]), .RECT3_HEIGHT(rectangle3_heights[618]), .RECT3_WEIGHT(rectangle3_weights[618]), .FEAT_THRES(feature_thresholds[618]), .FEAT_ABOVE(feature_aboves[618]), .FEAT_BELOW(feature_belows[618])) ac618(.scan_win(scan_win618), .scan_win_std_dev(scan_win_std_dev[618]), .feature_accum(feature_accums[618]));
  accum_calculator #(.RECT1_X(rectangle1_xs[619]), .RECT1_Y(rectangle1_ys[619]), .RECT1_WIDTH(rectangle1_widths[619]), .RECT1_HEIGHT(rectangle1_heights[619]), .RECT1_WEIGHT(rectangle1_weights[619]), .RECT2_X(rectangle2_xs[619]), .RECT2_Y(rectangle2_ys[619]), .RECT2_WIDTH(rectangle2_widths[619]), .RECT2_HEIGHT(rectangle2_heights[619]), .RECT2_WEIGHT(rectangle2_weights[619]), .RECT3_X(rectangle3_xs[619]), .RECT3_Y(rectangle3_ys[619]), .RECT3_WIDTH(rectangle3_widths[619]), .RECT3_HEIGHT(rectangle3_heights[619]), .RECT3_WEIGHT(rectangle3_weights[619]), .FEAT_THRES(feature_thresholds[619]), .FEAT_ABOVE(feature_aboves[619]), .FEAT_BELOW(feature_belows[619])) ac619(.scan_win(scan_win619), .scan_win_std_dev(scan_win_std_dev[619]), .feature_accum(feature_accums[619]));
  accum_calculator #(.RECT1_X(rectangle1_xs[620]), .RECT1_Y(rectangle1_ys[620]), .RECT1_WIDTH(rectangle1_widths[620]), .RECT1_HEIGHT(rectangle1_heights[620]), .RECT1_WEIGHT(rectangle1_weights[620]), .RECT2_X(rectangle2_xs[620]), .RECT2_Y(rectangle2_ys[620]), .RECT2_WIDTH(rectangle2_widths[620]), .RECT2_HEIGHT(rectangle2_heights[620]), .RECT2_WEIGHT(rectangle2_weights[620]), .RECT3_X(rectangle3_xs[620]), .RECT3_Y(rectangle3_ys[620]), .RECT3_WIDTH(rectangle3_widths[620]), .RECT3_HEIGHT(rectangle3_heights[620]), .RECT3_WEIGHT(rectangle3_weights[620]), .FEAT_THRES(feature_thresholds[620]), .FEAT_ABOVE(feature_aboves[620]), .FEAT_BELOW(feature_belows[620])) ac620(.scan_win(scan_win620), .scan_win_std_dev(scan_win_std_dev[620]), .feature_accum(feature_accums[620]));
  accum_calculator #(.RECT1_X(rectangle1_xs[621]), .RECT1_Y(rectangle1_ys[621]), .RECT1_WIDTH(rectangle1_widths[621]), .RECT1_HEIGHT(rectangle1_heights[621]), .RECT1_WEIGHT(rectangle1_weights[621]), .RECT2_X(rectangle2_xs[621]), .RECT2_Y(rectangle2_ys[621]), .RECT2_WIDTH(rectangle2_widths[621]), .RECT2_HEIGHT(rectangle2_heights[621]), .RECT2_WEIGHT(rectangle2_weights[621]), .RECT3_X(rectangle3_xs[621]), .RECT3_Y(rectangle3_ys[621]), .RECT3_WIDTH(rectangle3_widths[621]), .RECT3_HEIGHT(rectangle3_heights[621]), .RECT3_WEIGHT(rectangle3_weights[621]), .FEAT_THRES(feature_thresholds[621]), .FEAT_ABOVE(feature_aboves[621]), .FEAT_BELOW(feature_belows[621])) ac621(.scan_win(scan_win621), .scan_win_std_dev(scan_win_std_dev[621]), .feature_accum(feature_accums[621]));
  accum_calculator #(.RECT1_X(rectangle1_xs[622]), .RECT1_Y(rectangle1_ys[622]), .RECT1_WIDTH(rectangle1_widths[622]), .RECT1_HEIGHT(rectangle1_heights[622]), .RECT1_WEIGHT(rectangle1_weights[622]), .RECT2_X(rectangle2_xs[622]), .RECT2_Y(rectangle2_ys[622]), .RECT2_WIDTH(rectangle2_widths[622]), .RECT2_HEIGHT(rectangle2_heights[622]), .RECT2_WEIGHT(rectangle2_weights[622]), .RECT3_X(rectangle3_xs[622]), .RECT3_Y(rectangle3_ys[622]), .RECT3_WIDTH(rectangle3_widths[622]), .RECT3_HEIGHT(rectangle3_heights[622]), .RECT3_WEIGHT(rectangle3_weights[622]), .FEAT_THRES(feature_thresholds[622]), .FEAT_ABOVE(feature_aboves[622]), .FEAT_BELOW(feature_belows[622])) ac622(.scan_win(scan_win622), .scan_win_std_dev(scan_win_std_dev[622]), .feature_accum(feature_accums[622]));
  accum_calculator #(.RECT1_X(rectangle1_xs[623]), .RECT1_Y(rectangle1_ys[623]), .RECT1_WIDTH(rectangle1_widths[623]), .RECT1_HEIGHT(rectangle1_heights[623]), .RECT1_WEIGHT(rectangle1_weights[623]), .RECT2_X(rectangle2_xs[623]), .RECT2_Y(rectangle2_ys[623]), .RECT2_WIDTH(rectangle2_widths[623]), .RECT2_HEIGHT(rectangle2_heights[623]), .RECT2_WEIGHT(rectangle2_weights[623]), .RECT3_X(rectangle3_xs[623]), .RECT3_Y(rectangle3_ys[623]), .RECT3_WIDTH(rectangle3_widths[623]), .RECT3_HEIGHT(rectangle3_heights[623]), .RECT3_WEIGHT(rectangle3_weights[623]), .FEAT_THRES(feature_thresholds[623]), .FEAT_ABOVE(feature_aboves[623]), .FEAT_BELOW(feature_belows[623])) ac623(.scan_win(scan_win623), .scan_win_std_dev(scan_win_std_dev[623]), .feature_accum(feature_accums[623]));
  accum_calculator #(.RECT1_X(rectangle1_xs[624]), .RECT1_Y(rectangle1_ys[624]), .RECT1_WIDTH(rectangle1_widths[624]), .RECT1_HEIGHT(rectangle1_heights[624]), .RECT1_WEIGHT(rectangle1_weights[624]), .RECT2_X(rectangle2_xs[624]), .RECT2_Y(rectangle2_ys[624]), .RECT2_WIDTH(rectangle2_widths[624]), .RECT2_HEIGHT(rectangle2_heights[624]), .RECT2_WEIGHT(rectangle2_weights[624]), .RECT3_X(rectangle3_xs[624]), .RECT3_Y(rectangle3_ys[624]), .RECT3_WIDTH(rectangle3_widths[624]), .RECT3_HEIGHT(rectangle3_heights[624]), .RECT3_WEIGHT(rectangle3_weights[624]), .FEAT_THRES(feature_thresholds[624]), .FEAT_ABOVE(feature_aboves[624]), .FEAT_BELOW(feature_belows[624])) ac624(.scan_win(scan_win624), .scan_win_std_dev(scan_win_std_dev[624]), .feature_accum(feature_accums[624]));
  accum_calculator #(.RECT1_X(rectangle1_xs[625]), .RECT1_Y(rectangle1_ys[625]), .RECT1_WIDTH(rectangle1_widths[625]), .RECT1_HEIGHT(rectangle1_heights[625]), .RECT1_WEIGHT(rectangle1_weights[625]), .RECT2_X(rectangle2_xs[625]), .RECT2_Y(rectangle2_ys[625]), .RECT2_WIDTH(rectangle2_widths[625]), .RECT2_HEIGHT(rectangle2_heights[625]), .RECT2_WEIGHT(rectangle2_weights[625]), .RECT3_X(rectangle3_xs[625]), .RECT3_Y(rectangle3_ys[625]), .RECT3_WIDTH(rectangle3_widths[625]), .RECT3_HEIGHT(rectangle3_heights[625]), .RECT3_WEIGHT(rectangle3_weights[625]), .FEAT_THRES(feature_thresholds[625]), .FEAT_ABOVE(feature_aboves[625]), .FEAT_BELOW(feature_belows[625])) ac625(.scan_win(scan_win625), .scan_win_std_dev(scan_win_std_dev[625]), .feature_accum(feature_accums[625]));
  accum_calculator #(.RECT1_X(rectangle1_xs[626]), .RECT1_Y(rectangle1_ys[626]), .RECT1_WIDTH(rectangle1_widths[626]), .RECT1_HEIGHT(rectangle1_heights[626]), .RECT1_WEIGHT(rectangle1_weights[626]), .RECT2_X(rectangle2_xs[626]), .RECT2_Y(rectangle2_ys[626]), .RECT2_WIDTH(rectangle2_widths[626]), .RECT2_HEIGHT(rectangle2_heights[626]), .RECT2_WEIGHT(rectangle2_weights[626]), .RECT3_X(rectangle3_xs[626]), .RECT3_Y(rectangle3_ys[626]), .RECT3_WIDTH(rectangle3_widths[626]), .RECT3_HEIGHT(rectangle3_heights[626]), .RECT3_WEIGHT(rectangle3_weights[626]), .FEAT_THRES(feature_thresholds[626]), .FEAT_ABOVE(feature_aboves[626]), .FEAT_BELOW(feature_belows[626])) ac626(.scan_win(scan_win626), .scan_win_std_dev(scan_win_std_dev[626]), .feature_accum(feature_accums[626]));
  accum_calculator #(.RECT1_X(rectangle1_xs[627]), .RECT1_Y(rectangle1_ys[627]), .RECT1_WIDTH(rectangle1_widths[627]), .RECT1_HEIGHT(rectangle1_heights[627]), .RECT1_WEIGHT(rectangle1_weights[627]), .RECT2_X(rectangle2_xs[627]), .RECT2_Y(rectangle2_ys[627]), .RECT2_WIDTH(rectangle2_widths[627]), .RECT2_HEIGHT(rectangle2_heights[627]), .RECT2_WEIGHT(rectangle2_weights[627]), .RECT3_X(rectangle3_xs[627]), .RECT3_Y(rectangle3_ys[627]), .RECT3_WIDTH(rectangle3_widths[627]), .RECT3_HEIGHT(rectangle3_heights[627]), .RECT3_WEIGHT(rectangle3_weights[627]), .FEAT_THRES(feature_thresholds[627]), .FEAT_ABOVE(feature_aboves[627]), .FEAT_BELOW(feature_belows[627])) ac627(.scan_win(scan_win627), .scan_win_std_dev(scan_win_std_dev[627]), .feature_accum(feature_accums[627]));
  accum_calculator #(.RECT1_X(rectangle1_xs[628]), .RECT1_Y(rectangle1_ys[628]), .RECT1_WIDTH(rectangle1_widths[628]), .RECT1_HEIGHT(rectangle1_heights[628]), .RECT1_WEIGHT(rectangle1_weights[628]), .RECT2_X(rectangle2_xs[628]), .RECT2_Y(rectangle2_ys[628]), .RECT2_WIDTH(rectangle2_widths[628]), .RECT2_HEIGHT(rectangle2_heights[628]), .RECT2_WEIGHT(rectangle2_weights[628]), .RECT3_X(rectangle3_xs[628]), .RECT3_Y(rectangle3_ys[628]), .RECT3_WIDTH(rectangle3_widths[628]), .RECT3_HEIGHT(rectangle3_heights[628]), .RECT3_WEIGHT(rectangle3_weights[628]), .FEAT_THRES(feature_thresholds[628]), .FEAT_ABOVE(feature_aboves[628]), .FEAT_BELOW(feature_belows[628])) ac628(.scan_win(scan_win628), .scan_win_std_dev(scan_win_std_dev[628]), .feature_accum(feature_accums[628]));
  accum_calculator #(.RECT1_X(rectangle1_xs[629]), .RECT1_Y(rectangle1_ys[629]), .RECT1_WIDTH(rectangle1_widths[629]), .RECT1_HEIGHT(rectangle1_heights[629]), .RECT1_WEIGHT(rectangle1_weights[629]), .RECT2_X(rectangle2_xs[629]), .RECT2_Y(rectangle2_ys[629]), .RECT2_WIDTH(rectangle2_widths[629]), .RECT2_HEIGHT(rectangle2_heights[629]), .RECT2_WEIGHT(rectangle2_weights[629]), .RECT3_X(rectangle3_xs[629]), .RECT3_Y(rectangle3_ys[629]), .RECT3_WIDTH(rectangle3_widths[629]), .RECT3_HEIGHT(rectangle3_heights[629]), .RECT3_WEIGHT(rectangle3_weights[629]), .FEAT_THRES(feature_thresholds[629]), .FEAT_ABOVE(feature_aboves[629]), .FEAT_BELOW(feature_belows[629])) ac629(.scan_win(scan_win629), .scan_win_std_dev(scan_win_std_dev[629]), .feature_accum(feature_accums[629]));
  accum_calculator #(.RECT1_X(rectangle1_xs[630]), .RECT1_Y(rectangle1_ys[630]), .RECT1_WIDTH(rectangle1_widths[630]), .RECT1_HEIGHT(rectangle1_heights[630]), .RECT1_WEIGHT(rectangle1_weights[630]), .RECT2_X(rectangle2_xs[630]), .RECT2_Y(rectangle2_ys[630]), .RECT2_WIDTH(rectangle2_widths[630]), .RECT2_HEIGHT(rectangle2_heights[630]), .RECT2_WEIGHT(rectangle2_weights[630]), .RECT3_X(rectangle3_xs[630]), .RECT3_Y(rectangle3_ys[630]), .RECT3_WIDTH(rectangle3_widths[630]), .RECT3_HEIGHT(rectangle3_heights[630]), .RECT3_WEIGHT(rectangle3_weights[630]), .FEAT_THRES(feature_thresholds[630]), .FEAT_ABOVE(feature_aboves[630]), .FEAT_BELOW(feature_belows[630])) ac630(.scan_win(scan_win630), .scan_win_std_dev(scan_win_std_dev[630]), .feature_accum(feature_accums[630]));
  accum_calculator #(.RECT1_X(rectangle1_xs[631]), .RECT1_Y(rectangle1_ys[631]), .RECT1_WIDTH(rectangle1_widths[631]), .RECT1_HEIGHT(rectangle1_heights[631]), .RECT1_WEIGHT(rectangle1_weights[631]), .RECT2_X(rectangle2_xs[631]), .RECT2_Y(rectangle2_ys[631]), .RECT2_WIDTH(rectangle2_widths[631]), .RECT2_HEIGHT(rectangle2_heights[631]), .RECT2_WEIGHT(rectangle2_weights[631]), .RECT3_X(rectangle3_xs[631]), .RECT3_Y(rectangle3_ys[631]), .RECT3_WIDTH(rectangle3_widths[631]), .RECT3_HEIGHT(rectangle3_heights[631]), .RECT3_WEIGHT(rectangle3_weights[631]), .FEAT_THRES(feature_thresholds[631]), .FEAT_ABOVE(feature_aboves[631]), .FEAT_BELOW(feature_belows[631])) ac631(.scan_win(scan_win631), .scan_win_std_dev(scan_win_std_dev[631]), .feature_accum(feature_accums[631]));
  accum_calculator #(.RECT1_X(rectangle1_xs[632]), .RECT1_Y(rectangle1_ys[632]), .RECT1_WIDTH(rectangle1_widths[632]), .RECT1_HEIGHT(rectangle1_heights[632]), .RECT1_WEIGHT(rectangle1_weights[632]), .RECT2_X(rectangle2_xs[632]), .RECT2_Y(rectangle2_ys[632]), .RECT2_WIDTH(rectangle2_widths[632]), .RECT2_HEIGHT(rectangle2_heights[632]), .RECT2_WEIGHT(rectangle2_weights[632]), .RECT3_X(rectangle3_xs[632]), .RECT3_Y(rectangle3_ys[632]), .RECT3_WIDTH(rectangle3_widths[632]), .RECT3_HEIGHT(rectangle3_heights[632]), .RECT3_WEIGHT(rectangle3_weights[632]), .FEAT_THRES(feature_thresholds[632]), .FEAT_ABOVE(feature_aboves[632]), .FEAT_BELOW(feature_belows[632])) ac632(.scan_win(scan_win632), .scan_win_std_dev(scan_win_std_dev[632]), .feature_accum(feature_accums[632]));
  accum_calculator #(.RECT1_X(rectangle1_xs[633]), .RECT1_Y(rectangle1_ys[633]), .RECT1_WIDTH(rectangle1_widths[633]), .RECT1_HEIGHT(rectangle1_heights[633]), .RECT1_WEIGHT(rectangle1_weights[633]), .RECT2_X(rectangle2_xs[633]), .RECT2_Y(rectangle2_ys[633]), .RECT2_WIDTH(rectangle2_widths[633]), .RECT2_HEIGHT(rectangle2_heights[633]), .RECT2_WEIGHT(rectangle2_weights[633]), .RECT3_X(rectangle3_xs[633]), .RECT3_Y(rectangle3_ys[633]), .RECT3_WIDTH(rectangle3_widths[633]), .RECT3_HEIGHT(rectangle3_heights[633]), .RECT3_WEIGHT(rectangle3_weights[633]), .FEAT_THRES(feature_thresholds[633]), .FEAT_ABOVE(feature_aboves[633]), .FEAT_BELOW(feature_belows[633])) ac633(.scan_win(scan_win633), .scan_win_std_dev(scan_win_std_dev[633]), .feature_accum(feature_accums[633]));
  accum_calculator #(.RECT1_X(rectangle1_xs[634]), .RECT1_Y(rectangle1_ys[634]), .RECT1_WIDTH(rectangle1_widths[634]), .RECT1_HEIGHT(rectangle1_heights[634]), .RECT1_WEIGHT(rectangle1_weights[634]), .RECT2_X(rectangle2_xs[634]), .RECT2_Y(rectangle2_ys[634]), .RECT2_WIDTH(rectangle2_widths[634]), .RECT2_HEIGHT(rectangle2_heights[634]), .RECT2_WEIGHT(rectangle2_weights[634]), .RECT3_X(rectangle3_xs[634]), .RECT3_Y(rectangle3_ys[634]), .RECT3_WIDTH(rectangle3_widths[634]), .RECT3_HEIGHT(rectangle3_heights[634]), .RECT3_WEIGHT(rectangle3_weights[634]), .FEAT_THRES(feature_thresholds[634]), .FEAT_ABOVE(feature_aboves[634]), .FEAT_BELOW(feature_belows[634])) ac634(.scan_win(scan_win634), .scan_win_std_dev(scan_win_std_dev[634]), .feature_accum(feature_accums[634]));
  accum_calculator #(.RECT1_X(rectangle1_xs[635]), .RECT1_Y(rectangle1_ys[635]), .RECT1_WIDTH(rectangle1_widths[635]), .RECT1_HEIGHT(rectangle1_heights[635]), .RECT1_WEIGHT(rectangle1_weights[635]), .RECT2_X(rectangle2_xs[635]), .RECT2_Y(rectangle2_ys[635]), .RECT2_WIDTH(rectangle2_widths[635]), .RECT2_HEIGHT(rectangle2_heights[635]), .RECT2_WEIGHT(rectangle2_weights[635]), .RECT3_X(rectangle3_xs[635]), .RECT3_Y(rectangle3_ys[635]), .RECT3_WIDTH(rectangle3_widths[635]), .RECT3_HEIGHT(rectangle3_heights[635]), .RECT3_WEIGHT(rectangle3_weights[635]), .FEAT_THRES(feature_thresholds[635]), .FEAT_ABOVE(feature_aboves[635]), .FEAT_BELOW(feature_belows[635])) ac635(.scan_win(scan_win635), .scan_win_std_dev(scan_win_std_dev[635]), .feature_accum(feature_accums[635]));
  accum_calculator #(.RECT1_X(rectangle1_xs[636]), .RECT1_Y(rectangle1_ys[636]), .RECT1_WIDTH(rectangle1_widths[636]), .RECT1_HEIGHT(rectangle1_heights[636]), .RECT1_WEIGHT(rectangle1_weights[636]), .RECT2_X(rectangle2_xs[636]), .RECT2_Y(rectangle2_ys[636]), .RECT2_WIDTH(rectangle2_widths[636]), .RECT2_HEIGHT(rectangle2_heights[636]), .RECT2_WEIGHT(rectangle2_weights[636]), .RECT3_X(rectangle3_xs[636]), .RECT3_Y(rectangle3_ys[636]), .RECT3_WIDTH(rectangle3_widths[636]), .RECT3_HEIGHT(rectangle3_heights[636]), .RECT3_WEIGHT(rectangle3_weights[636]), .FEAT_THRES(feature_thresholds[636]), .FEAT_ABOVE(feature_aboves[636]), .FEAT_BELOW(feature_belows[636])) ac636(.scan_win(scan_win636), .scan_win_std_dev(scan_win_std_dev[636]), .feature_accum(feature_accums[636]));
  accum_calculator #(.RECT1_X(rectangle1_xs[637]), .RECT1_Y(rectangle1_ys[637]), .RECT1_WIDTH(rectangle1_widths[637]), .RECT1_HEIGHT(rectangle1_heights[637]), .RECT1_WEIGHT(rectangle1_weights[637]), .RECT2_X(rectangle2_xs[637]), .RECT2_Y(rectangle2_ys[637]), .RECT2_WIDTH(rectangle2_widths[637]), .RECT2_HEIGHT(rectangle2_heights[637]), .RECT2_WEIGHT(rectangle2_weights[637]), .RECT3_X(rectangle3_xs[637]), .RECT3_Y(rectangle3_ys[637]), .RECT3_WIDTH(rectangle3_widths[637]), .RECT3_HEIGHT(rectangle3_heights[637]), .RECT3_WEIGHT(rectangle3_weights[637]), .FEAT_THRES(feature_thresholds[637]), .FEAT_ABOVE(feature_aboves[637]), .FEAT_BELOW(feature_belows[637])) ac637(.scan_win(scan_win637), .scan_win_std_dev(scan_win_std_dev[637]), .feature_accum(feature_accums[637]));
  accum_calculator #(.RECT1_X(rectangle1_xs[638]), .RECT1_Y(rectangle1_ys[638]), .RECT1_WIDTH(rectangle1_widths[638]), .RECT1_HEIGHT(rectangle1_heights[638]), .RECT1_WEIGHT(rectangle1_weights[638]), .RECT2_X(rectangle2_xs[638]), .RECT2_Y(rectangle2_ys[638]), .RECT2_WIDTH(rectangle2_widths[638]), .RECT2_HEIGHT(rectangle2_heights[638]), .RECT2_WEIGHT(rectangle2_weights[638]), .RECT3_X(rectangle3_xs[638]), .RECT3_Y(rectangle3_ys[638]), .RECT3_WIDTH(rectangle3_widths[638]), .RECT3_HEIGHT(rectangle3_heights[638]), .RECT3_WEIGHT(rectangle3_weights[638]), .FEAT_THRES(feature_thresholds[638]), .FEAT_ABOVE(feature_aboves[638]), .FEAT_BELOW(feature_belows[638])) ac638(.scan_win(scan_win638), .scan_win_std_dev(scan_win_std_dev[638]), .feature_accum(feature_accums[638]));
  accum_calculator #(.RECT1_X(rectangle1_xs[639]), .RECT1_Y(rectangle1_ys[639]), .RECT1_WIDTH(rectangle1_widths[639]), .RECT1_HEIGHT(rectangle1_heights[639]), .RECT1_WEIGHT(rectangle1_weights[639]), .RECT2_X(rectangle2_xs[639]), .RECT2_Y(rectangle2_ys[639]), .RECT2_WIDTH(rectangle2_widths[639]), .RECT2_HEIGHT(rectangle2_heights[639]), .RECT2_WEIGHT(rectangle2_weights[639]), .RECT3_X(rectangle3_xs[639]), .RECT3_Y(rectangle3_ys[639]), .RECT3_WIDTH(rectangle3_widths[639]), .RECT3_HEIGHT(rectangle3_heights[639]), .RECT3_WEIGHT(rectangle3_weights[639]), .FEAT_THRES(feature_thresholds[639]), .FEAT_ABOVE(feature_aboves[639]), .FEAT_BELOW(feature_belows[639])) ac639(.scan_win(scan_win639), .scan_win_std_dev(scan_win_std_dev[639]), .feature_accum(feature_accums[639]));
  accum_calculator #(.RECT1_X(rectangle1_xs[640]), .RECT1_Y(rectangle1_ys[640]), .RECT1_WIDTH(rectangle1_widths[640]), .RECT1_HEIGHT(rectangle1_heights[640]), .RECT1_WEIGHT(rectangle1_weights[640]), .RECT2_X(rectangle2_xs[640]), .RECT2_Y(rectangle2_ys[640]), .RECT2_WIDTH(rectangle2_widths[640]), .RECT2_HEIGHT(rectangle2_heights[640]), .RECT2_WEIGHT(rectangle2_weights[640]), .RECT3_X(rectangle3_xs[640]), .RECT3_Y(rectangle3_ys[640]), .RECT3_WIDTH(rectangle3_widths[640]), .RECT3_HEIGHT(rectangle3_heights[640]), .RECT3_WEIGHT(rectangle3_weights[640]), .FEAT_THRES(feature_thresholds[640]), .FEAT_ABOVE(feature_aboves[640]), .FEAT_BELOW(feature_belows[640])) ac640(.scan_win(scan_win640), .scan_win_std_dev(scan_win_std_dev[640]), .feature_accum(feature_accums[640]));
  accum_calculator #(.RECT1_X(rectangle1_xs[641]), .RECT1_Y(rectangle1_ys[641]), .RECT1_WIDTH(rectangle1_widths[641]), .RECT1_HEIGHT(rectangle1_heights[641]), .RECT1_WEIGHT(rectangle1_weights[641]), .RECT2_X(rectangle2_xs[641]), .RECT2_Y(rectangle2_ys[641]), .RECT2_WIDTH(rectangle2_widths[641]), .RECT2_HEIGHT(rectangle2_heights[641]), .RECT2_WEIGHT(rectangle2_weights[641]), .RECT3_X(rectangle3_xs[641]), .RECT3_Y(rectangle3_ys[641]), .RECT3_WIDTH(rectangle3_widths[641]), .RECT3_HEIGHT(rectangle3_heights[641]), .RECT3_WEIGHT(rectangle3_weights[641]), .FEAT_THRES(feature_thresholds[641]), .FEAT_ABOVE(feature_aboves[641]), .FEAT_BELOW(feature_belows[641])) ac641(.scan_win(scan_win641), .scan_win_std_dev(scan_win_std_dev[641]), .feature_accum(feature_accums[641]));
  accum_calculator #(.RECT1_X(rectangle1_xs[642]), .RECT1_Y(rectangle1_ys[642]), .RECT1_WIDTH(rectangle1_widths[642]), .RECT1_HEIGHT(rectangle1_heights[642]), .RECT1_WEIGHT(rectangle1_weights[642]), .RECT2_X(rectangle2_xs[642]), .RECT2_Y(rectangle2_ys[642]), .RECT2_WIDTH(rectangle2_widths[642]), .RECT2_HEIGHT(rectangle2_heights[642]), .RECT2_WEIGHT(rectangle2_weights[642]), .RECT3_X(rectangle3_xs[642]), .RECT3_Y(rectangle3_ys[642]), .RECT3_WIDTH(rectangle3_widths[642]), .RECT3_HEIGHT(rectangle3_heights[642]), .RECT3_WEIGHT(rectangle3_weights[642]), .FEAT_THRES(feature_thresholds[642]), .FEAT_ABOVE(feature_aboves[642]), .FEAT_BELOW(feature_belows[642])) ac642(.scan_win(scan_win642), .scan_win_std_dev(scan_win_std_dev[642]), .feature_accum(feature_accums[642]));
  accum_calculator #(.RECT1_X(rectangle1_xs[643]), .RECT1_Y(rectangle1_ys[643]), .RECT1_WIDTH(rectangle1_widths[643]), .RECT1_HEIGHT(rectangle1_heights[643]), .RECT1_WEIGHT(rectangle1_weights[643]), .RECT2_X(rectangle2_xs[643]), .RECT2_Y(rectangle2_ys[643]), .RECT2_WIDTH(rectangle2_widths[643]), .RECT2_HEIGHT(rectangle2_heights[643]), .RECT2_WEIGHT(rectangle2_weights[643]), .RECT3_X(rectangle3_xs[643]), .RECT3_Y(rectangle3_ys[643]), .RECT3_WIDTH(rectangle3_widths[643]), .RECT3_HEIGHT(rectangle3_heights[643]), .RECT3_WEIGHT(rectangle3_weights[643]), .FEAT_THRES(feature_thresholds[643]), .FEAT_ABOVE(feature_aboves[643]), .FEAT_BELOW(feature_belows[643])) ac643(.scan_win(scan_win643), .scan_win_std_dev(scan_win_std_dev[643]), .feature_accum(feature_accums[643]));
  accum_calculator #(.RECT1_X(rectangle1_xs[644]), .RECT1_Y(rectangle1_ys[644]), .RECT1_WIDTH(rectangle1_widths[644]), .RECT1_HEIGHT(rectangle1_heights[644]), .RECT1_WEIGHT(rectangle1_weights[644]), .RECT2_X(rectangle2_xs[644]), .RECT2_Y(rectangle2_ys[644]), .RECT2_WIDTH(rectangle2_widths[644]), .RECT2_HEIGHT(rectangle2_heights[644]), .RECT2_WEIGHT(rectangle2_weights[644]), .RECT3_X(rectangle3_xs[644]), .RECT3_Y(rectangle3_ys[644]), .RECT3_WIDTH(rectangle3_widths[644]), .RECT3_HEIGHT(rectangle3_heights[644]), .RECT3_WEIGHT(rectangle3_weights[644]), .FEAT_THRES(feature_thresholds[644]), .FEAT_ABOVE(feature_aboves[644]), .FEAT_BELOW(feature_belows[644])) ac644(.scan_win(scan_win644), .scan_win_std_dev(scan_win_std_dev[644]), .feature_accum(feature_accums[644]));
  accum_calculator #(.RECT1_X(rectangle1_xs[645]), .RECT1_Y(rectangle1_ys[645]), .RECT1_WIDTH(rectangle1_widths[645]), .RECT1_HEIGHT(rectangle1_heights[645]), .RECT1_WEIGHT(rectangle1_weights[645]), .RECT2_X(rectangle2_xs[645]), .RECT2_Y(rectangle2_ys[645]), .RECT2_WIDTH(rectangle2_widths[645]), .RECT2_HEIGHT(rectangle2_heights[645]), .RECT2_WEIGHT(rectangle2_weights[645]), .RECT3_X(rectangle3_xs[645]), .RECT3_Y(rectangle3_ys[645]), .RECT3_WIDTH(rectangle3_widths[645]), .RECT3_HEIGHT(rectangle3_heights[645]), .RECT3_WEIGHT(rectangle3_weights[645]), .FEAT_THRES(feature_thresholds[645]), .FEAT_ABOVE(feature_aboves[645]), .FEAT_BELOW(feature_belows[645])) ac645(.scan_win(scan_win645), .scan_win_std_dev(scan_win_std_dev[645]), .feature_accum(feature_accums[645]));
  accum_calculator #(.RECT1_X(rectangle1_xs[646]), .RECT1_Y(rectangle1_ys[646]), .RECT1_WIDTH(rectangle1_widths[646]), .RECT1_HEIGHT(rectangle1_heights[646]), .RECT1_WEIGHT(rectangle1_weights[646]), .RECT2_X(rectangle2_xs[646]), .RECT2_Y(rectangle2_ys[646]), .RECT2_WIDTH(rectangle2_widths[646]), .RECT2_HEIGHT(rectangle2_heights[646]), .RECT2_WEIGHT(rectangle2_weights[646]), .RECT3_X(rectangle3_xs[646]), .RECT3_Y(rectangle3_ys[646]), .RECT3_WIDTH(rectangle3_widths[646]), .RECT3_HEIGHT(rectangle3_heights[646]), .RECT3_WEIGHT(rectangle3_weights[646]), .FEAT_THRES(feature_thresholds[646]), .FEAT_ABOVE(feature_aboves[646]), .FEAT_BELOW(feature_belows[646])) ac646(.scan_win(scan_win646), .scan_win_std_dev(scan_win_std_dev[646]), .feature_accum(feature_accums[646]));
  accum_calculator #(.RECT1_X(rectangle1_xs[647]), .RECT1_Y(rectangle1_ys[647]), .RECT1_WIDTH(rectangle1_widths[647]), .RECT1_HEIGHT(rectangle1_heights[647]), .RECT1_WEIGHT(rectangle1_weights[647]), .RECT2_X(rectangle2_xs[647]), .RECT2_Y(rectangle2_ys[647]), .RECT2_WIDTH(rectangle2_widths[647]), .RECT2_HEIGHT(rectangle2_heights[647]), .RECT2_WEIGHT(rectangle2_weights[647]), .RECT3_X(rectangle3_xs[647]), .RECT3_Y(rectangle3_ys[647]), .RECT3_WIDTH(rectangle3_widths[647]), .RECT3_HEIGHT(rectangle3_heights[647]), .RECT3_WEIGHT(rectangle3_weights[647]), .FEAT_THRES(feature_thresholds[647]), .FEAT_ABOVE(feature_aboves[647]), .FEAT_BELOW(feature_belows[647])) ac647(.scan_win(scan_win647), .scan_win_std_dev(scan_win_std_dev[647]), .feature_accum(feature_accums[647]));
  accum_calculator #(.RECT1_X(rectangle1_xs[648]), .RECT1_Y(rectangle1_ys[648]), .RECT1_WIDTH(rectangle1_widths[648]), .RECT1_HEIGHT(rectangle1_heights[648]), .RECT1_WEIGHT(rectangle1_weights[648]), .RECT2_X(rectangle2_xs[648]), .RECT2_Y(rectangle2_ys[648]), .RECT2_WIDTH(rectangle2_widths[648]), .RECT2_HEIGHT(rectangle2_heights[648]), .RECT2_WEIGHT(rectangle2_weights[648]), .RECT3_X(rectangle3_xs[648]), .RECT3_Y(rectangle3_ys[648]), .RECT3_WIDTH(rectangle3_widths[648]), .RECT3_HEIGHT(rectangle3_heights[648]), .RECT3_WEIGHT(rectangle3_weights[648]), .FEAT_THRES(feature_thresholds[648]), .FEAT_ABOVE(feature_aboves[648]), .FEAT_BELOW(feature_belows[648])) ac648(.scan_win(scan_win648), .scan_win_std_dev(scan_win_std_dev[648]), .feature_accum(feature_accums[648]));
  accum_calculator #(.RECT1_X(rectangle1_xs[649]), .RECT1_Y(rectangle1_ys[649]), .RECT1_WIDTH(rectangle1_widths[649]), .RECT1_HEIGHT(rectangle1_heights[649]), .RECT1_WEIGHT(rectangle1_weights[649]), .RECT2_X(rectangle2_xs[649]), .RECT2_Y(rectangle2_ys[649]), .RECT2_WIDTH(rectangle2_widths[649]), .RECT2_HEIGHT(rectangle2_heights[649]), .RECT2_WEIGHT(rectangle2_weights[649]), .RECT3_X(rectangle3_xs[649]), .RECT3_Y(rectangle3_ys[649]), .RECT3_WIDTH(rectangle3_widths[649]), .RECT3_HEIGHT(rectangle3_heights[649]), .RECT3_WEIGHT(rectangle3_weights[649]), .FEAT_THRES(feature_thresholds[649]), .FEAT_ABOVE(feature_aboves[649]), .FEAT_BELOW(feature_belows[649])) ac649(.scan_win(scan_win649), .scan_win_std_dev(scan_win_std_dev[649]), .feature_accum(feature_accums[649]));
  accum_calculator #(.RECT1_X(rectangle1_xs[650]), .RECT1_Y(rectangle1_ys[650]), .RECT1_WIDTH(rectangle1_widths[650]), .RECT1_HEIGHT(rectangle1_heights[650]), .RECT1_WEIGHT(rectangle1_weights[650]), .RECT2_X(rectangle2_xs[650]), .RECT2_Y(rectangle2_ys[650]), .RECT2_WIDTH(rectangle2_widths[650]), .RECT2_HEIGHT(rectangle2_heights[650]), .RECT2_WEIGHT(rectangle2_weights[650]), .RECT3_X(rectangle3_xs[650]), .RECT3_Y(rectangle3_ys[650]), .RECT3_WIDTH(rectangle3_widths[650]), .RECT3_HEIGHT(rectangle3_heights[650]), .RECT3_WEIGHT(rectangle3_weights[650]), .FEAT_THRES(feature_thresholds[650]), .FEAT_ABOVE(feature_aboves[650]), .FEAT_BELOW(feature_belows[650])) ac650(.scan_win(scan_win650), .scan_win_std_dev(scan_win_std_dev[650]), .feature_accum(feature_accums[650]));
  accum_calculator #(.RECT1_X(rectangle1_xs[651]), .RECT1_Y(rectangle1_ys[651]), .RECT1_WIDTH(rectangle1_widths[651]), .RECT1_HEIGHT(rectangle1_heights[651]), .RECT1_WEIGHT(rectangle1_weights[651]), .RECT2_X(rectangle2_xs[651]), .RECT2_Y(rectangle2_ys[651]), .RECT2_WIDTH(rectangle2_widths[651]), .RECT2_HEIGHT(rectangle2_heights[651]), .RECT2_WEIGHT(rectangle2_weights[651]), .RECT3_X(rectangle3_xs[651]), .RECT3_Y(rectangle3_ys[651]), .RECT3_WIDTH(rectangle3_widths[651]), .RECT3_HEIGHT(rectangle3_heights[651]), .RECT3_WEIGHT(rectangle3_weights[651]), .FEAT_THRES(feature_thresholds[651]), .FEAT_ABOVE(feature_aboves[651]), .FEAT_BELOW(feature_belows[651])) ac651(.scan_win(scan_win651), .scan_win_std_dev(scan_win_std_dev[651]), .feature_accum(feature_accums[651]));
  accum_calculator #(.RECT1_X(rectangle1_xs[652]), .RECT1_Y(rectangle1_ys[652]), .RECT1_WIDTH(rectangle1_widths[652]), .RECT1_HEIGHT(rectangle1_heights[652]), .RECT1_WEIGHT(rectangle1_weights[652]), .RECT2_X(rectangle2_xs[652]), .RECT2_Y(rectangle2_ys[652]), .RECT2_WIDTH(rectangle2_widths[652]), .RECT2_HEIGHT(rectangle2_heights[652]), .RECT2_WEIGHT(rectangle2_weights[652]), .RECT3_X(rectangle3_xs[652]), .RECT3_Y(rectangle3_ys[652]), .RECT3_WIDTH(rectangle3_widths[652]), .RECT3_HEIGHT(rectangle3_heights[652]), .RECT3_WEIGHT(rectangle3_weights[652]), .FEAT_THRES(feature_thresholds[652]), .FEAT_ABOVE(feature_aboves[652]), .FEAT_BELOW(feature_belows[652])) ac652(.scan_win(scan_win652), .scan_win_std_dev(scan_win_std_dev[652]), .feature_accum(feature_accums[652]));
  accum_calculator #(.RECT1_X(rectangle1_xs[653]), .RECT1_Y(rectangle1_ys[653]), .RECT1_WIDTH(rectangle1_widths[653]), .RECT1_HEIGHT(rectangle1_heights[653]), .RECT1_WEIGHT(rectangle1_weights[653]), .RECT2_X(rectangle2_xs[653]), .RECT2_Y(rectangle2_ys[653]), .RECT2_WIDTH(rectangle2_widths[653]), .RECT2_HEIGHT(rectangle2_heights[653]), .RECT2_WEIGHT(rectangle2_weights[653]), .RECT3_X(rectangle3_xs[653]), .RECT3_Y(rectangle3_ys[653]), .RECT3_WIDTH(rectangle3_widths[653]), .RECT3_HEIGHT(rectangle3_heights[653]), .RECT3_WEIGHT(rectangle3_weights[653]), .FEAT_THRES(feature_thresholds[653]), .FEAT_ABOVE(feature_aboves[653]), .FEAT_BELOW(feature_belows[653])) ac653(.scan_win(scan_win653), .scan_win_std_dev(scan_win_std_dev[653]), .feature_accum(feature_accums[653]));
  accum_calculator #(.RECT1_X(rectangle1_xs[654]), .RECT1_Y(rectangle1_ys[654]), .RECT1_WIDTH(rectangle1_widths[654]), .RECT1_HEIGHT(rectangle1_heights[654]), .RECT1_WEIGHT(rectangle1_weights[654]), .RECT2_X(rectangle2_xs[654]), .RECT2_Y(rectangle2_ys[654]), .RECT2_WIDTH(rectangle2_widths[654]), .RECT2_HEIGHT(rectangle2_heights[654]), .RECT2_WEIGHT(rectangle2_weights[654]), .RECT3_X(rectangle3_xs[654]), .RECT3_Y(rectangle3_ys[654]), .RECT3_WIDTH(rectangle3_widths[654]), .RECT3_HEIGHT(rectangle3_heights[654]), .RECT3_WEIGHT(rectangle3_weights[654]), .FEAT_THRES(feature_thresholds[654]), .FEAT_ABOVE(feature_aboves[654]), .FEAT_BELOW(feature_belows[654])) ac654(.scan_win(scan_win654), .scan_win_std_dev(scan_win_std_dev[654]), .feature_accum(feature_accums[654]));
  accum_calculator #(.RECT1_X(rectangle1_xs[655]), .RECT1_Y(rectangle1_ys[655]), .RECT1_WIDTH(rectangle1_widths[655]), .RECT1_HEIGHT(rectangle1_heights[655]), .RECT1_WEIGHT(rectangle1_weights[655]), .RECT2_X(rectangle2_xs[655]), .RECT2_Y(rectangle2_ys[655]), .RECT2_WIDTH(rectangle2_widths[655]), .RECT2_HEIGHT(rectangle2_heights[655]), .RECT2_WEIGHT(rectangle2_weights[655]), .RECT3_X(rectangle3_xs[655]), .RECT3_Y(rectangle3_ys[655]), .RECT3_WIDTH(rectangle3_widths[655]), .RECT3_HEIGHT(rectangle3_heights[655]), .RECT3_WEIGHT(rectangle3_weights[655]), .FEAT_THRES(feature_thresholds[655]), .FEAT_ABOVE(feature_aboves[655]), .FEAT_BELOW(feature_belows[655])) ac655(.scan_win(scan_win655), .scan_win_std_dev(scan_win_std_dev[655]), .feature_accum(feature_accums[655]));
  accum_calculator #(.RECT1_X(rectangle1_xs[656]), .RECT1_Y(rectangle1_ys[656]), .RECT1_WIDTH(rectangle1_widths[656]), .RECT1_HEIGHT(rectangle1_heights[656]), .RECT1_WEIGHT(rectangle1_weights[656]), .RECT2_X(rectangle2_xs[656]), .RECT2_Y(rectangle2_ys[656]), .RECT2_WIDTH(rectangle2_widths[656]), .RECT2_HEIGHT(rectangle2_heights[656]), .RECT2_WEIGHT(rectangle2_weights[656]), .RECT3_X(rectangle3_xs[656]), .RECT3_Y(rectangle3_ys[656]), .RECT3_WIDTH(rectangle3_widths[656]), .RECT3_HEIGHT(rectangle3_heights[656]), .RECT3_WEIGHT(rectangle3_weights[656]), .FEAT_THRES(feature_thresholds[656]), .FEAT_ABOVE(feature_aboves[656]), .FEAT_BELOW(feature_belows[656])) ac656(.scan_win(scan_win656), .scan_win_std_dev(scan_win_std_dev[656]), .feature_accum(feature_accums[656]));
  accum_calculator #(.RECT1_X(rectangle1_xs[657]), .RECT1_Y(rectangle1_ys[657]), .RECT1_WIDTH(rectangle1_widths[657]), .RECT1_HEIGHT(rectangle1_heights[657]), .RECT1_WEIGHT(rectangle1_weights[657]), .RECT2_X(rectangle2_xs[657]), .RECT2_Y(rectangle2_ys[657]), .RECT2_WIDTH(rectangle2_widths[657]), .RECT2_HEIGHT(rectangle2_heights[657]), .RECT2_WEIGHT(rectangle2_weights[657]), .RECT3_X(rectangle3_xs[657]), .RECT3_Y(rectangle3_ys[657]), .RECT3_WIDTH(rectangle3_widths[657]), .RECT3_HEIGHT(rectangle3_heights[657]), .RECT3_WEIGHT(rectangle3_weights[657]), .FEAT_THRES(feature_thresholds[657]), .FEAT_ABOVE(feature_aboves[657]), .FEAT_BELOW(feature_belows[657])) ac657(.scan_win(scan_win657), .scan_win_std_dev(scan_win_std_dev[657]), .feature_accum(feature_accums[657]));
  accum_calculator #(.RECT1_X(rectangle1_xs[658]), .RECT1_Y(rectangle1_ys[658]), .RECT1_WIDTH(rectangle1_widths[658]), .RECT1_HEIGHT(rectangle1_heights[658]), .RECT1_WEIGHT(rectangle1_weights[658]), .RECT2_X(rectangle2_xs[658]), .RECT2_Y(rectangle2_ys[658]), .RECT2_WIDTH(rectangle2_widths[658]), .RECT2_HEIGHT(rectangle2_heights[658]), .RECT2_WEIGHT(rectangle2_weights[658]), .RECT3_X(rectangle3_xs[658]), .RECT3_Y(rectangle3_ys[658]), .RECT3_WIDTH(rectangle3_widths[658]), .RECT3_HEIGHT(rectangle3_heights[658]), .RECT3_WEIGHT(rectangle3_weights[658]), .FEAT_THRES(feature_thresholds[658]), .FEAT_ABOVE(feature_aboves[658]), .FEAT_BELOW(feature_belows[658])) ac658(.scan_win(scan_win658), .scan_win_std_dev(scan_win_std_dev[658]), .feature_accum(feature_accums[658]));
  accum_calculator #(.RECT1_X(rectangle1_xs[659]), .RECT1_Y(rectangle1_ys[659]), .RECT1_WIDTH(rectangle1_widths[659]), .RECT1_HEIGHT(rectangle1_heights[659]), .RECT1_WEIGHT(rectangle1_weights[659]), .RECT2_X(rectangle2_xs[659]), .RECT2_Y(rectangle2_ys[659]), .RECT2_WIDTH(rectangle2_widths[659]), .RECT2_HEIGHT(rectangle2_heights[659]), .RECT2_WEIGHT(rectangle2_weights[659]), .RECT3_X(rectangle3_xs[659]), .RECT3_Y(rectangle3_ys[659]), .RECT3_WIDTH(rectangle3_widths[659]), .RECT3_HEIGHT(rectangle3_heights[659]), .RECT3_WEIGHT(rectangle3_weights[659]), .FEAT_THRES(feature_thresholds[659]), .FEAT_ABOVE(feature_aboves[659]), .FEAT_BELOW(feature_belows[659])) ac659(.scan_win(scan_win659), .scan_win_std_dev(scan_win_std_dev[659]), .feature_accum(feature_accums[659]));
  accum_calculator #(.RECT1_X(rectangle1_xs[660]), .RECT1_Y(rectangle1_ys[660]), .RECT1_WIDTH(rectangle1_widths[660]), .RECT1_HEIGHT(rectangle1_heights[660]), .RECT1_WEIGHT(rectangle1_weights[660]), .RECT2_X(rectangle2_xs[660]), .RECT2_Y(rectangle2_ys[660]), .RECT2_WIDTH(rectangle2_widths[660]), .RECT2_HEIGHT(rectangle2_heights[660]), .RECT2_WEIGHT(rectangle2_weights[660]), .RECT3_X(rectangle3_xs[660]), .RECT3_Y(rectangle3_ys[660]), .RECT3_WIDTH(rectangle3_widths[660]), .RECT3_HEIGHT(rectangle3_heights[660]), .RECT3_WEIGHT(rectangle3_weights[660]), .FEAT_THRES(feature_thresholds[660]), .FEAT_ABOVE(feature_aboves[660]), .FEAT_BELOW(feature_belows[660])) ac660(.scan_win(scan_win660), .scan_win_std_dev(scan_win_std_dev[660]), .feature_accum(feature_accums[660]));
  accum_calculator #(.RECT1_X(rectangle1_xs[661]), .RECT1_Y(rectangle1_ys[661]), .RECT1_WIDTH(rectangle1_widths[661]), .RECT1_HEIGHT(rectangle1_heights[661]), .RECT1_WEIGHT(rectangle1_weights[661]), .RECT2_X(rectangle2_xs[661]), .RECT2_Y(rectangle2_ys[661]), .RECT2_WIDTH(rectangle2_widths[661]), .RECT2_HEIGHT(rectangle2_heights[661]), .RECT2_WEIGHT(rectangle2_weights[661]), .RECT3_X(rectangle3_xs[661]), .RECT3_Y(rectangle3_ys[661]), .RECT3_WIDTH(rectangle3_widths[661]), .RECT3_HEIGHT(rectangle3_heights[661]), .RECT3_WEIGHT(rectangle3_weights[661]), .FEAT_THRES(feature_thresholds[661]), .FEAT_ABOVE(feature_aboves[661]), .FEAT_BELOW(feature_belows[661])) ac661(.scan_win(scan_win661), .scan_win_std_dev(scan_win_std_dev[661]), .feature_accum(feature_accums[661]));
  accum_calculator #(.RECT1_X(rectangle1_xs[662]), .RECT1_Y(rectangle1_ys[662]), .RECT1_WIDTH(rectangle1_widths[662]), .RECT1_HEIGHT(rectangle1_heights[662]), .RECT1_WEIGHT(rectangle1_weights[662]), .RECT2_X(rectangle2_xs[662]), .RECT2_Y(rectangle2_ys[662]), .RECT2_WIDTH(rectangle2_widths[662]), .RECT2_HEIGHT(rectangle2_heights[662]), .RECT2_WEIGHT(rectangle2_weights[662]), .RECT3_X(rectangle3_xs[662]), .RECT3_Y(rectangle3_ys[662]), .RECT3_WIDTH(rectangle3_widths[662]), .RECT3_HEIGHT(rectangle3_heights[662]), .RECT3_WEIGHT(rectangle3_weights[662]), .FEAT_THRES(feature_thresholds[662]), .FEAT_ABOVE(feature_aboves[662]), .FEAT_BELOW(feature_belows[662])) ac662(.scan_win(scan_win662), .scan_win_std_dev(scan_win_std_dev[662]), .feature_accum(feature_accums[662]));
  accum_calculator #(.RECT1_X(rectangle1_xs[663]), .RECT1_Y(rectangle1_ys[663]), .RECT1_WIDTH(rectangle1_widths[663]), .RECT1_HEIGHT(rectangle1_heights[663]), .RECT1_WEIGHT(rectangle1_weights[663]), .RECT2_X(rectangle2_xs[663]), .RECT2_Y(rectangle2_ys[663]), .RECT2_WIDTH(rectangle2_widths[663]), .RECT2_HEIGHT(rectangle2_heights[663]), .RECT2_WEIGHT(rectangle2_weights[663]), .RECT3_X(rectangle3_xs[663]), .RECT3_Y(rectangle3_ys[663]), .RECT3_WIDTH(rectangle3_widths[663]), .RECT3_HEIGHT(rectangle3_heights[663]), .RECT3_WEIGHT(rectangle3_weights[663]), .FEAT_THRES(feature_thresholds[663]), .FEAT_ABOVE(feature_aboves[663]), .FEAT_BELOW(feature_belows[663])) ac663(.scan_win(scan_win663), .scan_win_std_dev(scan_win_std_dev[663]), .feature_accum(feature_accums[663]));
  accum_calculator #(.RECT1_X(rectangle1_xs[664]), .RECT1_Y(rectangle1_ys[664]), .RECT1_WIDTH(rectangle1_widths[664]), .RECT1_HEIGHT(rectangle1_heights[664]), .RECT1_WEIGHT(rectangle1_weights[664]), .RECT2_X(rectangle2_xs[664]), .RECT2_Y(rectangle2_ys[664]), .RECT2_WIDTH(rectangle2_widths[664]), .RECT2_HEIGHT(rectangle2_heights[664]), .RECT2_WEIGHT(rectangle2_weights[664]), .RECT3_X(rectangle3_xs[664]), .RECT3_Y(rectangle3_ys[664]), .RECT3_WIDTH(rectangle3_widths[664]), .RECT3_HEIGHT(rectangle3_heights[664]), .RECT3_WEIGHT(rectangle3_weights[664]), .FEAT_THRES(feature_thresholds[664]), .FEAT_ABOVE(feature_aboves[664]), .FEAT_BELOW(feature_belows[664])) ac664(.scan_win(scan_win664), .scan_win_std_dev(scan_win_std_dev[664]), .feature_accum(feature_accums[664]));
  accum_calculator #(.RECT1_X(rectangle1_xs[665]), .RECT1_Y(rectangle1_ys[665]), .RECT1_WIDTH(rectangle1_widths[665]), .RECT1_HEIGHT(rectangle1_heights[665]), .RECT1_WEIGHT(rectangle1_weights[665]), .RECT2_X(rectangle2_xs[665]), .RECT2_Y(rectangle2_ys[665]), .RECT2_WIDTH(rectangle2_widths[665]), .RECT2_HEIGHT(rectangle2_heights[665]), .RECT2_WEIGHT(rectangle2_weights[665]), .RECT3_X(rectangle3_xs[665]), .RECT3_Y(rectangle3_ys[665]), .RECT3_WIDTH(rectangle3_widths[665]), .RECT3_HEIGHT(rectangle3_heights[665]), .RECT3_WEIGHT(rectangle3_weights[665]), .FEAT_THRES(feature_thresholds[665]), .FEAT_ABOVE(feature_aboves[665]), .FEAT_BELOW(feature_belows[665])) ac665(.scan_win(scan_win665), .scan_win_std_dev(scan_win_std_dev[665]), .feature_accum(feature_accums[665]));
  accum_calculator #(.RECT1_X(rectangle1_xs[666]), .RECT1_Y(rectangle1_ys[666]), .RECT1_WIDTH(rectangle1_widths[666]), .RECT1_HEIGHT(rectangle1_heights[666]), .RECT1_WEIGHT(rectangle1_weights[666]), .RECT2_X(rectangle2_xs[666]), .RECT2_Y(rectangle2_ys[666]), .RECT2_WIDTH(rectangle2_widths[666]), .RECT2_HEIGHT(rectangle2_heights[666]), .RECT2_WEIGHT(rectangle2_weights[666]), .RECT3_X(rectangle3_xs[666]), .RECT3_Y(rectangle3_ys[666]), .RECT3_WIDTH(rectangle3_widths[666]), .RECT3_HEIGHT(rectangle3_heights[666]), .RECT3_WEIGHT(rectangle3_weights[666]), .FEAT_THRES(feature_thresholds[666]), .FEAT_ABOVE(feature_aboves[666]), .FEAT_BELOW(feature_belows[666])) ac666(.scan_win(scan_win666), .scan_win_std_dev(scan_win_std_dev[666]), .feature_accum(feature_accums[666]));
  accum_calculator #(.RECT1_X(rectangle1_xs[667]), .RECT1_Y(rectangle1_ys[667]), .RECT1_WIDTH(rectangle1_widths[667]), .RECT1_HEIGHT(rectangle1_heights[667]), .RECT1_WEIGHT(rectangle1_weights[667]), .RECT2_X(rectangle2_xs[667]), .RECT2_Y(rectangle2_ys[667]), .RECT2_WIDTH(rectangle2_widths[667]), .RECT2_HEIGHT(rectangle2_heights[667]), .RECT2_WEIGHT(rectangle2_weights[667]), .RECT3_X(rectangle3_xs[667]), .RECT3_Y(rectangle3_ys[667]), .RECT3_WIDTH(rectangle3_widths[667]), .RECT3_HEIGHT(rectangle3_heights[667]), .RECT3_WEIGHT(rectangle3_weights[667]), .FEAT_THRES(feature_thresholds[667]), .FEAT_ABOVE(feature_aboves[667]), .FEAT_BELOW(feature_belows[667])) ac667(.scan_win(scan_win667), .scan_win_std_dev(scan_win_std_dev[667]), .feature_accum(feature_accums[667]));
  accum_calculator #(.RECT1_X(rectangle1_xs[668]), .RECT1_Y(rectangle1_ys[668]), .RECT1_WIDTH(rectangle1_widths[668]), .RECT1_HEIGHT(rectangle1_heights[668]), .RECT1_WEIGHT(rectangle1_weights[668]), .RECT2_X(rectangle2_xs[668]), .RECT2_Y(rectangle2_ys[668]), .RECT2_WIDTH(rectangle2_widths[668]), .RECT2_HEIGHT(rectangle2_heights[668]), .RECT2_WEIGHT(rectangle2_weights[668]), .RECT3_X(rectangle3_xs[668]), .RECT3_Y(rectangle3_ys[668]), .RECT3_WIDTH(rectangle3_widths[668]), .RECT3_HEIGHT(rectangle3_heights[668]), .RECT3_WEIGHT(rectangle3_weights[668]), .FEAT_THRES(feature_thresholds[668]), .FEAT_ABOVE(feature_aboves[668]), .FEAT_BELOW(feature_belows[668])) ac668(.scan_win(scan_win668), .scan_win_std_dev(scan_win_std_dev[668]), .feature_accum(feature_accums[668]));
  accum_calculator #(.RECT1_X(rectangle1_xs[669]), .RECT1_Y(rectangle1_ys[669]), .RECT1_WIDTH(rectangle1_widths[669]), .RECT1_HEIGHT(rectangle1_heights[669]), .RECT1_WEIGHT(rectangle1_weights[669]), .RECT2_X(rectangle2_xs[669]), .RECT2_Y(rectangle2_ys[669]), .RECT2_WIDTH(rectangle2_widths[669]), .RECT2_HEIGHT(rectangle2_heights[669]), .RECT2_WEIGHT(rectangle2_weights[669]), .RECT3_X(rectangle3_xs[669]), .RECT3_Y(rectangle3_ys[669]), .RECT3_WIDTH(rectangle3_widths[669]), .RECT3_HEIGHT(rectangle3_heights[669]), .RECT3_WEIGHT(rectangle3_weights[669]), .FEAT_THRES(feature_thresholds[669]), .FEAT_ABOVE(feature_aboves[669]), .FEAT_BELOW(feature_belows[669])) ac669(.scan_win(scan_win669), .scan_win_std_dev(scan_win_std_dev[669]), .feature_accum(feature_accums[669]));
  accum_calculator #(.RECT1_X(rectangle1_xs[670]), .RECT1_Y(rectangle1_ys[670]), .RECT1_WIDTH(rectangle1_widths[670]), .RECT1_HEIGHT(rectangle1_heights[670]), .RECT1_WEIGHT(rectangle1_weights[670]), .RECT2_X(rectangle2_xs[670]), .RECT2_Y(rectangle2_ys[670]), .RECT2_WIDTH(rectangle2_widths[670]), .RECT2_HEIGHT(rectangle2_heights[670]), .RECT2_WEIGHT(rectangle2_weights[670]), .RECT3_X(rectangle3_xs[670]), .RECT3_Y(rectangle3_ys[670]), .RECT3_WIDTH(rectangle3_widths[670]), .RECT3_HEIGHT(rectangle3_heights[670]), .RECT3_WEIGHT(rectangle3_weights[670]), .FEAT_THRES(feature_thresholds[670]), .FEAT_ABOVE(feature_aboves[670]), .FEAT_BELOW(feature_belows[670])) ac670(.scan_win(scan_win670), .scan_win_std_dev(scan_win_std_dev[670]), .feature_accum(feature_accums[670]));
  accum_calculator #(.RECT1_X(rectangle1_xs[671]), .RECT1_Y(rectangle1_ys[671]), .RECT1_WIDTH(rectangle1_widths[671]), .RECT1_HEIGHT(rectangle1_heights[671]), .RECT1_WEIGHT(rectangle1_weights[671]), .RECT2_X(rectangle2_xs[671]), .RECT2_Y(rectangle2_ys[671]), .RECT2_WIDTH(rectangle2_widths[671]), .RECT2_HEIGHT(rectangle2_heights[671]), .RECT2_WEIGHT(rectangle2_weights[671]), .RECT3_X(rectangle3_xs[671]), .RECT3_Y(rectangle3_ys[671]), .RECT3_WIDTH(rectangle3_widths[671]), .RECT3_HEIGHT(rectangle3_heights[671]), .RECT3_WEIGHT(rectangle3_weights[671]), .FEAT_THRES(feature_thresholds[671]), .FEAT_ABOVE(feature_aboves[671]), .FEAT_BELOW(feature_belows[671])) ac671(.scan_win(scan_win671), .scan_win_std_dev(scan_win_std_dev[671]), .feature_accum(feature_accums[671]));
  accum_calculator #(.RECT1_X(rectangle1_xs[672]), .RECT1_Y(rectangle1_ys[672]), .RECT1_WIDTH(rectangle1_widths[672]), .RECT1_HEIGHT(rectangle1_heights[672]), .RECT1_WEIGHT(rectangle1_weights[672]), .RECT2_X(rectangle2_xs[672]), .RECT2_Y(rectangle2_ys[672]), .RECT2_WIDTH(rectangle2_widths[672]), .RECT2_HEIGHT(rectangle2_heights[672]), .RECT2_WEIGHT(rectangle2_weights[672]), .RECT3_X(rectangle3_xs[672]), .RECT3_Y(rectangle3_ys[672]), .RECT3_WIDTH(rectangle3_widths[672]), .RECT3_HEIGHT(rectangle3_heights[672]), .RECT3_WEIGHT(rectangle3_weights[672]), .FEAT_THRES(feature_thresholds[672]), .FEAT_ABOVE(feature_aboves[672]), .FEAT_BELOW(feature_belows[672])) ac672(.scan_win(scan_win672), .scan_win_std_dev(scan_win_std_dev[672]), .feature_accum(feature_accums[672]));
  accum_calculator #(.RECT1_X(rectangle1_xs[673]), .RECT1_Y(rectangle1_ys[673]), .RECT1_WIDTH(rectangle1_widths[673]), .RECT1_HEIGHT(rectangle1_heights[673]), .RECT1_WEIGHT(rectangle1_weights[673]), .RECT2_X(rectangle2_xs[673]), .RECT2_Y(rectangle2_ys[673]), .RECT2_WIDTH(rectangle2_widths[673]), .RECT2_HEIGHT(rectangle2_heights[673]), .RECT2_WEIGHT(rectangle2_weights[673]), .RECT3_X(rectangle3_xs[673]), .RECT3_Y(rectangle3_ys[673]), .RECT3_WIDTH(rectangle3_widths[673]), .RECT3_HEIGHT(rectangle3_heights[673]), .RECT3_WEIGHT(rectangle3_weights[673]), .FEAT_THRES(feature_thresholds[673]), .FEAT_ABOVE(feature_aboves[673]), .FEAT_BELOW(feature_belows[673])) ac673(.scan_win(scan_win673), .scan_win_std_dev(scan_win_std_dev[673]), .feature_accum(feature_accums[673]));
  accum_calculator #(.RECT1_X(rectangle1_xs[674]), .RECT1_Y(rectangle1_ys[674]), .RECT1_WIDTH(rectangle1_widths[674]), .RECT1_HEIGHT(rectangle1_heights[674]), .RECT1_WEIGHT(rectangle1_weights[674]), .RECT2_X(rectangle2_xs[674]), .RECT2_Y(rectangle2_ys[674]), .RECT2_WIDTH(rectangle2_widths[674]), .RECT2_HEIGHT(rectangle2_heights[674]), .RECT2_WEIGHT(rectangle2_weights[674]), .RECT3_X(rectangle3_xs[674]), .RECT3_Y(rectangle3_ys[674]), .RECT3_WIDTH(rectangle3_widths[674]), .RECT3_HEIGHT(rectangle3_heights[674]), .RECT3_WEIGHT(rectangle3_weights[674]), .FEAT_THRES(feature_thresholds[674]), .FEAT_ABOVE(feature_aboves[674]), .FEAT_BELOW(feature_belows[674])) ac674(.scan_win(scan_win674), .scan_win_std_dev(scan_win_std_dev[674]), .feature_accum(feature_accums[674]));
  accum_calculator #(.RECT1_X(rectangle1_xs[675]), .RECT1_Y(rectangle1_ys[675]), .RECT1_WIDTH(rectangle1_widths[675]), .RECT1_HEIGHT(rectangle1_heights[675]), .RECT1_WEIGHT(rectangle1_weights[675]), .RECT2_X(rectangle2_xs[675]), .RECT2_Y(rectangle2_ys[675]), .RECT2_WIDTH(rectangle2_widths[675]), .RECT2_HEIGHT(rectangle2_heights[675]), .RECT2_WEIGHT(rectangle2_weights[675]), .RECT3_X(rectangle3_xs[675]), .RECT3_Y(rectangle3_ys[675]), .RECT3_WIDTH(rectangle3_widths[675]), .RECT3_HEIGHT(rectangle3_heights[675]), .RECT3_WEIGHT(rectangle3_weights[675]), .FEAT_THRES(feature_thresholds[675]), .FEAT_ABOVE(feature_aboves[675]), .FEAT_BELOW(feature_belows[675])) ac675(.scan_win(scan_win675), .scan_win_std_dev(scan_win_std_dev[675]), .feature_accum(feature_accums[675]));
  accum_calculator #(.RECT1_X(rectangle1_xs[676]), .RECT1_Y(rectangle1_ys[676]), .RECT1_WIDTH(rectangle1_widths[676]), .RECT1_HEIGHT(rectangle1_heights[676]), .RECT1_WEIGHT(rectangle1_weights[676]), .RECT2_X(rectangle2_xs[676]), .RECT2_Y(rectangle2_ys[676]), .RECT2_WIDTH(rectangle2_widths[676]), .RECT2_HEIGHT(rectangle2_heights[676]), .RECT2_WEIGHT(rectangle2_weights[676]), .RECT3_X(rectangle3_xs[676]), .RECT3_Y(rectangle3_ys[676]), .RECT3_WIDTH(rectangle3_widths[676]), .RECT3_HEIGHT(rectangle3_heights[676]), .RECT3_WEIGHT(rectangle3_weights[676]), .FEAT_THRES(feature_thresholds[676]), .FEAT_ABOVE(feature_aboves[676]), .FEAT_BELOW(feature_belows[676])) ac676(.scan_win(scan_win676), .scan_win_std_dev(scan_win_std_dev[676]), .feature_accum(feature_accums[676]));
  accum_calculator #(.RECT1_X(rectangle1_xs[677]), .RECT1_Y(rectangle1_ys[677]), .RECT1_WIDTH(rectangle1_widths[677]), .RECT1_HEIGHT(rectangle1_heights[677]), .RECT1_WEIGHT(rectangle1_weights[677]), .RECT2_X(rectangle2_xs[677]), .RECT2_Y(rectangle2_ys[677]), .RECT2_WIDTH(rectangle2_widths[677]), .RECT2_HEIGHT(rectangle2_heights[677]), .RECT2_WEIGHT(rectangle2_weights[677]), .RECT3_X(rectangle3_xs[677]), .RECT3_Y(rectangle3_ys[677]), .RECT3_WIDTH(rectangle3_widths[677]), .RECT3_HEIGHT(rectangle3_heights[677]), .RECT3_WEIGHT(rectangle3_weights[677]), .FEAT_THRES(feature_thresholds[677]), .FEAT_ABOVE(feature_aboves[677]), .FEAT_BELOW(feature_belows[677])) ac677(.scan_win(scan_win677), .scan_win_std_dev(scan_win_std_dev[677]), .feature_accum(feature_accums[677]));
  accum_calculator #(.RECT1_X(rectangle1_xs[678]), .RECT1_Y(rectangle1_ys[678]), .RECT1_WIDTH(rectangle1_widths[678]), .RECT1_HEIGHT(rectangle1_heights[678]), .RECT1_WEIGHT(rectangle1_weights[678]), .RECT2_X(rectangle2_xs[678]), .RECT2_Y(rectangle2_ys[678]), .RECT2_WIDTH(rectangle2_widths[678]), .RECT2_HEIGHT(rectangle2_heights[678]), .RECT2_WEIGHT(rectangle2_weights[678]), .RECT3_X(rectangle3_xs[678]), .RECT3_Y(rectangle3_ys[678]), .RECT3_WIDTH(rectangle3_widths[678]), .RECT3_HEIGHT(rectangle3_heights[678]), .RECT3_WEIGHT(rectangle3_weights[678]), .FEAT_THRES(feature_thresholds[678]), .FEAT_ABOVE(feature_aboves[678]), .FEAT_BELOW(feature_belows[678])) ac678(.scan_win(scan_win678), .scan_win_std_dev(scan_win_std_dev[678]), .feature_accum(feature_accums[678]));
  accum_calculator #(.RECT1_X(rectangle1_xs[679]), .RECT1_Y(rectangle1_ys[679]), .RECT1_WIDTH(rectangle1_widths[679]), .RECT1_HEIGHT(rectangle1_heights[679]), .RECT1_WEIGHT(rectangle1_weights[679]), .RECT2_X(rectangle2_xs[679]), .RECT2_Y(rectangle2_ys[679]), .RECT2_WIDTH(rectangle2_widths[679]), .RECT2_HEIGHT(rectangle2_heights[679]), .RECT2_WEIGHT(rectangle2_weights[679]), .RECT3_X(rectangle3_xs[679]), .RECT3_Y(rectangle3_ys[679]), .RECT3_WIDTH(rectangle3_widths[679]), .RECT3_HEIGHT(rectangle3_heights[679]), .RECT3_WEIGHT(rectangle3_weights[679]), .FEAT_THRES(feature_thresholds[679]), .FEAT_ABOVE(feature_aboves[679]), .FEAT_BELOW(feature_belows[679])) ac679(.scan_win(scan_win679), .scan_win_std_dev(scan_win_std_dev[679]), .feature_accum(feature_accums[679]));
  accum_calculator #(.RECT1_X(rectangle1_xs[680]), .RECT1_Y(rectangle1_ys[680]), .RECT1_WIDTH(rectangle1_widths[680]), .RECT1_HEIGHT(rectangle1_heights[680]), .RECT1_WEIGHT(rectangle1_weights[680]), .RECT2_X(rectangle2_xs[680]), .RECT2_Y(rectangle2_ys[680]), .RECT2_WIDTH(rectangle2_widths[680]), .RECT2_HEIGHT(rectangle2_heights[680]), .RECT2_WEIGHT(rectangle2_weights[680]), .RECT3_X(rectangle3_xs[680]), .RECT3_Y(rectangle3_ys[680]), .RECT3_WIDTH(rectangle3_widths[680]), .RECT3_HEIGHT(rectangle3_heights[680]), .RECT3_WEIGHT(rectangle3_weights[680]), .FEAT_THRES(feature_thresholds[680]), .FEAT_ABOVE(feature_aboves[680]), .FEAT_BELOW(feature_belows[680])) ac680(.scan_win(scan_win680), .scan_win_std_dev(scan_win_std_dev[680]), .feature_accum(feature_accums[680]));
  accum_calculator #(.RECT1_X(rectangle1_xs[681]), .RECT1_Y(rectangle1_ys[681]), .RECT1_WIDTH(rectangle1_widths[681]), .RECT1_HEIGHT(rectangle1_heights[681]), .RECT1_WEIGHT(rectangle1_weights[681]), .RECT2_X(rectangle2_xs[681]), .RECT2_Y(rectangle2_ys[681]), .RECT2_WIDTH(rectangle2_widths[681]), .RECT2_HEIGHT(rectangle2_heights[681]), .RECT2_WEIGHT(rectangle2_weights[681]), .RECT3_X(rectangle3_xs[681]), .RECT3_Y(rectangle3_ys[681]), .RECT3_WIDTH(rectangle3_widths[681]), .RECT3_HEIGHT(rectangle3_heights[681]), .RECT3_WEIGHT(rectangle3_weights[681]), .FEAT_THRES(feature_thresholds[681]), .FEAT_ABOVE(feature_aboves[681]), .FEAT_BELOW(feature_belows[681])) ac681(.scan_win(scan_win681), .scan_win_std_dev(scan_win_std_dev[681]), .feature_accum(feature_accums[681]));
  accum_calculator #(.RECT1_X(rectangle1_xs[682]), .RECT1_Y(rectangle1_ys[682]), .RECT1_WIDTH(rectangle1_widths[682]), .RECT1_HEIGHT(rectangle1_heights[682]), .RECT1_WEIGHT(rectangle1_weights[682]), .RECT2_X(rectangle2_xs[682]), .RECT2_Y(rectangle2_ys[682]), .RECT2_WIDTH(rectangle2_widths[682]), .RECT2_HEIGHT(rectangle2_heights[682]), .RECT2_WEIGHT(rectangle2_weights[682]), .RECT3_X(rectangle3_xs[682]), .RECT3_Y(rectangle3_ys[682]), .RECT3_WIDTH(rectangle3_widths[682]), .RECT3_HEIGHT(rectangle3_heights[682]), .RECT3_WEIGHT(rectangle3_weights[682]), .FEAT_THRES(feature_thresholds[682]), .FEAT_ABOVE(feature_aboves[682]), .FEAT_BELOW(feature_belows[682])) ac682(.scan_win(scan_win682), .scan_win_std_dev(scan_win_std_dev[682]), .feature_accum(feature_accums[682]));
  accum_calculator #(.RECT1_X(rectangle1_xs[683]), .RECT1_Y(rectangle1_ys[683]), .RECT1_WIDTH(rectangle1_widths[683]), .RECT1_HEIGHT(rectangle1_heights[683]), .RECT1_WEIGHT(rectangle1_weights[683]), .RECT2_X(rectangle2_xs[683]), .RECT2_Y(rectangle2_ys[683]), .RECT2_WIDTH(rectangle2_widths[683]), .RECT2_HEIGHT(rectangle2_heights[683]), .RECT2_WEIGHT(rectangle2_weights[683]), .RECT3_X(rectangle3_xs[683]), .RECT3_Y(rectangle3_ys[683]), .RECT3_WIDTH(rectangle3_widths[683]), .RECT3_HEIGHT(rectangle3_heights[683]), .RECT3_WEIGHT(rectangle3_weights[683]), .FEAT_THRES(feature_thresholds[683]), .FEAT_ABOVE(feature_aboves[683]), .FEAT_BELOW(feature_belows[683])) ac683(.scan_win(scan_win683), .scan_win_std_dev(scan_win_std_dev[683]), .feature_accum(feature_accums[683]));
  accum_calculator #(.RECT1_X(rectangle1_xs[684]), .RECT1_Y(rectangle1_ys[684]), .RECT1_WIDTH(rectangle1_widths[684]), .RECT1_HEIGHT(rectangle1_heights[684]), .RECT1_WEIGHT(rectangle1_weights[684]), .RECT2_X(rectangle2_xs[684]), .RECT2_Y(rectangle2_ys[684]), .RECT2_WIDTH(rectangle2_widths[684]), .RECT2_HEIGHT(rectangle2_heights[684]), .RECT2_WEIGHT(rectangle2_weights[684]), .RECT3_X(rectangle3_xs[684]), .RECT3_Y(rectangle3_ys[684]), .RECT3_WIDTH(rectangle3_widths[684]), .RECT3_HEIGHT(rectangle3_heights[684]), .RECT3_WEIGHT(rectangle3_weights[684]), .FEAT_THRES(feature_thresholds[684]), .FEAT_ABOVE(feature_aboves[684]), .FEAT_BELOW(feature_belows[684])) ac684(.scan_win(scan_win684), .scan_win_std_dev(scan_win_std_dev[684]), .feature_accum(feature_accums[684]));
  accum_calculator #(.RECT1_X(rectangle1_xs[685]), .RECT1_Y(rectangle1_ys[685]), .RECT1_WIDTH(rectangle1_widths[685]), .RECT1_HEIGHT(rectangle1_heights[685]), .RECT1_WEIGHT(rectangle1_weights[685]), .RECT2_X(rectangle2_xs[685]), .RECT2_Y(rectangle2_ys[685]), .RECT2_WIDTH(rectangle2_widths[685]), .RECT2_HEIGHT(rectangle2_heights[685]), .RECT2_WEIGHT(rectangle2_weights[685]), .RECT3_X(rectangle3_xs[685]), .RECT3_Y(rectangle3_ys[685]), .RECT3_WIDTH(rectangle3_widths[685]), .RECT3_HEIGHT(rectangle3_heights[685]), .RECT3_WEIGHT(rectangle3_weights[685]), .FEAT_THRES(feature_thresholds[685]), .FEAT_ABOVE(feature_aboves[685]), .FEAT_BELOW(feature_belows[685])) ac685(.scan_win(scan_win685), .scan_win_std_dev(scan_win_std_dev[685]), .feature_accum(feature_accums[685]));
  accum_calculator #(.RECT1_X(rectangle1_xs[686]), .RECT1_Y(rectangle1_ys[686]), .RECT1_WIDTH(rectangle1_widths[686]), .RECT1_HEIGHT(rectangle1_heights[686]), .RECT1_WEIGHT(rectangle1_weights[686]), .RECT2_X(rectangle2_xs[686]), .RECT2_Y(rectangle2_ys[686]), .RECT2_WIDTH(rectangle2_widths[686]), .RECT2_HEIGHT(rectangle2_heights[686]), .RECT2_WEIGHT(rectangle2_weights[686]), .RECT3_X(rectangle3_xs[686]), .RECT3_Y(rectangle3_ys[686]), .RECT3_WIDTH(rectangle3_widths[686]), .RECT3_HEIGHT(rectangle3_heights[686]), .RECT3_WEIGHT(rectangle3_weights[686]), .FEAT_THRES(feature_thresholds[686]), .FEAT_ABOVE(feature_aboves[686]), .FEAT_BELOW(feature_belows[686])) ac686(.scan_win(scan_win686), .scan_win_std_dev(scan_win_std_dev[686]), .feature_accum(feature_accums[686]));
  accum_calculator #(.RECT1_X(rectangle1_xs[687]), .RECT1_Y(rectangle1_ys[687]), .RECT1_WIDTH(rectangle1_widths[687]), .RECT1_HEIGHT(rectangle1_heights[687]), .RECT1_WEIGHT(rectangle1_weights[687]), .RECT2_X(rectangle2_xs[687]), .RECT2_Y(rectangle2_ys[687]), .RECT2_WIDTH(rectangle2_widths[687]), .RECT2_HEIGHT(rectangle2_heights[687]), .RECT2_WEIGHT(rectangle2_weights[687]), .RECT3_X(rectangle3_xs[687]), .RECT3_Y(rectangle3_ys[687]), .RECT3_WIDTH(rectangle3_widths[687]), .RECT3_HEIGHT(rectangle3_heights[687]), .RECT3_WEIGHT(rectangle3_weights[687]), .FEAT_THRES(feature_thresholds[687]), .FEAT_ABOVE(feature_aboves[687]), .FEAT_BELOW(feature_belows[687])) ac687(.scan_win(scan_win687), .scan_win_std_dev(scan_win_std_dev[687]), .feature_accum(feature_accums[687]));
  accum_calculator #(.RECT1_X(rectangle1_xs[688]), .RECT1_Y(rectangle1_ys[688]), .RECT1_WIDTH(rectangle1_widths[688]), .RECT1_HEIGHT(rectangle1_heights[688]), .RECT1_WEIGHT(rectangle1_weights[688]), .RECT2_X(rectangle2_xs[688]), .RECT2_Y(rectangle2_ys[688]), .RECT2_WIDTH(rectangle2_widths[688]), .RECT2_HEIGHT(rectangle2_heights[688]), .RECT2_WEIGHT(rectangle2_weights[688]), .RECT3_X(rectangle3_xs[688]), .RECT3_Y(rectangle3_ys[688]), .RECT3_WIDTH(rectangle3_widths[688]), .RECT3_HEIGHT(rectangle3_heights[688]), .RECT3_WEIGHT(rectangle3_weights[688]), .FEAT_THRES(feature_thresholds[688]), .FEAT_ABOVE(feature_aboves[688]), .FEAT_BELOW(feature_belows[688])) ac688(.scan_win(scan_win688), .scan_win_std_dev(scan_win_std_dev[688]), .feature_accum(feature_accums[688]));
  accum_calculator #(.RECT1_X(rectangle1_xs[689]), .RECT1_Y(rectangle1_ys[689]), .RECT1_WIDTH(rectangle1_widths[689]), .RECT1_HEIGHT(rectangle1_heights[689]), .RECT1_WEIGHT(rectangle1_weights[689]), .RECT2_X(rectangle2_xs[689]), .RECT2_Y(rectangle2_ys[689]), .RECT2_WIDTH(rectangle2_widths[689]), .RECT2_HEIGHT(rectangle2_heights[689]), .RECT2_WEIGHT(rectangle2_weights[689]), .RECT3_X(rectangle3_xs[689]), .RECT3_Y(rectangle3_ys[689]), .RECT3_WIDTH(rectangle3_widths[689]), .RECT3_HEIGHT(rectangle3_heights[689]), .RECT3_WEIGHT(rectangle3_weights[689]), .FEAT_THRES(feature_thresholds[689]), .FEAT_ABOVE(feature_aboves[689]), .FEAT_BELOW(feature_belows[689])) ac689(.scan_win(scan_win689), .scan_win_std_dev(scan_win_std_dev[689]), .feature_accum(feature_accums[689]));
  accum_calculator #(.RECT1_X(rectangle1_xs[690]), .RECT1_Y(rectangle1_ys[690]), .RECT1_WIDTH(rectangle1_widths[690]), .RECT1_HEIGHT(rectangle1_heights[690]), .RECT1_WEIGHT(rectangle1_weights[690]), .RECT2_X(rectangle2_xs[690]), .RECT2_Y(rectangle2_ys[690]), .RECT2_WIDTH(rectangle2_widths[690]), .RECT2_HEIGHT(rectangle2_heights[690]), .RECT2_WEIGHT(rectangle2_weights[690]), .RECT3_X(rectangle3_xs[690]), .RECT3_Y(rectangle3_ys[690]), .RECT3_WIDTH(rectangle3_widths[690]), .RECT3_HEIGHT(rectangle3_heights[690]), .RECT3_WEIGHT(rectangle3_weights[690]), .FEAT_THRES(feature_thresholds[690]), .FEAT_ABOVE(feature_aboves[690]), .FEAT_BELOW(feature_belows[690])) ac690(.scan_win(scan_win690), .scan_win_std_dev(scan_win_std_dev[690]), .feature_accum(feature_accums[690]));
  accum_calculator #(.RECT1_X(rectangle1_xs[691]), .RECT1_Y(rectangle1_ys[691]), .RECT1_WIDTH(rectangle1_widths[691]), .RECT1_HEIGHT(rectangle1_heights[691]), .RECT1_WEIGHT(rectangle1_weights[691]), .RECT2_X(rectangle2_xs[691]), .RECT2_Y(rectangle2_ys[691]), .RECT2_WIDTH(rectangle2_widths[691]), .RECT2_HEIGHT(rectangle2_heights[691]), .RECT2_WEIGHT(rectangle2_weights[691]), .RECT3_X(rectangle3_xs[691]), .RECT3_Y(rectangle3_ys[691]), .RECT3_WIDTH(rectangle3_widths[691]), .RECT3_HEIGHT(rectangle3_heights[691]), .RECT3_WEIGHT(rectangle3_weights[691]), .FEAT_THRES(feature_thresholds[691]), .FEAT_ABOVE(feature_aboves[691]), .FEAT_BELOW(feature_belows[691])) ac691(.scan_win(scan_win691), .scan_win_std_dev(scan_win_std_dev[691]), .feature_accum(feature_accums[691]));
  accum_calculator #(.RECT1_X(rectangle1_xs[692]), .RECT1_Y(rectangle1_ys[692]), .RECT1_WIDTH(rectangle1_widths[692]), .RECT1_HEIGHT(rectangle1_heights[692]), .RECT1_WEIGHT(rectangle1_weights[692]), .RECT2_X(rectangle2_xs[692]), .RECT2_Y(rectangle2_ys[692]), .RECT2_WIDTH(rectangle2_widths[692]), .RECT2_HEIGHT(rectangle2_heights[692]), .RECT2_WEIGHT(rectangle2_weights[692]), .RECT3_X(rectangle3_xs[692]), .RECT3_Y(rectangle3_ys[692]), .RECT3_WIDTH(rectangle3_widths[692]), .RECT3_HEIGHT(rectangle3_heights[692]), .RECT3_WEIGHT(rectangle3_weights[692]), .FEAT_THRES(feature_thresholds[692]), .FEAT_ABOVE(feature_aboves[692]), .FEAT_BELOW(feature_belows[692])) ac692(.scan_win(scan_win692), .scan_win_std_dev(scan_win_std_dev[692]), .feature_accum(feature_accums[692]));
  accum_calculator #(.RECT1_X(rectangle1_xs[693]), .RECT1_Y(rectangle1_ys[693]), .RECT1_WIDTH(rectangle1_widths[693]), .RECT1_HEIGHT(rectangle1_heights[693]), .RECT1_WEIGHT(rectangle1_weights[693]), .RECT2_X(rectangle2_xs[693]), .RECT2_Y(rectangle2_ys[693]), .RECT2_WIDTH(rectangle2_widths[693]), .RECT2_HEIGHT(rectangle2_heights[693]), .RECT2_WEIGHT(rectangle2_weights[693]), .RECT3_X(rectangle3_xs[693]), .RECT3_Y(rectangle3_ys[693]), .RECT3_WIDTH(rectangle3_widths[693]), .RECT3_HEIGHT(rectangle3_heights[693]), .RECT3_WEIGHT(rectangle3_weights[693]), .FEAT_THRES(feature_thresholds[693]), .FEAT_ABOVE(feature_aboves[693]), .FEAT_BELOW(feature_belows[693])) ac693(.scan_win(scan_win693), .scan_win_std_dev(scan_win_std_dev[693]), .feature_accum(feature_accums[693]));
  accum_calculator #(.RECT1_X(rectangle1_xs[694]), .RECT1_Y(rectangle1_ys[694]), .RECT1_WIDTH(rectangle1_widths[694]), .RECT1_HEIGHT(rectangle1_heights[694]), .RECT1_WEIGHT(rectangle1_weights[694]), .RECT2_X(rectangle2_xs[694]), .RECT2_Y(rectangle2_ys[694]), .RECT2_WIDTH(rectangle2_widths[694]), .RECT2_HEIGHT(rectangle2_heights[694]), .RECT2_WEIGHT(rectangle2_weights[694]), .RECT3_X(rectangle3_xs[694]), .RECT3_Y(rectangle3_ys[694]), .RECT3_WIDTH(rectangle3_widths[694]), .RECT3_HEIGHT(rectangle3_heights[694]), .RECT3_WEIGHT(rectangle3_weights[694]), .FEAT_THRES(feature_thresholds[694]), .FEAT_ABOVE(feature_aboves[694]), .FEAT_BELOW(feature_belows[694])) ac694(.scan_win(scan_win694), .scan_win_std_dev(scan_win_std_dev[694]), .feature_accum(feature_accums[694]));
  accum_calculator #(.RECT1_X(rectangle1_xs[695]), .RECT1_Y(rectangle1_ys[695]), .RECT1_WIDTH(rectangle1_widths[695]), .RECT1_HEIGHT(rectangle1_heights[695]), .RECT1_WEIGHT(rectangle1_weights[695]), .RECT2_X(rectangle2_xs[695]), .RECT2_Y(rectangle2_ys[695]), .RECT2_WIDTH(rectangle2_widths[695]), .RECT2_HEIGHT(rectangle2_heights[695]), .RECT2_WEIGHT(rectangle2_weights[695]), .RECT3_X(rectangle3_xs[695]), .RECT3_Y(rectangle3_ys[695]), .RECT3_WIDTH(rectangle3_widths[695]), .RECT3_HEIGHT(rectangle3_heights[695]), .RECT3_WEIGHT(rectangle3_weights[695]), .FEAT_THRES(feature_thresholds[695]), .FEAT_ABOVE(feature_aboves[695]), .FEAT_BELOW(feature_belows[695])) ac695(.scan_win(scan_win695), .scan_win_std_dev(scan_win_std_dev[695]), .feature_accum(feature_accums[695]));
  accum_calculator #(.RECT1_X(rectangle1_xs[696]), .RECT1_Y(rectangle1_ys[696]), .RECT1_WIDTH(rectangle1_widths[696]), .RECT1_HEIGHT(rectangle1_heights[696]), .RECT1_WEIGHT(rectangle1_weights[696]), .RECT2_X(rectangle2_xs[696]), .RECT2_Y(rectangle2_ys[696]), .RECT2_WIDTH(rectangle2_widths[696]), .RECT2_HEIGHT(rectangle2_heights[696]), .RECT2_WEIGHT(rectangle2_weights[696]), .RECT3_X(rectangle3_xs[696]), .RECT3_Y(rectangle3_ys[696]), .RECT3_WIDTH(rectangle3_widths[696]), .RECT3_HEIGHT(rectangle3_heights[696]), .RECT3_WEIGHT(rectangle3_weights[696]), .FEAT_THRES(feature_thresholds[696]), .FEAT_ABOVE(feature_aboves[696]), .FEAT_BELOW(feature_belows[696])) ac696(.scan_win(scan_win696), .scan_win_std_dev(scan_win_std_dev[696]), .feature_accum(feature_accums[696]));
  accum_calculator #(.RECT1_X(rectangle1_xs[697]), .RECT1_Y(rectangle1_ys[697]), .RECT1_WIDTH(rectangle1_widths[697]), .RECT1_HEIGHT(rectangle1_heights[697]), .RECT1_WEIGHT(rectangle1_weights[697]), .RECT2_X(rectangle2_xs[697]), .RECT2_Y(rectangle2_ys[697]), .RECT2_WIDTH(rectangle2_widths[697]), .RECT2_HEIGHT(rectangle2_heights[697]), .RECT2_WEIGHT(rectangle2_weights[697]), .RECT3_X(rectangle3_xs[697]), .RECT3_Y(rectangle3_ys[697]), .RECT3_WIDTH(rectangle3_widths[697]), .RECT3_HEIGHT(rectangle3_heights[697]), .RECT3_WEIGHT(rectangle3_weights[697]), .FEAT_THRES(feature_thresholds[697]), .FEAT_ABOVE(feature_aboves[697]), .FEAT_BELOW(feature_belows[697])) ac697(.scan_win(scan_win697), .scan_win_std_dev(scan_win_std_dev[697]), .feature_accum(feature_accums[697]));
  accum_calculator #(.RECT1_X(rectangle1_xs[698]), .RECT1_Y(rectangle1_ys[698]), .RECT1_WIDTH(rectangle1_widths[698]), .RECT1_HEIGHT(rectangle1_heights[698]), .RECT1_WEIGHT(rectangle1_weights[698]), .RECT2_X(rectangle2_xs[698]), .RECT2_Y(rectangle2_ys[698]), .RECT2_WIDTH(rectangle2_widths[698]), .RECT2_HEIGHT(rectangle2_heights[698]), .RECT2_WEIGHT(rectangle2_weights[698]), .RECT3_X(rectangle3_xs[698]), .RECT3_Y(rectangle3_ys[698]), .RECT3_WIDTH(rectangle3_widths[698]), .RECT3_HEIGHT(rectangle3_heights[698]), .RECT3_WEIGHT(rectangle3_weights[698]), .FEAT_THRES(feature_thresholds[698]), .FEAT_ABOVE(feature_aboves[698]), .FEAT_BELOW(feature_belows[698])) ac698(.scan_win(scan_win698), .scan_win_std_dev(scan_win_std_dev[698]), .feature_accum(feature_accums[698]));
  accum_calculator #(.RECT1_X(rectangle1_xs[699]), .RECT1_Y(rectangle1_ys[699]), .RECT1_WIDTH(rectangle1_widths[699]), .RECT1_HEIGHT(rectangle1_heights[699]), .RECT1_WEIGHT(rectangle1_weights[699]), .RECT2_X(rectangle2_xs[699]), .RECT2_Y(rectangle2_ys[699]), .RECT2_WIDTH(rectangle2_widths[699]), .RECT2_HEIGHT(rectangle2_heights[699]), .RECT2_WEIGHT(rectangle2_weights[699]), .RECT3_X(rectangle3_xs[699]), .RECT3_Y(rectangle3_ys[699]), .RECT3_WIDTH(rectangle3_widths[699]), .RECT3_HEIGHT(rectangle3_heights[699]), .RECT3_WEIGHT(rectangle3_weights[699]), .FEAT_THRES(feature_thresholds[699]), .FEAT_ABOVE(feature_aboves[699]), .FEAT_BELOW(feature_belows[699])) ac699(.scan_win(scan_win699), .scan_win_std_dev(scan_win_std_dev[699]), .feature_accum(feature_accums[699]));
  accum_calculator #(.RECT1_X(rectangle1_xs[700]), .RECT1_Y(rectangle1_ys[700]), .RECT1_WIDTH(rectangle1_widths[700]), .RECT1_HEIGHT(rectangle1_heights[700]), .RECT1_WEIGHT(rectangle1_weights[700]), .RECT2_X(rectangle2_xs[700]), .RECT2_Y(rectangle2_ys[700]), .RECT2_WIDTH(rectangle2_widths[700]), .RECT2_HEIGHT(rectangle2_heights[700]), .RECT2_WEIGHT(rectangle2_weights[700]), .RECT3_X(rectangle3_xs[700]), .RECT3_Y(rectangle3_ys[700]), .RECT3_WIDTH(rectangle3_widths[700]), .RECT3_HEIGHT(rectangle3_heights[700]), .RECT3_WEIGHT(rectangle3_weights[700]), .FEAT_THRES(feature_thresholds[700]), .FEAT_ABOVE(feature_aboves[700]), .FEAT_BELOW(feature_belows[700])) ac700(.scan_win(scan_win700), .scan_win_std_dev(scan_win_std_dev[700]), .feature_accum(feature_accums[700]));
  accum_calculator #(.RECT1_X(rectangle1_xs[701]), .RECT1_Y(rectangle1_ys[701]), .RECT1_WIDTH(rectangle1_widths[701]), .RECT1_HEIGHT(rectangle1_heights[701]), .RECT1_WEIGHT(rectangle1_weights[701]), .RECT2_X(rectangle2_xs[701]), .RECT2_Y(rectangle2_ys[701]), .RECT2_WIDTH(rectangle2_widths[701]), .RECT2_HEIGHT(rectangle2_heights[701]), .RECT2_WEIGHT(rectangle2_weights[701]), .RECT3_X(rectangle3_xs[701]), .RECT3_Y(rectangle3_ys[701]), .RECT3_WIDTH(rectangle3_widths[701]), .RECT3_HEIGHT(rectangle3_heights[701]), .RECT3_WEIGHT(rectangle3_weights[701]), .FEAT_THRES(feature_thresholds[701]), .FEAT_ABOVE(feature_aboves[701]), .FEAT_BELOW(feature_belows[701])) ac701(.scan_win(scan_win701), .scan_win_std_dev(scan_win_std_dev[701]), .feature_accum(feature_accums[701]));
  accum_calculator #(.RECT1_X(rectangle1_xs[702]), .RECT1_Y(rectangle1_ys[702]), .RECT1_WIDTH(rectangle1_widths[702]), .RECT1_HEIGHT(rectangle1_heights[702]), .RECT1_WEIGHT(rectangle1_weights[702]), .RECT2_X(rectangle2_xs[702]), .RECT2_Y(rectangle2_ys[702]), .RECT2_WIDTH(rectangle2_widths[702]), .RECT2_HEIGHT(rectangle2_heights[702]), .RECT2_WEIGHT(rectangle2_weights[702]), .RECT3_X(rectangle3_xs[702]), .RECT3_Y(rectangle3_ys[702]), .RECT3_WIDTH(rectangle3_widths[702]), .RECT3_HEIGHT(rectangle3_heights[702]), .RECT3_WEIGHT(rectangle3_weights[702]), .FEAT_THRES(feature_thresholds[702]), .FEAT_ABOVE(feature_aboves[702]), .FEAT_BELOW(feature_belows[702])) ac702(.scan_win(scan_win702), .scan_win_std_dev(scan_win_std_dev[702]), .feature_accum(feature_accums[702]));
  accum_calculator #(.RECT1_X(rectangle1_xs[703]), .RECT1_Y(rectangle1_ys[703]), .RECT1_WIDTH(rectangle1_widths[703]), .RECT1_HEIGHT(rectangle1_heights[703]), .RECT1_WEIGHT(rectangle1_weights[703]), .RECT2_X(rectangle2_xs[703]), .RECT2_Y(rectangle2_ys[703]), .RECT2_WIDTH(rectangle2_widths[703]), .RECT2_HEIGHT(rectangle2_heights[703]), .RECT2_WEIGHT(rectangle2_weights[703]), .RECT3_X(rectangle3_xs[703]), .RECT3_Y(rectangle3_ys[703]), .RECT3_WIDTH(rectangle3_widths[703]), .RECT3_HEIGHT(rectangle3_heights[703]), .RECT3_WEIGHT(rectangle3_weights[703]), .FEAT_THRES(feature_thresholds[703]), .FEAT_ABOVE(feature_aboves[703]), .FEAT_BELOW(feature_belows[703])) ac703(.scan_win(scan_win703), .scan_win_std_dev(scan_win_std_dev[703]), .feature_accum(feature_accums[703]));
  accum_calculator #(.RECT1_X(rectangle1_xs[704]), .RECT1_Y(rectangle1_ys[704]), .RECT1_WIDTH(rectangle1_widths[704]), .RECT1_HEIGHT(rectangle1_heights[704]), .RECT1_WEIGHT(rectangle1_weights[704]), .RECT2_X(rectangle2_xs[704]), .RECT2_Y(rectangle2_ys[704]), .RECT2_WIDTH(rectangle2_widths[704]), .RECT2_HEIGHT(rectangle2_heights[704]), .RECT2_WEIGHT(rectangle2_weights[704]), .RECT3_X(rectangle3_xs[704]), .RECT3_Y(rectangle3_ys[704]), .RECT3_WIDTH(rectangle3_widths[704]), .RECT3_HEIGHT(rectangle3_heights[704]), .RECT3_WEIGHT(rectangle3_weights[704]), .FEAT_THRES(feature_thresholds[704]), .FEAT_ABOVE(feature_aboves[704]), .FEAT_BELOW(feature_belows[704])) ac704(.scan_win(scan_win704), .scan_win_std_dev(scan_win_std_dev[704]), .feature_accum(feature_accums[704]));
  accum_calculator #(.RECT1_X(rectangle1_xs[705]), .RECT1_Y(rectangle1_ys[705]), .RECT1_WIDTH(rectangle1_widths[705]), .RECT1_HEIGHT(rectangle1_heights[705]), .RECT1_WEIGHT(rectangle1_weights[705]), .RECT2_X(rectangle2_xs[705]), .RECT2_Y(rectangle2_ys[705]), .RECT2_WIDTH(rectangle2_widths[705]), .RECT2_HEIGHT(rectangle2_heights[705]), .RECT2_WEIGHT(rectangle2_weights[705]), .RECT3_X(rectangle3_xs[705]), .RECT3_Y(rectangle3_ys[705]), .RECT3_WIDTH(rectangle3_widths[705]), .RECT3_HEIGHT(rectangle3_heights[705]), .RECT3_WEIGHT(rectangle3_weights[705]), .FEAT_THRES(feature_thresholds[705]), .FEAT_ABOVE(feature_aboves[705]), .FEAT_BELOW(feature_belows[705])) ac705(.scan_win(scan_win705), .scan_win_std_dev(scan_win_std_dev[705]), .feature_accum(feature_accums[705]));
  accum_calculator #(.RECT1_X(rectangle1_xs[706]), .RECT1_Y(rectangle1_ys[706]), .RECT1_WIDTH(rectangle1_widths[706]), .RECT1_HEIGHT(rectangle1_heights[706]), .RECT1_WEIGHT(rectangle1_weights[706]), .RECT2_X(rectangle2_xs[706]), .RECT2_Y(rectangle2_ys[706]), .RECT2_WIDTH(rectangle2_widths[706]), .RECT2_HEIGHT(rectangle2_heights[706]), .RECT2_WEIGHT(rectangle2_weights[706]), .RECT3_X(rectangle3_xs[706]), .RECT3_Y(rectangle3_ys[706]), .RECT3_WIDTH(rectangle3_widths[706]), .RECT3_HEIGHT(rectangle3_heights[706]), .RECT3_WEIGHT(rectangle3_weights[706]), .FEAT_THRES(feature_thresholds[706]), .FEAT_ABOVE(feature_aboves[706]), .FEAT_BELOW(feature_belows[706])) ac706(.scan_win(scan_win706), .scan_win_std_dev(scan_win_std_dev[706]), .feature_accum(feature_accums[706]));
  accum_calculator #(.RECT1_X(rectangle1_xs[707]), .RECT1_Y(rectangle1_ys[707]), .RECT1_WIDTH(rectangle1_widths[707]), .RECT1_HEIGHT(rectangle1_heights[707]), .RECT1_WEIGHT(rectangle1_weights[707]), .RECT2_X(rectangle2_xs[707]), .RECT2_Y(rectangle2_ys[707]), .RECT2_WIDTH(rectangle2_widths[707]), .RECT2_HEIGHT(rectangle2_heights[707]), .RECT2_WEIGHT(rectangle2_weights[707]), .RECT3_X(rectangle3_xs[707]), .RECT3_Y(rectangle3_ys[707]), .RECT3_WIDTH(rectangle3_widths[707]), .RECT3_HEIGHT(rectangle3_heights[707]), .RECT3_WEIGHT(rectangle3_weights[707]), .FEAT_THRES(feature_thresholds[707]), .FEAT_ABOVE(feature_aboves[707]), .FEAT_BELOW(feature_belows[707])) ac707(.scan_win(scan_win707), .scan_win_std_dev(scan_win_std_dev[707]), .feature_accum(feature_accums[707]));
  accum_calculator #(.RECT1_X(rectangle1_xs[708]), .RECT1_Y(rectangle1_ys[708]), .RECT1_WIDTH(rectangle1_widths[708]), .RECT1_HEIGHT(rectangle1_heights[708]), .RECT1_WEIGHT(rectangle1_weights[708]), .RECT2_X(rectangle2_xs[708]), .RECT2_Y(rectangle2_ys[708]), .RECT2_WIDTH(rectangle2_widths[708]), .RECT2_HEIGHT(rectangle2_heights[708]), .RECT2_WEIGHT(rectangle2_weights[708]), .RECT3_X(rectangle3_xs[708]), .RECT3_Y(rectangle3_ys[708]), .RECT3_WIDTH(rectangle3_widths[708]), .RECT3_HEIGHT(rectangle3_heights[708]), .RECT3_WEIGHT(rectangle3_weights[708]), .FEAT_THRES(feature_thresholds[708]), .FEAT_ABOVE(feature_aboves[708]), .FEAT_BELOW(feature_belows[708])) ac708(.scan_win(scan_win708), .scan_win_std_dev(scan_win_std_dev[708]), .feature_accum(feature_accums[708]));
  accum_calculator #(.RECT1_X(rectangle1_xs[709]), .RECT1_Y(rectangle1_ys[709]), .RECT1_WIDTH(rectangle1_widths[709]), .RECT1_HEIGHT(rectangle1_heights[709]), .RECT1_WEIGHT(rectangle1_weights[709]), .RECT2_X(rectangle2_xs[709]), .RECT2_Y(rectangle2_ys[709]), .RECT2_WIDTH(rectangle2_widths[709]), .RECT2_HEIGHT(rectangle2_heights[709]), .RECT2_WEIGHT(rectangle2_weights[709]), .RECT3_X(rectangle3_xs[709]), .RECT3_Y(rectangle3_ys[709]), .RECT3_WIDTH(rectangle3_widths[709]), .RECT3_HEIGHT(rectangle3_heights[709]), .RECT3_WEIGHT(rectangle3_weights[709]), .FEAT_THRES(feature_thresholds[709]), .FEAT_ABOVE(feature_aboves[709]), .FEAT_BELOW(feature_belows[709])) ac709(.scan_win(scan_win709), .scan_win_std_dev(scan_win_std_dev[709]), .feature_accum(feature_accums[709]));
  accum_calculator #(.RECT1_X(rectangle1_xs[710]), .RECT1_Y(rectangle1_ys[710]), .RECT1_WIDTH(rectangle1_widths[710]), .RECT1_HEIGHT(rectangle1_heights[710]), .RECT1_WEIGHT(rectangle1_weights[710]), .RECT2_X(rectangle2_xs[710]), .RECT2_Y(rectangle2_ys[710]), .RECT2_WIDTH(rectangle2_widths[710]), .RECT2_HEIGHT(rectangle2_heights[710]), .RECT2_WEIGHT(rectangle2_weights[710]), .RECT3_X(rectangle3_xs[710]), .RECT3_Y(rectangle3_ys[710]), .RECT3_WIDTH(rectangle3_widths[710]), .RECT3_HEIGHT(rectangle3_heights[710]), .RECT3_WEIGHT(rectangle3_weights[710]), .FEAT_THRES(feature_thresholds[710]), .FEAT_ABOVE(feature_aboves[710]), .FEAT_BELOW(feature_belows[710])) ac710(.scan_win(scan_win710), .scan_win_std_dev(scan_win_std_dev[710]), .feature_accum(feature_accums[710]));
  accum_calculator #(.RECT1_X(rectangle1_xs[711]), .RECT1_Y(rectangle1_ys[711]), .RECT1_WIDTH(rectangle1_widths[711]), .RECT1_HEIGHT(rectangle1_heights[711]), .RECT1_WEIGHT(rectangle1_weights[711]), .RECT2_X(rectangle2_xs[711]), .RECT2_Y(rectangle2_ys[711]), .RECT2_WIDTH(rectangle2_widths[711]), .RECT2_HEIGHT(rectangle2_heights[711]), .RECT2_WEIGHT(rectangle2_weights[711]), .RECT3_X(rectangle3_xs[711]), .RECT3_Y(rectangle3_ys[711]), .RECT3_WIDTH(rectangle3_widths[711]), .RECT3_HEIGHT(rectangle3_heights[711]), .RECT3_WEIGHT(rectangle3_weights[711]), .FEAT_THRES(feature_thresholds[711]), .FEAT_ABOVE(feature_aboves[711]), .FEAT_BELOW(feature_belows[711])) ac711(.scan_win(scan_win711), .scan_win_std_dev(scan_win_std_dev[711]), .feature_accum(feature_accums[711]));
  accum_calculator #(.RECT1_X(rectangle1_xs[712]), .RECT1_Y(rectangle1_ys[712]), .RECT1_WIDTH(rectangle1_widths[712]), .RECT1_HEIGHT(rectangle1_heights[712]), .RECT1_WEIGHT(rectangle1_weights[712]), .RECT2_X(rectangle2_xs[712]), .RECT2_Y(rectangle2_ys[712]), .RECT2_WIDTH(rectangle2_widths[712]), .RECT2_HEIGHT(rectangle2_heights[712]), .RECT2_WEIGHT(rectangle2_weights[712]), .RECT3_X(rectangle3_xs[712]), .RECT3_Y(rectangle3_ys[712]), .RECT3_WIDTH(rectangle3_widths[712]), .RECT3_HEIGHT(rectangle3_heights[712]), .RECT3_WEIGHT(rectangle3_weights[712]), .FEAT_THRES(feature_thresholds[712]), .FEAT_ABOVE(feature_aboves[712]), .FEAT_BELOW(feature_belows[712])) ac712(.scan_win(scan_win712), .scan_win_std_dev(scan_win_std_dev[712]), .feature_accum(feature_accums[712]));
  accum_calculator #(.RECT1_X(rectangle1_xs[713]), .RECT1_Y(rectangle1_ys[713]), .RECT1_WIDTH(rectangle1_widths[713]), .RECT1_HEIGHT(rectangle1_heights[713]), .RECT1_WEIGHT(rectangle1_weights[713]), .RECT2_X(rectangle2_xs[713]), .RECT2_Y(rectangle2_ys[713]), .RECT2_WIDTH(rectangle2_widths[713]), .RECT2_HEIGHT(rectangle2_heights[713]), .RECT2_WEIGHT(rectangle2_weights[713]), .RECT3_X(rectangle3_xs[713]), .RECT3_Y(rectangle3_ys[713]), .RECT3_WIDTH(rectangle3_widths[713]), .RECT3_HEIGHT(rectangle3_heights[713]), .RECT3_WEIGHT(rectangle3_weights[713]), .FEAT_THRES(feature_thresholds[713]), .FEAT_ABOVE(feature_aboves[713]), .FEAT_BELOW(feature_belows[713])) ac713(.scan_win(scan_win713), .scan_win_std_dev(scan_win_std_dev[713]), .feature_accum(feature_accums[713]));
  accum_calculator #(.RECT1_X(rectangle1_xs[714]), .RECT1_Y(rectangle1_ys[714]), .RECT1_WIDTH(rectangle1_widths[714]), .RECT1_HEIGHT(rectangle1_heights[714]), .RECT1_WEIGHT(rectangle1_weights[714]), .RECT2_X(rectangle2_xs[714]), .RECT2_Y(rectangle2_ys[714]), .RECT2_WIDTH(rectangle2_widths[714]), .RECT2_HEIGHT(rectangle2_heights[714]), .RECT2_WEIGHT(rectangle2_weights[714]), .RECT3_X(rectangle3_xs[714]), .RECT3_Y(rectangle3_ys[714]), .RECT3_WIDTH(rectangle3_widths[714]), .RECT3_HEIGHT(rectangle3_heights[714]), .RECT3_WEIGHT(rectangle3_weights[714]), .FEAT_THRES(feature_thresholds[714]), .FEAT_ABOVE(feature_aboves[714]), .FEAT_BELOW(feature_belows[714])) ac714(.scan_win(scan_win714), .scan_win_std_dev(scan_win_std_dev[714]), .feature_accum(feature_accums[714]));
  accum_calculator #(.RECT1_X(rectangle1_xs[715]), .RECT1_Y(rectangle1_ys[715]), .RECT1_WIDTH(rectangle1_widths[715]), .RECT1_HEIGHT(rectangle1_heights[715]), .RECT1_WEIGHT(rectangle1_weights[715]), .RECT2_X(rectangle2_xs[715]), .RECT2_Y(rectangle2_ys[715]), .RECT2_WIDTH(rectangle2_widths[715]), .RECT2_HEIGHT(rectangle2_heights[715]), .RECT2_WEIGHT(rectangle2_weights[715]), .RECT3_X(rectangle3_xs[715]), .RECT3_Y(rectangle3_ys[715]), .RECT3_WIDTH(rectangle3_widths[715]), .RECT3_HEIGHT(rectangle3_heights[715]), .RECT3_WEIGHT(rectangle3_weights[715]), .FEAT_THRES(feature_thresholds[715]), .FEAT_ABOVE(feature_aboves[715]), .FEAT_BELOW(feature_belows[715])) ac715(.scan_win(scan_win715), .scan_win_std_dev(scan_win_std_dev[715]), .feature_accum(feature_accums[715]));
  accum_calculator #(.RECT1_X(rectangle1_xs[716]), .RECT1_Y(rectangle1_ys[716]), .RECT1_WIDTH(rectangle1_widths[716]), .RECT1_HEIGHT(rectangle1_heights[716]), .RECT1_WEIGHT(rectangle1_weights[716]), .RECT2_X(rectangle2_xs[716]), .RECT2_Y(rectangle2_ys[716]), .RECT2_WIDTH(rectangle2_widths[716]), .RECT2_HEIGHT(rectangle2_heights[716]), .RECT2_WEIGHT(rectangle2_weights[716]), .RECT3_X(rectangle3_xs[716]), .RECT3_Y(rectangle3_ys[716]), .RECT3_WIDTH(rectangle3_widths[716]), .RECT3_HEIGHT(rectangle3_heights[716]), .RECT3_WEIGHT(rectangle3_weights[716]), .FEAT_THRES(feature_thresholds[716]), .FEAT_ABOVE(feature_aboves[716]), .FEAT_BELOW(feature_belows[716])) ac716(.scan_win(scan_win716), .scan_win_std_dev(scan_win_std_dev[716]), .feature_accum(feature_accums[716]));
  accum_calculator #(.RECT1_X(rectangle1_xs[717]), .RECT1_Y(rectangle1_ys[717]), .RECT1_WIDTH(rectangle1_widths[717]), .RECT1_HEIGHT(rectangle1_heights[717]), .RECT1_WEIGHT(rectangle1_weights[717]), .RECT2_X(rectangle2_xs[717]), .RECT2_Y(rectangle2_ys[717]), .RECT2_WIDTH(rectangle2_widths[717]), .RECT2_HEIGHT(rectangle2_heights[717]), .RECT2_WEIGHT(rectangle2_weights[717]), .RECT3_X(rectangle3_xs[717]), .RECT3_Y(rectangle3_ys[717]), .RECT3_WIDTH(rectangle3_widths[717]), .RECT3_HEIGHT(rectangle3_heights[717]), .RECT3_WEIGHT(rectangle3_weights[717]), .FEAT_THRES(feature_thresholds[717]), .FEAT_ABOVE(feature_aboves[717]), .FEAT_BELOW(feature_belows[717])) ac717(.scan_win(scan_win717), .scan_win_std_dev(scan_win_std_dev[717]), .feature_accum(feature_accums[717]));
  accum_calculator #(.RECT1_X(rectangle1_xs[718]), .RECT1_Y(rectangle1_ys[718]), .RECT1_WIDTH(rectangle1_widths[718]), .RECT1_HEIGHT(rectangle1_heights[718]), .RECT1_WEIGHT(rectangle1_weights[718]), .RECT2_X(rectangle2_xs[718]), .RECT2_Y(rectangle2_ys[718]), .RECT2_WIDTH(rectangle2_widths[718]), .RECT2_HEIGHT(rectangle2_heights[718]), .RECT2_WEIGHT(rectangle2_weights[718]), .RECT3_X(rectangle3_xs[718]), .RECT3_Y(rectangle3_ys[718]), .RECT3_WIDTH(rectangle3_widths[718]), .RECT3_HEIGHT(rectangle3_heights[718]), .RECT3_WEIGHT(rectangle3_weights[718]), .FEAT_THRES(feature_thresholds[718]), .FEAT_ABOVE(feature_aboves[718]), .FEAT_BELOW(feature_belows[718])) ac718(.scan_win(scan_win718), .scan_win_std_dev(scan_win_std_dev[718]), .feature_accum(feature_accums[718]));
  accum_calculator #(.RECT1_X(rectangle1_xs[719]), .RECT1_Y(rectangle1_ys[719]), .RECT1_WIDTH(rectangle1_widths[719]), .RECT1_HEIGHT(rectangle1_heights[719]), .RECT1_WEIGHT(rectangle1_weights[719]), .RECT2_X(rectangle2_xs[719]), .RECT2_Y(rectangle2_ys[719]), .RECT2_WIDTH(rectangle2_widths[719]), .RECT2_HEIGHT(rectangle2_heights[719]), .RECT2_WEIGHT(rectangle2_weights[719]), .RECT3_X(rectangle3_xs[719]), .RECT3_Y(rectangle3_ys[719]), .RECT3_WIDTH(rectangle3_widths[719]), .RECT3_HEIGHT(rectangle3_heights[719]), .RECT3_WEIGHT(rectangle3_weights[719]), .FEAT_THRES(feature_thresholds[719]), .FEAT_ABOVE(feature_aboves[719]), .FEAT_BELOW(feature_belows[719])) ac719(.scan_win(scan_win719), .scan_win_std_dev(scan_win_std_dev[719]), .feature_accum(feature_accums[719]));
  accum_calculator #(.RECT1_X(rectangle1_xs[720]), .RECT1_Y(rectangle1_ys[720]), .RECT1_WIDTH(rectangle1_widths[720]), .RECT1_HEIGHT(rectangle1_heights[720]), .RECT1_WEIGHT(rectangle1_weights[720]), .RECT2_X(rectangle2_xs[720]), .RECT2_Y(rectangle2_ys[720]), .RECT2_WIDTH(rectangle2_widths[720]), .RECT2_HEIGHT(rectangle2_heights[720]), .RECT2_WEIGHT(rectangle2_weights[720]), .RECT3_X(rectangle3_xs[720]), .RECT3_Y(rectangle3_ys[720]), .RECT3_WIDTH(rectangle3_widths[720]), .RECT3_HEIGHT(rectangle3_heights[720]), .RECT3_WEIGHT(rectangle3_weights[720]), .FEAT_THRES(feature_thresholds[720]), .FEAT_ABOVE(feature_aboves[720]), .FEAT_BELOW(feature_belows[720])) ac720(.scan_win(scan_win720), .scan_win_std_dev(scan_win_std_dev[720]), .feature_accum(feature_accums[720]));
  accum_calculator #(.RECT1_X(rectangle1_xs[721]), .RECT1_Y(rectangle1_ys[721]), .RECT1_WIDTH(rectangle1_widths[721]), .RECT1_HEIGHT(rectangle1_heights[721]), .RECT1_WEIGHT(rectangle1_weights[721]), .RECT2_X(rectangle2_xs[721]), .RECT2_Y(rectangle2_ys[721]), .RECT2_WIDTH(rectangle2_widths[721]), .RECT2_HEIGHT(rectangle2_heights[721]), .RECT2_WEIGHT(rectangle2_weights[721]), .RECT3_X(rectangle3_xs[721]), .RECT3_Y(rectangle3_ys[721]), .RECT3_WIDTH(rectangle3_widths[721]), .RECT3_HEIGHT(rectangle3_heights[721]), .RECT3_WEIGHT(rectangle3_weights[721]), .FEAT_THRES(feature_thresholds[721]), .FEAT_ABOVE(feature_aboves[721]), .FEAT_BELOW(feature_belows[721])) ac721(.scan_win(scan_win721), .scan_win_std_dev(scan_win_std_dev[721]), .feature_accum(feature_accums[721]));
  accum_calculator #(.RECT1_X(rectangle1_xs[722]), .RECT1_Y(rectangle1_ys[722]), .RECT1_WIDTH(rectangle1_widths[722]), .RECT1_HEIGHT(rectangle1_heights[722]), .RECT1_WEIGHT(rectangle1_weights[722]), .RECT2_X(rectangle2_xs[722]), .RECT2_Y(rectangle2_ys[722]), .RECT2_WIDTH(rectangle2_widths[722]), .RECT2_HEIGHT(rectangle2_heights[722]), .RECT2_WEIGHT(rectangle2_weights[722]), .RECT3_X(rectangle3_xs[722]), .RECT3_Y(rectangle3_ys[722]), .RECT3_WIDTH(rectangle3_widths[722]), .RECT3_HEIGHT(rectangle3_heights[722]), .RECT3_WEIGHT(rectangle3_weights[722]), .FEAT_THRES(feature_thresholds[722]), .FEAT_ABOVE(feature_aboves[722]), .FEAT_BELOW(feature_belows[722])) ac722(.scan_win(scan_win722), .scan_win_std_dev(scan_win_std_dev[722]), .feature_accum(feature_accums[722]));
  accum_calculator #(.RECT1_X(rectangle1_xs[723]), .RECT1_Y(rectangle1_ys[723]), .RECT1_WIDTH(rectangle1_widths[723]), .RECT1_HEIGHT(rectangle1_heights[723]), .RECT1_WEIGHT(rectangle1_weights[723]), .RECT2_X(rectangle2_xs[723]), .RECT2_Y(rectangle2_ys[723]), .RECT2_WIDTH(rectangle2_widths[723]), .RECT2_HEIGHT(rectangle2_heights[723]), .RECT2_WEIGHT(rectangle2_weights[723]), .RECT3_X(rectangle3_xs[723]), .RECT3_Y(rectangle3_ys[723]), .RECT3_WIDTH(rectangle3_widths[723]), .RECT3_HEIGHT(rectangle3_heights[723]), .RECT3_WEIGHT(rectangle3_weights[723]), .FEAT_THRES(feature_thresholds[723]), .FEAT_ABOVE(feature_aboves[723]), .FEAT_BELOW(feature_belows[723])) ac723(.scan_win(scan_win723), .scan_win_std_dev(scan_win_std_dev[723]), .feature_accum(feature_accums[723]));
  accum_calculator #(.RECT1_X(rectangle1_xs[724]), .RECT1_Y(rectangle1_ys[724]), .RECT1_WIDTH(rectangle1_widths[724]), .RECT1_HEIGHT(rectangle1_heights[724]), .RECT1_WEIGHT(rectangle1_weights[724]), .RECT2_X(rectangle2_xs[724]), .RECT2_Y(rectangle2_ys[724]), .RECT2_WIDTH(rectangle2_widths[724]), .RECT2_HEIGHT(rectangle2_heights[724]), .RECT2_WEIGHT(rectangle2_weights[724]), .RECT3_X(rectangle3_xs[724]), .RECT3_Y(rectangle3_ys[724]), .RECT3_WIDTH(rectangle3_widths[724]), .RECT3_HEIGHT(rectangle3_heights[724]), .RECT3_WEIGHT(rectangle3_weights[724]), .FEAT_THRES(feature_thresholds[724]), .FEAT_ABOVE(feature_aboves[724]), .FEAT_BELOW(feature_belows[724])) ac724(.scan_win(scan_win724), .scan_win_std_dev(scan_win_std_dev[724]), .feature_accum(feature_accums[724]));
  accum_calculator #(.RECT1_X(rectangle1_xs[725]), .RECT1_Y(rectangle1_ys[725]), .RECT1_WIDTH(rectangle1_widths[725]), .RECT1_HEIGHT(rectangle1_heights[725]), .RECT1_WEIGHT(rectangle1_weights[725]), .RECT2_X(rectangle2_xs[725]), .RECT2_Y(rectangle2_ys[725]), .RECT2_WIDTH(rectangle2_widths[725]), .RECT2_HEIGHT(rectangle2_heights[725]), .RECT2_WEIGHT(rectangle2_weights[725]), .RECT3_X(rectangle3_xs[725]), .RECT3_Y(rectangle3_ys[725]), .RECT3_WIDTH(rectangle3_widths[725]), .RECT3_HEIGHT(rectangle3_heights[725]), .RECT3_WEIGHT(rectangle3_weights[725]), .FEAT_THRES(feature_thresholds[725]), .FEAT_ABOVE(feature_aboves[725]), .FEAT_BELOW(feature_belows[725])) ac725(.scan_win(scan_win725), .scan_win_std_dev(scan_win_std_dev[725]), .feature_accum(feature_accums[725]));
  accum_calculator #(.RECT1_X(rectangle1_xs[726]), .RECT1_Y(rectangle1_ys[726]), .RECT1_WIDTH(rectangle1_widths[726]), .RECT1_HEIGHT(rectangle1_heights[726]), .RECT1_WEIGHT(rectangle1_weights[726]), .RECT2_X(rectangle2_xs[726]), .RECT2_Y(rectangle2_ys[726]), .RECT2_WIDTH(rectangle2_widths[726]), .RECT2_HEIGHT(rectangle2_heights[726]), .RECT2_WEIGHT(rectangle2_weights[726]), .RECT3_X(rectangle3_xs[726]), .RECT3_Y(rectangle3_ys[726]), .RECT3_WIDTH(rectangle3_widths[726]), .RECT3_HEIGHT(rectangle3_heights[726]), .RECT3_WEIGHT(rectangle3_weights[726]), .FEAT_THRES(feature_thresholds[726]), .FEAT_ABOVE(feature_aboves[726]), .FEAT_BELOW(feature_belows[726])) ac726(.scan_win(scan_win726), .scan_win_std_dev(scan_win_std_dev[726]), .feature_accum(feature_accums[726]));
  accum_calculator #(.RECT1_X(rectangle1_xs[727]), .RECT1_Y(rectangle1_ys[727]), .RECT1_WIDTH(rectangle1_widths[727]), .RECT1_HEIGHT(rectangle1_heights[727]), .RECT1_WEIGHT(rectangle1_weights[727]), .RECT2_X(rectangle2_xs[727]), .RECT2_Y(rectangle2_ys[727]), .RECT2_WIDTH(rectangle2_widths[727]), .RECT2_HEIGHT(rectangle2_heights[727]), .RECT2_WEIGHT(rectangle2_weights[727]), .RECT3_X(rectangle3_xs[727]), .RECT3_Y(rectangle3_ys[727]), .RECT3_WIDTH(rectangle3_widths[727]), .RECT3_HEIGHT(rectangle3_heights[727]), .RECT3_WEIGHT(rectangle3_weights[727]), .FEAT_THRES(feature_thresholds[727]), .FEAT_ABOVE(feature_aboves[727]), .FEAT_BELOW(feature_belows[727])) ac727(.scan_win(scan_win727), .scan_win_std_dev(scan_win_std_dev[727]), .feature_accum(feature_accums[727]));
  accum_calculator #(.RECT1_X(rectangle1_xs[728]), .RECT1_Y(rectangle1_ys[728]), .RECT1_WIDTH(rectangle1_widths[728]), .RECT1_HEIGHT(rectangle1_heights[728]), .RECT1_WEIGHT(rectangle1_weights[728]), .RECT2_X(rectangle2_xs[728]), .RECT2_Y(rectangle2_ys[728]), .RECT2_WIDTH(rectangle2_widths[728]), .RECT2_HEIGHT(rectangle2_heights[728]), .RECT2_WEIGHT(rectangle2_weights[728]), .RECT3_X(rectangle3_xs[728]), .RECT3_Y(rectangle3_ys[728]), .RECT3_WIDTH(rectangle3_widths[728]), .RECT3_HEIGHT(rectangle3_heights[728]), .RECT3_WEIGHT(rectangle3_weights[728]), .FEAT_THRES(feature_thresholds[728]), .FEAT_ABOVE(feature_aboves[728]), .FEAT_BELOW(feature_belows[728])) ac728(.scan_win(scan_win728), .scan_win_std_dev(scan_win_std_dev[728]), .feature_accum(feature_accums[728]));
  accum_calculator #(.RECT1_X(rectangle1_xs[729]), .RECT1_Y(rectangle1_ys[729]), .RECT1_WIDTH(rectangle1_widths[729]), .RECT1_HEIGHT(rectangle1_heights[729]), .RECT1_WEIGHT(rectangle1_weights[729]), .RECT2_X(rectangle2_xs[729]), .RECT2_Y(rectangle2_ys[729]), .RECT2_WIDTH(rectangle2_widths[729]), .RECT2_HEIGHT(rectangle2_heights[729]), .RECT2_WEIGHT(rectangle2_weights[729]), .RECT3_X(rectangle3_xs[729]), .RECT3_Y(rectangle3_ys[729]), .RECT3_WIDTH(rectangle3_widths[729]), .RECT3_HEIGHT(rectangle3_heights[729]), .RECT3_WEIGHT(rectangle3_weights[729]), .FEAT_THRES(feature_thresholds[729]), .FEAT_ABOVE(feature_aboves[729]), .FEAT_BELOW(feature_belows[729])) ac729(.scan_win(scan_win729), .scan_win_std_dev(scan_win_std_dev[729]), .feature_accum(feature_accums[729]));
  accum_calculator #(.RECT1_X(rectangle1_xs[730]), .RECT1_Y(rectangle1_ys[730]), .RECT1_WIDTH(rectangle1_widths[730]), .RECT1_HEIGHT(rectangle1_heights[730]), .RECT1_WEIGHT(rectangle1_weights[730]), .RECT2_X(rectangle2_xs[730]), .RECT2_Y(rectangle2_ys[730]), .RECT2_WIDTH(rectangle2_widths[730]), .RECT2_HEIGHT(rectangle2_heights[730]), .RECT2_WEIGHT(rectangle2_weights[730]), .RECT3_X(rectangle3_xs[730]), .RECT3_Y(rectangle3_ys[730]), .RECT3_WIDTH(rectangle3_widths[730]), .RECT3_HEIGHT(rectangle3_heights[730]), .RECT3_WEIGHT(rectangle3_weights[730]), .FEAT_THRES(feature_thresholds[730]), .FEAT_ABOVE(feature_aboves[730]), .FEAT_BELOW(feature_belows[730])) ac730(.scan_win(scan_win730), .scan_win_std_dev(scan_win_std_dev[730]), .feature_accum(feature_accums[730]));
  accum_calculator #(.RECT1_X(rectangle1_xs[731]), .RECT1_Y(rectangle1_ys[731]), .RECT1_WIDTH(rectangle1_widths[731]), .RECT1_HEIGHT(rectangle1_heights[731]), .RECT1_WEIGHT(rectangle1_weights[731]), .RECT2_X(rectangle2_xs[731]), .RECT2_Y(rectangle2_ys[731]), .RECT2_WIDTH(rectangle2_widths[731]), .RECT2_HEIGHT(rectangle2_heights[731]), .RECT2_WEIGHT(rectangle2_weights[731]), .RECT3_X(rectangle3_xs[731]), .RECT3_Y(rectangle3_ys[731]), .RECT3_WIDTH(rectangle3_widths[731]), .RECT3_HEIGHT(rectangle3_heights[731]), .RECT3_WEIGHT(rectangle3_weights[731]), .FEAT_THRES(feature_thresholds[731]), .FEAT_ABOVE(feature_aboves[731]), .FEAT_BELOW(feature_belows[731])) ac731(.scan_win(scan_win731), .scan_win_std_dev(scan_win_std_dev[731]), .feature_accum(feature_accums[731]));
  accum_calculator #(.RECT1_X(rectangle1_xs[732]), .RECT1_Y(rectangle1_ys[732]), .RECT1_WIDTH(rectangle1_widths[732]), .RECT1_HEIGHT(rectangle1_heights[732]), .RECT1_WEIGHT(rectangle1_weights[732]), .RECT2_X(rectangle2_xs[732]), .RECT2_Y(rectangle2_ys[732]), .RECT2_WIDTH(rectangle2_widths[732]), .RECT2_HEIGHT(rectangle2_heights[732]), .RECT2_WEIGHT(rectangle2_weights[732]), .RECT3_X(rectangle3_xs[732]), .RECT3_Y(rectangle3_ys[732]), .RECT3_WIDTH(rectangle3_widths[732]), .RECT3_HEIGHT(rectangle3_heights[732]), .RECT3_WEIGHT(rectangle3_weights[732]), .FEAT_THRES(feature_thresholds[732]), .FEAT_ABOVE(feature_aboves[732]), .FEAT_BELOW(feature_belows[732])) ac732(.scan_win(scan_win732), .scan_win_std_dev(scan_win_std_dev[732]), .feature_accum(feature_accums[732]));
  accum_calculator #(.RECT1_X(rectangle1_xs[733]), .RECT1_Y(rectangle1_ys[733]), .RECT1_WIDTH(rectangle1_widths[733]), .RECT1_HEIGHT(rectangle1_heights[733]), .RECT1_WEIGHT(rectangle1_weights[733]), .RECT2_X(rectangle2_xs[733]), .RECT2_Y(rectangle2_ys[733]), .RECT2_WIDTH(rectangle2_widths[733]), .RECT2_HEIGHT(rectangle2_heights[733]), .RECT2_WEIGHT(rectangle2_weights[733]), .RECT3_X(rectangle3_xs[733]), .RECT3_Y(rectangle3_ys[733]), .RECT3_WIDTH(rectangle3_widths[733]), .RECT3_HEIGHT(rectangle3_heights[733]), .RECT3_WEIGHT(rectangle3_weights[733]), .FEAT_THRES(feature_thresholds[733]), .FEAT_ABOVE(feature_aboves[733]), .FEAT_BELOW(feature_belows[733])) ac733(.scan_win(scan_win733), .scan_win_std_dev(scan_win_std_dev[733]), .feature_accum(feature_accums[733]));
  accum_calculator #(.RECT1_X(rectangle1_xs[734]), .RECT1_Y(rectangle1_ys[734]), .RECT1_WIDTH(rectangle1_widths[734]), .RECT1_HEIGHT(rectangle1_heights[734]), .RECT1_WEIGHT(rectangle1_weights[734]), .RECT2_X(rectangle2_xs[734]), .RECT2_Y(rectangle2_ys[734]), .RECT2_WIDTH(rectangle2_widths[734]), .RECT2_HEIGHT(rectangle2_heights[734]), .RECT2_WEIGHT(rectangle2_weights[734]), .RECT3_X(rectangle3_xs[734]), .RECT3_Y(rectangle3_ys[734]), .RECT3_WIDTH(rectangle3_widths[734]), .RECT3_HEIGHT(rectangle3_heights[734]), .RECT3_WEIGHT(rectangle3_weights[734]), .FEAT_THRES(feature_thresholds[734]), .FEAT_ABOVE(feature_aboves[734]), .FEAT_BELOW(feature_belows[734])) ac734(.scan_win(scan_win734), .scan_win_std_dev(scan_win_std_dev[734]), .feature_accum(feature_accums[734]));
  accum_calculator #(.RECT1_X(rectangle1_xs[735]), .RECT1_Y(rectangle1_ys[735]), .RECT1_WIDTH(rectangle1_widths[735]), .RECT1_HEIGHT(rectangle1_heights[735]), .RECT1_WEIGHT(rectangle1_weights[735]), .RECT2_X(rectangle2_xs[735]), .RECT2_Y(rectangle2_ys[735]), .RECT2_WIDTH(rectangle2_widths[735]), .RECT2_HEIGHT(rectangle2_heights[735]), .RECT2_WEIGHT(rectangle2_weights[735]), .RECT3_X(rectangle3_xs[735]), .RECT3_Y(rectangle3_ys[735]), .RECT3_WIDTH(rectangle3_widths[735]), .RECT3_HEIGHT(rectangle3_heights[735]), .RECT3_WEIGHT(rectangle3_weights[735]), .FEAT_THRES(feature_thresholds[735]), .FEAT_ABOVE(feature_aboves[735]), .FEAT_BELOW(feature_belows[735])) ac735(.scan_win(scan_win735), .scan_win_std_dev(scan_win_std_dev[735]), .feature_accum(feature_accums[735]));
  accum_calculator #(.RECT1_X(rectangle1_xs[736]), .RECT1_Y(rectangle1_ys[736]), .RECT1_WIDTH(rectangle1_widths[736]), .RECT1_HEIGHT(rectangle1_heights[736]), .RECT1_WEIGHT(rectangle1_weights[736]), .RECT2_X(rectangle2_xs[736]), .RECT2_Y(rectangle2_ys[736]), .RECT2_WIDTH(rectangle2_widths[736]), .RECT2_HEIGHT(rectangle2_heights[736]), .RECT2_WEIGHT(rectangle2_weights[736]), .RECT3_X(rectangle3_xs[736]), .RECT3_Y(rectangle3_ys[736]), .RECT3_WIDTH(rectangle3_widths[736]), .RECT3_HEIGHT(rectangle3_heights[736]), .RECT3_WEIGHT(rectangle3_weights[736]), .FEAT_THRES(feature_thresholds[736]), .FEAT_ABOVE(feature_aboves[736]), .FEAT_BELOW(feature_belows[736])) ac736(.scan_win(scan_win736), .scan_win_std_dev(scan_win_std_dev[736]), .feature_accum(feature_accums[736]));
  accum_calculator #(.RECT1_X(rectangle1_xs[737]), .RECT1_Y(rectangle1_ys[737]), .RECT1_WIDTH(rectangle1_widths[737]), .RECT1_HEIGHT(rectangle1_heights[737]), .RECT1_WEIGHT(rectangle1_weights[737]), .RECT2_X(rectangle2_xs[737]), .RECT2_Y(rectangle2_ys[737]), .RECT2_WIDTH(rectangle2_widths[737]), .RECT2_HEIGHT(rectangle2_heights[737]), .RECT2_WEIGHT(rectangle2_weights[737]), .RECT3_X(rectangle3_xs[737]), .RECT3_Y(rectangle3_ys[737]), .RECT3_WIDTH(rectangle3_widths[737]), .RECT3_HEIGHT(rectangle3_heights[737]), .RECT3_WEIGHT(rectangle3_weights[737]), .FEAT_THRES(feature_thresholds[737]), .FEAT_ABOVE(feature_aboves[737]), .FEAT_BELOW(feature_belows[737])) ac737(.scan_win(scan_win737), .scan_win_std_dev(scan_win_std_dev[737]), .feature_accum(feature_accums[737]));
  accum_calculator #(.RECT1_X(rectangle1_xs[738]), .RECT1_Y(rectangle1_ys[738]), .RECT1_WIDTH(rectangle1_widths[738]), .RECT1_HEIGHT(rectangle1_heights[738]), .RECT1_WEIGHT(rectangle1_weights[738]), .RECT2_X(rectangle2_xs[738]), .RECT2_Y(rectangle2_ys[738]), .RECT2_WIDTH(rectangle2_widths[738]), .RECT2_HEIGHT(rectangle2_heights[738]), .RECT2_WEIGHT(rectangle2_weights[738]), .RECT3_X(rectangle3_xs[738]), .RECT3_Y(rectangle3_ys[738]), .RECT3_WIDTH(rectangle3_widths[738]), .RECT3_HEIGHT(rectangle3_heights[738]), .RECT3_WEIGHT(rectangle3_weights[738]), .FEAT_THRES(feature_thresholds[738]), .FEAT_ABOVE(feature_aboves[738]), .FEAT_BELOW(feature_belows[738])) ac738(.scan_win(scan_win738), .scan_win_std_dev(scan_win_std_dev[738]), .feature_accum(feature_accums[738]));
  accum_calculator #(.RECT1_X(rectangle1_xs[739]), .RECT1_Y(rectangle1_ys[739]), .RECT1_WIDTH(rectangle1_widths[739]), .RECT1_HEIGHT(rectangle1_heights[739]), .RECT1_WEIGHT(rectangle1_weights[739]), .RECT2_X(rectangle2_xs[739]), .RECT2_Y(rectangle2_ys[739]), .RECT2_WIDTH(rectangle2_widths[739]), .RECT2_HEIGHT(rectangle2_heights[739]), .RECT2_WEIGHT(rectangle2_weights[739]), .RECT3_X(rectangle3_xs[739]), .RECT3_Y(rectangle3_ys[739]), .RECT3_WIDTH(rectangle3_widths[739]), .RECT3_HEIGHT(rectangle3_heights[739]), .RECT3_WEIGHT(rectangle3_weights[739]), .FEAT_THRES(feature_thresholds[739]), .FEAT_ABOVE(feature_aboves[739]), .FEAT_BELOW(feature_belows[739])) ac739(.scan_win(scan_win739), .scan_win_std_dev(scan_win_std_dev[739]), .feature_accum(feature_accums[739]));
  accum_calculator #(.RECT1_X(rectangle1_xs[740]), .RECT1_Y(rectangle1_ys[740]), .RECT1_WIDTH(rectangle1_widths[740]), .RECT1_HEIGHT(rectangle1_heights[740]), .RECT1_WEIGHT(rectangle1_weights[740]), .RECT2_X(rectangle2_xs[740]), .RECT2_Y(rectangle2_ys[740]), .RECT2_WIDTH(rectangle2_widths[740]), .RECT2_HEIGHT(rectangle2_heights[740]), .RECT2_WEIGHT(rectangle2_weights[740]), .RECT3_X(rectangle3_xs[740]), .RECT3_Y(rectangle3_ys[740]), .RECT3_WIDTH(rectangle3_widths[740]), .RECT3_HEIGHT(rectangle3_heights[740]), .RECT3_WEIGHT(rectangle3_weights[740]), .FEAT_THRES(feature_thresholds[740]), .FEAT_ABOVE(feature_aboves[740]), .FEAT_BELOW(feature_belows[740])) ac740(.scan_win(scan_win740), .scan_win_std_dev(scan_win_std_dev[740]), .feature_accum(feature_accums[740]));
  accum_calculator #(.RECT1_X(rectangle1_xs[741]), .RECT1_Y(rectangle1_ys[741]), .RECT1_WIDTH(rectangle1_widths[741]), .RECT1_HEIGHT(rectangle1_heights[741]), .RECT1_WEIGHT(rectangle1_weights[741]), .RECT2_X(rectangle2_xs[741]), .RECT2_Y(rectangle2_ys[741]), .RECT2_WIDTH(rectangle2_widths[741]), .RECT2_HEIGHT(rectangle2_heights[741]), .RECT2_WEIGHT(rectangle2_weights[741]), .RECT3_X(rectangle3_xs[741]), .RECT3_Y(rectangle3_ys[741]), .RECT3_WIDTH(rectangle3_widths[741]), .RECT3_HEIGHT(rectangle3_heights[741]), .RECT3_WEIGHT(rectangle3_weights[741]), .FEAT_THRES(feature_thresholds[741]), .FEAT_ABOVE(feature_aboves[741]), .FEAT_BELOW(feature_belows[741])) ac741(.scan_win(scan_win741), .scan_win_std_dev(scan_win_std_dev[741]), .feature_accum(feature_accums[741]));
  accum_calculator #(.RECT1_X(rectangle1_xs[742]), .RECT1_Y(rectangle1_ys[742]), .RECT1_WIDTH(rectangle1_widths[742]), .RECT1_HEIGHT(rectangle1_heights[742]), .RECT1_WEIGHT(rectangle1_weights[742]), .RECT2_X(rectangle2_xs[742]), .RECT2_Y(rectangle2_ys[742]), .RECT2_WIDTH(rectangle2_widths[742]), .RECT2_HEIGHT(rectangle2_heights[742]), .RECT2_WEIGHT(rectangle2_weights[742]), .RECT3_X(rectangle3_xs[742]), .RECT3_Y(rectangle3_ys[742]), .RECT3_WIDTH(rectangle3_widths[742]), .RECT3_HEIGHT(rectangle3_heights[742]), .RECT3_WEIGHT(rectangle3_weights[742]), .FEAT_THRES(feature_thresholds[742]), .FEAT_ABOVE(feature_aboves[742]), .FEAT_BELOW(feature_belows[742])) ac742(.scan_win(scan_win742), .scan_win_std_dev(scan_win_std_dev[742]), .feature_accum(feature_accums[742]));
  accum_calculator #(.RECT1_X(rectangle1_xs[743]), .RECT1_Y(rectangle1_ys[743]), .RECT1_WIDTH(rectangle1_widths[743]), .RECT1_HEIGHT(rectangle1_heights[743]), .RECT1_WEIGHT(rectangle1_weights[743]), .RECT2_X(rectangle2_xs[743]), .RECT2_Y(rectangle2_ys[743]), .RECT2_WIDTH(rectangle2_widths[743]), .RECT2_HEIGHT(rectangle2_heights[743]), .RECT2_WEIGHT(rectangle2_weights[743]), .RECT3_X(rectangle3_xs[743]), .RECT3_Y(rectangle3_ys[743]), .RECT3_WIDTH(rectangle3_widths[743]), .RECT3_HEIGHT(rectangle3_heights[743]), .RECT3_WEIGHT(rectangle3_weights[743]), .FEAT_THRES(feature_thresholds[743]), .FEAT_ABOVE(feature_aboves[743]), .FEAT_BELOW(feature_belows[743])) ac743(.scan_win(scan_win743), .scan_win_std_dev(scan_win_std_dev[743]), .feature_accum(feature_accums[743]));
  accum_calculator #(.RECT1_X(rectangle1_xs[744]), .RECT1_Y(rectangle1_ys[744]), .RECT1_WIDTH(rectangle1_widths[744]), .RECT1_HEIGHT(rectangle1_heights[744]), .RECT1_WEIGHT(rectangle1_weights[744]), .RECT2_X(rectangle2_xs[744]), .RECT2_Y(rectangle2_ys[744]), .RECT2_WIDTH(rectangle2_widths[744]), .RECT2_HEIGHT(rectangle2_heights[744]), .RECT2_WEIGHT(rectangle2_weights[744]), .RECT3_X(rectangle3_xs[744]), .RECT3_Y(rectangle3_ys[744]), .RECT3_WIDTH(rectangle3_widths[744]), .RECT3_HEIGHT(rectangle3_heights[744]), .RECT3_WEIGHT(rectangle3_weights[744]), .FEAT_THRES(feature_thresholds[744]), .FEAT_ABOVE(feature_aboves[744]), .FEAT_BELOW(feature_belows[744])) ac744(.scan_win(scan_win744), .scan_win_std_dev(scan_win_std_dev[744]), .feature_accum(feature_accums[744]));
  accum_calculator #(.RECT1_X(rectangle1_xs[745]), .RECT1_Y(rectangle1_ys[745]), .RECT1_WIDTH(rectangle1_widths[745]), .RECT1_HEIGHT(rectangle1_heights[745]), .RECT1_WEIGHT(rectangle1_weights[745]), .RECT2_X(rectangle2_xs[745]), .RECT2_Y(rectangle2_ys[745]), .RECT2_WIDTH(rectangle2_widths[745]), .RECT2_HEIGHT(rectangle2_heights[745]), .RECT2_WEIGHT(rectangle2_weights[745]), .RECT3_X(rectangle3_xs[745]), .RECT3_Y(rectangle3_ys[745]), .RECT3_WIDTH(rectangle3_widths[745]), .RECT3_HEIGHT(rectangle3_heights[745]), .RECT3_WEIGHT(rectangle3_weights[745]), .FEAT_THRES(feature_thresholds[745]), .FEAT_ABOVE(feature_aboves[745]), .FEAT_BELOW(feature_belows[745])) ac745(.scan_win(scan_win745), .scan_win_std_dev(scan_win_std_dev[745]), .feature_accum(feature_accums[745]));
  accum_calculator #(.RECT1_X(rectangle1_xs[746]), .RECT1_Y(rectangle1_ys[746]), .RECT1_WIDTH(rectangle1_widths[746]), .RECT1_HEIGHT(rectangle1_heights[746]), .RECT1_WEIGHT(rectangle1_weights[746]), .RECT2_X(rectangle2_xs[746]), .RECT2_Y(rectangle2_ys[746]), .RECT2_WIDTH(rectangle2_widths[746]), .RECT2_HEIGHT(rectangle2_heights[746]), .RECT2_WEIGHT(rectangle2_weights[746]), .RECT3_X(rectangle3_xs[746]), .RECT3_Y(rectangle3_ys[746]), .RECT3_WIDTH(rectangle3_widths[746]), .RECT3_HEIGHT(rectangle3_heights[746]), .RECT3_WEIGHT(rectangle3_weights[746]), .FEAT_THRES(feature_thresholds[746]), .FEAT_ABOVE(feature_aboves[746]), .FEAT_BELOW(feature_belows[746])) ac746(.scan_win(scan_win746), .scan_win_std_dev(scan_win_std_dev[746]), .feature_accum(feature_accums[746]));
  accum_calculator #(.RECT1_X(rectangle1_xs[747]), .RECT1_Y(rectangle1_ys[747]), .RECT1_WIDTH(rectangle1_widths[747]), .RECT1_HEIGHT(rectangle1_heights[747]), .RECT1_WEIGHT(rectangle1_weights[747]), .RECT2_X(rectangle2_xs[747]), .RECT2_Y(rectangle2_ys[747]), .RECT2_WIDTH(rectangle2_widths[747]), .RECT2_HEIGHT(rectangle2_heights[747]), .RECT2_WEIGHT(rectangle2_weights[747]), .RECT3_X(rectangle3_xs[747]), .RECT3_Y(rectangle3_ys[747]), .RECT3_WIDTH(rectangle3_widths[747]), .RECT3_HEIGHT(rectangle3_heights[747]), .RECT3_WEIGHT(rectangle3_weights[747]), .FEAT_THRES(feature_thresholds[747]), .FEAT_ABOVE(feature_aboves[747]), .FEAT_BELOW(feature_belows[747])) ac747(.scan_win(scan_win747), .scan_win_std_dev(scan_win_std_dev[747]), .feature_accum(feature_accums[747]));
  accum_calculator #(.RECT1_X(rectangle1_xs[748]), .RECT1_Y(rectangle1_ys[748]), .RECT1_WIDTH(rectangle1_widths[748]), .RECT1_HEIGHT(rectangle1_heights[748]), .RECT1_WEIGHT(rectangle1_weights[748]), .RECT2_X(rectangle2_xs[748]), .RECT2_Y(rectangle2_ys[748]), .RECT2_WIDTH(rectangle2_widths[748]), .RECT2_HEIGHT(rectangle2_heights[748]), .RECT2_WEIGHT(rectangle2_weights[748]), .RECT3_X(rectangle3_xs[748]), .RECT3_Y(rectangle3_ys[748]), .RECT3_WIDTH(rectangle3_widths[748]), .RECT3_HEIGHT(rectangle3_heights[748]), .RECT3_WEIGHT(rectangle3_weights[748]), .FEAT_THRES(feature_thresholds[748]), .FEAT_ABOVE(feature_aboves[748]), .FEAT_BELOW(feature_belows[748])) ac748(.scan_win(scan_win748), .scan_win_std_dev(scan_win_std_dev[748]), .feature_accum(feature_accums[748]));
  accum_calculator #(.RECT1_X(rectangle1_xs[749]), .RECT1_Y(rectangle1_ys[749]), .RECT1_WIDTH(rectangle1_widths[749]), .RECT1_HEIGHT(rectangle1_heights[749]), .RECT1_WEIGHT(rectangle1_weights[749]), .RECT2_X(rectangle2_xs[749]), .RECT2_Y(rectangle2_ys[749]), .RECT2_WIDTH(rectangle2_widths[749]), .RECT2_HEIGHT(rectangle2_heights[749]), .RECT2_WEIGHT(rectangle2_weights[749]), .RECT3_X(rectangle3_xs[749]), .RECT3_Y(rectangle3_ys[749]), .RECT3_WIDTH(rectangle3_widths[749]), .RECT3_HEIGHT(rectangle3_heights[749]), .RECT3_WEIGHT(rectangle3_weights[749]), .FEAT_THRES(feature_thresholds[749]), .FEAT_ABOVE(feature_aboves[749]), .FEAT_BELOW(feature_belows[749])) ac749(.scan_win(scan_win749), .scan_win_std_dev(scan_win_std_dev[749]), .feature_accum(feature_accums[749]));
  accum_calculator #(.RECT1_X(rectangle1_xs[750]), .RECT1_Y(rectangle1_ys[750]), .RECT1_WIDTH(rectangle1_widths[750]), .RECT1_HEIGHT(rectangle1_heights[750]), .RECT1_WEIGHT(rectangle1_weights[750]), .RECT2_X(rectangle2_xs[750]), .RECT2_Y(rectangle2_ys[750]), .RECT2_WIDTH(rectangle2_widths[750]), .RECT2_HEIGHT(rectangle2_heights[750]), .RECT2_WEIGHT(rectangle2_weights[750]), .RECT3_X(rectangle3_xs[750]), .RECT3_Y(rectangle3_ys[750]), .RECT3_WIDTH(rectangle3_widths[750]), .RECT3_HEIGHT(rectangle3_heights[750]), .RECT3_WEIGHT(rectangle3_weights[750]), .FEAT_THRES(feature_thresholds[750]), .FEAT_ABOVE(feature_aboves[750]), .FEAT_BELOW(feature_belows[750])) ac750(.scan_win(scan_win750), .scan_win_std_dev(scan_win_std_dev[750]), .feature_accum(feature_accums[750]));
  accum_calculator #(.RECT1_X(rectangle1_xs[751]), .RECT1_Y(rectangle1_ys[751]), .RECT1_WIDTH(rectangle1_widths[751]), .RECT1_HEIGHT(rectangle1_heights[751]), .RECT1_WEIGHT(rectangle1_weights[751]), .RECT2_X(rectangle2_xs[751]), .RECT2_Y(rectangle2_ys[751]), .RECT2_WIDTH(rectangle2_widths[751]), .RECT2_HEIGHT(rectangle2_heights[751]), .RECT2_WEIGHT(rectangle2_weights[751]), .RECT3_X(rectangle3_xs[751]), .RECT3_Y(rectangle3_ys[751]), .RECT3_WIDTH(rectangle3_widths[751]), .RECT3_HEIGHT(rectangle3_heights[751]), .RECT3_WEIGHT(rectangle3_weights[751]), .FEAT_THRES(feature_thresholds[751]), .FEAT_ABOVE(feature_aboves[751]), .FEAT_BELOW(feature_belows[751])) ac751(.scan_win(scan_win751), .scan_win_std_dev(scan_win_std_dev[751]), .feature_accum(feature_accums[751]));
  accum_calculator #(.RECT1_X(rectangle1_xs[752]), .RECT1_Y(rectangle1_ys[752]), .RECT1_WIDTH(rectangle1_widths[752]), .RECT1_HEIGHT(rectangle1_heights[752]), .RECT1_WEIGHT(rectangle1_weights[752]), .RECT2_X(rectangle2_xs[752]), .RECT2_Y(rectangle2_ys[752]), .RECT2_WIDTH(rectangle2_widths[752]), .RECT2_HEIGHT(rectangle2_heights[752]), .RECT2_WEIGHT(rectangle2_weights[752]), .RECT3_X(rectangle3_xs[752]), .RECT3_Y(rectangle3_ys[752]), .RECT3_WIDTH(rectangle3_widths[752]), .RECT3_HEIGHT(rectangle3_heights[752]), .RECT3_WEIGHT(rectangle3_weights[752]), .FEAT_THRES(feature_thresholds[752]), .FEAT_ABOVE(feature_aboves[752]), .FEAT_BELOW(feature_belows[752])) ac752(.scan_win(scan_win752), .scan_win_std_dev(scan_win_std_dev[752]), .feature_accum(feature_accums[752]));
  accum_calculator #(.RECT1_X(rectangle1_xs[753]), .RECT1_Y(rectangle1_ys[753]), .RECT1_WIDTH(rectangle1_widths[753]), .RECT1_HEIGHT(rectangle1_heights[753]), .RECT1_WEIGHT(rectangle1_weights[753]), .RECT2_X(rectangle2_xs[753]), .RECT2_Y(rectangle2_ys[753]), .RECT2_WIDTH(rectangle2_widths[753]), .RECT2_HEIGHT(rectangle2_heights[753]), .RECT2_WEIGHT(rectangle2_weights[753]), .RECT3_X(rectangle3_xs[753]), .RECT3_Y(rectangle3_ys[753]), .RECT3_WIDTH(rectangle3_widths[753]), .RECT3_HEIGHT(rectangle3_heights[753]), .RECT3_WEIGHT(rectangle3_weights[753]), .FEAT_THRES(feature_thresholds[753]), .FEAT_ABOVE(feature_aboves[753]), .FEAT_BELOW(feature_belows[753])) ac753(.scan_win(scan_win753), .scan_win_std_dev(scan_win_std_dev[753]), .feature_accum(feature_accums[753]));
  accum_calculator #(.RECT1_X(rectangle1_xs[754]), .RECT1_Y(rectangle1_ys[754]), .RECT1_WIDTH(rectangle1_widths[754]), .RECT1_HEIGHT(rectangle1_heights[754]), .RECT1_WEIGHT(rectangle1_weights[754]), .RECT2_X(rectangle2_xs[754]), .RECT2_Y(rectangle2_ys[754]), .RECT2_WIDTH(rectangle2_widths[754]), .RECT2_HEIGHT(rectangle2_heights[754]), .RECT2_WEIGHT(rectangle2_weights[754]), .RECT3_X(rectangle3_xs[754]), .RECT3_Y(rectangle3_ys[754]), .RECT3_WIDTH(rectangle3_widths[754]), .RECT3_HEIGHT(rectangle3_heights[754]), .RECT3_WEIGHT(rectangle3_weights[754]), .FEAT_THRES(feature_thresholds[754]), .FEAT_ABOVE(feature_aboves[754]), .FEAT_BELOW(feature_belows[754])) ac754(.scan_win(scan_win754), .scan_win_std_dev(scan_win_std_dev[754]), .feature_accum(feature_accums[754]));
  accum_calculator #(.RECT1_X(rectangle1_xs[755]), .RECT1_Y(rectangle1_ys[755]), .RECT1_WIDTH(rectangle1_widths[755]), .RECT1_HEIGHT(rectangle1_heights[755]), .RECT1_WEIGHT(rectangle1_weights[755]), .RECT2_X(rectangle2_xs[755]), .RECT2_Y(rectangle2_ys[755]), .RECT2_WIDTH(rectangle2_widths[755]), .RECT2_HEIGHT(rectangle2_heights[755]), .RECT2_WEIGHT(rectangle2_weights[755]), .RECT3_X(rectangle3_xs[755]), .RECT3_Y(rectangle3_ys[755]), .RECT3_WIDTH(rectangle3_widths[755]), .RECT3_HEIGHT(rectangle3_heights[755]), .RECT3_WEIGHT(rectangle3_weights[755]), .FEAT_THRES(feature_thresholds[755]), .FEAT_ABOVE(feature_aboves[755]), .FEAT_BELOW(feature_belows[755])) ac755(.scan_win(scan_win755), .scan_win_std_dev(scan_win_std_dev[755]), .feature_accum(feature_accums[755]));
  accum_calculator #(.RECT1_X(rectangle1_xs[756]), .RECT1_Y(rectangle1_ys[756]), .RECT1_WIDTH(rectangle1_widths[756]), .RECT1_HEIGHT(rectangle1_heights[756]), .RECT1_WEIGHT(rectangle1_weights[756]), .RECT2_X(rectangle2_xs[756]), .RECT2_Y(rectangle2_ys[756]), .RECT2_WIDTH(rectangle2_widths[756]), .RECT2_HEIGHT(rectangle2_heights[756]), .RECT2_WEIGHT(rectangle2_weights[756]), .RECT3_X(rectangle3_xs[756]), .RECT3_Y(rectangle3_ys[756]), .RECT3_WIDTH(rectangle3_widths[756]), .RECT3_HEIGHT(rectangle3_heights[756]), .RECT3_WEIGHT(rectangle3_weights[756]), .FEAT_THRES(feature_thresholds[756]), .FEAT_ABOVE(feature_aboves[756]), .FEAT_BELOW(feature_belows[756])) ac756(.scan_win(scan_win756), .scan_win_std_dev(scan_win_std_dev[756]), .feature_accum(feature_accums[756]));
  accum_calculator #(.RECT1_X(rectangle1_xs[757]), .RECT1_Y(rectangle1_ys[757]), .RECT1_WIDTH(rectangle1_widths[757]), .RECT1_HEIGHT(rectangle1_heights[757]), .RECT1_WEIGHT(rectangle1_weights[757]), .RECT2_X(rectangle2_xs[757]), .RECT2_Y(rectangle2_ys[757]), .RECT2_WIDTH(rectangle2_widths[757]), .RECT2_HEIGHT(rectangle2_heights[757]), .RECT2_WEIGHT(rectangle2_weights[757]), .RECT3_X(rectangle3_xs[757]), .RECT3_Y(rectangle3_ys[757]), .RECT3_WIDTH(rectangle3_widths[757]), .RECT3_HEIGHT(rectangle3_heights[757]), .RECT3_WEIGHT(rectangle3_weights[757]), .FEAT_THRES(feature_thresholds[757]), .FEAT_ABOVE(feature_aboves[757]), .FEAT_BELOW(feature_belows[757])) ac757(.scan_win(scan_win757), .scan_win_std_dev(scan_win_std_dev[757]), .feature_accum(feature_accums[757]));
  accum_calculator #(.RECT1_X(rectangle1_xs[758]), .RECT1_Y(rectangle1_ys[758]), .RECT1_WIDTH(rectangle1_widths[758]), .RECT1_HEIGHT(rectangle1_heights[758]), .RECT1_WEIGHT(rectangle1_weights[758]), .RECT2_X(rectangle2_xs[758]), .RECT2_Y(rectangle2_ys[758]), .RECT2_WIDTH(rectangle2_widths[758]), .RECT2_HEIGHT(rectangle2_heights[758]), .RECT2_WEIGHT(rectangle2_weights[758]), .RECT3_X(rectangle3_xs[758]), .RECT3_Y(rectangle3_ys[758]), .RECT3_WIDTH(rectangle3_widths[758]), .RECT3_HEIGHT(rectangle3_heights[758]), .RECT3_WEIGHT(rectangle3_weights[758]), .FEAT_THRES(feature_thresholds[758]), .FEAT_ABOVE(feature_aboves[758]), .FEAT_BELOW(feature_belows[758])) ac758(.scan_win(scan_win758), .scan_win_std_dev(scan_win_std_dev[758]), .feature_accum(feature_accums[758]));
  accum_calculator #(.RECT1_X(rectangle1_xs[759]), .RECT1_Y(rectangle1_ys[759]), .RECT1_WIDTH(rectangle1_widths[759]), .RECT1_HEIGHT(rectangle1_heights[759]), .RECT1_WEIGHT(rectangle1_weights[759]), .RECT2_X(rectangle2_xs[759]), .RECT2_Y(rectangle2_ys[759]), .RECT2_WIDTH(rectangle2_widths[759]), .RECT2_HEIGHT(rectangle2_heights[759]), .RECT2_WEIGHT(rectangle2_weights[759]), .RECT3_X(rectangle3_xs[759]), .RECT3_Y(rectangle3_ys[759]), .RECT3_WIDTH(rectangle3_widths[759]), .RECT3_HEIGHT(rectangle3_heights[759]), .RECT3_WEIGHT(rectangle3_weights[759]), .FEAT_THRES(feature_thresholds[759]), .FEAT_ABOVE(feature_aboves[759]), .FEAT_BELOW(feature_belows[759])) ac759(.scan_win(scan_win759), .scan_win_std_dev(scan_win_std_dev[759]), .feature_accum(feature_accums[759]));
  accum_calculator #(.RECT1_X(rectangle1_xs[760]), .RECT1_Y(rectangle1_ys[760]), .RECT1_WIDTH(rectangle1_widths[760]), .RECT1_HEIGHT(rectangle1_heights[760]), .RECT1_WEIGHT(rectangle1_weights[760]), .RECT2_X(rectangle2_xs[760]), .RECT2_Y(rectangle2_ys[760]), .RECT2_WIDTH(rectangle2_widths[760]), .RECT2_HEIGHT(rectangle2_heights[760]), .RECT2_WEIGHT(rectangle2_weights[760]), .RECT3_X(rectangle3_xs[760]), .RECT3_Y(rectangle3_ys[760]), .RECT3_WIDTH(rectangle3_widths[760]), .RECT3_HEIGHT(rectangle3_heights[760]), .RECT3_WEIGHT(rectangle3_weights[760]), .FEAT_THRES(feature_thresholds[760]), .FEAT_ABOVE(feature_aboves[760]), .FEAT_BELOW(feature_belows[760])) ac760(.scan_win(scan_win760), .scan_win_std_dev(scan_win_std_dev[760]), .feature_accum(feature_accums[760]));
  accum_calculator #(.RECT1_X(rectangle1_xs[761]), .RECT1_Y(rectangle1_ys[761]), .RECT1_WIDTH(rectangle1_widths[761]), .RECT1_HEIGHT(rectangle1_heights[761]), .RECT1_WEIGHT(rectangle1_weights[761]), .RECT2_X(rectangle2_xs[761]), .RECT2_Y(rectangle2_ys[761]), .RECT2_WIDTH(rectangle2_widths[761]), .RECT2_HEIGHT(rectangle2_heights[761]), .RECT2_WEIGHT(rectangle2_weights[761]), .RECT3_X(rectangle3_xs[761]), .RECT3_Y(rectangle3_ys[761]), .RECT3_WIDTH(rectangle3_widths[761]), .RECT3_HEIGHT(rectangle3_heights[761]), .RECT3_WEIGHT(rectangle3_weights[761]), .FEAT_THRES(feature_thresholds[761]), .FEAT_ABOVE(feature_aboves[761]), .FEAT_BELOW(feature_belows[761])) ac761(.scan_win(scan_win761), .scan_win_std_dev(scan_win_std_dev[761]), .feature_accum(feature_accums[761]));
  accum_calculator #(.RECT1_X(rectangle1_xs[762]), .RECT1_Y(rectangle1_ys[762]), .RECT1_WIDTH(rectangle1_widths[762]), .RECT1_HEIGHT(rectangle1_heights[762]), .RECT1_WEIGHT(rectangle1_weights[762]), .RECT2_X(rectangle2_xs[762]), .RECT2_Y(rectangle2_ys[762]), .RECT2_WIDTH(rectangle2_widths[762]), .RECT2_HEIGHT(rectangle2_heights[762]), .RECT2_WEIGHT(rectangle2_weights[762]), .RECT3_X(rectangle3_xs[762]), .RECT3_Y(rectangle3_ys[762]), .RECT3_WIDTH(rectangle3_widths[762]), .RECT3_HEIGHT(rectangle3_heights[762]), .RECT3_WEIGHT(rectangle3_weights[762]), .FEAT_THRES(feature_thresholds[762]), .FEAT_ABOVE(feature_aboves[762]), .FEAT_BELOW(feature_belows[762])) ac762(.scan_win(scan_win762), .scan_win_std_dev(scan_win_std_dev[762]), .feature_accum(feature_accums[762]));
  accum_calculator #(.RECT1_X(rectangle1_xs[763]), .RECT1_Y(rectangle1_ys[763]), .RECT1_WIDTH(rectangle1_widths[763]), .RECT1_HEIGHT(rectangle1_heights[763]), .RECT1_WEIGHT(rectangle1_weights[763]), .RECT2_X(rectangle2_xs[763]), .RECT2_Y(rectangle2_ys[763]), .RECT2_WIDTH(rectangle2_widths[763]), .RECT2_HEIGHT(rectangle2_heights[763]), .RECT2_WEIGHT(rectangle2_weights[763]), .RECT3_X(rectangle3_xs[763]), .RECT3_Y(rectangle3_ys[763]), .RECT3_WIDTH(rectangle3_widths[763]), .RECT3_HEIGHT(rectangle3_heights[763]), .RECT3_WEIGHT(rectangle3_weights[763]), .FEAT_THRES(feature_thresholds[763]), .FEAT_ABOVE(feature_aboves[763]), .FEAT_BELOW(feature_belows[763])) ac763(.scan_win(scan_win763), .scan_win_std_dev(scan_win_std_dev[763]), .feature_accum(feature_accums[763]));
  accum_calculator #(.RECT1_X(rectangle1_xs[764]), .RECT1_Y(rectangle1_ys[764]), .RECT1_WIDTH(rectangle1_widths[764]), .RECT1_HEIGHT(rectangle1_heights[764]), .RECT1_WEIGHT(rectangle1_weights[764]), .RECT2_X(rectangle2_xs[764]), .RECT2_Y(rectangle2_ys[764]), .RECT2_WIDTH(rectangle2_widths[764]), .RECT2_HEIGHT(rectangle2_heights[764]), .RECT2_WEIGHT(rectangle2_weights[764]), .RECT3_X(rectangle3_xs[764]), .RECT3_Y(rectangle3_ys[764]), .RECT3_WIDTH(rectangle3_widths[764]), .RECT3_HEIGHT(rectangle3_heights[764]), .RECT3_WEIGHT(rectangle3_weights[764]), .FEAT_THRES(feature_thresholds[764]), .FEAT_ABOVE(feature_aboves[764]), .FEAT_BELOW(feature_belows[764])) ac764(.scan_win(scan_win764), .scan_win_std_dev(scan_win_std_dev[764]), .feature_accum(feature_accums[764]));
  accum_calculator #(.RECT1_X(rectangle1_xs[765]), .RECT1_Y(rectangle1_ys[765]), .RECT1_WIDTH(rectangle1_widths[765]), .RECT1_HEIGHT(rectangle1_heights[765]), .RECT1_WEIGHT(rectangle1_weights[765]), .RECT2_X(rectangle2_xs[765]), .RECT2_Y(rectangle2_ys[765]), .RECT2_WIDTH(rectangle2_widths[765]), .RECT2_HEIGHT(rectangle2_heights[765]), .RECT2_WEIGHT(rectangle2_weights[765]), .RECT3_X(rectangle3_xs[765]), .RECT3_Y(rectangle3_ys[765]), .RECT3_WIDTH(rectangle3_widths[765]), .RECT3_HEIGHT(rectangle3_heights[765]), .RECT3_WEIGHT(rectangle3_weights[765]), .FEAT_THRES(feature_thresholds[765]), .FEAT_ABOVE(feature_aboves[765]), .FEAT_BELOW(feature_belows[765])) ac765(.scan_win(scan_win765), .scan_win_std_dev(scan_win_std_dev[765]), .feature_accum(feature_accums[765]));
  accum_calculator #(.RECT1_X(rectangle1_xs[766]), .RECT1_Y(rectangle1_ys[766]), .RECT1_WIDTH(rectangle1_widths[766]), .RECT1_HEIGHT(rectangle1_heights[766]), .RECT1_WEIGHT(rectangle1_weights[766]), .RECT2_X(rectangle2_xs[766]), .RECT2_Y(rectangle2_ys[766]), .RECT2_WIDTH(rectangle2_widths[766]), .RECT2_HEIGHT(rectangle2_heights[766]), .RECT2_WEIGHT(rectangle2_weights[766]), .RECT3_X(rectangle3_xs[766]), .RECT3_Y(rectangle3_ys[766]), .RECT3_WIDTH(rectangle3_widths[766]), .RECT3_HEIGHT(rectangle3_heights[766]), .RECT3_WEIGHT(rectangle3_weights[766]), .FEAT_THRES(feature_thresholds[766]), .FEAT_ABOVE(feature_aboves[766]), .FEAT_BELOW(feature_belows[766])) ac766(.scan_win(scan_win766), .scan_win_std_dev(scan_win_std_dev[766]), .feature_accum(feature_accums[766]));
  accum_calculator #(.RECT1_X(rectangle1_xs[767]), .RECT1_Y(rectangle1_ys[767]), .RECT1_WIDTH(rectangle1_widths[767]), .RECT1_HEIGHT(rectangle1_heights[767]), .RECT1_WEIGHT(rectangle1_weights[767]), .RECT2_X(rectangle2_xs[767]), .RECT2_Y(rectangle2_ys[767]), .RECT2_WIDTH(rectangle2_widths[767]), .RECT2_HEIGHT(rectangle2_heights[767]), .RECT2_WEIGHT(rectangle2_weights[767]), .RECT3_X(rectangle3_xs[767]), .RECT3_Y(rectangle3_ys[767]), .RECT3_WIDTH(rectangle3_widths[767]), .RECT3_HEIGHT(rectangle3_heights[767]), .RECT3_WEIGHT(rectangle3_weights[767]), .FEAT_THRES(feature_thresholds[767]), .FEAT_ABOVE(feature_aboves[767]), .FEAT_BELOW(feature_belows[767])) ac767(.scan_win(scan_win767), .scan_win_std_dev(scan_win_std_dev[767]), .feature_accum(feature_accums[767]));
  accum_calculator #(.RECT1_X(rectangle1_xs[768]), .RECT1_Y(rectangle1_ys[768]), .RECT1_WIDTH(rectangle1_widths[768]), .RECT1_HEIGHT(rectangle1_heights[768]), .RECT1_WEIGHT(rectangle1_weights[768]), .RECT2_X(rectangle2_xs[768]), .RECT2_Y(rectangle2_ys[768]), .RECT2_WIDTH(rectangle2_widths[768]), .RECT2_HEIGHT(rectangle2_heights[768]), .RECT2_WEIGHT(rectangle2_weights[768]), .RECT3_X(rectangle3_xs[768]), .RECT3_Y(rectangle3_ys[768]), .RECT3_WIDTH(rectangle3_widths[768]), .RECT3_HEIGHT(rectangle3_heights[768]), .RECT3_WEIGHT(rectangle3_weights[768]), .FEAT_THRES(feature_thresholds[768]), .FEAT_ABOVE(feature_aboves[768]), .FEAT_BELOW(feature_belows[768])) ac768(.scan_win(scan_win768), .scan_win_std_dev(scan_win_std_dev[768]), .feature_accum(feature_accums[768]));
  accum_calculator #(.RECT1_X(rectangle1_xs[769]), .RECT1_Y(rectangle1_ys[769]), .RECT1_WIDTH(rectangle1_widths[769]), .RECT1_HEIGHT(rectangle1_heights[769]), .RECT1_WEIGHT(rectangle1_weights[769]), .RECT2_X(rectangle2_xs[769]), .RECT2_Y(rectangle2_ys[769]), .RECT2_WIDTH(rectangle2_widths[769]), .RECT2_HEIGHT(rectangle2_heights[769]), .RECT2_WEIGHT(rectangle2_weights[769]), .RECT3_X(rectangle3_xs[769]), .RECT3_Y(rectangle3_ys[769]), .RECT3_WIDTH(rectangle3_widths[769]), .RECT3_HEIGHT(rectangle3_heights[769]), .RECT3_WEIGHT(rectangle3_weights[769]), .FEAT_THRES(feature_thresholds[769]), .FEAT_ABOVE(feature_aboves[769]), .FEAT_BELOW(feature_belows[769])) ac769(.scan_win(scan_win769), .scan_win_std_dev(scan_win_std_dev[769]), .feature_accum(feature_accums[769]));
  accum_calculator #(.RECT1_X(rectangle1_xs[770]), .RECT1_Y(rectangle1_ys[770]), .RECT1_WIDTH(rectangle1_widths[770]), .RECT1_HEIGHT(rectangle1_heights[770]), .RECT1_WEIGHT(rectangle1_weights[770]), .RECT2_X(rectangle2_xs[770]), .RECT2_Y(rectangle2_ys[770]), .RECT2_WIDTH(rectangle2_widths[770]), .RECT2_HEIGHT(rectangle2_heights[770]), .RECT2_WEIGHT(rectangle2_weights[770]), .RECT3_X(rectangle3_xs[770]), .RECT3_Y(rectangle3_ys[770]), .RECT3_WIDTH(rectangle3_widths[770]), .RECT3_HEIGHT(rectangle3_heights[770]), .RECT3_WEIGHT(rectangle3_weights[770]), .FEAT_THRES(feature_thresholds[770]), .FEAT_ABOVE(feature_aboves[770]), .FEAT_BELOW(feature_belows[770])) ac770(.scan_win(scan_win770), .scan_win_std_dev(scan_win_std_dev[770]), .feature_accum(feature_accums[770]));
  accum_calculator #(.RECT1_X(rectangle1_xs[771]), .RECT1_Y(rectangle1_ys[771]), .RECT1_WIDTH(rectangle1_widths[771]), .RECT1_HEIGHT(rectangle1_heights[771]), .RECT1_WEIGHT(rectangle1_weights[771]), .RECT2_X(rectangle2_xs[771]), .RECT2_Y(rectangle2_ys[771]), .RECT2_WIDTH(rectangle2_widths[771]), .RECT2_HEIGHT(rectangle2_heights[771]), .RECT2_WEIGHT(rectangle2_weights[771]), .RECT3_X(rectangle3_xs[771]), .RECT3_Y(rectangle3_ys[771]), .RECT3_WIDTH(rectangle3_widths[771]), .RECT3_HEIGHT(rectangle3_heights[771]), .RECT3_WEIGHT(rectangle3_weights[771]), .FEAT_THRES(feature_thresholds[771]), .FEAT_ABOVE(feature_aboves[771]), .FEAT_BELOW(feature_belows[771])) ac771(.scan_win(scan_win771), .scan_win_std_dev(scan_win_std_dev[771]), .feature_accum(feature_accums[771]));
  accum_calculator #(.RECT1_X(rectangle1_xs[772]), .RECT1_Y(rectangle1_ys[772]), .RECT1_WIDTH(rectangle1_widths[772]), .RECT1_HEIGHT(rectangle1_heights[772]), .RECT1_WEIGHT(rectangle1_weights[772]), .RECT2_X(rectangle2_xs[772]), .RECT2_Y(rectangle2_ys[772]), .RECT2_WIDTH(rectangle2_widths[772]), .RECT2_HEIGHT(rectangle2_heights[772]), .RECT2_WEIGHT(rectangle2_weights[772]), .RECT3_X(rectangle3_xs[772]), .RECT3_Y(rectangle3_ys[772]), .RECT3_WIDTH(rectangle3_widths[772]), .RECT3_HEIGHT(rectangle3_heights[772]), .RECT3_WEIGHT(rectangle3_weights[772]), .FEAT_THRES(feature_thresholds[772]), .FEAT_ABOVE(feature_aboves[772]), .FEAT_BELOW(feature_belows[772])) ac772(.scan_win(scan_win772), .scan_win_std_dev(scan_win_std_dev[772]), .feature_accum(feature_accums[772]));
  accum_calculator #(.RECT1_X(rectangle1_xs[773]), .RECT1_Y(rectangle1_ys[773]), .RECT1_WIDTH(rectangle1_widths[773]), .RECT1_HEIGHT(rectangle1_heights[773]), .RECT1_WEIGHT(rectangle1_weights[773]), .RECT2_X(rectangle2_xs[773]), .RECT2_Y(rectangle2_ys[773]), .RECT2_WIDTH(rectangle2_widths[773]), .RECT2_HEIGHT(rectangle2_heights[773]), .RECT2_WEIGHT(rectangle2_weights[773]), .RECT3_X(rectangle3_xs[773]), .RECT3_Y(rectangle3_ys[773]), .RECT3_WIDTH(rectangle3_widths[773]), .RECT3_HEIGHT(rectangle3_heights[773]), .RECT3_WEIGHT(rectangle3_weights[773]), .FEAT_THRES(feature_thresholds[773]), .FEAT_ABOVE(feature_aboves[773]), .FEAT_BELOW(feature_belows[773])) ac773(.scan_win(scan_win773), .scan_win_std_dev(scan_win_std_dev[773]), .feature_accum(feature_accums[773]));
  accum_calculator #(.RECT1_X(rectangle1_xs[774]), .RECT1_Y(rectangle1_ys[774]), .RECT1_WIDTH(rectangle1_widths[774]), .RECT1_HEIGHT(rectangle1_heights[774]), .RECT1_WEIGHT(rectangle1_weights[774]), .RECT2_X(rectangle2_xs[774]), .RECT2_Y(rectangle2_ys[774]), .RECT2_WIDTH(rectangle2_widths[774]), .RECT2_HEIGHT(rectangle2_heights[774]), .RECT2_WEIGHT(rectangle2_weights[774]), .RECT3_X(rectangle3_xs[774]), .RECT3_Y(rectangle3_ys[774]), .RECT3_WIDTH(rectangle3_widths[774]), .RECT3_HEIGHT(rectangle3_heights[774]), .RECT3_WEIGHT(rectangle3_weights[774]), .FEAT_THRES(feature_thresholds[774]), .FEAT_ABOVE(feature_aboves[774]), .FEAT_BELOW(feature_belows[774])) ac774(.scan_win(scan_win774), .scan_win_std_dev(scan_win_std_dev[774]), .feature_accum(feature_accums[774]));
  accum_calculator #(.RECT1_X(rectangle1_xs[775]), .RECT1_Y(rectangle1_ys[775]), .RECT1_WIDTH(rectangle1_widths[775]), .RECT1_HEIGHT(rectangle1_heights[775]), .RECT1_WEIGHT(rectangle1_weights[775]), .RECT2_X(rectangle2_xs[775]), .RECT2_Y(rectangle2_ys[775]), .RECT2_WIDTH(rectangle2_widths[775]), .RECT2_HEIGHT(rectangle2_heights[775]), .RECT2_WEIGHT(rectangle2_weights[775]), .RECT3_X(rectangle3_xs[775]), .RECT3_Y(rectangle3_ys[775]), .RECT3_WIDTH(rectangle3_widths[775]), .RECT3_HEIGHT(rectangle3_heights[775]), .RECT3_WEIGHT(rectangle3_weights[775]), .FEAT_THRES(feature_thresholds[775]), .FEAT_ABOVE(feature_aboves[775]), .FEAT_BELOW(feature_belows[775])) ac775(.scan_win(scan_win775), .scan_win_std_dev(scan_win_std_dev[775]), .feature_accum(feature_accums[775]));
  accum_calculator #(.RECT1_X(rectangle1_xs[776]), .RECT1_Y(rectangle1_ys[776]), .RECT1_WIDTH(rectangle1_widths[776]), .RECT1_HEIGHT(rectangle1_heights[776]), .RECT1_WEIGHT(rectangle1_weights[776]), .RECT2_X(rectangle2_xs[776]), .RECT2_Y(rectangle2_ys[776]), .RECT2_WIDTH(rectangle2_widths[776]), .RECT2_HEIGHT(rectangle2_heights[776]), .RECT2_WEIGHT(rectangle2_weights[776]), .RECT3_X(rectangle3_xs[776]), .RECT3_Y(rectangle3_ys[776]), .RECT3_WIDTH(rectangle3_widths[776]), .RECT3_HEIGHT(rectangle3_heights[776]), .RECT3_WEIGHT(rectangle3_weights[776]), .FEAT_THRES(feature_thresholds[776]), .FEAT_ABOVE(feature_aboves[776]), .FEAT_BELOW(feature_belows[776])) ac776(.scan_win(scan_win776), .scan_win_std_dev(scan_win_std_dev[776]), .feature_accum(feature_accums[776]));
  accum_calculator #(.RECT1_X(rectangle1_xs[777]), .RECT1_Y(rectangle1_ys[777]), .RECT1_WIDTH(rectangle1_widths[777]), .RECT1_HEIGHT(rectangle1_heights[777]), .RECT1_WEIGHT(rectangle1_weights[777]), .RECT2_X(rectangle2_xs[777]), .RECT2_Y(rectangle2_ys[777]), .RECT2_WIDTH(rectangle2_widths[777]), .RECT2_HEIGHT(rectangle2_heights[777]), .RECT2_WEIGHT(rectangle2_weights[777]), .RECT3_X(rectangle3_xs[777]), .RECT3_Y(rectangle3_ys[777]), .RECT3_WIDTH(rectangle3_widths[777]), .RECT3_HEIGHT(rectangle3_heights[777]), .RECT3_WEIGHT(rectangle3_weights[777]), .FEAT_THRES(feature_thresholds[777]), .FEAT_ABOVE(feature_aboves[777]), .FEAT_BELOW(feature_belows[777])) ac777(.scan_win(scan_win777), .scan_win_std_dev(scan_win_std_dev[777]), .feature_accum(feature_accums[777]));
  accum_calculator #(.RECT1_X(rectangle1_xs[778]), .RECT1_Y(rectangle1_ys[778]), .RECT1_WIDTH(rectangle1_widths[778]), .RECT1_HEIGHT(rectangle1_heights[778]), .RECT1_WEIGHT(rectangle1_weights[778]), .RECT2_X(rectangle2_xs[778]), .RECT2_Y(rectangle2_ys[778]), .RECT2_WIDTH(rectangle2_widths[778]), .RECT2_HEIGHT(rectangle2_heights[778]), .RECT2_WEIGHT(rectangle2_weights[778]), .RECT3_X(rectangle3_xs[778]), .RECT3_Y(rectangle3_ys[778]), .RECT3_WIDTH(rectangle3_widths[778]), .RECT3_HEIGHT(rectangle3_heights[778]), .RECT3_WEIGHT(rectangle3_weights[778]), .FEAT_THRES(feature_thresholds[778]), .FEAT_ABOVE(feature_aboves[778]), .FEAT_BELOW(feature_belows[778])) ac778(.scan_win(scan_win778), .scan_win_std_dev(scan_win_std_dev[778]), .feature_accum(feature_accums[778]));
  accum_calculator #(.RECT1_X(rectangle1_xs[779]), .RECT1_Y(rectangle1_ys[779]), .RECT1_WIDTH(rectangle1_widths[779]), .RECT1_HEIGHT(rectangle1_heights[779]), .RECT1_WEIGHT(rectangle1_weights[779]), .RECT2_X(rectangle2_xs[779]), .RECT2_Y(rectangle2_ys[779]), .RECT2_WIDTH(rectangle2_widths[779]), .RECT2_HEIGHT(rectangle2_heights[779]), .RECT2_WEIGHT(rectangle2_weights[779]), .RECT3_X(rectangle3_xs[779]), .RECT3_Y(rectangle3_ys[779]), .RECT3_WIDTH(rectangle3_widths[779]), .RECT3_HEIGHT(rectangle3_heights[779]), .RECT3_WEIGHT(rectangle3_weights[779]), .FEAT_THRES(feature_thresholds[779]), .FEAT_ABOVE(feature_aboves[779]), .FEAT_BELOW(feature_belows[779])) ac779(.scan_win(scan_win779), .scan_win_std_dev(scan_win_std_dev[779]), .feature_accum(feature_accums[779]));
  accum_calculator #(.RECT1_X(rectangle1_xs[780]), .RECT1_Y(rectangle1_ys[780]), .RECT1_WIDTH(rectangle1_widths[780]), .RECT1_HEIGHT(rectangle1_heights[780]), .RECT1_WEIGHT(rectangle1_weights[780]), .RECT2_X(rectangle2_xs[780]), .RECT2_Y(rectangle2_ys[780]), .RECT2_WIDTH(rectangle2_widths[780]), .RECT2_HEIGHT(rectangle2_heights[780]), .RECT2_WEIGHT(rectangle2_weights[780]), .RECT3_X(rectangle3_xs[780]), .RECT3_Y(rectangle3_ys[780]), .RECT3_WIDTH(rectangle3_widths[780]), .RECT3_HEIGHT(rectangle3_heights[780]), .RECT3_WEIGHT(rectangle3_weights[780]), .FEAT_THRES(feature_thresholds[780]), .FEAT_ABOVE(feature_aboves[780]), .FEAT_BELOW(feature_belows[780])) ac780(.scan_win(scan_win780), .scan_win_std_dev(scan_win_std_dev[780]), .feature_accum(feature_accums[780]));
  accum_calculator #(.RECT1_X(rectangle1_xs[781]), .RECT1_Y(rectangle1_ys[781]), .RECT1_WIDTH(rectangle1_widths[781]), .RECT1_HEIGHT(rectangle1_heights[781]), .RECT1_WEIGHT(rectangle1_weights[781]), .RECT2_X(rectangle2_xs[781]), .RECT2_Y(rectangle2_ys[781]), .RECT2_WIDTH(rectangle2_widths[781]), .RECT2_HEIGHT(rectangle2_heights[781]), .RECT2_WEIGHT(rectangle2_weights[781]), .RECT3_X(rectangle3_xs[781]), .RECT3_Y(rectangle3_ys[781]), .RECT3_WIDTH(rectangle3_widths[781]), .RECT3_HEIGHT(rectangle3_heights[781]), .RECT3_WEIGHT(rectangle3_weights[781]), .FEAT_THRES(feature_thresholds[781]), .FEAT_ABOVE(feature_aboves[781]), .FEAT_BELOW(feature_belows[781])) ac781(.scan_win(scan_win781), .scan_win_std_dev(scan_win_std_dev[781]), .feature_accum(feature_accums[781]));
  accum_calculator #(.RECT1_X(rectangle1_xs[782]), .RECT1_Y(rectangle1_ys[782]), .RECT1_WIDTH(rectangle1_widths[782]), .RECT1_HEIGHT(rectangle1_heights[782]), .RECT1_WEIGHT(rectangle1_weights[782]), .RECT2_X(rectangle2_xs[782]), .RECT2_Y(rectangle2_ys[782]), .RECT2_WIDTH(rectangle2_widths[782]), .RECT2_HEIGHT(rectangle2_heights[782]), .RECT2_WEIGHT(rectangle2_weights[782]), .RECT3_X(rectangle3_xs[782]), .RECT3_Y(rectangle3_ys[782]), .RECT3_WIDTH(rectangle3_widths[782]), .RECT3_HEIGHT(rectangle3_heights[782]), .RECT3_WEIGHT(rectangle3_weights[782]), .FEAT_THRES(feature_thresholds[782]), .FEAT_ABOVE(feature_aboves[782]), .FEAT_BELOW(feature_belows[782])) ac782(.scan_win(scan_win782), .scan_win_std_dev(scan_win_std_dev[782]), .feature_accum(feature_accums[782]));
  accum_calculator #(.RECT1_X(rectangle1_xs[783]), .RECT1_Y(rectangle1_ys[783]), .RECT1_WIDTH(rectangle1_widths[783]), .RECT1_HEIGHT(rectangle1_heights[783]), .RECT1_WEIGHT(rectangle1_weights[783]), .RECT2_X(rectangle2_xs[783]), .RECT2_Y(rectangle2_ys[783]), .RECT2_WIDTH(rectangle2_widths[783]), .RECT2_HEIGHT(rectangle2_heights[783]), .RECT2_WEIGHT(rectangle2_weights[783]), .RECT3_X(rectangle3_xs[783]), .RECT3_Y(rectangle3_ys[783]), .RECT3_WIDTH(rectangle3_widths[783]), .RECT3_HEIGHT(rectangle3_heights[783]), .RECT3_WEIGHT(rectangle3_weights[783]), .FEAT_THRES(feature_thresholds[783]), .FEAT_ABOVE(feature_aboves[783]), .FEAT_BELOW(feature_belows[783])) ac783(.scan_win(scan_win783), .scan_win_std_dev(scan_win_std_dev[783]), .feature_accum(feature_accums[783]));
  accum_calculator #(.RECT1_X(rectangle1_xs[784]), .RECT1_Y(rectangle1_ys[784]), .RECT1_WIDTH(rectangle1_widths[784]), .RECT1_HEIGHT(rectangle1_heights[784]), .RECT1_WEIGHT(rectangle1_weights[784]), .RECT2_X(rectangle2_xs[784]), .RECT2_Y(rectangle2_ys[784]), .RECT2_WIDTH(rectangle2_widths[784]), .RECT2_HEIGHT(rectangle2_heights[784]), .RECT2_WEIGHT(rectangle2_weights[784]), .RECT3_X(rectangle3_xs[784]), .RECT3_Y(rectangle3_ys[784]), .RECT3_WIDTH(rectangle3_widths[784]), .RECT3_HEIGHT(rectangle3_heights[784]), .RECT3_WEIGHT(rectangle3_weights[784]), .FEAT_THRES(feature_thresholds[784]), .FEAT_ABOVE(feature_aboves[784]), .FEAT_BELOW(feature_belows[784])) ac784(.scan_win(scan_win784), .scan_win_std_dev(scan_win_std_dev[784]), .feature_accum(feature_accums[784]));
  accum_calculator #(.RECT1_X(rectangle1_xs[785]), .RECT1_Y(rectangle1_ys[785]), .RECT1_WIDTH(rectangle1_widths[785]), .RECT1_HEIGHT(rectangle1_heights[785]), .RECT1_WEIGHT(rectangle1_weights[785]), .RECT2_X(rectangle2_xs[785]), .RECT2_Y(rectangle2_ys[785]), .RECT2_WIDTH(rectangle2_widths[785]), .RECT2_HEIGHT(rectangle2_heights[785]), .RECT2_WEIGHT(rectangle2_weights[785]), .RECT3_X(rectangle3_xs[785]), .RECT3_Y(rectangle3_ys[785]), .RECT3_WIDTH(rectangle3_widths[785]), .RECT3_HEIGHT(rectangle3_heights[785]), .RECT3_WEIGHT(rectangle3_weights[785]), .FEAT_THRES(feature_thresholds[785]), .FEAT_ABOVE(feature_aboves[785]), .FEAT_BELOW(feature_belows[785])) ac785(.scan_win(scan_win785), .scan_win_std_dev(scan_win_std_dev[785]), .feature_accum(feature_accums[785]));
  accum_calculator #(.RECT1_X(rectangle1_xs[786]), .RECT1_Y(rectangle1_ys[786]), .RECT1_WIDTH(rectangle1_widths[786]), .RECT1_HEIGHT(rectangle1_heights[786]), .RECT1_WEIGHT(rectangle1_weights[786]), .RECT2_X(rectangle2_xs[786]), .RECT2_Y(rectangle2_ys[786]), .RECT2_WIDTH(rectangle2_widths[786]), .RECT2_HEIGHT(rectangle2_heights[786]), .RECT2_WEIGHT(rectangle2_weights[786]), .RECT3_X(rectangle3_xs[786]), .RECT3_Y(rectangle3_ys[786]), .RECT3_WIDTH(rectangle3_widths[786]), .RECT3_HEIGHT(rectangle3_heights[786]), .RECT3_WEIGHT(rectangle3_weights[786]), .FEAT_THRES(feature_thresholds[786]), .FEAT_ABOVE(feature_aboves[786]), .FEAT_BELOW(feature_belows[786])) ac786(.scan_win(scan_win786), .scan_win_std_dev(scan_win_std_dev[786]), .feature_accum(feature_accums[786]));
  accum_calculator #(.RECT1_X(rectangle1_xs[787]), .RECT1_Y(rectangle1_ys[787]), .RECT1_WIDTH(rectangle1_widths[787]), .RECT1_HEIGHT(rectangle1_heights[787]), .RECT1_WEIGHT(rectangle1_weights[787]), .RECT2_X(rectangle2_xs[787]), .RECT2_Y(rectangle2_ys[787]), .RECT2_WIDTH(rectangle2_widths[787]), .RECT2_HEIGHT(rectangle2_heights[787]), .RECT2_WEIGHT(rectangle2_weights[787]), .RECT3_X(rectangle3_xs[787]), .RECT3_Y(rectangle3_ys[787]), .RECT3_WIDTH(rectangle3_widths[787]), .RECT3_HEIGHT(rectangle3_heights[787]), .RECT3_WEIGHT(rectangle3_weights[787]), .FEAT_THRES(feature_thresholds[787]), .FEAT_ABOVE(feature_aboves[787]), .FEAT_BELOW(feature_belows[787])) ac787(.scan_win(scan_win787), .scan_win_std_dev(scan_win_std_dev[787]), .feature_accum(feature_accums[787]));
  accum_calculator #(.RECT1_X(rectangle1_xs[788]), .RECT1_Y(rectangle1_ys[788]), .RECT1_WIDTH(rectangle1_widths[788]), .RECT1_HEIGHT(rectangle1_heights[788]), .RECT1_WEIGHT(rectangle1_weights[788]), .RECT2_X(rectangle2_xs[788]), .RECT2_Y(rectangle2_ys[788]), .RECT2_WIDTH(rectangle2_widths[788]), .RECT2_HEIGHT(rectangle2_heights[788]), .RECT2_WEIGHT(rectangle2_weights[788]), .RECT3_X(rectangle3_xs[788]), .RECT3_Y(rectangle3_ys[788]), .RECT3_WIDTH(rectangle3_widths[788]), .RECT3_HEIGHT(rectangle3_heights[788]), .RECT3_WEIGHT(rectangle3_weights[788]), .FEAT_THRES(feature_thresholds[788]), .FEAT_ABOVE(feature_aboves[788]), .FEAT_BELOW(feature_belows[788])) ac788(.scan_win(scan_win788), .scan_win_std_dev(scan_win_std_dev[788]), .feature_accum(feature_accums[788]));
  accum_calculator #(.RECT1_X(rectangle1_xs[789]), .RECT1_Y(rectangle1_ys[789]), .RECT1_WIDTH(rectangle1_widths[789]), .RECT1_HEIGHT(rectangle1_heights[789]), .RECT1_WEIGHT(rectangle1_weights[789]), .RECT2_X(rectangle2_xs[789]), .RECT2_Y(rectangle2_ys[789]), .RECT2_WIDTH(rectangle2_widths[789]), .RECT2_HEIGHT(rectangle2_heights[789]), .RECT2_WEIGHT(rectangle2_weights[789]), .RECT3_X(rectangle3_xs[789]), .RECT3_Y(rectangle3_ys[789]), .RECT3_WIDTH(rectangle3_widths[789]), .RECT3_HEIGHT(rectangle3_heights[789]), .RECT3_WEIGHT(rectangle3_weights[789]), .FEAT_THRES(feature_thresholds[789]), .FEAT_ABOVE(feature_aboves[789]), .FEAT_BELOW(feature_belows[789])) ac789(.scan_win(scan_win789), .scan_win_std_dev(scan_win_std_dev[789]), .feature_accum(feature_accums[789]));
  accum_calculator #(.RECT1_X(rectangle1_xs[790]), .RECT1_Y(rectangle1_ys[790]), .RECT1_WIDTH(rectangle1_widths[790]), .RECT1_HEIGHT(rectangle1_heights[790]), .RECT1_WEIGHT(rectangle1_weights[790]), .RECT2_X(rectangle2_xs[790]), .RECT2_Y(rectangle2_ys[790]), .RECT2_WIDTH(rectangle2_widths[790]), .RECT2_HEIGHT(rectangle2_heights[790]), .RECT2_WEIGHT(rectangle2_weights[790]), .RECT3_X(rectangle3_xs[790]), .RECT3_Y(rectangle3_ys[790]), .RECT3_WIDTH(rectangle3_widths[790]), .RECT3_HEIGHT(rectangle3_heights[790]), .RECT3_WEIGHT(rectangle3_weights[790]), .FEAT_THRES(feature_thresholds[790]), .FEAT_ABOVE(feature_aboves[790]), .FEAT_BELOW(feature_belows[790])) ac790(.scan_win(scan_win790), .scan_win_std_dev(scan_win_std_dev[790]), .feature_accum(feature_accums[790]));
  accum_calculator #(.RECT1_X(rectangle1_xs[791]), .RECT1_Y(rectangle1_ys[791]), .RECT1_WIDTH(rectangle1_widths[791]), .RECT1_HEIGHT(rectangle1_heights[791]), .RECT1_WEIGHT(rectangle1_weights[791]), .RECT2_X(rectangle2_xs[791]), .RECT2_Y(rectangle2_ys[791]), .RECT2_WIDTH(rectangle2_widths[791]), .RECT2_HEIGHT(rectangle2_heights[791]), .RECT2_WEIGHT(rectangle2_weights[791]), .RECT3_X(rectangle3_xs[791]), .RECT3_Y(rectangle3_ys[791]), .RECT3_WIDTH(rectangle3_widths[791]), .RECT3_HEIGHT(rectangle3_heights[791]), .RECT3_WEIGHT(rectangle3_weights[791]), .FEAT_THRES(feature_thresholds[791]), .FEAT_ABOVE(feature_aboves[791]), .FEAT_BELOW(feature_belows[791])) ac791(.scan_win(scan_win791), .scan_win_std_dev(scan_win_std_dev[791]), .feature_accum(feature_accums[791]));
  accum_calculator #(.RECT1_X(rectangle1_xs[792]), .RECT1_Y(rectangle1_ys[792]), .RECT1_WIDTH(rectangle1_widths[792]), .RECT1_HEIGHT(rectangle1_heights[792]), .RECT1_WEIGHT(rectangle1_weights[792]), .RECT2_X(rectangle2_xs[792]), .RECT2_Y(rectangle2_ys[792]), .RECT2_WIDTH(rectangle2_widths[792]), .RECT2_HEIGHT(rectangle2_heights[792]), .RECT2_WEIGHT(rectangle2_weights[792]), .RECT3_X(rectangle3_xs[792]), .RECT3_Y(rectangle3_ys[792]), .RECT3_WIDTH(rectangle3_widths[792]), .RECT3_HEIGHT(rectangle3_heights[792]), .RECT3_WEIGHT(rectangle3_weights[792]), .FEAT_THRES(feature_thresholds[792]), .FEAT_ABOVE(feature_aboves[792]), .FEAT_BELOW(feature_belows[792])) ac792(.scan_win(scan_win792), .scan_win_std_dev(scan_win_std_dev[792]), .feature_accum(feature_accums[792]));
  accum_calculator #(.RECT1_X(rectangle1_xs[793]), .RECT1_Y(rectangle1_ys[793]), .RECT1_WIDTH(rectangle1_widths[793]), .RECT1_HEIGHT(rectangle1_heights[793]), .RECT1_WEIGHT(rectangle1_weights[793]), .RECT2_X(rectangle2_xs[793]), .RECT2_Y(rectangle2_ys[793]), .RECT2_WIDTH(rectangle2_widths[793]), .RECT2_HEIGHT(rectangle2_heights[793]), .RECT2_WEIGHT(rectangle2_weights[793]), .RECT3_X(rectangle3_xs[793]), .RECT3_Y(rectangle3_ys[793]), .RECT3_WIDTH(rectangle3_widths[793]), .RECT3_HEIGHT(rectangle3_heights[793]), .RECT3_WEIGHT(rectangle3_weights[793]), .FEAT_THRES(feature_thresholds[793]), .FEAT_ABOVE(feature_aboves[793]), .FEAT_BELOW(feature_belows[793])) ac793(.scan_win(scan_win793), .scan_win_std_dev(scan_win_std_dev[793]), .feature_accum(feature_accums[793]));
  accum_calculator #(.RECT1_X(rectangle1_xs[794]), .RECT1_Y(rectangle1_ys[794]), .RECT1_WIDTH(rectangle1_widths[794]), .RECT1_HEIGHT(rectangle1_heights[794]), .RECT1_WEIGHT(rectangle1_weights[794]), .RECT2_X(rectangle2_xs[794]), .RECT2_Y(rectangle2_ys[794]), .RECT2_WIDTH(rectangle2_widths[794]), .RECT2_HEIGHT(rectangle2_heights[794]), .RECT2_WEIGHT(rectangle2_weights[794]), .RECT3_X(rectangle3_xs[794]), .RECT3_Y(rectangle3_ys[794]), .RECT3_WIDTH(rectangle3_widths[794]), .RECT3_HEIGHT(rectangle3_heights[794]), .RECT3_WEIGHT(rectangle3_weights[794]), .FEAT_THRES(feature_thresholds[794]), .FEAT_ABOVE(feature_aboves[794]), .FEAT_BELOW(feature_belows[794])) ac794(.scan_win(scan_win794), .scan_win_std_dev(scan_win_std_dev[794]), .feature_accum(feature_accums[794]));
  accum_calculator #(.RECT1_X(rectangle1_xs[795]), .RECT1_Y(rectangle1_ys[795]), .RECT1_WIDTH(rectangle1_widths[795]), .RECT1_HEIGHT(rectangle1_heights[795]), .RECT1_WEIGHT(rectangle1_weights[795]), .RECT2_X(rectangle2_xs[795]), .RECT2_Y(rectangle2_ys[795]), .RECT2_WIDTH(rectangle2_widths[795]), .RECT2_HEIGHT(rectangle2_heights[795]), .RECT2_WEIGHT(rectangle2_weights[795]), .RECT3_X(rectangle3_xs[795]), .RECT3_Y(rectangle3_ys[795]), .RECT3_WIDTH(rectangle3_widths[795]), .RECT3_HEIGHT(rectangle3_heights[795]), .RECT3_WEIGHT(rectangle3_weights[795]), .FEAT_THRES(feature_thresholds[795]), .FEAT_ABOVE(feature_aboves[795]), .FEAT_BELOW(feature_belows[795])) ac795(.scan_win(scan_win795), .scan_win_std_dev(scan_win_std_dev[795]), .feature_accum(feature_accums[795]));
  accum_calculator #(.RECT1_X(rectangle1_xs[796]), .RECT1_Y(rectangle1_ys[796]), .RECT1_WIDTH(rectangle1_widths[796]), .RECT1_HEIGHT(rectangle1_heights[796]), .RECT1_WEIGHT(rectangle1_weights[796]), .RECT2_X(rectangle2_xs[796]), .RECT2_Y(rectangle2_ys[796]), .RECT2_WIDTH(rectangle2_widths[796]), .RECT2_HEIGHT(rectangle2_heights[796]), .RECT2_WEIGHT(rectangle2_weights[796]), .RECT3_X(rectangle3_xs[796]), .RECT3_Y(rectangle3_ys[796]), .RECT3_WIDTH(rectangle3_widths[796]), .RECT3_HEIGHT(rectangle3_heights[796]), .RECT3_WEIGHT(rectangle3_weights[796]), .FEAT_THRES(feature_thresholds[796]), .FEAT_ABOVE(feature_aboves[796]), .FEAT_BELOW(feature_belows[796])) ac796(.scan_win(scan_win796), .scan_win_std_dev(scan_win_std_dev[796]), .feature_accum(feature_accums[796]));
  accum_calculator #(.RECT1_X(rectangle1_xs[797]), .RECT1_Y(rectangle1_ys[797]), .RECT1_WIDTH(rectangle1_widths[797]), .RECT1_HEIGHT(rectangle1_heights[797]), .RECT1_WEIGHT(rectangle1_weights[797]), .RECT2_X(rectangle2_xs[797]), .RECT2_Y(rectangle2_ys[797]), .RECT2_WIDTH(rectangle2_widths[797]), .RECT2_HEIGHT(rectangle2_heights[797]), .RECT2_WEIGHT(rectangle2_weights[797]), .RECT3_X(rectangle3_xs[797]), .RECT3_Y(rectangle3_ys[797]), .RECT3_WIDTH(rectangle3_widths[797]), .RECT3_HEIGHT(rectangle3_heights[797]), .RECT3_WEIGHT(rectangle3_weights[797]), .FEAT_THRES(feature_thresholds[797]), .FEAT_ABOVE(feature_aboves[797]), .FEAT_BELOW(feature_belows[797])) ac797(.scan_win(scan_win797), .scan_win_std_dev(scan_win_std_dev[797]), .feature_accum(feature_accums[797]));
  accum_calculator #(.RECT1_X(rectangle1_xs[798]), .RECT1_Y(rectangle1_ys[798]), .RECT1_WIDTH(rectangle1_widths[798]), .RECT1_HEIGHT(rectangle1_heights[798]), .RECT1_WEIGHT(rectangle1_weights[798]), .RECT2_X(rectangle2_xs[798]), .RECT2_Y(rectangle2_ys[798]), .RECT2_WIDTH(rectangle2_widths[798]), .RECT2_HEIGHT(rectangle2_heights[798]), .RECT2_WEIGHT(rectangle2_weights[798]), .RECT3_X(rectangle3_xs[798]), .RECT3_Y(rectangle3_ys[798]), .RECT3_WIDTH(rectangle3_widths[798]), .RECT3_HEIGHT(rectangle3_heights[798]), .RECT3_WEIGHT(rectangle3_weights[798]), .FEAT_THRES(feature_thresholds[798]), .FEAT_ABOVE(feature_aboves[798]), .FEAT_BELOW(feature_belows[798])) ac798(.scan_win(scan_win798), .scan_win_std_dev(scan_win_std_dev[798]), .feature_accum(feature_accums[798]));
  accum_calculator #(.RECT1_X(rectangle1_xs[799]), .RECT1_Y(rectangle1_ys[799]), .RECT1_WIDTH(rectangle1_widths[799]), .RECT1_HEIGHT(rectangle1_heights[799]), .RECT1_WEIGHT(rectangle1_weights[799]), .RECT2_X(rectangle2_xs[799]), .RECT2_Y(rectangle2_ys[799]), .RECT2_WIDTH(rectangle2_widths[799]), .RECT2_HEIGHT(rectangle2_heights[799]), .RECT2_WEIGHT(rectangle2_weights[799]), .RECT3_X(rectangle3_xs[799]), .RECT3_Y(rectangle3_ys[799]), .RECT3_WIDTH(rectangle3_widths[799]), .RECT3_HEIGHT(rectangle3_heights[799]), .RECT3_WEIGHT(rectangle3_weights[799]), .FEAT_THRES(feature_thresholds[799]), .FEAT_ABOVE(feature_aboves[799]), .FEAT_BELOW(feature_belows[799])) ac799(.scan_win(scan_win799), .scan_win_std_dev(scan_win_std_dev[799]), .feature_accum(feature_accums[799]));
  accum_calculator #(.RECT1_X(rectangle1_xs[800]), .RECT1_Y(rectangle1_ys[800]), .RECT1_WIDTH(rectangle1_widths[800]), .RECT1_HEIGHT(rectangle1_heights[800]), .RECT1_WEIGHT(rectangle1_weights[800]), .RECT2_X(rectangle2_xs[800]), .RECT2_Y(rectangle2_ys[800]), .RECT2_WIDTH(rectangle2_widths[800]), .RECT2_HEIGHT(rectangle2_heights[800]), .RECT2_WEIGHT(rectangle2_weights[800]), .RECT3_X(rectangle3_xs[800]), .RECT3_Y(rectangle3_ys[800]), .RECT3_WIDTH(rectangle3_widths[800]), .RECT3_HEIGHT(rectangle3_heights[800]), .RECT3_WEIGHT(rectangle3_weights[800]), .FEAT_THRES(feature_thresholds[800]), .FEAT_ABOVE(feature_aboves[800]), .FEAT_BELOW(feature_belows[800])) ac800(.scan_win(scan_win800), .scan_win_std_dev(scan_win_std_dev[800]), .feature_accum(feature_accums[800]));
  accum_calculator #(.RECT1_X(rectangle1_xs[801]), .RECT1_Y(rectangle1_ys[801]), .RECT1_WIDTH(rectangle1_widths[801]), .RECT1_HEIGHT(rectangle1_heights[801]), .RECT1_WEIGHT(rectangle1_weights[801]), .RECT2_X(rectangle2_xs[801]), .RECT2_Y(rectangle2_ys[801]), .RECT2_WIDTH(rectangle2_widths[801]), .RECT2_HEIGHT(rectangle2_heights[801]), .RECT2_WEIGHT(rectangle2_weights[801]), .RECT3_X(rectangle3_xs[801]), .RECT3_Y(rectangle3_ys[801]), .RECT3_WIDTH(rectangle3_widths[801]), .RECT3_HEIGHT(rectangle3_heights[801]), .RECT3_WEIGHT(rectangle3_weights[801]), .FEAT_THRES(feature_thresholds[801]), .FEAT_ABOVE(feature_aboves[801]), .FEAT_BELOW(feature_belows[801])) ac801(.scan_win(scan_win801), .scan_win_std_dev(scan_win_std_dev[801]), .feature_accum(feature_accums[801]));
  accum_calculator #(.RECT1_X(rectangle1_xs[802]), .RECT1_Y(rectangle1_ys[802]), .RECT1_WIDTH(rectangle1_widths[802]), .RECT1_HEIGHT(rectangle1_heights[802]), .RECT1_WEIGHT(rectangle1_weights[802]), .RECT2_X(rectangle2_xs[802]), .RECT2_Y(rectangle2_ys[802]), .RECT2_WIDTH(rectangle2_widths[802]), .RECT2_HEIGHT(rectangle2_heights[802]), .RECT2_WEIGHT(rectangle2_weights[802]), .RECT3_X(rectangle3_xs[802]), .RECT3_Y(rectangle3_ys[802]), .RECT3_WIDTH(rectangle3_widths[802]), .RECT3_HEIGHT(rectangle3_heights[802]), .RECT3_WEIGHT(rectangle3_weights[802]), .FEAT_THRES(feature_thresholds[802]), .FEAT_ABOVE(feature_aboves[802]), .FEAT_BELOW(feature_belows[802])) ac802(.scan_win(scan_win802), .scan_win_std_dev(scan_win_std_dev[802]), .feature_accum(feature_accums[802]));
  accum_calculator #(.RECT1_X(rectangle1_xs[803]), .RECT1_Y(rectangle1_ys[803]), .RECT1_WIDTH(rectangle1_widths[803]), .RECT1_HEIGHT(rectangle1_heights[803]), .RECT1_WEIGHT(rectangle1_weights[803]), .RECT2_X(rectangle2_xs[803]), .RECT2_Y(rectangle2_ys[803]), .RECT2_WIDTH(rectangle2_widths[803]), .RECT2_HEIGHT(rectangle2_heights[803]), .RECT2_WEIGHT(rectangle2_weights[803]), .RECT3_X(rectangle3_xs[803]), .RECT3_Y(rectangle3_ys[803]), .RECT3_WIDTH(rectangle3_widths[803]), .RECT3_HEIGHT(rectangle3_heights[803]), .RECT3_WEIGHT(rectangle3_weights[803]), .FEAT_THRES(feature_thresholds[803]), .FEAT_ABOVE(feature_aboves[803]), .FEAT_BELOW(feature_belows[803])) ac803(.scan_win(scan_win803), .scan_win_std_dev(scan_win_std_dev[803]), .feature_accum(feature_accums[803]));
  accum_calculator #(.RECT1_X(rectangle1_xs[804]), .RECT1_Y(rectangle1_ys[804]), .RECT1_WIDTH(rectangle1_widths[804]), .RECT1_HEIGHT(rectangle1_heights[804]), .RECT1_WEIGHT(rectangle1_weights[804]), .RECT2_X(rectangle2_xs[804]), .RECT2_Y(rectangle2_ys[804]), .RECT2_WIDTH(rectangle2_widths[804]), .RECT2_HEIGHT(rectangle2_heights[804]), .RECT2_WEIGHT(rectangle2_weights[804]), .RECT3_X(rectangle3_xs[804]), .RECT3_Y(rectangle3_ys[804]), .RECT3_WIDTH(rectangle3_widths[804]), .RECT3_HEIGHT(rectangle3_heights[804]), .RECT3_WEIGHT(rectangle3_weights[804]), .FEAT_THRES(feature_thresholds[804]), .FEAT_ABOVE(feature_aboves[804]), .FEAT_BELOW(feature_belows[804])) ac804(.scan_win(scan_win804), .scan_win_std_dev(scan_win_std_dev[804]), .feature_accum(feature_accums[804]));
  accum_calculator #(.RECT1_X(rectangle1_xs[805]), .RECT1_Y(rectangle1_ys[805]), .RECT1_WIDTH(rectangle1_widths[805]), .RECT1_HEIGHT(rectangle1_heights[805]), .RECT1_WEIGHT(rectangle1_weights[805]), .RECT2_X(rectangle2_xs[805]), .RECT2_Y(rectangle2_ys[805]), .RECT2_WIDTH(rectangle2_widths[805]), .RECT2_HEIGHT(rectangle2_heights[805]), .RECT2_WEIGHT(rectangle2_weights[805]), .RECT3_X(rectangle3_xs[805]), .RECT3_Y(rectangle3_ys[805]), .RECT3_WIDTH(rectangle3_widths[805]), .RECT3_HEIGHT(rectangle3_heights[805]), .RECT3_WEIGHT(rectangle3_weights[805]), .FEAT_THRES(feature_thresholds[805]), .FEAT_ABOVE(feature_aboves[805]), .FEAT_BELOW(feature_belows[805])) ac805(.scan_win(scan_win805), .scan_win_std_dev(scan_win_std_dev[805]), .feature_accum(feature_accums[805]));
  accum_calculator #(.RECT1_X(rectangle1_xs[806]), .RECT1_Y(rectangle1_ys[806]), .RECT1_WIDTH(rectangle1_widths[806]), .RECT1_HEIGHT(rectangle1_heights[806]), .RECT1_WEIGHT(rectangle1_weights[806]), .RECT2_X(rectangle2_xs[806]), .RECT2_Y(rectangle2_ys[806]), .RECT2_WIDTH(rectangle2_widths[806]), .RECT2_HEIGHT(rectangle2_heights[806]), .RECT2_WEIGHT(rectangle2_weights[806]), .RECT3_X(rectangle3_xs[806]), .RECT3_Y(rectangle3_ys[806]), .RECT3_WIDTH(rectangle3_widths[806]), .RECT3_HEIGHT(rectangle3_heights[806]), .RECT3_WEIGHT(rectangle3_weights[806]), .FEAT_THRES(feature_thresholds[806]), .FEAT_ABOVE(feature_aboves[806]), .FEAT_BELOW(feature_belows[806])) ac806(.scan_win(scan_win806), .scan_win_std_dev(scan_win_std_dev[806]), .feature_accum(feature_accums[806]));
  accum_calculator #(.RECT1_X(rectangle1_xs[807]), .RECT1_Y(rectangle1_ys[807]), .RECT1_WIDTH(rectangle1_widths[807]), .RECT1_HEIGHT(rectangle1_heights[807]), .RECT1_WEIGHT(rectangle1_weights[807]), .RECT2_X(rectangle2_xs[807]), .RECT2_Y(rectangle2_ys[807]), .RECT2_WIDTH(rectangle2_widths[807]), .RECT2_HEIGHT(rectangle2_heights[807]), .RECT2_WEIGHT(rectangle2_weights[807]), .RECT3_X(rectangle3_xs[807]), .RECT3_Y(rectangle3_ys[807]), .RECT3_WIDTH(rectangle3_widths[807]), .RECT3_HEIGHT(rectangle3_heights[807]), .RECT3_WEIGHT(rectangle3_weights[807]), .FEAT_THRES(feature_thresholds[807]), .FEAT_ABOVE(feature_aboves[807]), .FEAT_BELOW(feature_belows[807])) ac807(.scan_win(scan_win807), .scan_win_std_dev(scan_win_std_dev[807]), .feature_accum(feature_accums[807]));
  accum_calculator #(.RECT1_X(rectangle1_xs[808]), .RECT1_Y(rectangle1_ys[808]), .RECT1_WIDTH(rectangle1_widths[808]), .RECT1_HEIGHT(rectangle1_heights[808]), .RECT1_WEIGHT(rectangle1_weights[808]), .RECT2_X(rectangle2_xs[808]), .RECT2_Y(rectangle2_ys[808]), .RECT2_WIDTH(rectangle2_widths[808]), .RECT2_HEIGHT(rectangle2_heights[808]), .RECT2_WEIGHT(rectangle2_weights[808]), .RECT3_X(rectangle3_xs[808]), .RECT3_Y(rectangle3_ys[808]), .RECT3_WIDTH(rectangle3_widths[808]), .RECT3_HEIGHT(rectangle3_heights[808]), .RECT3_WEIGHT(rectangle3_weights[808]), .FEAT_THRES(feature_thresholds[808]), .FEAT_ABOVE(feature_aboves[808]), .FEAT_BELOW(feature_belows[808])) ac808(.scan_win(scan_win808), .scan_win_std_dev(scan_win_std_dev[808]), .feature_accum(feature_accums[808]));
  accum_calculator #(.RECT1_X(rectangle1_xs[809]), .RECT1_Y(rectangle1_ys[809]), .RECT1_WIDTH(rectangle1_widths[809]), .RECT1_HEIGHT(rectangle1_heights[809]), .RECT1_WEIGHT(rectangle1_weights[809]), .RECT2_X(rectangle2_xs[809]), .RECT2_Y(rectangle2_ys[809]), .RECT2_WIDTH(rectangle2_widths[809]), .RECT2_HEIGHT(rectangle2_heights[809]), .RECT2_WEIGHT(rectangle2_weights[809]), .RECT3_X(rectangle3_xs[809]), .RECT3_Y(rectangle3_ys[809]), .RECT3_WIDTH(rectangle3_widths[809]), .RECT3_HEIGHT(rectangle3_heights[809]), .RECT3_WEIGHT(rectangle3_weights[809]), .FEAT_THRES(feature_thresholds[809]), .FEAT_ABOVE(feature_aboves[809]), .FEAT_BELOW(feature_belows[809])) ac809(.scan_win(scan_win809), .scan_win_std_dev(scan_win_std_dev[809]), .feature_accum(feature_accums[809]));
  accum_calculator #(.RECT1_X(rectangle1_xs[810]), .RECT1_Y(rectangle1_ys[810]), .RECT1_WIDTH(rectangle1_widths[810]), .RECT1_HEIGHT(rectangle1_heights[810]), .RECT1_WEIGHT(rectangle1_weights[810]), .RECT2_X(rectangle2_xs[810]), .RECT2_Y(rectangle2_ys[810]), .RECT2_WIDTH(rectangle2_widths[810]), .RECT2_HEIGHT(rectangle2_heights[810]), .RECT2_WEIGHT(rectangle2_weights[810]), .RECT3_X(rectangle3_xs[810]), .RECT3_Y(rectangle3_ys[810]), .RECT3_WIDTH(rectangle3_widths[810]), .RECT3_HEIGHT(rectangle3_heights[810]), .RECT3_WEIGHT(rectangle3_weights[810]), .FEAT_THRES(feature_thresholds[810]), .FEAT_ABOVE(feature_aboves[810]), .FEAT_BELOW(feature_belows[810])) ac810(.scan_win(scan_win810), .scan_win_std_dev(scan_win_std_dev[810]), .feature_accum(feature_accums[810]));
  accum_calculator #(.RECT1_X(rectangle1_xs[811]), .RECT1_Y(rectangle1_ys[811]), .RECT1_WIDTH(rectangle1_widths[811]), .RECT1_HEIGHT(rectangle1_heights[811]), .RECT1_WEIGHT(rectangle1_weights[811]), .RECT2_X(rectangle2_xs[811]), .RECT2_Y(rectangle2_ys[811]), .RECT2_WIDTH(rectangle2_widths[811]), .RECT2_HEIGHT(rectangle2_heights[811]), .RECT2_WEIGHT(rectangle2_weights[811]), .RECT3_X(rectangle3_xs[811]), .RECT3_Y(rectangle3_ys[811]), .RECT3_WIDTH(rectangle3_widths[811]), .RECT3_HEIGHT(rectangle3_heights[811]), .RECT3_WEIGHT(rectangle3_weights[811]), .FEAT_THRES(feature_thresholds[811]), .FEAT_ABOVE(feature_aboves[811]), .FEAT_BELOW(feature_belows[811])) ac811(.scan_win(scan_win811), .scan_win_std_dev(scan_win_std_dev[811]), .feature_accum(feature_accums[811]));
  accum_calculator #(.RECT1_X(rectangle1_xs[812]), .RECT1_Y(rectangle1_ys[812]), .RECT1_WIDTH(rectangle1_widths[812]), .RECT1_HEIGHT(rectangle1_heights[812]), .RECT1_WEIGHT(rectangle1_weights[812]), .RECT2_X(rectangle2_xs[812]), .RECT2_Y(rectangle2_ys[812]), .RECT2_WIDTH(rectangle2_widths[812]), .RECT2_HEIGHT(rectangle2_heights[812]), .RECT2_WEIGHT(rectangle2_weights[812]), .RECT3_X(rectangle3_xs[812]), .RECT3_Y(rectangle3_ys[812]), .RECT3_WIDTH(rectangle3_widths[812]), .RECT3_HEIGHT(rectangle3_heights[812]), .RECT3_WEIGHT(rectangle3_weights[812]), .FEAT_THRES(feature_thresholds[812]), .FEAT_ABOVE(feature_aboves[812]), .FEAT_BELOW(feature_belows[812])) ac812(.scan_win(scan_win812), .scan_win_std_dev(scan_win_std_dev[812]), .feature_accum(feature_accums[812]));
  accum_calculator #(.RECT1_X(rectangle1_xs[813]), .RECT1_Y(rectangle1_ys[813]), .RECT1_WIDTH(rectangle1_widths[813]), .RECT1_HEIGHT(rectangle1_heights[813]), .RECT1_WEIGHT(rectangle1_weights[813]), .RECT2_X(rectangle2_xs[813]), .RECT2_Y(rectangle2_ys[813]), .RECT2_WIDTH(rectangle2_widths[813]), .RECT2_HEIGHT(rectangle2_heights[813]), .RECT2_WEIGHT(rectangle2_weights[813]), .RECT3_X(rectangle3_xs[813]), .RECT3_Y(rectangle3_ys[813]), .RECT3_WIDTH(rectangle3_widths[813]), .RECT3_HEIGHT(rectangle3_heights[813]), .RECT3_WEIGHT(rectangle3_weights[813]), .FEAT_THRES(feature_thresholds[813]), .FEAT_ABOVE(feature_aboves[813]), .FEAT_BELOW(feature_belows[813])) ac813(.scan_win(scan_win813), .scan_win_std_dev(scan_win_std_dev[813]), .feature_accum(feature_accums[813]));
  accum_calculator #(.RECT1_X(rectangle1_xs[814]), .RECT1_Y(rectangle1_ys[814]), .RECT1_WIDTH(rectangle1_widths[814]), .RECT1_HEIGHT(rectangle1_heights[814]), .RECT1_WEIGHT(rectangle1_weights[814]), .RECT2_X(rectangle2_xs[814]), .RECT2_Y(rectangle2_ys[814]), .RECT2_WIDTH(rectangle2_widths[814]), .RECT2_HEIGHT(rectangle2_heights[814]), .RECT2_WEIGHT(rectangle2_weights[814]), .RECT3_X(rectangle3_xs[814]), .RECT3_Y(rectangle3_ys[814]), .RECT3_WIDTH(rectangle3_widths[814]), .RECT3_HEIGHT(rectangle3_heights[814]), .RECT3_WEIGHT(rectangle3_weights[814]), .FEAT_THRES(feature_thresholds[814]), .FEAT_ABOVE(feature_aboves[814]), .FEAT_BELOW(feature_belows[814])) ac814(.scan_win(scan_win814), .scan_win_std_dev(scan_win_std_dev[814]), .feature_accum(feature_accums[814]));
  accum_calculator #(.RECT1_X(rectangle1_xs[815]), .RECT1_Y(rectangle1_ys[815]), .RECT1_WIDTH(rectangle1_widths[815]), .RECT1_HEIGHT(rectangle1_heights[815]), .RECT1_WEIGHT(rectangle1_weights[815]), .RECT2_X(rectangle2_xs[815]), .RECT2_Y(rectangle2_ys[815]), .RECT2_WIDTH(rectangle2_widths[815]), .RECT2_HEIGHT(rectangle2_heights[815]), .RECT2_WEIGHT(rectangle2_weights[815]), .RECT3_X(rectangle3_xs[815]), .RECT3_Y(rectangle3_ys[815]), .RECT3_WIDTH(rectangle3_widths[815]), .RECT3_HEIGHT(rectangle3_heights[815]), .RECT3_WEIGHT(rectangle3_weights[815]), .FEAT_THRES(feature_thresholds[815]), .FEAT_ABOVE(feature_aboves[815]), .FEAT_BELOW(feature_belows[815])) ac815(.scan_win(scan_win815), .scan_win_std_dev(scan_win_std_dev[815]), .feature_accum(feature_accums[815]));
  accum_calculator #(.RECT1_X(rectangle1_xs[816]), .RECT1_Y(rectangle1_ys[816]), .RECT1_WIDTH(rectangle1_widths[816]), .RECT1_HEIGHT(rectangle1_heights[816]), .RECT1_WEIGHT(rectangle1_weights[816]), .RECT2_X(rectangle2_xs[816]), .RECT2_Y(rectangle2_ys[816]), .RECT2_WIDTH(rectangle2_widths[816]), .RECT2_HEIGHT(rectangle2_heights[816]), .RECT2_WEIGHT(rectangle2_weights[816]), .RECT3_X(rectangle3_xs[816]), .RECT3_Y(rectangle3_ys[816]), .RECT3_WIDTH(rectangle3_widths[816]), .RECT3_HEIGHT(rectangle3_heights[816]), .RECT3_WEIGHT(rectangle3_weights[816]), .FEAT_THRES(feature_thresholds[816]), .FEAT_ABOVE(feature_aboves[816]), .FEAT_BELOW(feature_belows[816])) ac816(.scan_win(scan_win816), .scan_win_std_dev(scan_win_std_dev[816]), .feature_accum(feature_accums[816]));
  accum_calculator #(.RECT1_X(rectangle1_xs[817]), .RECT1_Y(rectangle1_ys[817]), .RECT1_WIDTH(rectangle1_widths[817]), .RECT1_HEIGHT(rectangle1_heights[817]), .RECT1_WEIGHT(rectangle1_weights[817]), .RECT2_X(rectangle2_xs[817]), .RECT2_Y(rectangle2_ys[817]), .RECT2_WIDTH(rectangle2_widths[817]), .RECT2_HEIGHT(rectangle2_heights[817]), .RECT2_WEIGHT(rectangle2_weights[817]), .RECT3_X(rectangle3_xs[817]), .RECT3_Y(rectangle3_ys[817]), .RECT3_WIDTH(rectangle3_widths[817]), .RECT3_HEIGHT(rectangle3_heights[817]), .RECT3_WEIGHT(rectangle3_weights[817]), .FEAT_THRES(feature_thresholds[817]), .FEAT_ABOVE(feature_aboves[817]), .FEAT_BELOW(feature_belows[817])) ac817(.scan_win(scan_win817), .scan_win_std_dev(scan_win_std_dev[817]), .feature_accum(feature_accums[817]));
  accum_calculator #(.RECT1_X(rectangle1_xs[818]), .RECT1_Y(rectangle1_ys[818]), .RECT1_WIDTH(rectangle1_widths[818]), .RECT1_HEIGHT(rectangle1_heights[818]), .RECT1_WEIGHT(rectangle1_weights[818]), .RECT2_X(rectangle2_xs[818]), .RECT2_Y(rectangle2_ys[818]), .RECT2_WIDTH(rectangle2_widths[818]), .RECT2_HEIGHT(rectangle2_heights[818]), .RECT2_WEIGHT(rectangle2_weights[818]), .RECT3_X(rectangle3_xs[818]), .RECT3_Y(rectangle3_ys[818]), .RECT3_WIDTH(rectangle3_widths[818]), .RECT3_HEIGHT(rectangle3_heights[818]), .RECT3_WEIGHT(rectangle3_weights[818]), .FEAT_THRES(feature_thresholds[818]), .FEAT_ABOVE(feature_aboves[818]), .FEAT_BELOW(feature_belows[818])) ac818(.scan_win(scan_win818), .scan_win_std_dev(scan_win_std_dev[818]), .feature_accum(feature_accums[818]));
  accum_calculator #(.RECT1_X(rectangle1_xs[819]), .RECT1_Y(rectangle1_ys[819]), .RECT1_WIDTH(rectangle1_widths[819]), .RECT1_HEIGHT(rectangle1_heights[819]), .RECT1_WEIGHT(rectangle1_weights[819]), .RECT2_X(rectangle2_xs[819]), .RECT2_Y(rectangle2_ys[819]), .RECT2_WIDTH(rectangle2_widths[819]), .RECT2_HEIGHT(rectangle2_heights[819]), .RECT2_WEIGHT(rectangle2_weights[819]), .RECT3_X(rectangle3_xs[819]), .RECT3_Y(rectangle3_ys[819]), .RECT3_WIDTH(rectangle3_widths[819]), .RECT3_HEIGHT(rectangle3_heights[819]), .RECT3_WEIGHT(rectangle3_weights[819]), .FEAT_THRES(feature_thresholds[819]), .FEAT_ABOVE(feature_aboves[819]), .FEAT_BELOW(feature_belows[819])) ac819(.scan_win(scan_win819), .scan_win_std_dev(scan_win_std_dev[819]), .feature_accum(feature_accums[819]));
  accum_calculator #(.RECT1_X(rectangle1_xs[820]), .RECT1_Y(rectangle1_ys[820]), .RECT1_WIDTH(rectangle1_widths[820]), .RECT1_HEIGHT(rectangle1_heights[820]), .RECT1_WEIGHT(rectangle1_weights[820]), .RECT2_X(rectangle2_xs[820]), .RECT2_Y(rectangle2_ys[820]), .RECT2_WIDTH(rectangle2_widths[820]), .RECT2_HEIGHT(rectangle2_heights[820]), .RECT2_WEIGHT(rectangle2_weights[820]), .RECT3_X(rectangle3_xs[820]), .RECT3_Y(rectangle3_ys[820]), .RECT3_WIDTH(rectangle3_widths[820]), .RECT3_HEIGHT(rectangle3_heights[820]), .RECT3_WEIGHT(rectangle3_weights[820]), .FEAT_THRES(feature_thresholds[820]), .FEAT_ABOVE(feature_aboves[820]), .FEAT_BELOW(feature_belows[820])) ac820(.scan_win(scan_win820), .scan_win_std_dev(scan_win_std_dev[820]), .feature_accum(feature_accums[820]));
  accum_calculator #(.RECT1_X(rectangle1_xs[821]), .RECT1_Y(rectangle1_ys[821]), .RECT1_WIDTH(rectangle1_widths[821]), .RECT1_HEIGHT(rectangle1_heights[821]), .RECT1_WEIGHT(rectangle1_weights[821]), .RECT2_X(rectangle2_xs[821]), .RECT2_Y(rectangle2_ys[821]), .RECT2_WIDTH(rectangle2_widths[821]), .RECT2_HEIGHT(rectangle2_heights[821]), .RECT2_WEIGHT(rectangle2_weights[821]), .RECT3_X(rectangle3_xs[821]), .RECT3_Y(rectangle3_ys[821]), .RECT3_WIDTH(rectangle3_widths[821]), .RECT3_HEIGHT(rectangle3_heights[821]), .RECT3_WEIGHT(rectangle3_weights[821]), .FEAT_THRES(feature_thresholds[821]), .FEAT_ABOVE(feature_aboves[821]), .FEAT_BELOW(feature_belows[821])) ac821(.scan_win(scan_win821), .scan_win_std_dev(scan_win_std_dev[821]), .feature_accum(feature_accums[821]));
  accum_calculator #(.RECT1_X(rectangle1_xs[822]), .RECT1_Y(rectangle1_ys[822]), .RECT1_WIDTH(rectangle1_widths[822]), .RECT1_HEIGHT(rectangle1_heights[822]), .RECT1_WEIGHT(rectangle1_weights[822]), .RECT2_X(rectangle2_xs[822]), .RECT2_Y(rectangle2_ys[822]), .RECT2_WIDTH(rectangle2_widths[822]), .RECT2_HEIGHT(rectangle2_heights[822]), .RECT2_WEIGHT(rectangle2_weights[822]), .RECT3_X(rectangle3_xs[822]), .RECT3_Y(rectangle3_ys[822]), .RECT3_WIDTH(rectangle3_widths[822]), .RECT3_HEIGHT(rectangle3_heights[822]), .RECT3_WEIGHT(rectangle3_weights[822]), .FEAT_THRES(feature_thresholds[822]), .FEAT_ABOVE(feature_aboves[822]), .FEAT_BELOW(feature_belows[822])) ac822(.scan_win(scan_win822), .scan_win_std_dev(scan_win_std_dev[822]), .feature_accum(feature_accums[822]));
  accum_calculator #(.RECT1_X(rectangle1_xs[823]), .RECT1_Y(rectangle1_ys[823]), .RECT1_WIDTH(rectangle1_widths[823]), .RECT1_HEIGHT(rectangle1_heights[823]), .RECT1_WEIGHT(rectangle1_weights[823]), .RECT2_X(rectangle2_xs[823]), .RECT2_Y(rectangle2_ys[823]), .RECT2_WIDTH(rectangle2_widths[823]), .RECT2_HEIGHT(rectangle2_heights[823]), .RECT2_WEIGHT(rectangle2_weights[823]), .RECT3_X(rectangle3_xs[823]), .RECT3_Y(rectangle3_ys[823]), .RECT3_WIDTH(rectangle3_widths[823]), .RECT3_HEIGHT(rectangle3_heights[823]), .RECT3_WEIGHT(rectangle3_weights[823]), .FEAT_THRES(feature_thresholds[823]), .FEAT_ABOVE(feature_aboves[823]), .FEAT_BELOW(feature_belows[823])) ac823(.scan_win(scan_win823), .scan_win_std_dev(scan_win_std_dev[823]), .feature_accum(feature_accums[823]));
  accum_calculator #(.RECT1_X(rectangle1_xs[824]), .RECT1_Y(rectangle1_ys[824]), .RECT1_WIDTH(rectangle1_widths[824]), .RECT1_HEIGHT(rectangle1_heights[824]), .RECT1_WEIGHT(rectangle1_weights[824]), .RECT2_X(rectangle2_xs[824]), .RECT2_Y(rectangle2_ys[824]), .RECT2_WIDTH(rectangle2_widths[824]), .RECT2_HEIGHT(rectangle2_heights[824]), .RECT2_WEIGHT(rectangle2_weights[824]), .RECT3_X(rectangle3_xs[824]), .RECT3_Y(rectangle3_ys[824]), .RECT3_WIDTH(rectangle3_widths[824]), .RECT3_HEIGHT(rectangle3_heights[824]), .RECT3_WEIGHT(rectangle3_weights[824]), .FEAT_THRES(feature_thresholds[824]), .FEAT_ABOVE(feature_aboves[824]), .FEAT_BELOW(feature_belows[824])) ac824(.scan_win(scan_win824), .scan_win_std_dev(scan_win_std_dev[824]), .feature_accum(feature_accums[824]));
  accum_calculator #(.RECT1_X(rectangle1_xs[825]), .RECT1_Y(rectangle1_ys[825]), .RECT1_WIDTH(rectangle1_widths[825]), .RECT1_HEIGHT(rectangle1_heights[825]), .RECT1_WEIGHT(rectangle1_weights[825]), .RECT2_X(rectangle2_xs[825]), .RECT2_Y(rectangle2_ys[825]), .RECT2_WIDTH(rectangle2_widths[825]), .RECT2_HEIGHT(rectangle2_heights[825]), .RECT2_WEIGHT(rectangle2_weights[825]), .RECT3_X(rectangle3_xs[825]), .RECT3_Y(rectangle3_ys[825]), .RECT3_WIDTH(rectangle3_widths[825]), .RECT3_HEIGHT(rectangle3_heights[825]), .RECT3_WEIGHT(rectangle3_weights[825]), .FEAT_THRES(feature_thresholds[825]), .FEAT_ABOVE(feature_aboves[825]), .FEAT_BELOW(feature_belows[825])) ac825(.scan_win(scan_win825), .scan_win_std_dev(scan_win_std_dev[825]), .feature_accum(feature_accums[825]));
  accum_calculator #(.RECT1_X(rectangle1_xs[826]), .RECT1_Y(rectangle1_ys[826]), .RECT1_WIDTH(rectangle1_widths[826]), .RECT1_HEIGHT(rectangle1_heights[826]), .RECT1_WEIGHT(rectangle1_weights[826]), .RECT2_X(rectangle2_xs[826]), .RECT2_Y(rectangle2_ys[826]), .RECT2_WIDTH(rectangle2_widths[826]), .RECT2_HEIGHT(rectangle2_heights[826]), .RECT2_WEIGHT(rectangle2_weights[826]), .RECT3_X(rectangle3_xs[826]), .RECT3_Y(rectangle3_ys[826]), .RECT3_WIDTH(rectangle3_widths[826]), .RECT3_HEIGHT(rectangle3_heights[826]), .RECT3_WEIGHT(rectangle3_weights[826]), .FEAT_THRES(feature_thresholds[826]), .FEAT_ABOVE(feature_aboves[826]), .FEAT_BELOW(feature_belows[826])) ac826(.scan_win(scan_win826), .scan_win_std_dev(scan_win_std_dev[826]), .feature_accum(feature_accums[826]));
  accum_calculator #(.RECT1_X(rectangle1_xs[827]), .RECT1_Y(rectangle1_ys[827]), .RECT1_WIDTH(rectangle1_widths[827]), .RECT1_HEIGHT(rectangle1_heights[827]), .RECT1_WEIGHT(rectangle1_weights[827]), .RECT2_X(rectangle2_xs[827]), .RECT2_Y(rectangle2_ys[827]), .RECT2_WIDTH(rectangle2_widths[827]), .RECT2_HEIGHT(rectangle2_heights[827]), .RECT2_WEIGHT(rectangle2_weights[827]), .RECT3_X(rectangle3_xs[827]), .RECT3_Y(rectangle3_ys[827]), .RECT3_WIDTH(rectangle3_widths[827]), .RECT3_HEIGHT(rectangle3_heights[827]), .RECT3_WEIGHT(rectangle3_weights[827]), .FEAT_THRES(feature_thresholds[827]), .FEAT_ABOVE(feature_aboves[827]), .FEAT_BELOW(feature_belows[827])) ac827(.scan_win(scan_win827), .scan_win_std_dev(scan_win_std_dev[827]), .feature_accum(feature_accums[827]));
  accum_calculator #(.RECT1_X(rectangle1_xs[828]), .RECT1_Y(rectangle1_ys[828]), .RECT1_WIDTH(rectangle1_widths[828]), .RECT1_HEIGHT(rectangle1_heights[828]), .RECT1_WEIGHT(rectangle1_weights[828]), .RECT2_X(rectangle2_xs[828]), .RECT2_Y(rectangle2_ys[828]), .RECT2_WIDTH(rectangle2_widths[828]), .RECT2_HEIGHT(rectangle2_heights[828]), .RECT2_WEIGHT(rectangle2_weights[828]), .RECT3_X(rectangle3_xs[828]), .RECT3_Y(rectangle3_ys[828]), .RECT3_WIDTH(rectangle3_widths[828]), .RECT3_HEIGHT(rectangle3_heights[828]), .RECT3_WEIGHT(rectangle3_weights[828]), .FEAT_THRES(feature_thresholds[828]), .FEAT_ABOVE(feature_aboves[828]), .FEAT_BELOW(feature_belows[828])) ac828(.scan_win(scan_win828), .scan_win_std_dev(scan_win_std_dev[828]), .feature_accum(feature_accums[828]));
  accum_calculator #(.RECT1_X(rectangle1_xs[829]), .RECT1_Y(rectangle1_ys[829]), .RECT1_WIDTH(rectangle1_widths[829]), .RECT1_HEIGHT(rectangle1_heights[829]), .RECT1_WEIGHT(rectangle1_weights[829]), .RECT2_X(rectangle2_xs[829]), .RECT2_Y(rectangle2_ys[829]), .RECT2_WIDTH(rectangle2_widths[829]), .RECT2_HEIGHT(rectangle2_heights[829]), .RECT2_WEIGHT(rectangle2_weights[829]), .RECT3_X(rectangle3_xs[829]), .RECT3_Y(rectangle3_ys[829]), .RECT3_WIDTH(rectangle3_widths[829]), .RECT3_HEIGHT(rectangle3_heights[829]), .RECT3_WEIGHT(rectangle3_weights[829]), .FEAT_THRES(feature_thresholds[829]), .FEAT_ABOVE(feature_aboves[829]), .FEAT_BELOW(feature_belows[829])) ac829(.scan_win(scan_win829), .scan_win_std_dev(scan_win_std_dev[829]), .feature_accum(feature_accums[829]));
  accum_calculator #(.RECT1_X(rectangle1_xs[830]), .RECT1_Y(rectangle1_ys[830]), .RECT1_WIDTH(rectangle1_widths[830]), .RECT1_HEIGHT(rectangle1_heights[830]), .RECT1_WEIGHT(rectangle1_weights[830]), .RECT2_X(rectangle2_xs[830]), .RECT2_Y(rectangle2_ys[830]), .RECT2_WIDTH(rectangle2_widths[830]), .RECT2_HEIGHT(rectangle2_heights[830]), .RECT2_WEIGHT(rectangle2_weights[830]), .RECT3_X(rectangle3_xs[830]), .RECT3_Y(rectangle3_ys[830]), .RECT3_WIDTH(rectangle3_widths[830]), .RECT3_HEIGHT(rectangle3_heights[830]), .RECT3_WEIGHT(rectangle3_weights[830]), .FEAT_THRES(feature_thresholds[830]), .FEAT_ABOVE(feature_aboves[830]), .FEAT_BELOW(feature_belows[830])) ac830(.scan_win(scan_win830), .scan_win_std_dev(scan_win_std_dev[830]), .feature_accum(feature_accums[830]));
  accum_calculator #(.RECT1_X(rectangle1_xs[831]), .RECT1_Y(rectangle1_ys[831]), .RECT1_WIDTH(rectangle1_widths[831]), .RECT1_HEIGHT(rectangle1_heights[831]), .RECT1_WEIGHT(rectangle1_weights[831]), .RECT2_X(rectangle2_xs[831]), .RECT2_Y(rectangle2_ys[831]), .RECT2_WIDTH(rectangle2_widths[831]), .RECT2_HEIGHT(rectangle2_heights[831]), .RECT2_WEIGHT(rectangle2_weights[831]), .RECT3_X(rectangle3_xs[831]), .RECT3_Y(rectangle3_ys[831]), .RECT3_WIDTH(rectangle3_widths[831]), .RECT3_HEIGHT(rectangle3_heights[831]), .RECT3_WEIGHT(rectangle3_weights[831]), .FEAT_THRES(feature_thresholds[831]), .FEAT_ABOVE(feature_aboves[831]), .FEAT_BELOW(feature_belows[831])) ac831(.scan_win(scan_win831), .scan_win_std_dev(scan_win_std_dev[831]), .feature_accum(feature_accums[831]));
  accum_calculator #(.RECT1_X(rectangle1_xs[832]), .RECT1_Y(rectangle1_ys[832]), .RECT1_WIDTH(rectangle1_widths[832]), .RECT1_HEIGHT(rectangle1_heights[832]), .RECT1_WEIGHT(rectangle1_weights[832]), .RECT2_X(rectangle2_xs[832]), .RECT2_Y(rectangle2_ys[832]), .RECT2_WIDTH(rectangle2_widths[832]), .RECT2_HEIGHT(rectangle2_heights[832]), .RECT2_WEIGHT(rectangle2_weights[832]), .RECT3_X(rectangle3_xs[832]), .RECT3_Y(rectangle3_ys[832]), .RECT3_WIDTH(rectangle3_widths[832]), .RECT3_HEIGHT(rectangle3_heights[832]), .RECT3_WEIGHT(rectangle3_weights[832]), .FEAT_THRES(feature_thresholds[832]), .FEAT_ABOVE(feature_aboves[832]), .FEAT_BELOW(feature_belows[832])) ac832(.scan_win(scan_win832), .scan_win_std_dev(scan_win_std_dev[832]), .feature_accum(feature_accums[832]));
  accum_calculator #(.RECT1_X(rectangle1_xs[833]), .RECT1_Y(rectangle1_ys[833]), .RECT1_WIDTH(rectangle1_widths[833]), .RECT1_HEIGHT(rectangle1_heights[833]), .RECT1_WEIGHT(rectangle1_weights[833]), .RECT2_X(rectangle2_xs[833]), .RECT2_Y(rectangle2_ys[833]), .RECT2_WIDTH(rectangle2_widths[833]), .RECT2_HEIGHT(rectangle2_heights[833]), .RECT2_WEIGHT(rectangle2_weights[833]), .RECT3_X(rectangle3_xs[833]), .RECT3_Y(rectangle3_ys[833]), .RECT3_WIDTH(rectangle3_widths[833]), .RECT3_HEIGHT(rectangle3_heights[833]), .RECT3_WEIGHT(rectangle3_weights[833]), .FEAT_THRES(feature_thresholds[833]), .FEAT_ABOVE(feature_aboves[833]), .FEAT_BELOW(feature_belows[833])) ac833(.scan_win(scan_win833), .scan_win_std_dev(scan_win_std_dev[833]), .feature_accum(feature_accums[833]));
  accum_calculator #(.RECT1_X(rectangle1_xs[834]), .RECT1_Y(rectangle1_ys[834]), .RECT1_WIDTH(rectangle1_widths[834]), .RECT1_HEIGHT(rectangle1_heights[834]), .RECT1_WEIGHT(rectangle1_weights[834]), .RECT2_X(rectangle2_xs[834]), .RECT2_Y(rectangle2_ys[834]), .RECT2_WIDTH(rectangle2_widths[834]), .RECT2_HEIGHT(rectangle2_heights[834]), .RECT2_WEIGHT(rectangle2_weights[834]), .RECT3_X(rectangle3_xs[834]), .RECT3_Y(rectangle3_ys[834]), .RECT3_WIDTH(rectangle3_widths[834]), .RECT3_HEIGHT(rectangle3_heights[834]), .RECT3_WEIGHT(rectangle3_weights[834]), .FEAT_THRES(feature_thresholds[834]), .FEAT_ABOVE(feature_aboves[834]), .FEAT_BELOW(feature_belows[834])) ac834(.scan_win(scan_win834), .scan_win_std_dev(scan_win_std_dev[834]), .feature_accum(feature_accums[834]));
  accum_calculator #(.RECT1_X(rectangle1_xs[835]), .RECT1_Y(rectangle1_ys[835]), .RECT1_WIDTH(rectangle1_widths[835]), .RECT1_HEIGHT(rectangle1_heights[835]), .RECT1_WEIGHT(rectangle1_weights[835]), .RECT2_X(rectangle2_xs[835]), .RECT2_Y(rectangle2_ys[835]), .RECT2_WIDTH(rectangle2_widths[835]), .RECT2_HEIGHT(rectangle2_heights[835]), .RECT2_WEIGHT(rectangle2_weights[835]), .RECT3_X(rectangle3_xs[835]), .RECT3_Y(rectangle3_ys[835]), .RECT3_WIDTH(rectangle3_widths[835]), .RECT3_HEIGHT(rectangle3_heights[835]), .RECT3_WEIGHT(rectangle3_weights[835]), .FEAT_THRES(feature_thresholds[835]), .FEAT_ABOVE(feature_aboves[835]), .FEAT_BELOW(feature_belows[835])) ac835(.scan_win(scan_win835), .scan_win_std_dev(scan_win_std_dev[835]), .feature_accum(feature_accums[835]));
  accum_calculator #(.RECT1_X(rectangle1_xs[836]), .RECT1_Y(rectangle1_ys[836]), .RECT1_WIDTH(rectangle1_widths[836]), .RECT1_HEIGHT(rectangle1_heights[836]), .RECT1_WEIGHT(rectangle1_weights[836]), .RECT2_X(rectangle2_xs[836]), .RECT2_Y(rectangle2_ys[836]), .RECT2_WIDTH(rectangle2_widths[836]), .RECT2_HEIGHT(rectangle2_heights[836]), .RECT2_WEIGHT(rectangle2_weights[836]), .RECT3_X(rectangle3_xs[836]), .RECT3_Y(rectangle3_ys[836]), .RECT3_WIDTH(rectangle3_widths[836]), .RECT3_HEIGHT(rectangle3_heights[836]), .RECT3_WEIGHT(rectangle3_weights[836]), .FEAT_THRES(feature_thresholds[836]), .FEAT_ABOVE(feature_aboves[836]), .FEAT_BELOW(feature_belows[836])) ac836(.scan_win(scan_win836), .scan_win_std_dev(scan_win_std_dev[836]), .feature_accum(feature_accums[836]));
  accum_calculator #(.RECT1_X(rectangle1_xs[837]), .RECT1_Y(rectangle1_ys[837]), .RECT1_WIDTH(rectangle1_widths[837]), .RECT1_HEIGHT(rectangle1_heights[837]), .RECT1_WEIGHT(rectangle1_weights[837]), .RECT2_X(rectangle2_xs[837]), .RECT2_Y(rectangle2_ys[837]), .RECT2_WIDTH(rectangle2_widths[837]), .RECT2_HEIGHT(rectangle2_heights[837]), .RECT2_WEIGHT(rectangle2_weights[837]), .RECT3_X(rectangle3_xs[837]), .RECT3_Y(rectangle3_ys[837]), .RECT3_WIDTH(rectangle3_widths[837]), .RECT3_HEIGHT(rectangle3_heights[837]), .RECT3_WEIGHT(rectangle3_weights[837]), .FEAT_THRES(feature_thresholds[837]), .FEAT_ABOVE(feature_aboves[837]), .FEAT_BELOW(feature_belows[837])) ac837(.scan_win(scan_win837), .scan_win_std_dev(scan_win_std_dev[837]), .feature_accum(feature_accums[837]));
  accum_calculator #(.RECT1_X(rectangle1_xs[838]), .RECT1_Y(rectangle1_ys[838]), .RECT1_WIDTH(rectangle1_widths[838]), .RECT1_HEIGHT(rectangle1_heights[838]), .RECT1_WEIGHT(rectangle1_weights[838]), .RECT2_X(rectangle2_xs[838]), .RECT2_Y(rectangle2_ys[838]), .RECT2_WIDTH(rectangle2_widths[838]), .RECT2_HEIGHT(rectangle2_heights[838]), .RECT2_WEIGHT(rectangle2_weights[838]), .RECT3_X(rectangle3_xs[838]), .RECT3_Y(rectangle3_ys[838]), .RECT3_WIDTH(rectangle3_widths[838]), .RECT3_HEIGHT(rectangle3_heights[838]), .RECT3_WEIGHT(rectangle3_weights[838]), .FEAT_THRES(feature_thresholds[838]), .FEAT_ABOVE(feature_aboves[838]), .FEAT_BELOW(feature_belows[838])) ac838(.scan_win(scan_win838), .scan_win_std_dev(scan_win_std_dev[838]), .feature_accum(feature_accums[838]));
  accum_calculator #(.RECT1_X(rectangle1_xs[839]), .RECT1_Y(rectangle1_ys[839]), .RECT1_WIDTH(rectangle1_widths[839]), .RECT1_HEIGHT(rectangle1_heights[839]), .RECT1_WEIGHT(rectangle1_weights[839]), .RECT2_X(rectangle2_xs[839]), .RECT2_Y(rectangle2_ys[839]), .RECT2_WIDTH(rectangle2_widths[839]), .RECT2_HEIGHT(rectangle2_heights[839]), .RECT2_WEIGHT(rectangle2_weights[839]), .RECT3_X(rectangle3_xs[839]), .RECT3_Y(rectangle3_ys[839]), .RECT3_WIDTH(rectangle3_widths[839]), .RECT3_HEIGHT(rectangle3_heights[839]), .RECT3_WEIGHT(rectangle3_weights[839]), .FEAT_THRES(feature_thresholds[839]), .FEAT_ABOVE(feature_aboves[839]), .FEAT_BELOW(feature_belows[839])) ac839(.scan_win(scan_win839), .scan_win_std_dev(scan_win_std_dev[839]), .feature_accum(feature_accums[839]));
  accum_calculator #(.RECT1_X(rectangle1_xs[840]), .RECT1_Y(rectangle1_ys[840]), .RECT1_WIDTH(rectangle1_widths[840]), .RECT1_HEIGHT(rectangle1_heights[840]), .RECT1_WEIGHT(rectangle1_weights[840]), .RECT2_X(rectangle2_xs[840]), .RECT2_Y(rectangle2_ys[840]), .RECT2_WIDTH(rectangle2_widths[840]), .RECT2_HEIGHT(rectangle2_heights[840]), .RECT2_WEIGHT(rectangle2_weights[840]), .RECT3_X(rectangle3_xs[840]), .RECT3_Y(rectangle3_ys[840]), .RECT3_WIDTH(rectangle3_widths[840]), .RECT3_HEIGHT(rectangle3_heights[840]), .RECT3_WEIGHT(rectangle3_weights[840]), .FEAT_THRES(feature_thresholds[840]), .FEAT_ABOVE(feature_aboves[840]), .FEAT_BELOW(feature_belows[840])) ac840(.scan_win(scan_win840), .scan_win_std_dev(scan_win_std_dev[840]), .feature_accum(feature_accums[840]));
  accum_calculator #(.RECT1_X(rectangle1_xs[841]), .RECT1_Y(rectangle1_ys[841]), .RECT1_WIDTH(rectangle1_widths[841]), .RECT1_HEIGHT(rectangle1_heights[841]), .RECT1_WEIGHT(rectangle1_weights[841]), .RECT2_X(rectangle2_xs[841]), .RECT2_Y(rectangle2_ys[841]), .RECT2_WIDTH(rectangle2_widths[841]), .RECT2_HEIGHT(rectangle2_heights[841]), .RECT2_WEIGHT(rectangle2_weights[841]), .RECT3_X(rectangle3_xs[841]), .RECT3_Y(rectangle3_ys[841]), .RECT3_WIDTH(rectangle3_widths[841]), .RECT3_HEIGHT(rectangle3_heights[841]), .RECT3_WEIGHT(rectangle3_weights[841]), .FEAT_THRES(feature_thresholds[841]), .FEAT_ABOVE(feature_aboves[841]), .FEAT_BELOW(feature_belows[841])) ac841(.scan_win(scan_win841), .scan_win_std_dev(scan_win_std_dev[841]), .feature_accum(feature_accums[841]));
  accum_calculator #(.RECT1_X(rectangle1_xs[842]), .RECT1_Y(rectangle1_ys[842]), .RECT1_WIDTH(rectangle1_widths[842]), .RECT1_HEIGHT(rectangle1_heights[842]), .RECT1_WEIGHT(rectangle1_weights[842]), .RECT2_X(rectangle2_xs[842]), .RECT2_Y(rectangle2_ys[842]), .RECT2_WIDTH(rectangle2_widths[842]), .RECT2_HEIGHT(rectangle2_heights[842]), .RECT2_WEIGHT(rectangle2_weights[842]), .RECT3_X(rectangle3_xs[842]), .RECT3_Y(rectangle3_ys[842]), .RECT3_WIDTH(rectangle3_widths[842]), .RECT3_HEIGHT(rectangle3_heights[842]), .RECT3_WEIGHT(rectangle3_weights[842]), .FEAT_THRES(feature_thresholds[842]), .FEAT_ABOVE(feature_aboves[842]), .FEAT_BELOW(feature_belows[842])) ac842(.scan_win(scan_win842), .scan_win_std_dev(scan_win_std_dev[842]), .feature_accum(feature_accums[842]));
  accum_calculator #(.RECT1_X(rectangle1_xs[843]), .RECT1_Y(rectangle1_ys[843]), .RECT1_WIDTH(rectangle1_widths[843]), .RECT1_HEIGHT(rectangle1_heights[843]), .RECT1_WEIGHT(rectangle1_weights[843]), .RECT2_X(rectangle2_xs[843]), .RECT2_Y(rectangle2_ys[843]), .RECT2_WIDTH(rectangle2_widths[843]), .RECT2_HEIGHT(rectangle2_heights[843]), .RECT2_WEIGHT(rectangle2_weights[843]), .RECT3_X(rectangle3_xs[843]), .RECT3_Y(rectangle3_ys[843]), .RECT3_WIDTH(rectangle3_widths[843]), .RECT3_HEIGHT(rectangle3_heights[843]), .RECT3_WEIGHT(rectangle3_weights[843]), .FEAT_THRES(feature_thresholds[843]), .FEAT_ABOVE(feature_aboves[843]), .FEAT_BELOW(feature_belows[843])) ac843(.scan_win(scan_win843), .scan_win_std_dev(scan_win_std_dev[843]), .feature_accum(feature_accums[843]));
  accum_calculator #(.RECT1_X(rectangle1_xs[844]), .RECT1_Y(rectangle1_ys[844]), .RECT1_WIDTH(rectangle1_widths[844]), .RECT1_HEIGHT(rectangle1_heights[844]), .RECT1_WEIGHT(rectangle1_weights[844]), .RECT2_X(rectangle2_xs[844]), .RECT2_Y(rectangle2_ys[844]), .RECT2_WIDTH(rectangle2_widths[844]), .RECT2_HEIGHT(rectangle2_heights[844]), .RECT2_WEIGHT(rectangle2_weights[844]), .RECT3_X(rectangle3_xs[844]), .RECT3_Y(rectangle3_ys[844]), .RECT3_WIDTH(rectangle3_widths[844]), .RECT3_HEIGHT(rectangle3_heights[844]), .RECT3_WEIGHT(rectangle3_weights[844]), .FEAT_THRES(feature_thresholds[844]), .FEAT_ABOVE(feature_aboves[844]), .FEAT_BELOW(feature_belows[844])) ac844(.scan_win(scan_win844), .scan_win_std_dev(scan_win_std_dev[844]), .feature_accum(feature_accums[844]));
  accum_calculator #(.RECT1_X(rectangle1_xs[845]), .RECT1_Y(rectangle1_ys[845]), .RECT1_WIDTH(rectangle1_widths[845]), .RECT1_HEIGHT(rectangle1_heights[845]), .RECT1_WEIGHT(rectangle1_weights[845]), .RECT2_X(rectangle2_xs[845]), .RECT2_Y(rectangle2_ys[845]), .RECT2_WIDTH(rectangle2_widths[845]), .RECT2_HEIGHT(rectangle2_heights[845]), .RECT2_WEIGHT(rectangle2_weights[845]), .RECT3_X(rectangle3_xs[845]), .RECT3_Y(rectangle3_ys[845]), .RECT3_WIDTH(rectangle3_widths[845]), .RECT3_HEIGHT(rectangle3_heights[845]), .RECT3_WEIGHT(rectangle3_weights[845]), .FEAT_THRES(feature_thresholds[845]), .FEAT_ABOVE(feature_aboves[845]), .FEAT_BELOW(feature_belows[845])) ac845(.scan_win(scan_win845), .scan_win_std_dev(scan_win_std_dev[845]), .feature_accum(feature_accums[845]));
  accum_calculator #(.RECT1_X(rectangle1_xs[846]), .RECT1_Y(rectangle1_ys[846]), .RECT1_WIDTH(rectangle1_widths[846]), .RECT1_HEIGHT(rectangle1_heights[846]), .RECT1_WEIGHT(rectangle1_weights[846]), .RECT2_X(rectangle2_xs[846]), .RECT2_Y(rectangle2_ys[846]), .RECT2_WIDTH(rectangle2_widths[846]), .RECT2_HEIGHT(rectangle2_heights[846]), .RECT2_WEIGHT(rectangle2_weights[846]), .RECT3_X(rectangle3_xs[846]), .RECT3_Y(rectangle3_ys[846]), .RECT3_WIDTH(rectangle3_widths[846]), .RECT3_HEIGHT(rectangle3_heights[846]), .RECT3_WEIGHT(rectangle3_weights[846]), .FEAT_THRES(feature_thresholds[846]), .FEAT_ABOVE(feature_aboves[846]), .FEAT_BELOW(feature_belows[846])) ac846(.scan_win(scan_win846), .scan_win_std_dev(scan_win_std_dev[846]), .feature_accum(feature_accums[846]));
  accum_calculator #(.RECT1_X(rectangle1_xs[847]), .RECT1_Y(rectangle1_ys[847]), .RECT1_WIDTH(rectangle1_widths[847]), .RECT1_HEIGHT(rectangle1_heights[847]), .RECT1_WEIGHT(rectangle1_weights[847]), .RECT2_X(rectangle2_xs[847]), .RECT2_Y(rectangle2_ys[847]), .RECT2_WIDTH(rectangle2_widths[847]), .RECT2_HEIGHT(rectangle2_heights[847]), .RECT2_WEIGHT(rectangle2_weights[847]), .RECT3_X(rectangle3_xs[847]), .RECT3_Y(rectangle3_ys[847]), .RECT3_WIDTH(rectangle3_widths[847]), .RECT3_HEIGHT(rectangle3_heights[847]), .RECT3_WEIGHT(rectangle3_weights[847]), .FEAT_THRES(feature_thresholds[847]), .FEAT_ABOVE(feature_aboves[847]), .FEAT_BELOW(feature_belows[847])) ac847(.scan_win(scan_win847), .scan_win_std_dev(scan_win_std_dev[847]), .feature_accum(feature_accums[847]));
  accum_calculator #(.RECT1_X(rectangle1_xs[848]), .RECT1_Y(rectangle1_ys[848]), .RECT1_WIDTH(rectangle1_widths[848]), .RECT1_HEIGHT(rectangle1_heights[848]), .RECT1_WEIGHT(rectangle1_weights[848]), .RECT2_X(rectangle2_xs[848]), .RECT2_Y(rectangle2_ys[848]), .RECT2_WIDTH(rectangle2_widths[848]), .RECT2_HEIGHT(rectangle2_heights[848]), .RECT2_WEIGHT(rectangle2_weights[848]), .RECT3_X(rectangle3_xs[848]), .RECT3_Y(rectangle3_ys[848]), .RECT3_WIDTH(rectangle3_widths[848]), .RECT3_HEIGHT(rectangle3_heights[848]), .RECT3_WEIGHT(rectangle3_weights[848]), .FEAT_THRES(feature_thresholds[848]), .FEAT_ABOVE(feature_aboves[848]), .FEAT_BELOW(feature_belows[848])) ac848(.scan_win(scan_win848), .scan_win_std_dev(scan_win_std_dev[848]), .feature_accum(feature_accums[848]));
  accum_calculator #(.RECT1_X(rectangle1_xs[849]), .RECT1_Y(rectangle1_ys[849]), .RECT1_WIDTH(rectangle1_widths[849]), .RECT1_HEIGHT(rectangle1_heights[849]), .RECT1_WEIGHT(rectangle1_weights[849]), .RECT2_X(rectangle2_xs[849]), .RECT2_Y(rectangle2_ys[849]), .RECT2_WIDTH(rectangle2_widths[849]), .RECT2_HEIGHT(rectangle2_heights[849]), .RECT2_WEIGHT(rectangle2_weights[849]), .RECT3_X(rectangle3_xs[849]), .RECT3_Y(rectangle3_ys[849]), .RECT3_WIDTH(rectangle3_widths[849]), .RECT3_HEIGHT(rectangle3_heights[849]), .RECT3_WEIGHT(rectangle3_weights[849]), .FEAT_THRES(feature_thresholds[849]), .FEAT_ABOVE(feature_aboves[849]), .FEAT_BELOW(feature_belows[849])) ac849(.scan_win(scan_win849), .scan_win_std_dev(scan_win_std_dev[849]), .feature_accum(feature_accums[849]));
  accum_calculator #(.RECT1_X(rectangle1_xs[850]), .RECT1_Y(rectangle1_ys[850]), .RECT1_WIDTH(rectangle1_widths[850]), .RECT1_HEIGHT(rectangle1_heights[850]), .RECT1_WEIGHT(rectangle1_weights[850]), .RECT2_X(rectangle2_xs[850]), .RECT2_Y(rectangle2_ys[850]), .RECT2_WIDTH(rectangle2_widths[850]), .RECT2_HEIGHT(rectangle2_heights[850]), .RECT2_WEIGHT(rectangle2_weights[850]), .RECT3_X(rectangle3_xs[850]), .RECT3_Y(rectangle3_ys[850]), .RECT3_WIDTH(rectangle3_widths[850]), .RECT3_HEIGHT(rectangle3_heights[850]), .RECT3_WEIGHT(rectangle3_weights[850]), .FEAT_THRES(feature_thresholds[850]), .FEAT_ABOVE(feature_aboves[850]), .FEAT_BELOW(feature_belows[850])) ac850(.scan_win(scan_win850), .scan_win_std_dev(scan_win_std_dev[850]), .feature_accum(feature_accums[850]));
  accum_calculator #(.RECT1_X(rectangle1_xs[851]), .RECT1_Y(rectangle1_ys[851]), .RECT1_WIDTH(rectangle1_widths[851]), .RECT1_HEIGHT(rectangle1_heights[851]), .RECT1_WEIGHT(rectangle1_weights[851]), .RECT2_X(rectangle2_xs[851]), .RECT2_Y(rectangle2_ys[851]), .RECT2_WIDTH(rectangle2_widths[851]), .RECT2_HEIGHT(rectangle2_heights[851]), .RECT2_WEIGHT(rectangle2_weights[851]), .RECT3_X(rectangle3_xs[851]), .RECT3_Y(rectangle3_ys[851]), .RECT3_WIDTH(rectangle3_widths[851]), .RECT3_HEIGHT(rectangle3_heights[851]), .RECT3_WEIGHT(rectangle3_weights[851]), .FEAT_THRES(feature_thresholds[851]), .FEAT_ABOVE(feature_aboves[851]), .FEAT_BELOW(feature_belows[851])) ac851(.scan_win(scan_win851), .scan_win_std_dev(scan_win_std_dev[851]), .feature_accum(feature_accums[851]));
  accum_calculator #(.RECT1_X(rectangle1_xs[852]), .RECT1_Y(rectangle1_ys[852]), .RECT1_WIDTH(rectangle1_widths[852]), .RECT1_HEIGHT(rectangle1_heights[852]), .RECT1_WEIGHT(rectangle1_weights[852]), .RECT2_X(rectangle2_xs[852]), .RECT2_Y(rectangle2_ys[852]), .RECT2_WIDTH(rectangle2_widths[852]), .RECT2_HEIGHT(rectangle2_heights[852]), .RECT2_WEIGHT(rectangle2_weights[852]), .RECT3_X(rectangle3_xs[852]), .RECT3_Y(rectangle3_ys[852]), .RECT3_WIDTH(rectangle3_widths[852]), .RECT3_HEIGHT(rectangle3_heights[852]), .RECT3_WEIGHT(rectangle3_weights[852]), .FEAT_THRES(feature_thresholds[852]), .FEAT_ABOVE(feature_aboves[852]), .FEAT_BELOW(feature_belows[852])) ac852(.scan_win(scan_win852), .scan_win_std_dev(scan_win_std_dev[852]), .feature_accum(feature_accums[852]));
  accum_calculator #(.RECT1_X(rectangle1_xs[853]), .RECT1_Y(rectangle1_ys[853]), .RECT1_WIDTH(rectangle1_widths[853]), .RECT1_HEIGHT(rectangle1_heights[853]), .RECT1_WEIGHT(rectangle1_weights[853]), .RECT2_X(rectangle2_xs[853]), .RECT2_Y(rectangle2_ys[853]), .RECT2_WIDTH(rectangle2_widths[853]), .RECT2_HEIGHT(rectangle2_heights[853]), .RECT2_WEIGHT(rectangle2_weights[853]), .RECT3_X(rectangle3_xs[853]), .RECT3_Y(rectangle3_ys[853]), .RECT3_WIDTH(rectangle3_widths[853]), .RECT3_HEIGHT(rectangle3_heights[853]), .RECT3_WEIGHT(rectangle3_weights[853]), .FEAT_THRES(feature_thresholds[853]), .FEAT_ABOVE(feature_aboves[853]), .FEAT_BELOW(feature_belows[853])) ac853(.scan_win(scan_win853), .scan_win_std_dev(scan_win_std_dev[853]), .feature_accum(feature_accums[853]));
  accum_calculator #(.RECT1_X(rectangle1_xs[854]), .RECT1_Y(rectangle1_ys[854]), .RECT1_WIDTH(rectangle1_widths[854]), .RECT1_HEIGHT(rectangle1_heights[854]), .RECT1_WEIGHT(rectangle1_weights[854]), .RECT2_X(rectangle2_xs[854]), .RECT2_Y(rectangle2_ys[854]), .RECT2_WIDTH(rectangle2_widths[854]), .RECT2_HEIGHT(rectangle2_heights[854]), .RECT2_WEIGHT(rectangle2_weights[854]), .RECT3_X(rectangle3_xs[854]), .RECT3_Y(rectangle3_ys[854]), .RECT3_WIDTH(rectangle3_widths[854]), .RECT3_HEIGHT(rectangle3_heights[854]), .RECT3_WEIGHT(rectangle3_weights[854]), .FEAT_THRES(feature_thresholds[854]), .FEAT_ABOVE(feature_aboves[854]), .FEAT_BELOW(feature_belows[854])) ac854(.scan_win(scan_win854), .scan_win_std_dev(scan_win_std_dev[854]), .feature_accum(feature_accums[854]));
  accum_calculator #(.RECT1_X(rectangle1_xs[855]), .RECT1_Y(rectangle1_ys[855]), .RECT1_WIDTH(rectangle1_widths[855]), .RECT1_HEIGHT(rectangle1_heights[855]), .RECT1_WEIGHT(rectangle1_weights[855]), .RECT2_X(rectangle2_xs[855]), .RECT2_Y(rectangle2_ys[855]), .RECT2_WIDTH(rectangle2_widths[855]), .RECT2_HEIGHT(rectangle2_heights[855]), .RECT2_WEIGHT(rectangle2_weights[855]), .RECT3_X(rectangle3_xs[855]), .RECT3_Y(rectangle3_ys[855]), .RECT3_WIDTH(rectangle3_widths[855]), .RECT3_HEIGHT(rectangle3_heights[855]), .RECT3_WEIGHT(rectangle3_weights[855]), .FEAT_THRES(feature_thresholds[855]), .FEAT_ABOVE(feature_aboves[855]), .FEAT_BELOW(feature_belows[855])) ac855(.scan_win(scan_win855), .scan_win_std_dev(scan_win_std_dev[855]), .feature_accum(feature_accums[855]));
  accum_calculator #(.RECT1_X(rectangle1_xs[856]), .RECT1_Y(rectangle1_ys[856]), .RECT1_WIDTH(rectangle1_widths[856]), .RECT1_HEIGHT(rectangle1_heights[856]), .RECT1_WEIGHT(rectangle1_weights[856]), .RECT2_X(rectangle2_xs[856]), .RECT2_Y(rectangle2_ys[856]), .RECT2_WIDTH(rectangle2_widths[856]), .RECT2_HEIGHT(rectangle2_heights[856]), .RECT2_WEIGHT(rectangle2_weights[856]), .RECT3_X(rectangle3_xs[856]), .RECT3_Y(rectangle3_ys[856]), .RECT3_WIDTH(rectangle3_widths[856]), .RECT3_HEIGHT(rectangle3_heights[856]), .RECT3_WEIGHT(rectangle3_weights[856]), .FEAT_THRES(feature_thresholds[856]), .FEAT_ABOVE(feature_aboves[856]), .FEAT_BELOW(feature_belows[856])) ac856(.scan_win(scan_win856), .scan_win_std_dev(scan_win_std_dev[856]), .feature_accum(feature_accums[856]));
  accum_calculator #(.RECT1_X(rectangle1_xs[857]), .RECT1_Y(rectangle1_ys[857]), .RECT1_WIDTH(rectangle1_widths[857]), .RECT1_HEIGHT(rectangle1_heights[857]), .RECT1_WEIGHT(rectangle1_weights[857]), .RECT2_X(rectangle2_xs[857]), .RECT2_Y(rectangle2_ys[857]), .RECT2_WIDTH(rectangle2_widths[857]), .RECT2_HEIGHT(rectangle2_heights[857]), .RECT2_WEIGHT(rectangle2_weights[857]), .RECT3_X(rectangle3_xs[857]), .RECT3_Y(rectangle3_ys[857]), .RECT3_WIDTH(rectangle3_widths[857]), .RECT3_HEIGHT(rectangle3_heights[857]), .RECT3_WEIGHT(rectangle3_weights[857]), .FEAT_THRES(feature_thresholds[857]), .FEAT_ABOVE(feature_aboves[857]), .FEAT_BELOW(feature_belows[857])) ac857(.scan_win(scan_win857), .scan_win_std_dev(scan_win_std_dev[857]), .feature_accum(feature_accums[857]));
  accum_calculator #(.RECT1_X(rectangle1_xs[858]), .RECT1_Y(rectangle1_ys[858]), .RECT1_WIDTH(rectangle1_widths[858]), .RECT1_HEIGHT(rectangle1_heights[858]), .RECT1_WEIGHT(rectangle1_weights[858]), .RECT2_X(rectangle2_xs[858]), .RECT2_Y(rectangle2_ys[858]), .RECT2_WIDTH(rectangle2_widths[858]), .RECT2_HEIGHT(rectangle2_heights[858]), .RECT2_WEIGHT(rectangle2_weights[858]), .RECT3_X(rectangle3_xs[858]), .RECT3_Y(rectangle3_ys[858]), .RECT3_WIDTH(rectangle3_widths[858]), .RECT3_HEIGHT(rectangle3_heights[858]), .RECT3_WEIGHT(rectangle3_weights[858]), .FEAT_THRES(feature_thresholds[858]), .FEAT_ABOVE(feature_aboves[858]), .FEAT_BELOW(feature_belows[858])) ac858(.scan_win(scan_win858), .scan_win_std_dev(scan_win_std_dev[858]), .feature_accum(feature_accums[858]));
  accum_calculator #(.RECT1_X(rectangle1_xs[859]), .RECT1_Y(rectangle1_ys[859]), .RECT1_WIDTH(rectangle1_widths[859]), .RECT1_HEIGHT(rectangle1_heights[859]), .RECT1_WEIGHT(rectangle1_weights[859]), .RECT2_X(rectangle2_xs[859]), .RECT2_Y(rectangle2_ys[859]), .RECT2_WIDTH(rectangle2_widths[859]), .RECT2_HEIGHT(rectangle2_heights[859]), .RECT2_WEIGHT(rectangle2_weights[859]), .RECT3_X(rectangle3_xs[859]), .RECT3_Y(rectangle3_ys[859]), .RECT3_WIDTH(rectangle3_widths[859]), .RECT3_HEIGHT(rectangle3_heights[859]), .RECT3_WEIGHT(rectangle3_weights[859]), .FEAT_THRES(feature_thresholds[859]), .FEAT_ABOVE(feature_aboves[859]), .FEAT_BELOW(feature_belows[859])) ac859(.scan_win(scan_win859), .scan_win_std_dev(scan_win_std_dev[859]), .feature_accum(feature_accums[859]));
  accum_calculator #(.RECT1_X(rectangle1_xs[860]), .RECT1_Y(rectangle1_ys[860]), .RECT1_WIDTH(rectangle1_widths[860]), .RECT1_HEIGHT(rectangle1_heights[860]), .RECT1_WEIGHT(rectangle1_weights[860]), .RECT2_X(rectangle2_xs[860]), .RECT2_Y(rectangle2_ys[860]), .RECT2_WIDTH(rectangle2_widths[860]), .RECT2_HEIGHT(rectangle2_heights[860]), .RECT2_WEIGHT(rectangle2_weights[860]), .RECT3_X(rectangle3_xs[860]), .RECT3_Y(rectangle3_ys[860]), .RECT3_WIDTH(rectangle3_widths[860]), .RECT3_HEIGHT(rectangle3_heights[860]), .RECT3_WEIGHT(rectangle3_weights[860]), .FEAT_THRES(feature_thresholds[860]), .FEAT_ABOVE(feature_aboves[860]), .FEAT_BELOW(feature_belows[860])) ac860(.scan_win(scan_win860), .scan_win_std_dev(scan_win_std_dev[860]), .feature_accum(feature_accums[860]));
  accum_calculator #(.RECT1_X(rectangle1_xs[861]), .RECT1_Y(rectangle1_ys[861]), .RECT1_WIDTH(rectangle1_widths[861]), .RECT1_HEIGHT(rectangle1_heights[861]), .RECT1_WEIGHT(rectangle1_weights[861]), .RECT2_X(rectangle2_xs[861]), .RECT2_Y(rectangle2_ys[861]), .RECT2_WIDTH(rectangle2_widths[861]), .RECT2_HEIGHT(rectangle2_heights[861]), .RECT2_WEIGHT(rectangle2_weights[861]), .RECT3_X(rectangle3_xs[861]), .RECT3_Y(rectangle3_ys[861]), .RECT3_WIDTH(rectangle3_widths[861]), .RECT3_HEIGHT(rectangle3_heights[861]), .RECT3_WEIGHT(rectangle3_weights[861]), .FEAT_THRES(feature_thresholds[861]), .FEAT_ABOVE(feature_aboves[861]), .FEAT_BELOW(feature_belows[861])) ac861(.scan_win(scan_win861), .scan_win_std_dev(scan_win_std_dev[861]), .feature_accum(feature_accums[861]));
  accum_calculator #(.RECT1_X(rectangle1_xs[862]), .RECT1_Y(rectangle1_ys[862]), .RECT1_WIDTH(rectangle1_widths[862]), .RECT1_HEIGHT(rectangle1_heights[862]), .RECT1_WEIGHT(rectangle1_weights[862]), .RECT2_X(rectangle2_xs[862]), .RECT2_Y(rectangle2_ys[862]), .RECT2_WIDTH(rectangle2_widths[862]), .RECT2_HEIGHT(rectangle2_heights[862]), .RECT2_WEIGHT(rectangle2_weights[862]), .RECT3_X(rectangle3_xs[862]), .RECT3_Y(rectangle3_ys[862]), .RECT3_WIDTH(rectangle3_widths[862]), .RECT3_HEIGHT(rectangle3_heights[862]), .RECT3_WEIGHT(rectangle3_weights[862]), .FEAT_THRES(feature_thresholds[862]), .FEAT_ABOVE(feature_aboves[862]), .FEAT_BELOW(feature_belows[862])) ac862(.scan_win(scan_win862), .scan_win_std_dev(scan_win_std_dev[862]), .feature_accum(feature_accums[862]));
  accum_calculator #(.RECT1_X(rectangle1_xs[863]), .RECT1_Y(rectangle1_ys[863]), .RECT1_WIDTH(rectangle1_widths[863]), .RECT1_HEIGHT(rectangle1_heights[863]), .RECT1_WEIGHT(rectangle1_weights[863]), .RECT2_X(rectangle2_xs[863]), .RECT2_Y(rectangle2_ys[863]), .RECT2_WIDTH(rectangle2_widths[863]), .RECT2_HEIGHT(rectangle2_heights[863]), .RECT2_WEIGHT(rectangle2_weights[863]), .RECT3_X(rectangle3_xs[863]), .RECT3_Y(rectangle3_ys[863]), .RECT3_WIDTH(rectangle3_widths[863]), .RECT3_HEIGHT(rectangle3_heights[863]), .RECT3_WEIGHT(rectangle3_weights[863]), .FEAT_THRES(feature_thresholds[863]), .FEAT_ABOVE(feature_aboves[863]), .FEAT_BELOW(feature_belows[863])) ac863(.scan_win(scan_win863), .scan_win_std_dev(scan_win_std_dev[863]), .feature_accum(feature_accums[863]));
  accum_calculator #(.RECT1_X(rectangle1_xs[864]), .RECT1_Y(rectangle1_ys[864]), .RECT1_WIDTH(rectangle1_widths[864]), .RECT1_HEIGHT(rectangle1_heights[864]), .RECT1_WEIGHT(rectangle1_weights[864]), .RECT2_X(rectangle2_xs[864]), .RECT2_Y(rectangle2_ys[864]), .RECT2_WIDTH(rectangle2_widths[864]), .RECT2_HEIGHT(rectangle2_heights[864]), .RECT2_WEIGHT(rectangle2_weights[864]), .RECT3_X(rectangle3_xs[864]), .RECT3_Y(rectangle3_ys[864]), .RECT3_WIDTH(rectangle3_widths[864]), .RECT3_HEIGHT(rectangle3_heights[864]), .RECT3_WEIGHT(rectangle3_weights[864]), .FEAT_THRES(feature_thresholds[864]), .FEAT_ABOVE(feature_aboves[864]), .FEAT_BELOW(feature_belows[864])) ac864(.scan_win(scan_win864), .scan_win_std_dev(scan_win_std_dev[864]), .feature_accum(feature_accums[864]));
  accum_calculator #(.RECT1_X(rectangle1_xs[865]), .RECT1_Y(rectangle1_ys[865]), .RECT1_WIDTH(rectangle1_widths[865]), .RECT1_HEIGHT(rectangle1_heights[865]), .RECT1_WEIGHT(rectangle1_weights[865]), .RECT2_X(rectangle2_xs[865]), .RECT2_Y(rectangle2_ys[865]), .RECT2_WIDTH(rectangle2_widths[865]), .RECT2_HEIGHT(rectangle2_heights[865]), .RECT2_WEIGHT(rectangle2_weights[865]), .RECT3_X(rectangle3_xs[865]), .RECT3_Y(rectangle3_ys[865]), .RECT3_WIDTH(rectangle3_widths[865]), .RECT3_HEIGHT(rectangle3_heights[865]), .RECT3_WEIGHT(rectangle3_weights[865]), .FEAT_THRES(feature_thresholds[865]), .FEAT_ABOVE(feature_aboves[865]), .FEAT_BELOW(feature_belows[865])) ac865(.scan_win(scan_win865), .scan_win_std_dev(scan_win_std_dev[865]), .feature_accum(feature_accums[865]));
  accum_calculator #(.RECT1_X(rectangle1_xs[866]), .RECT1_Y(rectangle1_ys[866]), .RECT1_WIDTH(rectangle1_widths[866]), .RECT1_HEIGHT(rectangle1_heights[866]), .RECT1_WEIGHT(rectangle1_weights[866]), .RECT2_X(rectangle2_xs[866]), .RECT2_Y(rectangle2_ys[866]), .RECT2_WIDTH(rectangle2_widths[866]), .RECT2_HEIGHT(rectangle2_heights[866]), .RECT2_WEIGHT(rectangle2_weights[866]), .RECT3_X(rectangle3_xs[866]), .RECT3_Y(rectangle3_ys[866]), .RECT3_WIDTH(rectangle3_widths[866]), .RECT3_HEIGHT(rectangle3_heights[866]), .RECT3_WEIGHT(rectangle3_weights[866]), .FEAT_THRES(feature_thresholds[866]), .FEAT_ABOVE(feature_aboves[866]), .FEAT_BELOW(feature_belows[866])) ac866(.scan_win(scan_win866), .scan_win_std_dev(scan_win_std_dev[866]), .feature_accum(feature_accums[866]));
  accum_calculator #(.RECT1_X(rectangle1_xs[867]), .RECT1_Y(rectangle1_ys[867]), .RECT1_WIDTH(rectangle1_widths[867]), .RECT1_HEIGHT(rectangle1_heights[867]), .RECT1_WEIGHT(rectangle1_weights[867]), .RECT2_X(rectangle2_xs[867]), .RECT2_Y(rectangle2_ys[867]), .RECT2_WIDTH(rectangle2_widths[867]), .RECT2_HEIGHT(rectangle2_heights[867]), .RECT2_WEIGHT(rectangle2_weights[867]), .RECT3_X(rectangle3_xs[867]), .RECT3_Y(rectangle3_ys[867]), .RECT3_WIDTH(rectangle3_widths[867]), .RECT3_HEIGHT(rectangle3_heights[867]), .RECT3_WEIGHT(rectangle3_weights[867]), .FEAT_THRES(feature_thresholds[867]), .FEAT_ABOVE(feature_aboves[867]), .FEAT_BELOW(feature_belows[867])) ac867(.scan_win(scan_win867), .scan_win_std_dev(scan_win_std_dev[867]), .feature_accum(feature_accums[867]));
  accum_calculator #(.RECT1_X(rectangle1_xs[868]), .RECT1_Y(rectangle1_ys[868]), .RECT1_WIDTH(rectangle1_widths[868]), .RECT1_HEIGHT(rectangle1_heights[868]), .RECT1_WEIGHT(rectangle1_weights[868]), .RECT2_X(rectangle2_xs[868]), .RECT2_Y(rectangle2_ys[868]), .RECT2_WIDTH(rectangle2_widths[868]), .RECT2_HEIGHT(rectangle2_heights[868]), .RECT2_WEIGHT(rectangle2_weights[868]), .RECT3_X(rectangle3_xs[868]), .RECT3_Y(rectangle3_ys[868]), .RECT3_WIDTH(rectangle3_widths[868]), .RECT3_HEIGHT(rectangle3_heights[868]), .RECT3_WEIGHT(rectangle3_weights[868]), .FEAT_THRES(feature_thresholds[868]), .FEAT_ABOVE(feature_aboves[868]), .FEAT_BELOW(feature_belows[868])) ac868(.scan_win(scan_win868), .scan_win_std_dev(scan_win_std_dev[868]), .feature_accum(feature_accums[868]));
  accum_calculator #(.RECT1_X(rectangle1_xs[869]), .RECT1_Y(rectangle1_ys[869]), .RECT1_WIDTH(rectangle1_widths[869]), .RECT1_HEIGHT(rectangle1_heights[869]), .RECT1_WEIGHT(rectangle1_weights[869]), .RECT2_X(rectangle2_xs[869]), .RECT2_Y(rectangle2_ys[869]), .RECT2_WIDTH(rectangle2_widths[869]), .RECT2_HEIGHT(rectangle2_heights[869]), .RECT2_WEIGHT(rectangle2_weights[869]), .RECT3_X(rectangle3_xs[869]), .RECT3_Y(rectangle3_ys[869]), .RECT3_WIDTH(rectangle3_widths[869]), .RECT3_HEIGHT(rectangle3_heights[869]), .RECT3_WEIGHT(rectangle3_weights[869]), .FEAT_THRES(feature_thresholds[869]), .FEAT_ABOVE(feature_aboves[869]), .FEAT_BELOW(feature_belows[869])) ac869(.scan_win(scan_win869), .scan_win_std_dev(scan_win_std_dev[869]), .feature_accum(feature_accums[869]));
  accum_calculator #(.RECT1_X(rectangle1_xs[870]), .RECT1_Y(rectangle1_ys[870]), .RECT1_WIDTH(rectangle1_widths[870]), .RECT1_HEIGHT(rectangle1_heights[870]), .RECT1_WEIGHT(rectangle1_weights[870]), .RECT2_X(rectangle2_xs[870]), .RECT2_Y(rectangle2_ys[870]), .RECT2_WIDTH(rectangle2_widths[870]), .RECT2_HEIGHT(rectangle2_heights[870]), .RECT2_WEIGHT(rectangle2_weights[870]), .RECT3_X(rectangle3_xs[870]), .RECT3_Y(rectangle3_ys[870]), .RECT3_WIDTH(rectangle3_widths[870]), .RECT3_HEIGHT(rectangle3_heights[870]), .RECT3_WEIGHT(rectangle3_weights[870]), .FEAT_THRES(feature_thresholds[870]), .FEAT_ABOVE(feature_aboves[870]), .FEAT_BELOW(feature_belows[870])) ac870(.scan_win(scan_win870), .scan_win_std_dev(scan_win_std_dev[870]), .feature_accum(feature_accums[870]));
  accum_calculator #(.RECT1_X(rectangle1_xs[871]), .RECT1_Y(rectangle1_ys[871]), .RECT1_WIDTH(rectangle1_widths[871]), .RECT1_HEIGHT(rectangle1_heights[871]), .RECT1_WEIGHT(rectangle1_weights[871]), .RECT2_X(rectangle2_xs[871]), .RECT2_Y(rectangle2_ys[871]), .RECT2_WIDTH(rectangle2_widths[871]), .RECT2_HEIGHT(rectangle2_heights[871]), .RECT2_WEIGHT(rectangle2_weights[871]), .RECT3_X(rectangle3_xs[871]), .RECT3_Y(rectangle3_ys[871]), .RECT3_WIDTH(rectangle3_widths[871]), .RECT3_HEIGHT(rectangle3_heights[871]), .RECT3_WEIGHT(rectangle3_weights[871]), .FEAT_THRES(feature_thresholds[871]), .FEAT_ABOVE(feature_aboves[871]), .FEAT_BELOW(feature_belows[871])) ac871(.scan_win(scan_win871), .scan_win_std_dev(scan_win_std_dev[871]), .feature_accum(feature_accums[871]));
  accum_calculator #(.RECT1_X(rectangle1_xs[872]), .RECT1_Y(rectangle1_ys[872]), .RECT1_WIDTH(rectangle1_widths[872]), .RECT1_HEIGHT(rectangle1_heights[872]), .RECT1_WEIGHT(rectangle1_weights[872]), .RECT2_X(rectangle2_xs[872]), .RECT2_Y(rectangle2_ys[872]), .RECT2_WIDTH(rectangle2_widths[872]), .RECT2_HEIGHT(rectangle2_heights[872]), .RECT2_WEIGHT(rectangle2_weights[872]), .RECT3_X(rectangle3_xs[872]), .RECT3_Y(rectangle3_ys[872]), .RECT3_WIDTH(rectangle3_widths[872]), .RECT3_HEIGHT(rectangle3_heights[872]), .RECT3_WEIGHT(rectangle3_weights[872]), .FEAT_THRES(feature_thresholds[872]), .FEAT_ABOVE(feature_aboves[872]), .FEAT_BELOW(feature_belows[872])) ac872(.scan_win(scan_win872), .scan_win_std_dev(scan_win_std_dev[872]), .feature_accum(feature_accums[872]));
  accum_calculator #(.RECT1_X(rectangle1_xs[873]), .RECT1_Y(rectangle1_ys[873]), .RECT1_WIDTH(rectangle1_widths[873]), .RECT1_HEIGHT(rectangle1_heights[873]), .RECT1_WEIGHT(rectangle1_weights[873]), .RECT2_X(rectangle2_xs[873]), .RECT2_Y(rectangle2_ys[873]), .RECT2_WIDTH(rectangle2_widths[873]), .RECT2_HEIGHT(rectangle2_heights[873]), .RECT2_WEIGHT(rectangle2_weights[873]), .RECT3_X(rectangle3_xs[873]), .RECT3_Y(rectangle3_ys[873]), .RECT3_WIDTH(rectangle3_widths[873]), .RECT3_HEIGHT(rectangle3_heights[873]), .RECT3_WEIGHT(rectangle3_weights[873]), .FEAT_THRES(feature_thresholds[873]), .FEAT_ABOVE(feature_aboves[873]), .FEAT_BELOW(feature_belows[873])) ac873(.scan_win(scan_win873), .scan_win_std_dev(scan_win_std_dev[873]), .feature_accum(feature_accums[873]));
  accum_calculator #(.RECT1_X(rectangle1_xs[874]), .RECT1_Y(rectangle1_ys[874]), .RECT1_WIDTH(rectangle1_widths[874]), .RECT1_HEIGHT(rectangle1_heights[874]), .RECT1_WEIGHT(rectangle1_weights[874]), .RECT2_X(rectangle2_xs[874]), .RECT2_Y(rectangle2_ys[874]), .RECT2_WIDTH(rectangle2_widths[874]), .RECT2_HEIGHT(rectangle2_heights[874]), .RECT2_WEIGHT(rectangle2_weights[874]), .RECT3_X(rectangle3_xs[874]), .RECT3_Y(rectangle3_ys[874]), .RECT3_WIDTH(rectangle3_widths[874]), .RECT3_HEIGHT(rectangle3_heights[874]), .RECT3_WEIGHT(rectangle3_weights[874]), .FEAT_THRES(feature_thresholds[874]), .FEAT_ABOVE(feature_aboves[874]), .FEAT_BELOW(feature_belows[874])) ac874(.scan_win(scan_win874), .scan_win_std_dev(scan_win_std_dev[874]), .feature_accum(feature_accums[874]));
  accum_calculator #(.RECT1_X(rectangle1_xs[875]), .RECT1_Y(rectangle1_ys[875]), .RECT1_WIDTH(rectangle1_widths[875]), .RECT1_HEIGHT(rectangle1_heights[875]), .RECT1_WEIGHT(rectangle1_weights[875]), .RECT2_X(rectangle2_xs[875]), .RECT2_Y(rectangle2_ys[875]), .RECT2_WIDTH(rectangle2_widths[875]), .RECT2_HEIGHT(rectangle2_heights[875]), .RECT2_WEIGHT(rectangle2_weights[875]), .RECT3_X(rectangle3_xs[875]), .RECT3_Y(rectangle3_ys[875]), .RECT3_WIDTH(rectangle3_widths[875]), .RECT3_HEIGHT(rectangle3_heights[875]), .RECT3_WEIGHT(rectangle3_weights[875]), .FEAT_THRES(feature_thresholds[875]), .FEAT_ABOVE(feature_aboves[875]), .FEAT_BELOW(feature_belows[875])) ac875(.scan_win(scan_win875), .scan_win_std_dev(scan_win_std_dev[875]), .feature_accum(feature_accums[875]));
  accum_calculator #(.RECT1_X(rectangle1_xs[876]), .RECT1_Y(rectangle1_ys[876]), .RECT1_WIDTH(rectangle1_widths[876]), .RECT1_HEIGHT(rectangle1_heights[876]), .RECT1_WEIGHT(rectangle1_weights[876]), .RECT2_X(rectangle2_xs[876]), .RECT2_Y(rectangle2_ys[876]), .RECT2_WIDTH(rectangle2_widths[876]), .RECT2_HEIGHT(rectangle2_heights[876]), .RECT2_WEIGHT(rectangle2_weights[876]), .RECT3_X(rectangle3_xs[876]), .RECT3_Y(rectangle3_ys[876]), .RECT3_WIDTH(rectangle3_widths[876]), .RECT3_HEIGHT(rectangle3_heights[876]), .RECT3_WEIGHT(rectangle3_weights[876]), .FEAT_THRES(feature_thresholds[876]), .FEAT_ABOVE(feature_aboves[876]), .FEAT_BELOW(feature_belows[876])) ac876(.scan_win(scan_win876), .scan_win_std_dev(scan_win_std_dev[876]), .feature_accum(feature_accums[876]));
  accum_calculator #(.RECT1_X(rectangle1_xs[877]), .RECT1_Y(rectangle1_ys[877]), .RECT1_WIDTH(rectangle1_widths[877]), .RECT1_HEIGHT(rectangle1_heights[877]), .RECT1_WEIGHT(rectangle1_weights[877]), .RECT2_X(rectangle2_xs[877]), .RECT2_Y(rectangle2_ys[877]), .RECT2_WIDTH(rectangle2_widths[877]), .RECT2_HEIGHT(rectangle2_heights[877]), .RECT2_WEIGHT(rectangle2_weights[877]), .RECT3_X(rectangle3_xs[877]), .RECT3_Y(rectangle3_ys[877]), .RECT3_WIDTH(rectangle3_widths[877]), .RECT3_HEIGHT(rectangle3_heights[877]), .RECT3_WEIGHT(rectangle3_weights[877]), .FEAT_THRES(feature_thresholds[877]), .FEAT_ABOVE(feature_aboves[877]), .FEAT_BELOW(feature_belows[877])) ac877(.scan_win(scan_win877), .scan_win_std_dev(scan_win_std_dev[877]), .feature_accum(feature_accums[877]));
  accum_calculator #(.RECT1_X(rectangle1_xs[878]), .RECT1_Y(rectangle1_ys[878]), .RECT1_WIDTH(rectangle1_widths[878]), .RECT1_HEIGHT(rectangle1_heights[878]), .RECT1_WEIGHT(rectangle1_weights[878]), .RECT2_X(rectangle2_xs[878]), .RECT2_Y(rectangle2_ys[878]), .RECT2_WIDTH(rectangle2_widths[878]), .RECT2_HEIGHT(rectangle2_heights[878]), .RECT2_WEIGHT(rectangle2_weights[878]), .RECT3_X(rectangle3_xs[878]), .RECT3_Y(rectangle3_ys[878]), .RECT3_WIDTH(rectangle3_widths[878]), .RECT3_HEIGHT(rectangle3_heights[878]), .RECT3_WEIGHT(rectangle3_weights[878]), .FEAT_THRES(feature_thresholds[878]), .FEAT_ABOVE(feature_aboves[878]), .FEAT_BELOW(feature_belows[878])) ac878(.scan_win(scan_win878), .scan_win_std_dev(scan_win_std_dev[878]), .feature_accum(feature_accums[878]));
  accum_calculator #(.RECT1_X(rectangle1_xs[879]), .RECT1_Y(rectangle1_ys[879]), .RECT1_WIDTH(rectangle1_widths[879]), .RECT1_HEIGHT(rectangle1_heights[879]), .RECT1_WEIGHT(rectangle1_weights[879]), .RECT2_X(rectangle2_xs[879]), .RECT2_Y(rectangle2_ys[879]), .RECT2_WIDTH(rectangle2_widths[879]), .RECT2_HEIGHT(rectangle2_heights[879]), .RECT2_WEIGHT(rectangle2_weights[879]), .RECT3_X(rectangle3_xs[879]), .RECT3_Y(rectangle3_ys[879]), .RECT3_WIDTH(rectangle3_widths[879]), .RECT3_HEIGHT(rectangle3_heights[879]), .RECT3_WEIGHT(rectangle3_weights[879]), .FEAT_THRES(feature_thresholds[879]), .FEAT_ABOVE(feature_aboves[879]), .FEAT_BELOW(feature_belows[879])) ac879(.scan_win(scan_win879), .scan_win_std_dev(scan_win_std_dev[879]), .feature_accum(feature_accums[879]));
  accum_calculator #(.RECT1_X(rectangle1_xs[880]), .RECT1_Y(rectangle1_ys[880]), .RECT1_WIDTH(rectangle1_widths[880]), .RECT1_HEIGHT(rectangle1_heights[880]), .RECT1_WEIGHT(rectangle1_weights[880]), .RECT2_X(rectangle2_xs[880]), .RECT2_Y(rectangle2_ys[880]), .RECT2_WIDTH(rectangle2_widths[880]), .RECT2_HEIGHT(rectangle2_heights[880]), .RECT2_WEIGHT(rectangle2_weights[880]), .RECT3_X(rectangle3_xs[880]), .RECT3_Y(rectangle3_ys[880]), .RECT3_WIDTH(rectangle3_widths[880]), .RECT3_HEIGHT(rectangle3_heights[880]), .RECT3_WEIGHT(rectangle3_weights[880]), .FEAT_THRES(feature_thresholds[880]), .FEAT_ABOVE(feature_aboves[880]), .FEAT_BELOW(feature_belows[880])) ac880(.scan_win(scan_win880), .scan_win_std_dev(scan_win_std_dev[880]), .feature_accum(feature_accums[880]));
  accum_calculator #(.RECT1_X(rectangle1_xs[881]), .RECT1_Y(rectangle1_ys[881]), .RECT1_WIDTH(rectangle1_widths[881]), .RECT1_HEIGHT(rectangle1_heights[881]), .RECT1_WEIGHT(rectangle1_weights[881]), .RECT2_X(rectangle2_xs[881]), .RECT2_Y(rectangle2_ys[881]), .RECT2_WIDTH(rectangle2_widths[881]), .RECT2_HEIGHT(rectangle2_heights[881]), .RECT2_WEIGHT(rectangle2_weights[881]), .RECT3_X(rectangle3_xs[881]), .RECT3_Y(rectangle3_ys[881]), .RECT3_WIDTH(rectangle3_widths[881]), .RECT3_HEIGHT(rectangle3_heights[881]), .RECT3_WEIGHT(rectangle3_weights[881]), .FEAT_THRES(feature_thresholds[881]), .FEAT_ABOVE(feature_aboves[881]), .FEAT_BELOW(feature_belows[881])) ac881(.scan_win(scan_win881), .scan_win_std_dev(scan_win_std_dev[881]), .feature_accum(feature_accums[881]));
  accum_calculator #(.RECT1_X(rectangle1_xs[882]), .RECT1_Y(rectangle1_ys[882]), .RECT1_WIDTH(rectangle1_widths[882]), .RECT1_HEIGHT(rectangle1_heights[882]), .RECT1_WEIGHT(rectangle1_weights[882]), .RECT2_X(rectangle2_xs[882]), .RECT2_Y(rectangle2_ys[882]), .RECT2_WIDTH(rectangle2_widths[882]), .RECT2_HEIGHT(rectangle2_heights[882]), .RECT2_WEIGHT(rectangle2_weights[882]), .RECT3_X(rectangle3_xs[882]), .RECT3_Y(rectangle3_ys[882]), .RECT3_WIDTH(rectangle3_widths[882]), .RECT3_HEIGHT(rectangle3_heights[882]), .RECT3_WEIGHT(rectangle3_weights[882]), .FEAT_THRES(feature_thresholds[882]), .FEAT_ABOVE(feature_aboves[882]), .FEAT_BELOW(feature_belows[882])) ac882(.scan_win(scan_win882), .scan_win_std_dev(scan_win_std_dev[882]), .feature_accum(feature_accums[882]));
  accum_calculator #(.RECT1_X(rectangle1_xs[883]), .RECT1_Y(rectangle1_ys[883]), .RECT1_WIDTH(rectangle1_widths[883]), .RECT1_HEIGHT(rectangle1_heights[883]), .RECT1_WEIGHT(rectangle1_weights[883]), .RECT2_X(rectangle2_xs[883]), .RECT2_Y(rectangle2_ys[883]), .RECT2_WIDTH(rectangle2_widths[883]), .RECT2_HEIGHT(rectangle2_heights[883]), .RECT2_WEIGHT(rectangle2_weights[883]), .RECT3_X(rectangle3_xs[883]), .RECT3_Y(rectangle3_ys[883]), .RECT3_WIDTH(rectangle3_widths[883]), .RECT3_HEIGHT(rectangle3_heights[883]), .RECT3_WEIGHT(rectangle3_weights[883]), .FEAT_THRES(feature_thresholds[883]), .FEAT_ABOVE(feature_aboves[883]), .FEAT_BELOW(feature_belows[883])) ac883(.scan_win(scan_win883), .scan_win_std_dev(scan_win_std_dev[883]), .feature_accum(feature_accums[883]));
  accum_calculator #(.RECT1_X(rectangle1_xs[884]), .RECT1_Y(rectangle1_ys[884]), .RECT1_WIDTH(rectangle1_widths[884]), .RECT1_HEIGHT(rectangle1_heights[884]), .RECT1_WEIGHT(rectangle1_weights[884]), .RECT2_X(rectangle2_xs[884]), .RECT2_Y(rectangle2_ys[884]), .RECT2_WIDTH(rectangle2_widths[884]), .RECT2_HEIGHT(rectangle2_heights[884]), .RECT2_WEIGHT(rectangle2_weights[884]), .RECT3_X(rectangle3_xs[884]), .RECT3_Y(rectangle3_ys[884]), .RECT3_WIDTH(rectangle3_widths[884]), .RECT3_HEIGHT(rectangle3_heights[884]), .RECT3_WEIGHT(rectangle3_weights[884]), .FEAT_THRES(feature_thresholds[884]), .FEAT_ABOVE(feature_aboves[884]), .FEAT_BELOW(feature_belows[884])) ac884(.scan_win(scan_win884), .scan_win_std_dev(scan_win_std_dev[884]), .feature_accum(feature_accums[884]));
  accum_calculator #(.RECT1_X(rectangle1_xs[885]), .RECT1_Y(rectangle1_ys[885]), .RECT1_WIDTH(rectangle1_widths[885]), .RECT1_HEIGHT(rectangle1_heights[885]), .RECT1_WEIGHT(rectangle1_weights[885]), .RECT2_X(rectangle2_xs[885]), .RECT2_Y(rectangle2_ys[885]), .RECT2_WIDTH(rectangle2_widths[885]), .RECT2_HEIGHT(rectangle2_heights[885]), .RECT2_WEIGHT(rectangle2_weights[885]), .RECT3_X(rectangle3_xs[885]), .RECT3_Y(rectangle3_ys[885]), .RECT3_WIDTH(rectangle3_widths[885]), .RECT3_HEIGHT(rectangle3_heights[885]), .RECT3_WEIGHT(rectangle3_weights[885]), .FEAT_THRES(feature_thresholds[885]), .FEAT_ABOVE(feature_aboves[885]), .FEAT_BELOW(feature_belows[885])) ac885(.scan_win(scan_win885), .scan_win_std_dev(scan_win_std_dev[885]), .feature_accum(feature_accums[885]));
  accum_calculator #(.RECT1_X(rectangle1_xs[886]), .RECT1_Y(rectangle1_ys[886]), .RECT1_WIDTH(rectangle1_widths[886]), .RECT1_HEIGHT(rectangle1_heights[886]), .RECT1_WEIGHT(rectangle1_weights[886]), .RECT2_X(rectangle2_xs[886]), .RECT2_Y(rectangle2_ys[886]), .RECT2_WIDTH(rectangle2_widths[886]), .RECT2_HEIGHT(rectangle2_heights[886]), .RECT2_WEIGHT(rectangle2_weights[886]), .RECT3_X(rectangle3_xs[886]), .RECT3_Y(rectangle3_ys[886]), .RECT3_WIDTH(rectangle3_widths[886]), .RECT3_HEIGHT(rectangle3_heights[886]), .RECT3_WEIGHT(rectangle3_weights[886]), .FEAT_THRES(feature_thresholds[886]), .FEAT_ABOVE(feature_aboves[886]), .FEAT_BELOW(feature_belows[886])) ac886(.scan_win(scan_win886), .scan_win_std_dev(scan_win_std_dev[886]), .feature_accum(feature_accums[886]));
  accum_calculator #(.RECT1_X(rectangle1_xs[887]), .RECT1_Y(rectangle1_ys[887]), .RECT1_WIDTH(rectangle1_widths[887]), .RECT1_HEIGHT(rectangle1_heights[887]), .RECT1_WEIGHT(rectangle1_weights[887]), .RECT2_X(rectangle2_xs[887]), .RECT2_Y(rectangle2_ys[887]), .RECT2_WIDTH(rectangle2_widths[887]), .RECT2_HEIGHT(rectangle2_heights[887]), .RECT2_WEIGHT(rectangle2_weights[887]), .RECT3_X(rectangle3_xs[887]), .RECT3_Y(rectangle3_ys[887]), .RECT3_WIDTH(rectangle3_widths[887]), .RECT3_HEIGHT(rectangle3_heights[887]), .RECT3_WEIGHT(rectangle3_weights[887]), .FEAT_THRES(feature_thresholds[887]), .FEAT_ABOVE(feature_aboves[887]), .FEAT_BELOW(feature_belows[887])) ac887(.scan_win(scan_win887), .scan_win_std_dev(scan_win_std_dev[887]), .feature_accum(feature_accums[887]));
  accum_calculator #(.RECT1_X(rectangle1_xs[888]), .RECT1_Y(rectangle1_ys[888]), .RECT1_WIDTH(rectangle1_widths[888]), .RECT1_HEIGHT(rectangle1_heights[888]), .RECT1_WEIGHT(rectangle1_weights[888]), .RECT2_X(rectangle2_xs[888]), .RECT2_Y(rectangle2_ys[888]), .RECT2_WIDTH(rectangle2_widths[888]), .RECT2_HEIGHT(rectangle2_heights[888]), .RECT2_WEIGHT(rectangle2_weights[888]), .RECT3_X(rectangle3_xs[888]), .RECT3_Y(rectangle3_ys[888]), .RECT3_WIDTH(rectangle3_widths[888]), .RECT3_HEIGHT(rectangle3_heights[888]), .RECT3_WEIGHT(rectangle3_weights[888]), .FEAT_THRES(feature_thresholds[888]), .FEAT_ABOVE(feature_aboves[888]), .FEAT_BELOW(feature_belows[888])) ac888(.scan_win(scan_win888), .scan_win_std_dev(scan_win_std_dev[888]), .feature_accum(feature_accums[888]));
  accum_calculator #(.RECT1_X(rectangle1_xs[889]), .RECT1_Y(rectangle1_ys[889]), .RECT1_WIDTH(rectangle1_widths[889]), .RECT1_HEIGHT(rectangle1_heights[889]), .RECT1_WEIGHT(rectangle1_weights[889]), .RECT2_X(rectangle2_xs[889]), .RECT2_Y(rectangle2_ys[889]), .RECT2_WIDTH(rectangle2_widths[889]), .RECT2_HEIGHT(rectangle2_heights[889]), .RECT2_WEIGHT(rectangle2_weights[889]), .RECT3_X(rectangle3_xs[889]), .RECT3_Y(rectangle3_ys[889]), .RECT3_WIDTH(rectangle3_widths[889]), .RECT3_HEIGHT(rectangle3_heights[889]), .RECT3_WEIGHT(rectangle3_weights[889]), .FEAT_THRES(feature_thresholds[889]), .FEAT_ABOVE(feature_aboves[889]), .FEAT_BELOW(feature_belows[889])) ac889(.scan_win(scan_win889), .scan_win_std_dev(scan_win_std_dev[889]), .feature_accum(feature_accums[889]));
  accum_calculator #(.RECT1_X(rectangle1_xs[890]), .RECT1_Y(rectangle1_ys[890]), .RECT1_WIDTH(rectangle1_widths[890]), .RECT1_HEIGHT(rectangle1_heights[890]), .RECT1_WEIGHT(rectangle1_weights[890]), .RECT2_X(rectangle2_xs[890]), .RECT2_Y(rectangle2_ys[890]), .RECT2_WIDTH(rectangle2_widths[890]), .RECT2_HEIGHT(rectangle2_heights[890]), .RECT2_WEIGHT(rectangle2_weights[890]), .RECT3_X(rectangle3_xs[890]), .RECT3_Y(rectangle3_ys[890]), .RECT3_WIDTH(rectangle3_widths[890]), .RECT3_HEIGHT(rectangle3_heights[890]), .RECT3_WEIGHT(rectangle3_weights[890]), .FEAT_THRES(feature_thresholds[890]), .FEAT_ABOVE(feature_aboves[890]), .FEAT_BELOW(feature_belows[890])) ac890(.scan_win(scan_win890), .scan_win_std_dev(scan_win_std_dev[890]), .feature_accum(feature_accums[890]));
  accum_calculator #(.RECT1_X(rectangle1_xs[891]), .RECT1_Y(rectangle1_ys[891]), .RECT1_WIDTH(rectangle1_widths[891]), .RECT1_HEIGHT(rectangle1_heights[891]), .RECT1_WEIGHT(rectangle1_weights[891]), .RECT2_X(rectangle2_xs[891]), .RECT2_Y(rectangle2_ys[891]), .RECT2_WIDTH(rectangle2_widths[891]), .RECT2_HEIGHT(rectangle2_heights[891]), .RECT2_WEIGHT(rectangle2_weights[891]), .RECT3_X(rectangle3_xs[891]), .RECT3_Y(rectangle3_ys[891]), .RECT3_WIDTH(rectangle3_widths[891]), .RECT3_HEIGHT(rectangle3_heights[891]), .RECT3_WEIGHT(rectangle3_weights[891]), .FEAT_THRES(feature_thresholds[891]), .FEAT_ABOVE(feature_aboves[891]), .FEAT_BELOW(feature_belows[891])) ac891(.scan_win(scan_win891), .scan_win_std_dev(scan_win_std_dev[891]), .feature_accum(feature_accums[891]));
  accum_calculator #(.RECT1_X(rectangle1_xs[892]), .RECT1_Y(rectangle1_ys[892]), .RECT1_WIDTH(rectangle1_widths[892]), .RECT1_HEIGHT(rectangle1_heights[892]), .RECT1_WEIGHT(rectangle1_weights[892]), .RECT2_X(rectangle2_xs[892]), .RECT2_Y(rectangle2_ys[892]), .RECT2_WIDTH(rectangle2_widths[892]), .RECT2_HEIGHT(rectangle2_heights[892]), .RECT2_WEIGHT(rectangle2_weights[892]), .RECT3_X(rectangle3_xs[892]), .RECT3_Y(rectangle3_ys[892]), .RECT3_WIDTH(rectangle3_widths[892]), .RECT3_HEIGHT(rectangle3_heights[892]), .RECT3_WEIGHT(rectangle3_weights[892]), .FEAT_THRES(feature_thresholds[892]), .FEAT_ABOVE(feature_aboves[892]), .FEAT_BELOW(feature_belows[892])) ac892(.scan_win(scan_win892), .scan_win_std_dev(scan_win_std_dev[892]), .feature_accum(feature_accums[892]));
  accum_calculator #(.RECT1_X(rectangle1_xs[893]), .RECT1_Y(rectangle1_ys[893]), .RECT1_WIDTH(rectangle1_widths[893]), .RECT1_HEIGHT(rectangle1_heights[893]), .RECT1_WEIGHT(rectangle1_weights[893]), .RECT2_X(rectangle2_xs[893]), .RECT2_Y(rectangle2_ys[893]), .RECT2_WIDTH(rectangle2_widths[893]), .RECT2_HEIGHT(rectangle2_heights[893]), .RECT2_WEIGHT(rectangle2_weights[893]), .RECT3_X(rectangle3_xs[893]), .RECT3_Y(rectangle3_ys[893]), .RECT3_WIDTH(rectangle3_widths[893]), .RECT3_HEIGHT(rectangle3_heights[893]), .RECT3_WEIGHT(rectangle3_weights[893]), .FEAT_THRES(feature_thresholds[893]), .FEAT_ABOVE(feature_aboves[893]), .FEAT_BELOW(feature_belows[893])) ac893(.scan_win(scan_win893), .scan_win_std_dev(scan_win_std_dev[893]), .feature_accum(feature_accums[893]));
  accum_calculator #(.RECT1_X(rectangle1_xs[894]), .RECT1_Y(rectangle1_ys[894]), .RECT1_WIDTH(rectangle1_widths[894]), .RECT1_HEIGHT(rectangle1_heights[894]), .RECT1_WEIGHT(rectangle1_weights[894]), .RECT2_X(rectangle2_xs[894]), .RECT2_Y(rectangle2_ys[894]), .RECT2_WIDTH(rectangle2_widths[894]), .RECT2_HEIGHT(rectangle2_heights[894]), .RECT2_WEIGHT(rectangle2_weights[894]), .RECT3_X(rectangle3_xs[894]), .RECT3_Y(rectangle3_ys[894]), .RECT3_WIDTH(rectangle3_widths[894]), .RECT3_HEIGHT(rectangle3_heights[894]), .RECT3_WEIGHT(rectangle3_weights[894]), .FEAT_THRES(feature_thresholds[894]), .FEAT_ABOVE(feature_aboves[894]), .FEAT_BELOW(feature_belows[894])) ac894(.scan_win(scan_win894), .scan_win_std_dev(scan_win_std_dev[894]), .feature_accum(feature_accums[894]));
  accum_calculator #(.RECT1_X(rectangle1_xs[895]), .RECT1_Y(rectangle1_ys[895]), .RECT1_WIDTH(rectangle1_widths[895]), .RECT1_HEIGHT(rectangle1_heights[895]), .RECT1_WEIGHT(rectangle1_weights[895]), .RECT2_X(rectangle2_xs[895]), .RECT2_Y(rectangle2_ys[895]), .RECT2_WIDTH(rectangle2_widths[895]), .RECT2_HEIGHT(rectangle2_heights[895]), .RECT2_WEIGHT(rectangle2_weights[895]), .RECT3_X(rectangle3_xs[895]), .RECT3_Y(rectangle3_ys[895]), .RECT3_WIDTH(rectangle3_widths[895]), .RECT3_HEIGHT(rectangle3_heights[895]), .RECT3_WEIGHT(rectangle3_weights[895]), .FEAT_THRES(feature_thresholds[895]), .FEAT_ABOVE(feature_aboves[895]), .FEAT_BELOW(feature_belows[895])) ac895(.scan_win(scan_win895), .scan_win_std_dev(scan_win_std_dev[895]), .feature_accum(feature_accums[895]));
  accum_calculator #(.RECT1_X(rectangle1_xs[896]), .RECT1_Y(rectangle1_ys[896]), .RECT1_WIDTH(rectangle1_widths[896]), .RECT1_HEIGHT(rectangle1_heights[896]), .RECT1_WEIGHT(rectangle1_weights[896]), .RECT2_X(rectangle2_xs[896]), .RECT2_Y(rectangle2_ys[896]), .RECT2_WIDTH(rectangle2_widths[896]), .RECT2_HEIGHT(rectangle2_heights[896]), .RECT2_WEIGHT(rectangle2_weights[896]), .RECT3_X(rectangle3_xs[896]), .RECT3_Y(rectangle3_ys[896]), .RECT3_WIDTH(rectangle3_widths[896]), .RECT3_HEIGHT(rectangle3_heights[896]), .RECT3_WEIGHT(rectangle3_weights[896]), .FEAT_THRES(feature_thresholds[896]), .FEAT_ABOVE(feature_aboves[896]), .FEAT_BELOW(feature_belows[896])) ac896(.scan_win(scan_win896), .scan_win_std_dev(scan_win_std_dev[896]), .feature_accum(feature_accums[896]));
  accum_calculator #(.RECT1_X(rectangle1_xs[897]), .RECT1_Y(rectangle1_ys[897]), .RECT1_WIDTH(rectangle1_widths[897]), .RECT1_HEIGHT(rectangle1_heights[897]), .RECT1_WEIGHT(rectangle1_weights[897]), .RECT2_X(rectangle2_xs[897]), .RECT2_Y(rectangle2_ys[897]), .RECT2_WIDTH(rectangle2_widths[897]), .RECT2_HEIGHT(rectangle2_heights[897]), .RECT2_WEIGHT(rectangle2_weights[897]), .RECT3_X(rectangle3_xs[897]), .RECT3_Y(rectangle3_ys[897]), .RECT3_WIDTH(rectangle3_widths[897]), .RECT3_HEIGHT(rectangle3_heights[897]), .RECT3_WEIGHT(rectangle3_weights[897]), .FEAT_THRES(feature_thresholds[897]), .FEAT_ABOVE(feature_aboves[897]), .FEAT_BELOW(feature_belows[897])) ac897(.scan_win(scan_win897), .scan_win_std_dev(scan_win_std_dev[897]), .feature_accum(feature_accums[897]));
  accum_calculator #(.RECT1_X(rectangle1_xs[898]), .RECT1_Y(rectangle1_ys[898]), .RECT1_WIDTH(rectangle1_widths[898]), .RECT1_HEIGHT(rectangle1_heights[898]), .RECT1_WEIGHT(rectangle1_weights[898]), .RECT2_X(rectangle2_xs[898]), .RECT2_Y(rectangle2_ys[898]), .RECT2_WIDTH(rectangle2_widths[898]), .RECT2_HEIGHT(rectangle2_heights[898]), .RECT2_WEIGHT(rectangle2_weights[898]), .RECT3_X(rectangle3_xs[898]), .RECT3_Y(rectangle3_ys[898]), .RECT3_WIDTH(rectangle3_widths[898]), .RECT3_HEIGHT(rectangle3_heights[898]), .RECT3_WEIGHT(rectangle3_weights[898]), .FEAT_THRES(feature_thresholds[898]), .FEAT_ABOVE(feature_aboves[898]), .FEAT_BELOW(feature_belows[898])) ac898(.scan_win(scan_win898), .scan_win_std_dev(scan_win_std_dev[898]), .feature_accum(feature_accums[898]));
  accum_calculator #(.RECT1_X(rectangle1_xs[899]), .RECT1_Y(rectangle1_ys[899]), .RECT1_WIDTH(rectangle1_widths[899]), .RECT1_HEIGHT(rectangle1_heights[899]), .RECT1_WEIGHT(rectangle1_weights[899]), .RECT2_X(rectangle2_xs[899]), .RECT2_Y(rectangle2_ys[899]), .RECT2_WIDTH(rectangle2_widths[899]), .RECT2_HEIGHT(rectangle2_heights[899]), .RECT2_WEIGHT(rectangle2_weights[899]), .RECT3_X(rectangle3_xs[899]), .RECT3_Y(rectangle3_ys[899]), .RECT3_WIDTH(rectangle3_widths[899]), .RECT3_HEIGHT(rectangle3_heights[899]), .RECT3_WEIGHT(rectangle3_weights[899]), .FEAT_THRES(feature_thresholds[899]), .FEAT_ABOVE(feature_aboves[899]), .FEAT_BELOW(feature_belows[899])) ac899(.scan_win(scan_win899), .scan_win_std_dev(scan_win_std_dev[899]), .feature_accum(feature_accums[899]));
  accum_calculator #(.RECT1_X(rectangle1_xs[900]), .RECT1_Y(rectangle1_ys[900]), .RECT1_WIDTH(rectangle1_widths[900]), .RECT1_HEIGHT(rectangle1_heights[900]), .RECT1_WEIGHT(rectangle1_weights[900]), .RECT2_X(rectangle2_xs[900]), .RECT2_Y(rectangle2_ys[900]), .RECT2_WIDTH(rectangle2_widths[900]), .RECT2_HEIGHT(rectangle2_heights[900]), .RECT2_WEIGHT(rectangle2_weights[900]), .RECT3_X(rectangle3_xs[900]), .RECT3_Y(rectangle3_ys[900]), .RECT3_WIDTH(rectangle3_widths[900]), .RECT3_HEIGHT(rectangle3_heights[900]), .RECT3_WEIGHT(rectangle3_weights[900]), .FEAT_THRES(feature_thresholds[900]), .FEAT_ABOVE(feature_aboves[900]), .FEAT_BELOW(feature_belows[900])) ac900(.scan_win(scan_win900), .scan_win_std_dev(scan_win_std_dev[900]), .feature_accum(feature_accums[900]));
  accum_calculator #(.RECT1_X(rectangle1_xs[901]), .RECT1_Y(rectangle1_ys[901]), .RECT1_WIDTH(rectangle1_widths[901]), .RECT1_HEIGHT(rectangle1_heights[901]), .RECT1_WEIGHT(rectangle1_weights[901]), .RECT2_X(rectangle2_xs[901]), .RECT2_Y(rectangle2_ys[901]), .RECT2_WIDTH(rectangle2_widths[901]), .RECT2_HEIGHT(rectangle2_heights[901]), .RECT2_WEIGHT(rectangle2_weights[901]), .RECT3_X(rectangle3_xs[901]), .RECT3_Y(rectangle3_ys[901]), .RECT3_WIDTH(rectangle3_widths[901]), .RECT3_HEIGHT(rectangle3_heights[901]), .RECT3_WEIGHT(rectangle3_weights[901]), .FEAT_THRES(feature_thresholds[901]), .FEAT_ABOVE(feature_aboves[901]), .FEAT_BELOW(feature_belows[901])) ac901(.scan_win(scan_win901), .scan_win_std_dev(scan_win_std_dev[901]), .feature_accum(feature_accums[901]));
  accum_calculator #(.RECT1_X(rectangle1_xs[902]), .RECT1_Y(rectangle1_ys[902]), .RECT1_WIDTH(rectangle1_widths[902]), .RECT1_HEIGHT(rectangle1_heights[902]), .RECT1_WEIGHT(rectangle1_weights[902]), .RECT2_X(rectangle2_xs[902]), .RECT2_Y(rectangle2_ys[902]), .RECT2_WIDTH(rectangle2_widths[902]), .RECT2_HEIGHT(rectangle2_heights[902]), .RECT2_WEIGHT(rectangle2_weights[902]), .RECT3_X(rectangle3_xs[902]), .RECT3_Y(rectangle3_ys[902]), .RECT3_WIDTH(rectangle3_widths[902]), .RECT3_HEIGHT(rectangle3_heights[902]), .RECT3_WEIGHT(rectangle3_weights[902]), .FEAT_THRES(feature_thresholds[902]), .FEAT_ABOVE(feature_aboves[902]), .FEAT_BELOW(feature_belows[902])) ac902(.scan_win(scan_win902), .scan_win_std_dev(scan_win_std_dev[902]), .feature_accum(feature_accums[902]));
  accum_calculator #(.RECT1_X(rectangle1_xs[903]), .RECT1_Y(rectangle1_ys[903]), .RECT1_WIDTH(rectangle1_widths[903]), .RECT1_HEIGHT(rectangle1_heights[903]), .RECT1_WEIGHT(rectangle1_weights[903]), .RECT2_X(rectangle2_xs[903]), .RECT2_Y(rectangle2_ys[903]), .RECT2_WIDTH(rectangle2_widths[903]), .RECT2_HEIGHT(rectangle2_heights[903]), .RECT2_WEIGHT(rectangle2_weights[903]), .RECT3_X(rectangle3_xs[903]), .RECT3_Y(rectangle3_ys[903]), .RECT3_WIDTH(rectangle3_widths[903]), .RECT3_HEIGHT(rectangle3_heights[903]), .RECT3_WEIGHT(rectangle3_weights[903]), .FEAT_THRES(feature_thresholds[903]), .FEAT_ABOVE(feature_aboves[903]), .FEAT_BELOW(feature_belows[903])) ac903(.scan_win(scan_win903), .scan_win_std_dev(scan_win_std_dev[903]), .feature_accum(feature_accums[903]));
  accum_calculator #(.RECT1_X(rectangle1_xs[904]), .RECT1_Y(rectangle1_ys[904]), .RECT1_WIDTH(rectangle1_widths[904]), .RECT1_HEIGHT(rectangle1_heights[904]), .RECT1_WEIGHT(rectangle1_weights[904]), .RECT2_X(rectangle2_xs[904]), .RECT2_Y(rectangle2_ys[904]), .RECT2_WIDTH(rectangle2_widths[904]), .RECT2_HEIGHT(rectangle2_heights[904]), .RECT2_WEIGHT(rectangle2_weights[904]), .RECT3_X(rectangle3_xs[904]), .RECT3_Y(rectangle3_ys[904]), .RECT3_WIDTH(rectangle3_widths[904]), .RECT3_HEIGHT(rectangle3_heights[904]), .RECT3_WEIGHT(rectangle3_weights[904]), .FEAT_THRES(feature_thresholds[904]), .FEAT_ABOVE(feature_aboves[904]), .FEAT_BELOW(feature_belows[904])) ac904(.scan_win(scan_win904), .scan_win_std_dev(scan_win_std_dev[904]), .feature_accum(feature_accums[904]));
  accum_calculator #(.RECT1_X(rectangle1_xs[905]), .RECT1_Y(rectangle1_ys[905]), .RECT1_WIDTH(rectangle1_widths[905]), .RECT1_HEIGHT(rectangle1_heights[905]), .RECT1_WEIGHT(rectangle1_weights[905]), .RECT2_X(rectangle2_xs[905]), .RECT2_Y(rectangle2_ys[905]), .RECT2_WIDTH(rectangle2_widths[905]), .RECT2_HEIGHT(rectangle2_heights[905]), .RECT2_WEIGHT(rectangle2_weights[905]), .RECT3_X(rectangle3_xs[905]), .RECT3_Y(rectangle3_ys[905]), .RECT3_WIDTH(rectangle3_widths[905]), .RECT3_HEIGHT(rectangle3_heights[905]), .RECT3_WEIGHT(rectangle3_weights[905]), .FEAT_THRES(feature_thresholds[905]), .FEAT_ABOVE(feature_aboves[905]), .FEAT_BELOW(feature_belows[905])) ac905(.scan_win(scan_win905), .scan_win_std_dev(scan_win_std_dev[905]), .feature_accum(feature_accums[905]));
  accum_calculator #(.RECT1_X(rectangle1_xs[906]), .RECT1_Y(rectangle1_ys[906]), .RECT1_WIDTH(rectangle1_widths[906]), .RECT1_HEIGHT(rectangle1_heights[906]), .RECT1_WEIGHT(rectangle1_weights[906]), .RECT2_X(rectangle2_xs[906]), .RECT2_Y(rectangle2_ys[906]), .RECT2_WIDTH(rectangle2_widths[906]), .RECT2_HEIGHT(rectangle2_heights[906]), .RECT2_WEIGHT(rectangle2_weights[906]), .RECT3_X(rectangle3_xs[906]), .RECT3_Y(rectangle3_ys[906]), .RECT3_WIDTH(rectangle3_widths[906]), .RECT3_HEIGHT(rectangle3_heights[906]), .RECT3_WEIGHT(rectangle3_weights[906]), .FEAT_THRES(feature_thresholds[906]), .FEAT_ABOVE(feature_aboves[906]), .FEAT_BELOW(feature_belows[906])) ac906(.scan_win(scan_win906), .scan_win_std_dev(scan_win_std_dev[906]), .feature_accum(feature_accums[906]));
  accum_calculator #(.RECT1_X(rectangle1_xs[907]), .RECT1_Y(rectangle1_ys[907]), .RECT1_WIDTH(rectangle1_widths[907]), .RECT1_HEIGHT(rectangle1_heights[907]), .RECT1_WEIGHT(rectangle1_weights[907]), .RECT2_X(rectangle2_xs[907]), .RECT2_Y(rectangle2_ys[907]), .RECT2_WIDTH(rectangle2_widths[907]), .RECT2_HEIGHT(rectangle2_heights[907]), .RECT2_WEIGHT(rectangle2_weights[907]), .RECT3_X(rectangle3_xs[907]), .RECT3_Y(rectangle3_ys[907]), .RECT3_WIDTH(rectangle3_widths[907]), .RECT3_HEIGHT(rectangle3_heights[907]), .RECT3_WEIGHT(rectangle3_weights[907]), .FEAT_THRES(feature_thresholds[907]), .FEAT_ABOVE(feature_aboves[907]), .FEAT_BELOW(feature_belows[907])) ac907(.scan_win(scan_win907), .scan_win_std_dev(scan_win_std_dev[907]), .feature_accum(feature_accums[907]));
  accum_calculator #(.RECT1_X(rectangle1_xs[908]), .RECT1_Y(rectangle1_ys[908]), .RECT1_WIDTH(rectangle1_widths[908]), .RECT1_HEIGHT(rectangle1_heights[908]), .RECT1_WEIGHT(rectangle1_weights[908]), .RECT2_X(rectangle2_xs[908]), .RECT2_Y(rectangle2_ys[908]), .RECT2_WIDTH(rectangle2_widths[908]), .RECT2_HEIGHT(rectangle2_heights[908]), .RECT2_WEIGHT(rectangle2_weights[908]), .RECT3_X(rectangle3_xs[908]), .RECT3_Y(rectangle3_ys[908]), .RECT3_WIDTH(rectangle3_widths[908]), .RECT3_HEIGHT(rectangle3_heights[908]), .RECT3_WEIGHT(rectangle3_weights[908]), .FEAT_THRES(feature_thresholds[908]), .FEAT_ABOVE(feature_aboves[908]), .FEAT_BELOW(feature_belows[908])) ac908(.scan_win(scan_win908), .scan_win_std_dev(scan_win_std_dev[908]), .feature_accum(feature_accums[908]));
  accum_calculator #(.RECT1_X(rectangle1_xs[909]), .RECT1_Y(rectangle1_ys[909]), .RECT1_WIDTH(rectangle1_widths[909]), .RECT1_HEIGHT(rectangle1_heights[909]), .RECT1_WEIGHT(rectangle1_weights[909]), .RECT2_X(rectangle2_xs[909]), .RECT2_Y(rectangle2_ys[909]), .RECT2_WIDTH(rectangle2_widths[909]), .RECT2_HEIGHT(rectangle2_heights[909]), .RECT2_WEIGHT(rectangle2_weights[909]), .RECT3_X(rectangle3_xs[909]), .RECT3_Y(rectangle3_ys[909]), .RECT3_WIDTH(rectangle3_widths[909]), .RECT3_HEIGHT(rectangle3_heights[909]), .RECT3_WEIGHT(rectangle3_weights[909]), .FEAT_THRES(feature_thresholds[909]), .FEAT_ABOVE(feature_aboves[909]), .FEAT_BELOW(feature_belows[909])) ac909(.scan_win(scan_win909), .scan_win_std_dev(scan_win_std_dev[909]), .feature_accum(feature_accums[909]));
  accum_calculator #(.RECT1_X(rectangle1_xs[910]), .RECT1_Y(rectangle1_ys[910]), .RECT1_WIDTH(rectangle1_widths[910]), .RECT1_HEIGHT(rectangle1_heights[910]), .RECT1_WEIGHT(rectangle1_weights[910]), .RECT2_X(rectangle2_xs[910]), .RECT2_Y(rectangle2_ys[910]), .RECT2_WIDTH(rectangle2_widths[910]), .RECT2_HEIGHT(rectangle2_heights[910]), .RECT2_WEIGHT(rectangle2_weights[910]), .RECT3_X(rectangle3_xs[910]), .RECT3_Y(rectangle3_ys[910]), .RECT3_WIDTH(rectangle3_widths[910]), .RECT3_HEIGHT(rectangle3_heights[910]), .RECT3_WEIGHT(rectangle3_weights[910]), .FEAT_THRES(feature_thresholds[910]), .FEAT_ABOVE(feature_aboves[910]), .FEAT_BELOW(feature_belows[910])) ac910(.scan_win(scan_win910), .scan_win_std_dev(scan_win_std_dev[910]), .feature_accum(feature_accums[910]));
  accum_calculator #(.RECT1_X(rectangle1_xs[911]), .RECT1_Y(rectangle1_ys[911]), .RECT1_WIDTH(rectangle1_widths[911]), .RECT1_HEIGHT(rectangle1_heights[911]), .RECT1_WEIGHT(rectangle1_weights[911]), .RECT2_X(rectangle2_xs[911]), .RECT2_Y(rectangle2_ys[911]), .RECT2_WIDTH(rectangle2_widths[911]), .RECT2_HEIGHT(rectangle2_heights[911]), .RECT2_WEIGHT(rectangle2_weights[911]), .RECT3_X(rectangle3_xs[911]), .RECT3_Y(rectangle3_ys[911]), .RECT3_WIDTH(rectangle3_widths[911]), .RECT3_HEIGHT(rectangle3_heights[911]), .RECT3_WEIGHT(rectangle3_weights[911]), .FEAT_THRES(feature_thresholds[911]), .FEAT_ABOVE(feature_aboves[911]), .FEAT_BELOW(feature_belows[911])) ac911(.scan_win(scan_win911), .scan_win_std_dev(scan_win_std_dev[911]), .feature_accum(feature_accums[911]));
  accum_calculator #(.RECT1_X(rectangle1_xs[912]), .RECT1_Y(rectangle1_ys[912]), .RECT1_WIDTH(rectangle1_widths[912]), .RECT1_HEIGHT(rectangle1_heights[912]), .RECT1_WEIGHT(rectangle1_weights[912]), .RECT2_X(rectangle2_xs[912]), .RECT2_Y(rectangle2_ys[912]), .RECT2_WIDTH(rectangle2_widths[912]), .RECT2_HEIGHT(rectangle2_heights[912]), .RECT2_WEIGHT(rectangle2_weights[912]), .RECT3_X(rectangle3_xs[912]), .RECT3_Y(rectangle3_ys[912]), .RECT3_WIDTH(rectangle3_widths[912]), .RECT3_HEIGHT(rectangle3_heights[912]), .RECT3_WEIGHT(rectangle3_weights[912]), .FEAT_THRES(feature_thresholds[912]), .FEAT_ABOVE(feature_aboves[912]), .FEAT_BELOW(feature_belows[912])) ac912(.scan_win(scan_win912), .scan_win_std_dev(scan_win_std_dev[912]), .feature_accum(feature_accums[912]));
  accum_calculator #(.RECT1_X(rectangle1_xs[913]), .RECT1_Y(rectangle1_ys[913]), .RECT1_WIDTH(rectangle1_widths[913]), .RECT1_HEIGHT(rectangle1_heights[913]), .RECT1_WEIGHT(rectangle1_weights[913]), .RECT2_X(rectangle2_xs[913]), .RECT2_Y(rectangle2_ys[913]), .RECT2_WIDTH(rectangle2_widths[913]), .RECT2_HEIGHT(rectangle2_heights[913]), .RECT2_WEIGHT(rectangle2_weights[913]), .RECT3_X(rectangle3_xs[913]), .RECT3_Y(rectangle3_ys[913]), .RECT3_WIDTH(rectangle3_widths[913]), .RECT3_HEIGHT(rectangle3_heights[913]), .RECT3_WEIGHT(rectangle3_weights[913]), .FEAT_THRES(feature_thresholds[913]), .FEAT_ABOVE(feature_aboves[913]), .FEAT_BELOW(feature_belows[913])) ac913(.scan_win(scan_win913), .scan_win_std_dev(scan_win_std_dev[913]), .feature_accum(feature_accums[913]));
  accum_calculator #(.RECT1_X(rectangle1_xs[914]), .RECT1_Y(rectangle1_ys[914]), .RECT1_WIDTH(rectangle1_widths[914]), .RECT1_HEIGHT(rectangle1_heights[914]), .RECT1_WEIGHT(rectangle1_weights[914]), .RECT2_X(rectangle2_xs[914]), .RECT2_Y(rectangle2_ys[914]), .RECT2_WIDTH(rectangle2_widths[914]), .RECT2_HEIGHT(rectangle2_heights[914]), .RECT2_WEIGHT(rectangle2_weights[914]), .RECT3_X(rectangle3_xs[914]), .RECT3_Y(rectangle3_ys[914]), .RECT3_WIDTH(rectangle3_widths[914]), .RECT3_HEIGHT(rectangle3_heights[914]), .RECT3_WEIGHT(rectangle3_weights[914]), .FEAT_THRES(feature_thresholds[914]), .FEAT_ABOVE(feature_aboves[914]), .FEAT_BELOW(feature_belows[914])) ac914(.scan_win(scan_win914), .scan_win_std_dev(scan_win_std_dev[914]), .feature_accum(feature_accums[914]));
  accum_calculator #(.RECT1_X(rectangle1_xs[915]), .RECT1_Y(rectangle1_ys[915]), .RECT1_WIDTH(rectangle1_widths[915]), .RECT1_HEIGHT(rectangle1_heights[915]), .RECT1_WEIGHT(rectangle1_weights[915]), .RECT2_X(rectangle2_xs[915]), .RECT2_Y(rectangle2_ys[915]), .RECT2_WIDTH(rectangle2_widths[915]), .RECT2_HEIGHT(rectangle2_heights[915]), .RECT2_WEIGHT(rectangle2_weights[915]), .RECT3_X(rectangle3_xs[915]), .RECT3_Y(rectangle3_ys[915]), .RECT3_WIDTH(rectangle3_widths[915]), .RECT3_HEIGHT(rectangle3_heights[915]), .RECT3_WEIGHT(rectangle3_weights[915]), .FEAT_THRES(feature_thresholds[915]), .FEAT_ABOVE(feature_aboves[915]), .FEAT_BELOW(feature_belows[915])) ac915(.scan_win(scan_win915), .scan_win_std_dev(scan_win_std_dev[915]), .feature_accum(feature_accums[915]));
  accum_calculator #(.RECT1_X(rectangle1_xs[916]), .RECT1_Y(rectangle1_ys[916]), .RECT1_WIDTH(rectangle1_widths[916]), .RECT1_HEIGHT(rectangle1_heights[916]), .RECT1_WEIGHT(rectangle1_weights[916]), .RECT2_X(rectangle2_xs[916]), .RECT2_Y(rectangle2_ys[916]), .RECT2_WIDTH(rectangle2_widths[916]), .RECT2_HEIGHT(rectangle2_heights[916]), .RECT2_WEIGHT(rectangle2_weights[916]), .RECT3_X(rectangle3_xs[916]), .RECT3_Y(rectangle3_ys[916]), .RECT3_WIDTH(rectangle3_widths[916]), .RECT3_HEIGHT(rectangle3_heights[916]), .RECT3_WEIGHT(rectangle3_weights[916]), .FEAT_THRES(feature_thresholds[916]), .FEAT_ABOVE(feature_aboves[916]), .FEAT_BELOW(feature_belows[916])) ac916(.scan_win(scan_win916), .scan_win_std_dev(scan_win_std_dev[916]), .feature_accum(feature_accums[916]));
  accum_calculator #(.RECT1_X(rectangle1_xs[917]), .RECT1_Y(rectangle1_ys[917]), .RECT1_WIDTH(rectangle1_widths[917]), .RECT1_HEIGHT(rectangle1_heights[917]), .RECT1_WEIGHT(rectangle1_weights[917]), .RECT2_X(rectangle2_xs[917]), .RECT2_Y(rectangle2_ys[917]), .RECT2_WIDTH(rectangle2_widths[917]), .RECT2_HEIGHT(rectangle2_heights[917]), .RECT2_WEIGHT(rectangle2_weights[917]), .RECT3_X(rectangle3_xs[917]), .RECT3_Y(rectangle3_ys[917]), .RECT3_WIDTH(rectangle3_widths[917]), .RECT3_HEIGHT(rectangle3_heights[917]), .RECT3_WEIGHT(rectangle3_weights[917]), .FEAT_THRES(feature_thresholds[917]), .FEAT_ABOVE(feature_aboves[917]), .FEAT_BELOW(feature_belows[917])) ac917(.scan_win(scan_win917), .scan_win_std_dev(scan_win_std_dev[917]), .feature_accum(feature_accums[917]));
  accum_calculator #(.RECT1_X(rectangle1_xs[918]), .RECT1_Y(rectangle1_ys[918]), .RECT1_WIDTH(rectangle1_widths[918]), .RECT1_HEIGHT(rectangle1_heights[918]), .RECT1_WEIGHT(rectangle1_weights[918]), .RECT2_X(rectangle2_xs[918]), .RECT2_Y(rectangle2_ys[918]), .RECT2_WIDTH(rectangle2_widths[918]), .RECT2_HEIGHT(rectangle2_heights[918]), .RECT2_WEIGHT(rectangle2_weights[918]), .RECT3_X(rectangle3_xs[918]), .RECT3_Y(rectangle3_ys[918]), .RECT3_WIDTH(rectangle3_widths[918]), .RECT3_HEIGHT(rectangle3_heights[918]), .RECT3_WEIGHT(rectangle3_weights[918]), .FEAT_THRES(feature_thresholds[918]), .FEAT_ABOVE(feature_aboves[918]), .FEAT_BELOW(feature_belows[918])) ac918(.scan_win(scan_win918), .scan_win_std_dev(scan_win_std_dev[918]), .feature_accum(feature_accums[918]));
  accum_calculator #(.RECT1_X(rectangle1_xs[919]), .RECT1_Y(rectangle1_ys[919]), .RECT1_WIDTH(rectangle1_widths[919]), .RECT1_HEIGHT(rectangle1_heights[919]), .RECT1_WEIGHT(rectangle1_weights[919]), .RECT2_X(rectangle2_xs[919]), .RECT2_Y(rectangle2_ys[919]), .RECT2_WIDTH(rectangle2_widths[919]), .RECT2_HEIGHT(rectangle2_heights[919]), .RECT2_WEIGHT(rectangle2_weights[919]), .RECT3_X(rectangle3_xs[919]), .RECT3_Y(rectangle3_ys[919]), .RECT3_WIDTH(rectangle3_widths[919]), .RECT3_HEIGHT(rectangle3_heights[919]), .RECT3_WEIGHT(rectangle3_weights[919]), .FEAT_THRES(feature_thresholds[919]), .FEAT_ABOVE(feature_aboves[919]), .FEAT_BELOW(feature_belows[919])) ac919(.scan_win(scan_win919), .scan_win_std_dev(scan_win_std_dev[919]), .feature_accum(feature_accums[919]));
  accum_calculator #(.RECT1_X(rectangle1_xs[920]), .RECT1_Y(rectangle1_ys[920]), .RECT1_WIDTH(rectangle1_widths[920]), .RECT1_HEIGHT(rectangle1_heights[920]), .RECT1_WEIGHT(rectangle1_weights[920]), .RECT2_X(rectangle2_xs[920]), .RECT2_Y(rectangle2_ys[920]), .RECT2_WIDTH(rectangle2_widths[920]), .RECT2_HEIGHT(rectangle2_heights[920]), .RECT2_WEIGHT(rectangle2_weights[920]), .RECT3_X(rectangle3_xs[920]), .RECT3_Y(rectangle3_ys[920]), .RECT3_WIDTH(rectangle3_widths[920]), .RECT3_HEIGHT(rectangle3_heights[920]), .RECT3_WEIGHT(rectangle3_weights[920]), .FEAT_THRES(feature_thresholds[920]), .FEAT_ABOVE(feature_aboves[920]), .FEAT_BELOW(feature_belows[920])) ac920(.scan_win(scan_win920), .scan_win_std_dev(scan_win_std_dev[920]), .feature_accum(feature_accums[920]));
  accum_calculator #(.RECT1_X(rectangle1_xs[921]), .RECT1_Y(rectangle1_ys[921]), .RECT1_WIDTH(rectangle1_widths[921]), .RECT1_HEIGHT(rectangle1_heights[921]), .RECT1_WEIGHT(rectangle1_weights[921]), .RECT2_X(rectangle2_xs[921]), .RECT2_Y(rectangle2_ys[921]), .RECT2_WIDTH(rectangle2_widths[921]), .RECT2_HEIGHT(rectangle2_heights[921]), .RECT2_WEIGHT(rectangle2_weights[921]), .RECT3_X(rectangle3_xs[921]), .RECT3_Y(rectangle3_ys[921]), .RECT3_WIDTH(rectangle3_widths[921]), .RECT3_HEIGHT(rectangle3_heights[921]), .RECT3_WEIGHT(rectangle3_weights[921]), .FEAT_THRES(feature_thresholds[921]), .FEAT_ABOVE(feature_aboves[921]), .FEAT_BELOW(feature_belows[921])) ac921(.scan_win(scan_win921), .scan_win_std_dev(scan_win_std_dev[921]), .feature_accum(feature_accums[921]));
  accum_calculator #(.RECT1_X(rectangle1_xs[922]), .RECT1_Y(rectangle1_ys[922]), .RECT1_WIDTH(rectangle1_widths[922]), .RECT1_HEIGHT(rectangle1_heights[922]), .RECT1_WEIGHT(rectangle1_weights[922]), .RECT2_X(rectangle2_xs[922]), .RECT2_Y(rectangle2_ys[922]), .RECT2_WIDTH(rectangle2_widths[922]), .RECT2_HEIGHT(rectangle2_heights[922]), .RECT2_WEIGHT(rectangle2_weights[922]), .RECT3_X(rectangle3_xs[922]), .RECT3_Y(rectangle3_ys[922]), .RECT3_WIDTH(rectangle3_widths[922]), .RECT3_HEIGHT(rectangle3_heights[922]), .RECT3_WEIGHT(rectangle3_weights[922]), .FEAT_THRES(feature_thresholds[922]), .FEAT_ABOVE(feature_aboves[922]), .FEAT_BELOW(feature_belows[922])) ac922(.scan_win(scan_win922), .scan_win_std_dev(scan_win_std_dev[922]), .feature_accum(feature_accums[922]));
  accum_calculator #(.RECT1_X(rectangle1_xs[923]), .RECT1_Y(rectangle1_ys[923]), .RECT1_WIDTH(rectangle1_widths[923]), .RECT1_HEIGHT(rectangle1_heights[923]), .RECT1_WEIGHT(rectangle1_weights[923]), .RECT2_X(rectangle2_xs[923]), .RECT2_Y(rectangle2_ys[923]), .RECT2_WIDTH(rectangle2_widths[923]), .RECT2_HEIGHT(rectangle2_heights[923]), .RECT2_WEIGHT(rectangle2_weights[923]), .RECT3_X(rectangle3_xs[923]), .RECT3_Y(rectangle3_ys[923]), .RECT3_WIDTH(rectangle3_widths[923]), .RECT3_HEIGHT(rectangle3_heights[923]), .RECT3_WEIGHT(rectangle3_weights[923]), .FEAT_THRES(feature_thresholds[923]), .FEAT_ABOVE(feature_aboves[923]), .FEAT_BELOW(feature_belows[923])) ac923(.scan_win(scan_win923), .scan_win_std_dev(scan_win_std_dev[923]), .feature_accum(feature_accums[923]));
  accum_calculator #(.RECT1_X(rectangle1_xs[924]), .RECT1_Y(rectangle1_ys[924]), .RECT1_WIDTH(rectangle1_widths[924]), .RECT1_HEIGHT(rectangle1_heights[924]), .RECT1_WEIGHT(rectangle1_weights[924]), .RECT2_X(rectangle2_xs[924]), .RECT2_Y(rectangle2_ys[924]), .RECT2_WIDTH(rectangle2_widths[924]), .RECT2_HEIGHT(rectangle2_heights[924]), .RECT2_WEIGHT(rectangle2_weights[924]), .RECT3_X(rectangle3_xs[924]), .RECT3_Y(rectangle3_ys[924]), .RECT3_WIDTH(rectangle3_widths[924]), .RECT3_HEIGHT(rectangle3_heights[924]), .RECT3_WEIGHT(rectangle3_weights[924]), .FEAT_THRES(feature_thresholds[924]), .FEAT_ABOVE(feature_aboves[924]), .FEAT_BELOW(feature_belows[924])) ac924(.scan_win(scan_win924), .scan_win_std_dev(scan_win_std_dev[924]), .feature_accum(feature_accums[924]));
  accum_calculator #(.RECT1_X(rectangle1_xs[925]), .RECT1_Y(rectangle1_ys[925]), .RECT1_WIDTH(rectangle1_widths[925]), .RECT1_HEIGHT(rectangle1_heights[925]), .RECT1_WEIGHT(rectangle1_weights[925]), .RECT2_X(rectangle2_xs[925]), .RECT2_Y(rectangle2_ys[925]), .RECT2_WIDTH(rectangle2_widths[925]), .RECT2_HEIGHT(rectangle2_heights[925]), .RECT2_WEIGHT(rectangle2_weights[925]), .RECT3_X(rectangle3_xs[925]), .RECT3_Y(rectangle3_ys[925]), .RECT3_WIDTH(rectangle3_widths[925]), .RECT3_HEIGHT(rectangle3_heights[925]), .RECT3_WEIGHT(rectangle3_weights[925]), .FEAT_THRES(feature_thresholds[925]), .FEAT_ABOVE(feature_aboves[925]), .FEAT_BELOW(feature_belows[925])) ac925(.scan_win(scan_win925), .scan_win_std_dev(scan_win_std_dev[925]), .feature_accum(feature_accums[925]));
  accum_calculator #(.RECT1_X(rectangle1_xs[926]), .RECT1_Y(rectangle1_ys[926]), .RECT1_WIDTH(rectangle1_widths[926]), .RECT1_HEIGHT(rectangle1_heights[926]), .RECT1_WEIGHT(rectangle1_weights[926]), .RECT2_X(rectangle2_xs[926]), .RECT2_Y(rectangle2_ys[926]), .RECT2_WIDTH(rectangle2_widths[926]), .RECT2_HEIGHT(rectangle2_heights[926]), .RECT2_WEIGHT(rectangle2_weights[926]), .RECT3_X(rectangle3_xs[926]), .RECT3_Y(rectangle3_ys[926]), .RECT3_WIDTH(rectangle3_widths[926]), .RECT3_HEIGHT(rectangle3_heights[926]), .RECT3_WEIGHT(rectangle3_weights[926]), .FEAT_THRES(feature_thresholds[926]), .FEAT_ABOVE(feature_aboves[926]), .FEAT_BELOW(feature_belows[926])) ac926(.scan_win(scan_win926), .scan_win_std_dev(scan_win_std_dev[926]), .feature_accum(feature_accums[926]));
  accum_calculator #(.RECT1_X(rectangle1_xs[927]), .RECT1_Y(rectangle1_ys[927]), .RECT1_WIDTH(rectangle1_widths[927]), .RECT1_HEIGHT(rectangle1_heights[927]), .RECT1_WEIGHT(rectangle1_weights[927]), .RECT2_X(rectangle2_xs[927]), .RECT2_Y(rectangle2_ys[927]), .RECT2_WIDTH(rectangle2_widths[927]), .RECT2_HEIGHT(rectangle2_heights[927]), .RECT2_WEIGHT(rectangle2_weights[927]), .RECT3_X(rectangle3_xs[927]), .RECT3_Y(rectangle3_ys[927]), .RECT3_WIDTH(rectangle3_widths[927]), .RECT3_HEIGHT(rectangle3_heights[927]), .RECT3_WEIGHT(rectangle3_weights[927]), .FEAT_THRES(feature_thresholds[927]), .FEAT_ABOVE(feature_aboves[927]), .FEAT_BELOW(feature_belows[927])) ac927(.scan_win(scan_win927), .scan_win_std_dev(scan_win_std_dev[927]), .feature_accum(feature_accums[927]));
  accum_calculator #(.RECT1_X(rectangle1_xs[928]), .RECT1_Y(rectangle1_ys[928]), .RECT1_WIDTH(rectangle1_widths[928]), .RECT1_HEIGHT(rectangle1_heights[928]), .RECT1_WEIGHT(rectangle1_weights[928]), .RECT2_X(rectangle2_xs[928]), .RECT2_Y(rectangle2_ys[928]), .RECT2_WIDTH(rectangle2_widths[928]), .RECT2_HEIGHT(rectangle2_heights[928]), .RECT2_WEIGHT(rectangle2_weights[928]), .RECT3_X(rectangle3_xs[928]), .RECT3_Y(rectangle3_ys[928]), .RECT3_WIDTH(rectangle3_widths[928]), .RECT3_HEIGHT(rectangle3_heights[928]), .RECT3_WEIGHT(rectangle3_weights[928]), .FEAT_THRES(feature_thresholds[928]), .FEAT_ABOVE(feature_aboves[928]), .FEAT_BELOW(feature_belows[928])) ac928(.scan_win(scan_win928), .scan_win_std_dev(scan_win_std_dev[928]), .feature_accum(feature_accums[928]));
  accum_calculator #(.RECT1_X(rectangle1_xs[929]), .RECT1_Y(rectangle1_ys[929]), .RECT1_WIDTH(rectangle1_widths[929]), .RECT1_HEIGHT(rectangle1_heights[929]), .RECT1_WEIGHT(rectangle1_weights[929]), .RECT2_X(rectangle2_xs[929]), .RECT2_Y(rectangle2_ys[929]), .RECT2_WIDTH(rectangle2_widths[929]), .RECT2_HEIGHT(rectangle2_heights[929]), .RECT2_WEIGHT(rectangle2_weights[929]), .RECT3_X(rectangle3_xs[929]), .RECT3_Y(rectangle3_ys[929]), .RECT3_WIDTH(rectangle3_widths[929]), .RECT3_HEIGHT(rectangle3_heights[929]), .RECT3_WEIGHT(rectangle3_weights[929]), .FEAT_THRES(feature_thresholds[929]), .FEAT_ABOVE(feature_aboves[929]), .FEAT_BELOW(feature_belows[929])) ac929(.scan_win(scan_win929), .scan_win_std_dev(scan_win_std_dev[929]), .feature_accum(feature_accums[929]));
  accum_calculator #(.RECT1_X(rectangle1_xs[930]), .RECT1_Y(rectangle1_ys[930]), .RECT1_WIDTH(rectangle1_widths[930]), .RECT1_HEIGHT(rectangle1_heights[930]), .RECT1_WEIGHT(rectangle1_weights[930]), .RECT2_X(rectangle2_xs[930]), .RECT2_Y(rectangle2_ys[930]), .RECT2_WIDTH(rectangle2_widths[930]), .RECT2_HEIGHT(rectangle2_heights[930]), .RECT2_WEIGHT(rectangle2_weights[930]), .RECT3_X(rectangle3_xs[930]), .RECT3_Y(rectangle3_ys[930]), .RECT3_WIDTH(rectangle3_widths[930]), .RECT3_HEIGHT(rectangle3_heights[930]), .RECT3_WEIGHT(rectangle3_weights[930]), .FEAT_THRES(feature_thresholds[930]), .FEAT_ABOVE(feature_aboves[930]), .FEAT_BELOW(feature_belows[930])) ac930(.scan_win(scan_win930), .scan_win_std_dev(scan_win_std_dev[930]), .feature_accum(feature_accums[930]));
  accum_calculator #(.RECT1_X(rectangle1_xs[931]), .RECT1_Y(rectangle1_ys[931]), .RECT1_WIDTH(rectangle1_widths[931]), .RECT1_HEIGHT(rectangle1_heights[931]), .RECT1_WEIGHT(rectangle1_weights[931]), .RECT2_X(rectangle2_xs[931]), .RECT2_Y(rectangle2_ys[931]), .RECT2_WIDTH(rectangle2_widths[931]), .RECT2_HEIGHT(rectangle2_heights[931]), .RECT2_WEIGHT(rectangle2_weights[931]), .RECT3_X(rectangle3_xs[931]), .RECT3_Y(rectangle3_ys[931]), .RECT3_WIDTH(rectangle3_widths[931]), .RECT3_HEIGHT(rectangle3_heights[931]), .RECT3_WEIGHT(rectangle3_weights[931]), .FEAT_THRES(feature_thresholds[931]), .FEAT_ABOVE(feature_aboves[931]), .FEAT_BELOW(feature_belows[931])) ac931(.scan_win(scan_win931), .scan_win_std_dev(scan_win_std_dev[931]), .feature_accum(feature_accums[931]));
  accum_calculator #(.RECT1_X(rectangle1_xs[932]), .RECT1_Y(rectangle1_ys[932]), .RECT1_WIDTH(rectangle1_widths[932]), .RECT1_HEIGHT(rectangle1_heights[932]), .RECT1_WEIGHT(rectangle1_weights[932]), .RECT2_X(rectangle2_xs[932]), .RECT2_Y(rectangle2_ys[932]), .RECT2_WIDTH(rectangle2_widths[932]), .RECT2_HEIGHT(rectangle2_heights[932]), .RECT2_WEIGHT(rectangle2_weights[932]), .RECT3_X(rectangle3_xs[932]), .RECT3_Y(rectangle3_ys[932]), .RECT3_WIDTH(rectangle3_widths[932]), .RECT3_HEIGHT(rectangle3_heights[932]), .RECT3_WEIGHT(rectangle3_weights[932]), .FEAT_THRES(feature_thresholds[932]), .FEAT_ABOVE(feature_aboves[932]), .FEAT_BELOW(feature_belows[932])) ac932(.scan_win(scan_win932), .scan_win_std_dev(scan_win_std_dev[932]), .feature_accum(feature_accums[932]));
  accum_calculator #(.RECT1_X(rectangle1_xs[933]), .RECT1_Y(rectangle1_ys[933]), .RECT1_WIDTH(rectangle1_widths[933]), .RECT1_HEIGHT(rectangle1_heights[933]), .RECT1_WEIGHT(rectangle1_weights[933]), .RECT2_X(rectangle2_xs[933]), .RECT2_Y(rectangle2_ys[933]), .RECT2_WIDTH(rectangle2_widths[933]), .RECT2_HEIGHT(rectangle2_heights[933]), .RECT2_WEIGHT(rectangle2_weights[933]), .RECT3_X(rectangle3_xs[933]), .RECT3_Y(rectangle3_ys[933]), .RECT3_WIDTH(rectangle3_widths[933]), .RECT3_HEIGHT(rectangle3_heights[933]), .RECT3_WEIGHT(rectangle3_weights[933]), .FEAT_THRES(feature_thresholds[933]), .FEAT_ABOVE(feature_aboves[933]), .FEAT_BELOW(feature_belows[933])) ac933(.scan_win(scan_win933), .scan_win_std_dev(scan_win_std_dev[933]), .feature_accum(feature_accums[933]));
  accum_calculator #(.RECT1_X(rectangle1_xs[934]), .RECT1_Y(rectangle1_ys[934]), .RECT1_WIDTH(rectangle1_widths[934]), .RECT1_HEIGHT(rectangle1_heights[934]), .RECT1_WEIGHT(rectangle1_weights[934]), .RECT2_X(rectangle2_xs[934]), .RECT2_Y(rectangle2_ys[934]), .RECT2_WIDTH(rectangle2_widths[934]), .RECT2_HEIGHT(rectangle2_heights[934]), .RECT2_WEIGHT(rectangle2_weights[934]), .RECT3_X(rectangle3_xs[934]), .RECT3_Y(rectangle3_ys[934]), .RECT3_WIDTH(rectangle3_widths[934]), .RECT3_HEIGHT(rectangle3_heights[934]), .RECT3_WEIGHT(rectangle3_weights[934]), .FEAT_THRES(feature_thresholds[934]), .FEAT_ABOVE(feature_aboves[934]), .FEAT_BELOW(feature_belows[934])) ac934(.scan_win(scan_win934), .scan_win_std_dev(scan_win_std_dev[934]), .feature_accum(feature_accums[934]));
  accum_calculator #(.RECT1_X(rectangle1_xs[935]), .RECT1_Y(rectangle1_ys[935]), .RECT1_WIDTH(rectangle1_widths[935]), .RECT1_HEIGHT(rectangle1_heights[935]), .RECT1_WEIGHT(rectangle1_weights[935]), .RECT2_X(rectangle2_xs[935]), .RECT2_Y(rectangle2_ys[935]), .RECT2_WIDTH(rectangle2_widths[935]), .RECT2_HEIGHT(rectangle2_heights[935]), .RECT2_WEIGHT(rectangle2_weights[935]), .RECT3_X(rectangle3_xs[935]), .RECT3_Y(rectangle3_ys[935]), .RECT3_WIDTH(rectangle3_widths[935]), .RECT3_HEIGHT(rectangle3_heights[935]), .RECT3_WEIGHT(rectangle3_weights[935]), .FEAT_THRES(feature_thresholds[935]), .FEAT_ABOVE(feature_aboves[935]), .FEAT_BELOW(feature_belows[935])) ac935(.scan_win(scan_win935), .scan_win_std_dev(scan_win_std_dev[935]), .feature_accum(feature_accums[935]));
  accum_calculator #(.RECT1_X(rectangle1_xs[936]), .RECT1_Y(rectangle1_ys[936]), .RECT1_WIDTH(rectangle1_widths[936]), .RECT1_HEIGHT(rectangle1_heights[936]), .RECT1_WEIGHT(rectangle1_weights[936]), .RECT2_X(rectangle2_xs[936]), .RECT2_Y(rectangle2_ys[936]), .RECT2_WIDTH(rectangle2_widths[936]), .RECT2_HEIGHT(rectangle2_heights[936]), .RECT2_WEIGHT(rectangle2_weights[936]), .RECT3_X(rectangle3_xs[936]), .RECT3_Y(rectangle3_ys[936]), .RECT3_WIDTH(rectangle3_widths[936]), .RECT3_HEIGHT(rectangle3_heights[936]), .RECT3_WEIGHT(rectangle3_weights[936]), .FEAT_THRES(feature_thresholds[936]), .FEAT_ABOVE(feature_aboves[936]), .FEAT_BELOW(feature_belows[936])) ac936(.scan_win(scan_win936), .scan_win_std_dev(scan_win_std_dev[936]), .feature_accum(feature_accums[936]));
  accum_calculator #(.RECT1_X(rectangle1_xs[937]), .RECT1_Y(rectangle1_ys[937]), .RECT1_WIDTH(rectangle1_widths[937]), .RECT1_HEIGHT(rectangle1_heights[937]), .RECT1_WEIGHT(rectangle1_weights[937]), .RECT2_X(rectangle2_xs[937]), .RECT2_Y(rectangle2_ys[937]), .RECT2_WIDTH(rectangle2_widths[937]), .RECT2_HEIGHT(rectangle2_heights[937]), .RECT2_WEIGHT(rectangle2_weights[937]), .RECT3_X(rectangle3_xs[937]), .RECT3_Y(rectangle3_ys[937]), .RECT3_WIDTH(rectangle3_widths[937]), .RECT3_HEIGHT(rectangle3_heights[937]), .RECT3_WEIGHT(rectangle3_weights[937]), .FEAT_THRES(feature_thresholds[937]), .FEAT_ABOVE(feature_aboves[937]), .FEAT_BELOW(feature_belows[937])) ac937(.scan_win(scan_win937), .scan_win_std_dev(scan_win_std_dev[937]), .feature_accum(feature_accums[937]));
  accum_calculator #(.RECT1_X(rectangle1_xs[938]), .RECT1_Y(rectangle1_ys[938]), .RECT1_WIDTH(rectangle1_widths[938]), .RECT1_HEIGHT(rectangle1_heights[938]), .RECT1_WEIGHT(rectangle1_weights[938]), .RECT2_X(rectangle2_xs[938]), .RECT2_Y(rectangle2_ys[938]), .RECT2_WIDTH(rectangle2_widths[938]), .RECT2_HEIGHT(rectangle2_heights[938]), .RECT2_WEIGHT(rectangle2_weights[938]), .RECT3_X(rectangle3_xs[938]), .RECT3_Y(rectangle3_ys[938]), .RECT3_WIDTH(rectangle3_widths[938]), .RECT3_HEIGHT(rectangle3_heights[938]), .RECT3_WEIGHT(rectangle3_weights[938]), .FEAT_THRES(feature_thresholds[938]), .FEAT_ABOVE(feature_aboves[938]), .FEAT_BELOW(feature_belows[938])) ac938(.scan_win(scan_win938), .scan_win_std_dev(scan_win_std_dev[938]), .feature_accum(feature_accums[938]));
  accum_calculator #(.RECT1_X(rectangle1_xs[939]), .RECT1_Y(rectangle1_ys[939]), .RECT1_WIDTH(rectangle1_widths[939]), .RECT1_HEIGHT(rectangle1_heights[939]), .RECT1_WEIGHT(rectangle1_weights[939]), .RECT2_X(rectangle2_xs[939]), .RECT2_Y(rectangle2_ys[939]), .RECT2_WIDTH(rectangle2_widths[939]), .RECT2_HEIGHT(rectangle2_heights[939]), .RECT2_WEIGHT(rectangle2_weights[939]), .RECT3_X(rectangle3_xs[939]), .RECT3_Y(rectangle3_ys[939]), .RECT3_WIDTH(rectangle3_widths[939]), .RECT3_HEIGHT(rectangle3_heights[939]), .RECT3_WEIGHT(rectangle3_weights[939]), .FEAT_THRES(feature_thresholds[939]), .FEAT_ABOVE(feature_aboves[939]), .FEAT_BELOW(feature_belows[939])) ac939(.scan_win(scan_win939), .scan_win_std_dev(scan_win_std_dev[939]), .feature_accum(feature_accums[939]));
  accum_calculator #(.RECT1_X(rectangle1_xs[940]), .RECT1_Y(rectangle1_ys[940]), .RECT1_WIDTH(rectangle1_widths[940]), .RECT1_HEIGHT(rectangle1_heights[940]), .RECT1_WEIGHT(rectangle1_weights[940]), .RECT2_X(rectangle2_xs[940]), .RECT2_Y(rectangle2_ys[940]), .RECT2_WIDTH(rectangle2_widths[940]), .RECT2_HEIGHT(rectangle2_heights[940]), .RECT2_WEIGHT(rectangle2_weights[940]), .RECT3_X(rectangle3_xs[940]), .RECT3_Y(rectangle3_ys[940]), .RECT3_WIDTH(rectangle3_widths[940]), .RECT3_HEIGHT(rectangle3_heights[940]), .RECT3_WEIGHT(rectangle3_weights[940]), .FEAT_THRES(feature_thresholds[940]), .FEAT_ABOVE(feature_aboves[940]), .FEAT_BELOW(feature_belows[940])) ac940(.scan_win(scan_win940), .scan_win_std_dev(scan_win_std_dev[940]), .feature_accum(feature_accums[940]));
  accum_calculator #(.RECT1_X(rectangle1_xs[941]), .RECT1_Y(rectangle1_ys[941]), .RECT1_WIDTH(rectangle1_widths[941]), .RECT1_HEIGHT(rectangle1_heights[941]), .RECT1_WEIGHT(rectangle1_weights[941]), .RECT2_X(rectangle2_xs[941]), .RECT2_Y(rectangle2_ys[941]), .RECT2_WIDTH(rectangle2_widths[941]), .RECT2_HEIGHT(rectangle2_heights[941]), .RECT2_WEIGHT(rectangle2_weights[941]), .RECT3_X(rectangle3_xs[941]), .RECT3_Y(rectangle3_ys[941]), .RECT3_WIDTH(rectangle3_widths[941]), .RECT3_HEIGHT(rectangle3_heights[941]), .RECT3_WEIGHT(rectangle3_weights[941]), .FEAT_THRES(feature_thresholds[941]), .FEAT_ABOVE(feature_aboves[941]), .FEAT_BELOW(feature_belows[941])) ac941(.scan_win(scan_win941), .scan_win_std_dev(scan_win_std_dev[941]), .feature_accum(feature_accums[941]));
  accum_calculator #(.RECT1_X(rectangle1_xs[942]), .RECT1_Y(rectangle1_ys[942]), .RECT1_WIDTH(rectangle1_widths[942]), .RECT1_HEIGHT(rectangle1_heights[942]), .RECT1_WEIGHT(rectangle1_weights[942]), .RECT2_X(rectangle2_xs[942]), .RECT2_Y(rectangle2_ys[942]), .RECT2_WIDTH(rectangle2_widths[942]), .RECT2_HEIGHT(rectangle2_heights[942]), .RECT2_WEIGHT(rectangle2_weights[942]), .RECT3_X(rectangle3_xs[942]), .RECT3_Y(rectangle3_ys[942]), .RECT3_WIDTH(rectangle3_widths[942]), .RECT3_HEIGHT(rectangle3_heights[942]), .RECT3_WEIGHT(rectangle3_weights[942]), .FEAT_THRES(feature_thresholds[942]), .FEAT_ABOVE(feature_aboves[942]), .FEAT_BELOW(feature_belows[942])) ac942(.scan_win(scan_win942), .scan_win_std_dev(scan_win_std_dev[942]), .feature_accum(feature_accums[942]));
  accum_calculator #(.RECT1_X(rectangle1_xs[943]), .RECT1_Y(rectangle1_ys[943]), .RECT1_WIDTH(rectangle1_widths[943]), .RECT1_HEIGHT(rectangle1_heights[943]), .RECT1_WEIGHT(rectangle1_weights[943]), .RECT2_X(rectangle2_xs[943]), .RECT2_Y(rectangle2_ys[943]), .RECT2_WIDTH(rectangle2_widths[943]), .RECT2_HEIGHT(rectangle2_heights[943]), .RECT2_WEIGHT(rectangle2_weights[943]), .RECT3_X(rectangle3_xs[943]), .RECT3_Y(rectangle3_ys[943]), .RECT3_WIDTH(rectangle3_widths[943]), .RECT3_HEIGHT(rectangle3_heights[943]), .RECT3_WEIGHT(rectangle3_weights[943]), .FEAT_THRES(feature_thresholds[943]), .FEAT_ABOVE(feature_aboves[943]), .FEAT_BELOW(feature_belows[943])) ac943(.scan_win(scan_win943), .scan_win_std_dev(scan_win_std_dev[943]), .feature_accum(feature_accums[943]));
  accum_calculator #(.RECT1_X(rectangle1_xs[944]), .RECT1_Y(rectangle1_ys[944]), .RECT1_WIDTH(rectangle1_widths[944]), .RECT1_HEIGHT(rectangle1_heights[944]), .RECT1_WEIGHT(rectangle1_weights[944]), .RECT2_X(rectangle2_xs[944]), .RECT2_Y(rectangle2_ys[944]), .RECT2_WIDTH(rectangle2_widths[944]), .RECT2_HEIGHT(rectangle2_heights[944]), .RECT2_WEIGHT(rectangle2_weights[944]), .RECT3_X(rectangle3_xs[944]), .RECT3_Y(rectangle3_ys[944]), .RECT3_WIDTH(rectangle3_widths[944]), .RECT3_HEIGHT(rectangle3_heights[944]), .RECT3_WEIGHT(rectangle3_weights[944]), .FEAT_THRES(feature_thresholds[944]), .FEAT_ABOVE(feature_aboves[944]), .FEAT_BELOW(feature_belows[944])) ac944(.scan_win(scan_win944), .scan_win_std_dev(scan_win_std_dev[944]), .feature_accum(feature_accums[944]));
  accum_calculator #(.RECT1_X(rectangle1_xs[945]), .RECT1_Y(rectangle1_ys[945]), .RECT1_WIDTH(rectangle1_widths[945]), .RECT1_HEIGHT(rectangle1_heights[945]), .RECT1_WEIGHT(rectangle1_weights[945]), .RECT2_X(rectangle2_xs[945]), .RECT2_Y(rectangle2_ys[945]), .RECT2_WIDTH(rectangle2_widths[945]), .RECT2_HEIGHT(rectangle2_heights[945]), .RECT2_WEIGHT(rectangle2_weights[945]), .RECT3_X(rectangle3_xs[945]), .RECT3_Y(rectangle3_ys[945]), .RECT3_WIDTH(rectangle3_widths[945]), .RECT3_HEIGHT(rectangle3_heights[945]), .RECT3_WEIGHT(rectangle3_weights[945]), .FEAT_THRES(feature_thresholds[945]), .FEAT_ABOVE(feature_aboves[945]), .FEAT_BELOW(feature_belows[945])) ac945(.scan_win(scan_win945), .scan_win_std_dev(scan_win_std_dev[945]), .feature_accum(feature_accums[945]));
  accum_calculator #(.RECT1_X(rectangle1_xs[946]), .RECT1_Y(rectangle1_ys[946]), .RECT1_WIDTH(rectangle1_widths[946]), .RECT1_HEIGHT(rectangle1_heights[946]), .RECT1_WEIGHT(rectangle1_weights[946]), .RECT2_X(rectangle2_xs[946]), .RECT2_Y(rectangle2_ys[946]), .RECT2_WIDTH(rectangle2_widths[946]), .RECT2_HEIGHT(rectangle2_heights[946]), .RECT2_WEIGHT(rectangle2_weights[946]), .RECT3_X(rectangle3_xs[946]), .RECT3_Y(rectangle3_ys[946]), .RECT3_WIDTH(rectangle3_widths[946]), .RECT3_HEIGHT(rectangle3_heights[946]), .RECT3_WEIGHT(rectangle3_weights[946]), .FEAT_THRES(feature_thresholds[946]), .FEAT_ABOVE(feature_aboves[946]), .FEAT_BELOW(feature_belows[946])) ac946(.scan_win(scan_win946), .scan_win_std_dev(scan_win_std_dev[946]), .feature_accum(feature_accums[946]));
  accum_calculator #(.RECT1_X(rectangle1_xs[947]), .RECT1_Y(rectangle1_ys[947]), .RECT1_WIDTH(rectangle1_widths[947]), .RECT1_HEIGHT(rectangle1_heights[947]), .RECT1_WEIGHT(rectangle1_weights[947]), .RECT2_X(rectangle2_xs[947]), .RECT2_Y(rectangle2_ys[947]), .RECT2_WIDTH(rectangle2_widths[947]), .RECT2_HEIGHT(rectangle2_heights[947]), .RECT2_WEIGHT(rectangle2_weights[947]), .RECT3_X(rectangle3_xs[947]), .RECT3_Y(rectangle3_ys[947]), .RECT3_WIDTH(rectangle3_widths[947]), .RECT3_HEIGHT(rectangle3_heights[947]), .RECT3_WEIGHT(rectangle3_weights[947]), .FEAT_THRES(feature_thresholds[947]), .FEAT_ABOVE(feature_aboves[947]), .FEAT_BELOW(feature_belows[947])) ac947(.scan_win(scan_win947), .scan_win_std_dev(scan_win_std_dev[947]), .feature_accum(feature_accums[947]));
  accum_calculator #(.RECT1_X(rectangle1_xs[948]), .RECT1_Y(rectangle1_ys[948]), .RECT1_WIDTH(rectangle1_widths[948]), .RECT1_HEIGHT(rectangle1_heights[948]), .RECT1_WEIGHT(rectangle1_weights[948]), .RECT2_X(rectangle2_xs[948]), .RECT2_Y(rectangle2_ys[948]), .RECT2_WIDTH(rectangle2_widths[948]), .RECT2_HEIGHT(rectangle2_heights[948]), .RECT2_WEIGHT(rectangle2_weights[948]), .RECT3_X(rectangle3_xs[948]), .RECT3_Y(rectangle3_ys[948]), .RECT3_WIDTH(rectangle3_widths[948]), .RECT3_HEIGHT(rectangle3_heights[948]), .RECT3_WEIGHT(rectangle3_weights[948]), .FEAT_THRES(feature_thresholds[948]), .FEAT_ABOVE(feature_aboves[948]), .FEAT_BELOW(feature_belows[948])) ac948(.scan_win(scan_win948), .scan_win_std_dev(scan_win_std_dev[948]), .feature_accum(feature_accums[948]));
  accum_calculator #(.RECT1_X(rectangle1_xs[949]), .RECT1_Y(rectangle1_ys[949]), .RECT1_WIDTH(rectangle1_widths[949]), .RECT1_HEIGHT(rectangle1_heights[949]), .RECT1_WEIGHT(rectangle1_weights[949]), .RECT2_X(rectangle2_xs[949]), .RECT2_Y(rectangle2_ys[949]), .RECT2_WIDTH(rectangle2_widths[949]), .RECT2_HEIGHT(rectangle2_heights[949]), .RECT2_WEIGHT(rectangle2_weights[949]), .RECT3_X(rectangle3_xs[949]), .RECT3_Y(rectangle3_ys[949]), .RECT3_WIDTH(rectangle3_widths[949]), .RECT3_HEIGHT(rectangle3_heights[949]), .RECT3_WEIGHT(rectangle3_weights[949]), .FEAT_THRES(feature_thresholds[949]), .FEAT_ABOVE(feature_aboves[949]), .FEAT_BELOW(feature_belows[949])) ac949(.scan_win(scan_win949), .scan_win_std_dev(scan_win_std_dev[949]), .feature_accum(feature_accums[949]));
  accum_calculator #(.RECT1_X(rectangle1_xs[950]), .RECT1_Y(rectangle1_ys[950]), .RECT1_WIDTH(rectangle1_widths[950]), .RECT1_HEIGHT(rectangle1_heights[950]), .RECT1_WEIGHT(rectangle1_weights[950]), .RECT2_X(rectangle2_xs[950]), .RECT2_Y(rectangle2_ys[950]), .RECT2_WIDTH(rectangle2_widths[950]), .RECT2_HEIGHT(rectangle2_heights[950]), .RECT2_WEIGHT(rectangle2_weights[950]), .RECT3_X(rectangle3_xs[950]), .RECT3_Y(rectangle3_ys[950]), .RECT3_WIDTH(rectangle3_widths[950]), .RECT3_HEIGHT(rectangle3_heights[950]), .RECT3_WEIGHT(rectangle3_weights[950]), .FEAT_THRES(feature_thresholds[950]), .FEAT_ABOVE(feature_aboves[950]), .FEAT_BELOW(feature_belows[950])) ac950(.scan_win(scan_win950), .scan_win_std_dev(scan_win_std_dev[950]), .feature_accum(feature_accums[950]));
  accum_calculator #(.RECT1_X(rectangle1_xs[951]), .RECT1_Y(rectangle1_ys[951]), .RECT1_WIDTH(rectangle1_widths[951]), .RECT1_HEIGHT(rectangle1_heights[951]), .RECT1_WEIGHT(rectangle1_weights[951]), .RECT2_X(rectangle2_xs[951]), .RECT2_Y(rectangle2_ys[951]), .RECT2_WIDTH(rectangle2_widths[951]), .RECT2_HEIGHT(rectangle2_heights[951]), .RECT2_WEIGHT(rectangle2_weights[951]), .RECT3_X(rectangle3_xs[951]), .RECT3_Y(rectangle3_ys[951]), .RECT3_WIDTH(rectangle3_widths[951]), .RECT3_HEIGHT(rectangle3_heights[951]), .RECT3_WEIGHT(rectangle3_weights[951]), .FEAT_THRES(feature_thresholds[951]), .FEAT_ABOVE(feature_aboves[951]), .FEAT_BELOW(feature_belows[951])) ac951(.scan_win(scan_win951), .scan_win_std_dev(scan_win_std_dev[951]), .feature_accum(feature_accums[951]));
  accum_calculator #(.RECT1_X(rectangle1_xs[952]), .RECT1_Y(rectangle1_ys[952]), .RECT1_WIDTH(rectangle1_widths[952]), .RECT1_HEIGHT(rectangle1_heights[952]), .RECT1_WEIGHT(rectangle1_weights[952]), .RECT2_X(rectangle2_xs[952]), .RECT2_Y(rectangle2_ys[952]), .RECT2_WIDTH(rectangle2_widths[952]), .RECT2_HEIGHT(rectangle2_heights[952]), .RECT2_WEIGHT(rectangle2_weights[952]), .RECT3_X(rectangle3_xs[952]), .RECT3_Y(rectangle3_ys[952]), .RECT3_WIDTH(rectangle3_widths[952]), .RECT3_HEIGHT(rectangle3_heights[952]), .RECT3_WEIGHT(rectangle3_weights[952]), .FEAT_THRES(feature_thresholds[952]), .FEAT_ABOVE(feature_aboves[952]), .FEAT_BELOW(feature_belows[952])) ac952(.scan_win(scan_win952), .scan_win_std_dev(scan_win_std_dev[952]), .feature_accum(feature_accums[952]));
  accum_calculator #(.RECT1_X(rectangle1_xs[953]), .RECT1_Y(rectangle1_ys[953]), .RECT1_WIDTH(rectangle1_widths[953]), .RECT1_HEIGHT(rectangle1_heights[953]), .RECT1_WEIGHT(rectangle1_weights[953]), .RECT2_X(rectangle2_xs[953]), .RECT2_Y(rectangle2_ys[953]), .RECT2_WIDTH(rectangle2_widths[953]), .RECT2_HEIGHT(rectangle2_heights[953]), .RECT2_WEIGHT(rectangle2_weights[953]), .RECT3_X(rectangle3_xs[953]), .RECT3_Y(rectangle3_ys[953]), .RECT3_WIDTH(rectangle3_widths[953]), .RECT3_HEIGHT(rectangle3_heights[953]), .RECT3_WEIGHT(rectangle3_weights[953]), .FEAT_THRES(feature_thresholds[953]), .FEAT_ABOVE(feature_aboves[953]), .FEAT_BELOW(feature_belows[953])) ac953(.scan_win(scan_win953), .scan_win_std_dev(scan_win_std_dev[953]), .feature_accum(feature_accums[953]));
  accum_calculator #(.RECT1_X(rectangle1_xs[954]), .RECT1_Y(rectangle1_ys[954]), .RECT1_WIDTH(rectangle1_widths[954]), .RECT1_HEIGHT(rectangle1_heights[954]), .RECT1_WEIGHT(rectangle1_weights[954]), .RECT2_X(rectangle2_xs[954]), .RECT2_Y(rectangle2_ys[954]), .RECT2_WIDTH(rectangle2_widths[954]), .RECT2_HEIGHT(rectangle2_heights[954]), .RECT2_WEIGHT(rectangle2_weights[954]), .RECT3_X(rectangle3_xs[954]), .RECT3_Y(rectangle3_ys[954]), .RECT3_WIDTH(rectangle3_widths[954]), .RECT3_HEIGHT(rectangle3_heights[954]), .RECT3_WEIGHT(rectangle3_weights[954]), .FEAT_THRES(feature_thresholds[954]), .FEAT_ABOVE(feature_aboves[954]), .FEAT_BELOW(feature_belows[954])) ac954(.scan_win(scan_win954), .scan_win_std_dev(scan_win_std_dev[954]), .feature_accum(feature_accums[954]));
  accum_calculator #(.RECT1_X(rectangle1_xs[955]), .RECT1_Y(rectangle1_ys[955]), .RECT1_WIDTH(rectangle1_widths[955]), .RECT1_HEIGHT(rectangle1_heights[955]), .RECT1_WEIGHT(rectangle1_weights[955]), .RECT2_X(rectangle2_xs[955]), .RECT2_Y(rectangle2_ys[955]), .RECT2_WIDTH(rectangle2_widths[955]), .RECT2_HEIGHT(rectangle2_heights[955]), .RECT2_WEIGHT(rectangle2_weights[955]), .RECT3_X(rectangle3_xs[955]), .RECT3_Y(rectangle3_ys[955]), .RECT3_WIDTH(rectangle3_widths[955]), .RECT3_HEIGHT(rectangle3_heights[955]), .RECT3_WEIGHT(rectangle3_weights[955]), .FEAT_THRES(feature_thresholds[955]), .FEAT_ABOVE(feature_aboves[955]), .FEAT_BELOW(feature_belows[955])) ac955(.scan_win(scan_win955), .scan_win_std_dev(scan_win_std_dev[955]), .feature_accum(feature_accums[955]));
  accum_calculator #(.RECT1_X(rectangle1_xs[956]), .RECT1_Y(rectangle1_ys[956]), .RECT1_WIDTH(rectangle1_widths[956]), .RECT1_HEIGHT(rectangle1_heights[956]), .RECT1_WEIGHT(rectangle1_weights[956]), .RECT2_X(rectangle2_xs[956]), .RECT2_Y(rectangle2_ys[956]), .RECT2_WIDTH(rectangle2_widths[956]), .RECT2_HEIGHT(rectangle2_heights[956]), .RECT2_WEIGHT(rectangle2_weights[956]), .RECT3_X(rectangle3_xs[956]), .RECT3_Y(rectangle3_ys[956]), .RECT3_WIDTH(rectangle3_widths[956]), .RECT3_HEIGHT(rectangle3_heights[956]), .RECT3_WEIGHT(rectangle3_weights[956]), .FEAT_THRES(feature_thresholds[956]), .FEAT_ABOVE(feature_aboves[956]), .FEAT_BELOW(feature_belows[956])) ac956(.scan_win(scan_win956), .scan_win_std_dev(scan_win_std_dev[956]), .feature_accum(feature_accums[956]));
  accum_calculator #(.RECT1_X(rectangle1_xs[957]), .RECT1_Y(rectangle1_ys[957]), .RECT1_WIDTH(rectangle1_widths[957]), .RECT1_HEIGHT(rectangle1_heights[957]), .RECT1_WEIGHT(rectangle1_weights[957]), .RECT2_X(rectangle2_xs[957]), .RECT2_Y(rectangle2_ys[957]), .RECT2_WIDTH(rectangle2_widths[957]), .RECT2_HEIGHT(rectangle2_heights[957]), .RECT2_WEIGHT(rectangle2_weights[957]), .RECT3_X(rectangle3_xs[957]), .RECT3_Y(rectangle3_ys[957]), .RECT3_WIDTH(rectangle3_widths[957]), .RECT3_HEIGHT(rectangle3_heights[957]), .RECT3_WEIGHT(rectangle3_weights[957]), .FEAT_THRES(feature_thresholds[957]), .FEAT_ABOVE(feature_aboves[957]), .FEAT_BELOW(feature_belows[957])) ac957(.scan_win(scan_win957), .scan_win_std_dev(scan_win_std_dev[957]), .feature_accum(feature_accums[957]));
  accum_calculator #(.RECT1_X(rectangle1_xs[958]), .RECT1_Y(rectangle1_ys[958]), .RECT1_WIDTH(rectangle1_widths[958]), .RECT1_HEIGHT(rectangle1_heights[958]), .RECT1_WEIGHT(rectangle1_weights[958]), .RECT2_X(rectangle2_xs[958]), .RECT2_Y(rectangle2_ys[958]), .RECT2_WIDTH(rectangle2_widths[958]), .RECT2_HEIGHT(rectangle2_heights[958]), .RECT2_WEIGHT(rectangle2_weights[958]), .RECT3_X(rectangle3_xs[958]), .RECT3_Y(rectangle3_ys[958]), .RECT3_WIDTH(rectangle3_widths[958]), .RECT3_HEIGHT(rectangle3_heights[958]), .RECT3_WEIGHT(rectangle3_weights[958]), .FEAT_THRES(feature_thresholds[958]), .FEAT_ABOVE(feature_aboves[958]), .FEAT_BELOW(feature_belows[958])) ac958(.scan_win(scan_win958), .scan_win_std_dev(scan_win_std_dev[958]), .feature_accum(feature_accums[958]));
  accum_calculator #(.RECT1_X(rectangle1_xs[959]), .RECT1_Y(rectangle1_ys[959]), .RECT1_WIDTH(rectangle1_widths[959]), .RECT1_HEIGHT(rectangle1_heights[959]), .RECT1_WEIGHT(rectangle1_weights[959]), .RECT2_X(rectangle2_xs[959]), .RECT2_Y(rectangle2_ys[959]), .RECT2_WIDTH(rectangle2_widths[959]), .RECT2_HEIGHT(rectangle2_heights[959]), .RECT2_WEIGHT(rectangle2_weights[959]), .RECT3_X(rectangle3_xs[959]), .RECT3_Y(rectangle3_ys[959]), .RECT3_WIDTH(rectangle3_widths[959]), .RECT3_HEIGHT(rectangle3_heights[959]), .RECT3_WEIGHT(rectangle3_weights[959]), .FEAT_THRES(feature_thresholds[959]), .FEAT_ABOVE(feature_aboves[959]), .FEAT_BELOW(feature_belows[959])) ac959(.scan_win(scan_win959), .scan_win_std_dev(scan_win_std_dev[959]), .feature_accum(feature_accums[959]));
  accum_calculator #(.RECT1_X(rectangle1_xs[960]), .RECT1_Y(rectangle1_ys[960]), .RECT1_WIDTH(rectangle1_widths[960]), .RECT1_HEIGHT(rectangle1_heights[960]), .RECT1_WEIGHT(rectangle1_weights[960]), .RECT2_X(rectangle2_xs[960]), .RECT2_Y(rectangle2_ys[960]), .RECT2_WIDTH(rectangle2_widths[960]), .RECT2_HEIGHT(rectangle2_heights[960]), .RECT2_WEIGHT(rectangle2_weights[960]), .RECT3_X(rectangle3_xs[960]), .RECT3_Y(rectangle3_ys[960]), .RECT3_WIDTH(rectangle3_widths[960]), .RECT3_HEIGHT(rectangle3_heights[960]), .RECT3_WEIGHT(rectangle3_weights[960]), .FEAT_THRES(feature_thresholds[960]), .FEAT_ABOVE(feature_aboves[960]), .FEAT_BELOW(feature_belows[960])) ac960(.scan_win(scan_win960), .scan_win_std_dev(scan_win_std_dev[960]), .feature_accum(feature_accums[960]));
  accum_calculator #(.RECT1_X(rectangle1_xs[961]), .RECT1_Y(rectangle1_ys[961]), .RECT1_WIDTH(rectangle1_widths[961]), .RECT1_HEIGHT(rectangle1_heights[961]), .RECT1_WEIGHT(rectangle1_weights[961]), .RECT2_X(rectangle2_xs[961]), .RECT2_Y(rectangle2_ys[961]), .RECT2_WIDTH(rectangle2_widths[961]), .RECT2_HEIGHT(rectangle2_heights[961]), .RECT2_WEIGHT(rectangle2_weights[961]), .RECT3_X(rectangle3_xs[961]), .RECT3_Y(rectangle3_ys[961]), .RECT3_WIDTH(rectangle3_widths[961]), .RECT3_HEIGHT(rectangle3_heights[961]), .RECT3_WEIGHT(rectangle3_weights[961]), .FEAT_THRES(feature_thresholds[961]), .FEAT_ABOVE(feature_aboves[961]), .FEAT_BELOW(feature_belows[961])) ac961(.scan_win(scan_win961), .scan_win_std_dev(scan_win_std_dev[961]), .feature_accum(feature_accums[961]));
  accum_calculator #(.RECT1_X(rectangle1_xs[962]), .RECT1_Y(rectangle1_ys[962]), .RECT1_WIDTH(rectangle1_widths[962]), .RECT1_HEIGHT(rectangle1_heights[962]), .RECT1_WEIGHT(rectangle1_weights[962]), .RECT2_X(rectangle2_xs[962]), .RECT2_Y(rectangle2_ys[962]), .RECT2_WIDTH(rectangle2_widths[962]), .RECT2_HEIGHT(rectangle2_heights[962]), .RECT2_WEIGHT(rectangle2_weights[962]), .RECT3_X(rectangle3_xs[962]), .RECT3_Y(rectangle3_ys[962]), .RECT3_WIDTH(rectangle3_widths[962]), .RECT3_HEIGHT(rectangle3_heights[962]), .RECT3_WEIGHT(rectangle3_weights[962]), .FEAT_THRES(feature_thresholds[962]), .FEAT_ABOVE(feature_aboves[962]), .FEAT_BELOW(feature_belows[962])) ac962(.scan_win(scan_win962), .scan_win_std_dev(scan_win_std_dev[962]), .feature_accum(feature_accums[962]));
  accum_calculator #(.RECT1_X(rectangle1_xs[963]), .RECT1_Y(rectangle1_ys[963]), .RECT1_WIDTH(rectangle1_widths[963]), .RECT1_HEIGHT(rectangle1_heights[963]), .RECT1_WEIGHT(rectangle1_weights[963]), .RECT2_X(rectangle2_xs[963]), .RECT2_Y(rectangle2_ys[963]), .RECT2_WIDTH(rectangle2_widths[963]), .RECT2_HEIGHT(rectangle2_heights[963]), .RECT2_WEIGHT(rectangle2_weights[963]), .RECT3_X(rectangle3_xs[963]), .RECT3_Y(rectangle3_ys[963]), .RECT3_WIDTH(rectangle3_widths[963]), .RECT3_HEIGHT(rectangle3_heights[963]), .RECT3_WEIGHT(rectangle3_weights[963]), .FEAT_THRES(feature_thresholds[963]), .FEAT_ABOVE(feature_aboves[963]), .FEAT_BELOW(feature_belows[963])) ac963(.scan_win(scan_win963), .scan_win_std_dev(scan_win_std_dev[963]), .feature_accum(feature_accums[963]));
  accum_calculator #(.RECT1_X(rectangle1_xs[964]), .RECT1_Y(rectangle1_ys[964]), .RECT1_WIDTH(rectangle1_widths[964]), .RECT1_HEIGHT(rectangle1_heights[964]), .RECT1_WEIGHT(rectangle1_weights[964]), .RECT2_X(rectangle2_xs[964]), .RECT2_Y(rectangle2_ys[964]), .RECT2_WIDTH(rectangle2_widths[964]), .RECT2_HEIGHT(rectangle2_heights[964]), .RECT2_WEIGHT(rectangle2_weights[964]), .RECT3_X(rectangle3_xs[964]), .RECT3_Y(rectangle3_ys[964]), .RECT3_WIDTH(rectangle3_widths[964]), .RECT3_HEIGHT(rectangle3_heights[964]), .RECT3_WEIGHT(rectangle3_weights[964]), .FEAT_THRES(feature_thresholds[964]), .FEAT_ABOVE(feature_aboves[964]), .FEAT_BELOW(feature_belows[964])) ac964(.scan_win(scan_win964), .scan_win_std_dev(scan_win_std_dev[964]), .feature_accum(feature_accums[964]));
  accum_calculator #(.RECT1_X(rectangle1_xs[965]), .RECT1_Y(rectangle1_ys[965]), .RECT1_WIDTH(rectangle1_widths[965]), .RECT1_HEIGHT(rectangle1_heights[965]), .RECT1_WEIGHT(rectangle1_weights[965]), .RECT2_X(rectangle2_xs[965]), .RECT2_Y(rectangle2_ys[965]), .RECT2_WIDTH(rectangle2_widths[965]), .RECT2_HEIGHT(rectangle2_heights[965]), .RECT2_WEIGHT(rectangle2_weights[965]), .RECT3_X(rectangle3_xs[965]), .RECT3_Y(rectangle3_ys[965]), .RECT3_WIDTH(rectangle3_widths[965]), .RECT3_HEIGHT(rectangle3_heights[965]), .RECT3_WEIGHT(rectangle3_weights[965]), .FEAT_THRES(feature_thresholds[965]), .FEAT_ABOVE(feature_aboves[965]), .FEAT_BELOW(feature_belows[965])) ac965(.scan_win(scan_win965), .scan_win_std_dev(scan_win_std_dev[965]), .feature_accum(feature_accums[965]));
  accum_calculator #(.RECT1_X(rectangle1_xs[966]), .RECT1_Y(rectangle1_ys[966]), .RECT1_WIDTH(rectangle1_widths[966]), .RECT1_HEIGHT(rectangle1_heights[966]), .RECT1_WEIGHT(rectangle1_weights[966]), .RECT2_X(rectangle2_xs[966]), .RECT2_Y(rectangle2_ys[966]), .RECT2_WIDTH(rectangle2_widths[966]), .RECT2_HEIGHT(rectangle2_heights[966]), .RECT2_WEIGHT(rectangle2_weights[966]), .RECT3_X(rectangle3_xs[966]), .RECT3_Y(rectangle3_ys[966]), .RECT3_WIDTH(rectangle3_widths[966]), .RECT3_HEIGHT(rectangle3_heights[966]), .RECT3_WEIGHT(rectangle3_weights[966]), .FEAT_THRES(feature_thresholds[966]), .FEAT_ABOVE(feature_aboves[966]), .FEAT_BELOW(feature_belows[966])) ac966(.scan_win(scan_win966), .scan_win_std_dev(scan_win_std_dev[966]), .feature_accum(feature_accums[966]));
  accum_calculator #(.RECT1_X(rectangle1_xs[967]), .RECT1_Y(rectangle1_ys[967]), .RECT1_WIDTH(rectangle1_widths[967]), .RECT1_HEIGHT(rectangle1_heights[967]), .RECT1_WEIGHT(rectangle1_weights[967]), .RECT2_X(rectangle2_xs[967]), .RECT2_Y(rectangle2_ys[967]), .RECT2_WIDTH(rectangle2_widths[967]), .RECT2_HEIGHT(rectangle2_heights[967]), .RECT2_WEIGHT(rectangle2_weights[967]), .RECT3_X(rectangle3_xs[967]), .RECT3_Y(rectangle3_ys[967]), .RECT3_WIDTH(rectangle3_widths[967]), .RECT3_HEIGHT(rectangle3_heights[967]), .RECT3_WEIGHT(rectangle3_weights[967]), .FEAT_THRES(feature_thresholds[967]), .FEAT_ABOVE(feature_aboves[967]), .FEAT_BELOW(feature_belows[967])) ac967(.scan_win(scan_win967), .scan_win_std_dev(scan_win_std_dev[967]), .feature_accum(feature_accums[967]));
  accum_calculator #(.RECT1_X(rectangle1_xs[968]), .RECT1_Y(rectangle1_ys[968]), .RECT1_WIDTH(rectangle1_widths[968]), .RECT1_HEIGHT(rectangle1_heights[968]), .RECT1_WEIGHT(rectangle1_weights[968]), .RECT2_X(rectangle2_xs[968]), .RECT2_Y(rectangle2_ys[968]), .RECT2_WIDTH(rectangle2_widths[968]), .RECT2_HEIGHT(rectangle2_heights[968]), .RECT2_WEIGHT(rectangle2_weights[968]), .RECT3_X(rectangle3_xs[968]), .RECT3_Y(rectangle3_ys[968]), .RECT3_WIDTH(rectangle3_widths[968]), .RECT3_HEIGHT(rectangle3_heights[968]), .RECT3_WEIGHT(rectangle3_weights[968]), .FEAT_THRES(feature_thresholds[968]), .FEAT_ABOVE(feature_aboves[968]), .FEAT_BELOW(feature_belows[968])) ac968(.scan_win(scan_win968), .scan_win_std_dev(scan_win_std_dev[968]), .feature_accum(feature_accums[968]));
  accum_calculator #(.RECT1_X(rectangle1_xs[969]), .RECT1_Y(rectangle1_ys[969]), .RECT1_WIDTH(rectangle1_widths[969]), .RECT1_HEIGHT(rectangle1_heights[969]), .RECT1_WEIGHT(rectangle1_weights[969]), .RECT2_X(rectangle2_xs[969]), .RECT2_Y(rectangle2_ys[969]), .RECT2_WIDTH(rectangle2_widths[969]), .RECT2_HEIGHT(rectangle2_heights[969]), .RECT2_WEIGHT(rectangle2_weights[969]), .RECT3_X(rectangle3_xs[969]), .RECT3_Y(rectangle3_ys[969]), .RECT3_WIDTH(rectangle3_widths[969]), .RECT3_HEIGHT(rectangle3_heights[969]), .RECT3_WEIGHT(rectangle3_weights[969]), .FEAT_THRES(feature_thresholds[969]), .FEAT_ABOVE(feature_aboves[969]), .FEAT_BELOW(feature_belows[969])) ac969(.scan_win(scan_win969), .scan_win_std_dev(scan_win_std_dev[969]), .feature_accum(feature_accums[969]));
  accum_calculator #(.RECT1_X(rectangle1_xs[970]), .RECT1_Y(rectangle1_ys[970]), .RECT1_WIDTH(rectangle1_widths[970]), .RECT1_HEIGHT(rectangle1_heights[970]), .RECT1_WEIGHT(rectangle1_weights[970]), .RECT2_X(rectangle2_xs[970]), .RECT2_Y(rectangle2_ys[970]), .RECT2_WIDTH(rectangle2_widths[970]), .RECT2_HEIGHT(rectangle2_heights[970]), .RECT2_WEIGHT(rectangle2_weights[970]), .RECT3_X(rectangle3_xs[970]), .RECT3_Y(rectangle3_ys[970]), .RECT3_WIDTH(rectangle3_widths[970]), .RECT3_HEIGHT(rectangle3_heights[970]), .RECT3_WEIGHT(rectangle3_weights[970]), .FEAT_THRES(feature_thresholds[970]), .FEAT_ABOVE(feature_aboves[970]), .FEAT_BELOW(feature_belows[970])) ac970(.scan_win(scan_win970), .scan_win_std_dev(scan_win_std_dev[970]), .feature_accum(feature_accums[970]));
  accum_calculator #(.RECT1_X(rectangle1_xs[971]), .RECT1_Y(rectangle1_ys[971]), .RECT1_WIDTH(rectangle1_widths[971]), .RECT1_HEIGHT(rectangle1_heights[971]), .RECT1_WEIGHT(rectangle1_weights[971]), .RECT2_X(rectangle2_xs[971]), .RECT2_Y(rectangle2_ys[971]), .RECT2_WIDTH(rectangle2_widths[971]), .RECT2_HEIGHT(rectangle2_heights[971]), .RECT2_WEIGHT(rectangle2_weights[971]), .RECT3_X(rectangle3_xs[971]), .RECT3_Y(rectangle3_ys[971]), .RECT3_WIDTH(rectangle3_widths[971]), .RECT3_HEIGHT(rectangle3_heights[971]), .RECT3_WEIGHT(rectangle3_weights[971]), .FEAT_THRES(feature_thresholds[971]), .FEAT_ABOVE(feature_aboves[971]), .FEAT_BELOW(feature_belows[971])) ac971(.scan_win(scan_win971), .scan_win_std_dev(scan_win_std_dev[971]), .feature_accum(feature_accums[971]));
  accum_calculator #(.RECT1_X(rectangle1_xs[972]), .RECT1_Y(rectangle1_ys[972]), .RECT1_WIDTH(rectangle1_widths[972]), .RECT1_HEIGHT(rectangle1_heights[972]), .RECT1_WEIGHT(rectangle1_weights[972]), .RECT2_X(rectangle2_xs[972]), .RECT2_Y(rectangle2_ys[972]), .RECT2_WIDTH(rectangle2_widths[972]), .RECT2_HEIGHT(rectangle2_heights[972]), .RECT2_WEIGHT(rectangle2_weights[972]), .RECT3_X(rectangle3_xs[972]), .RECT3_Y(rectangle3_ys[972]), .RECT3_WIDTH(rectangle3_widths[972]), .RECT3_HEIGHT(rectangle3_heights[972]), .RECT3_WEIGHT(rectangle3_weights[972]), .FEAT_THRES(feature_thresholds[972]), .FEAT_ABOVE(feature_aboves[972]), .FEAT_BELOW(feature_belows[972])) ac972(.scan_win(scan_win972), .scan_win_std_dev(scan_win_std_dev[972]), .feature_accum(feature_accums[972]));
  accum_calculator #(.RECT1_X(rectangle1_xs[973]), .RECT1_Y(rectangle1_ys[973]), .RECT1_WIDTH(rectangle1_widths[973]), .RECT1_HEIGHT(rectangle1_heights[973]), .RECT1_WEIGHT(rectangle1_weights[973]), .RECT2_X(rectangle2_xs[973]), .RECT2_Y(rectangle2_ys[973]), .RECT2_WIDTH(rectangle2_widths[973]), .RECT2_HEIGHT(rectangle2_heights[973]), .RECT2_WEIGHT(rectangle2_weights[973]), .RECT3_X(rectangle3_xs[973]), .RECT3_Y(rectangle3_ys[973]), .RECT3_WIDTH(rectangle3_widths[973]), .RECT3_HEIGHT(rectangle3_heights[973]), .RECT3_WEIGHT(rectangle3_weights[973]), .FEAT_THRES(feature_thresholds[973]), .FEAT_ABOVE(feature_aboves[973]), .FEAT_BELOW(feature_belows[973])) ac973(.scan_win(scan_win973), .scan_win_std_dev(scan_win_std_dev[973]), .feature_accum(feature_accums[973]));
  accum_calculator #(.RECT1_X(rectangle1_xs[974]), .RECT1_Y(rectangle1_ys[974]), .RECT1_WIDTH(rectangle1_widths[974]), .RECT1_HEIGHT(rectangle1_heights[974]), .RECT1_WEIGHT(rectangle1_weights[974]), .RECT2_X(rectangle2_xs[974]), .RECT2_Y(rectangle2_ys[974]), .RECT2_WIDTH(rectangle2_widths[974]), .RECT2_HEIGHT(rectangle2_heights[974]), .RECT2_WEIGHT(rectangle2_weights[974]), .RECT3_X(rectangle3_xs[974]), .RECT3_Y(rectangle3_ys[974]), .RECT3_WIDTH(rectangle3_widths[974]), .RECT3_HEIGHT(rectangle3_heights[974]), .RECT3_WEIGHT(rectangle3_weights[974]), .FEAT_THRES(feature_thresholds[974]), .FEAT_ABOVE(feature_aboves[974]), .FEAT_BELOW(feature_belows[974])) ac974(.scan_win(scan_win974), .scan_win_std_dev(scan_win_std_dev[974]), .feature_accum(feature_accums[974]));
  accum_calculator #(.RECT1_X(rectangle1_xs[975]), .RECT1_Y(rectangle1_ys[975]), .RECT1_WIDTH(rectangle1_widths[975]), .RECT1_HEIGHT(rectangle1_heights[975]), .RECT1_WEIGHT(rectangle1_weights[975]), .RECT2_X(rectangle2_xs[975]), .RECT2_Y(rectangle2_ys[975]), .RECT2_WIDTH(rectangle2_widths[975]), .RECT2_HEIGHT(rectangle2_heights[975]), .RECT2_WEIGHT(rectangle2_weights[975]), .RECT3_X(rectangle3_xs[975]), .RECT3_Y(rectangle3_ys[975]), .RECT3_WIDTH(rectangle3_widths[975]), .RECT3_HEIGHT(rectangle3_heights[975]), .RECT3_WEIGHT(rectangle3_weights[975]), .FEAT_THRES(feature_thresholds[975]), .FEAT_ABOVE(feature_aboves[975]), .FEAT_BELOW(feature_belows[975])) ac975(.scan_win(scan_win975), .scan_win_std_dev(scan_win_std_dev[975]), .feature_accum(feature_accums[975]));
  accum_calculator #(.RECT1_X(rectangle1_xs[976]), .RECT1_Y(rectangle1_ys[976]), .RECT1_WIDTH(rectangle1_widths[976]), .RECT1_HEIGHT(rectangle1_heights[976]), .RECT1_WEIGHT(rectangle1_weights[976]), .RECT2_X(rectangle2_xs[976]), .RECT2_Y(rectangle2_ys[976]), .RECT2_WIDTH(rectangle2_widths[976]), .RECT2_HEIGHT(rectangle2_heights[976]), .RECT2_WEIGHT(rectangle2_weights[976]), .RECT3_X(rectangle3_xs[976]), .RECT3_Y(rectangle3_ys[976]), .RECT3_WIDTH(rectangle3_widths[976]), .RECT3_HEIGHT(rectangle3_heights[976]), .RECT3_WEIGHT(rectangle3_weights[976]), .FEAT_THRES(feature_thresholds[976]), .FEAT_ABOVE(feature_aboves[976]), .FEAT_BELOW(feature_belows[976])) ac976(.scan_win(scan_win976), .scan_win_std_dev(scan_win_std_dev[976]), .feature_accum(feature_accums[976]));
  accum_calculator #(.RECT1_X(rectangle1_xs[977]), .RECT1_Y(rectangle1_ys[977]), .RECT1_WIDTH(rectangle1_widths[977]), .RECT1_HEIGHT(rectangle1_heights[977]), .RECT1_WEIGHT(rectangle1_weights[977]), .RECT2_X(rectangle2_xs[977]), .RECT2_Y(rectangle2_ys[977]), .RECT2_WIDTH(rectangle2_widths[977]), .RECT2_HEIGHT(rectangle2_heights[977]), .RECT2_WEIGHT(rectangle2_weights[977]), .RECT3_X(rectangle3_xs[977]), .RECT3_Y(rectangle3_ys[977]), .RECT3_WIDTH(rectangle3_widths[977]), .RECT3_HEIGHT(rectangle3_heights[977]), .RECT3_WEIGHT(rectangle3_weights[977]), .FEAT_THRES(feature_thresholds[977]), .FEAT_ABOVE(feature_aboves[977]), .FEAT_BELOW(feature_belows[977])) ac977(.scan_win(scan_win977), .scan_win_std_dev(scan_win_std_dev[977]), .feature_accum(feature_accums[977]));
  accum_calculator #(.RECT1_X(rectangle1_xs[978]), .RECT1_Y(rectangle1_ys[978]), .RECT1_WIDTH(rectangle1_widths[978]), .RECT1_HEIGHT(rectangle1_heights[978]), .RECT1_WEIGHT(rectangle1_weights[978]), .RECT2_X(rectangle2_xs[978]), .RECT2_Y(rectangle2_ys[978]), .RECT2_WIDTH(rectangle2_widths[978]), .RECT2_HEIGHT(rectangle2_heights[978]), .RECT2_WEIGHT(rectangle2_weights[978]), .RECT3_X(rectangle3_xs[978]), .RECT3_Y(rectangle3_ys[978]), .RECT3_WIDTH(rectangle3_widths[978]), .RECT3_HEIGHT(rectangle3_heights[978]), .RECT3_WEIGHT(rectangle3_weights[978]), .FEAT_THRES(feature_thresholds[978]), .FEAT_ABOVE(feature_aboves[978]), .FEAT_BELOW(feature_belows[978])) ac978(.scan_win(scan_win978), .scan_win_std_dev(scan_win_std_dev[978]), .feature_accum(feature_accums[978]));
  accum_calculator #(.RECT1_X(rectangle1_xs[979]), .RECT1_Y(rectangle1_ys[979]), .RECT1_WIDTH(rectangle1_widths[979]), .RECT1_HEIGHT(rectangle1_heights[979]), .RECT1_WEIGHT(rectangle1_weights[979]), .RECT2_X(rectangle2_xs[979]), .RECT2_Y(rectangle2_ys[979]), .RECT2_WIDTH(rectangle2_widths[979]), .RECT2_HEIGHT(rectangle2_heights[979]), .RECT2_WEIGHT(rectangle2_weights[979]), .RECT3_X(rectangle3_xs[979]), .RECT3_Y(rectangle3_ys[979]), .RECT3_WIDTH(rectangle3_widths[979]), .RECT3_HEIGHT(rectangle3_heights[979]), .RECT3_WEIGHT(rectangle3_weights[979]), .FEAT_THRES(feature_thresholds[979]), .FEAT_ABOVE(feature_aboves[979]), .FEAT_BELOW(feature_belows[979])) ac979(.scan_win(scan_win979), .scan_win_std_dev(scan_win_std_dev[979]), .feature_accum(feature_accums[979]));
  accum_calculator #(.RECT1_X(rectangle1_xs[980]), .RECT1_Y(rectangle1_ys[980]), .RECT1_WIDTH(rectangle1_widths[980]), .RECT1_HEIGHT(rectangle1_heights[980]), .RECT1_WEIGHT(rectangle1_weights[980]), .RECT2_X(rectangle2_xs[980]), .RECT2_Y(rectangle2_ys[980]), .RECT2_WIDTH(rectangle2_widths[980]), .RECT2_HEIGHT(rectangle2_heights[980]), .RECT2_WEIGHT(rectangle2_weights[980]), .RECT3_X(rectangle3_xs[980]), .RECT3_Y(rectangle3_ys[980]), .RECT3_WIDTH(rectangle3_widths[980]), .RECT3_HEIGHT(rectangle3_heights[980]), .RECT3_WEIGHT(rectangle3_weights[980]), .FEAT_THRES(feature_thresholds[980]), .FEAT_ABOVE(feature_aboves[980]), .FEAT_BELOW(feature_belows[980])) ac980(.scan_win(scan_win980), .scan_win_std_dev(scan_win_std_dev[980]), .feature_accum(feature_accums[980]));
  accum_calculator #(.RECT1_X(rectangle1_xs[981]), .RECT1_Y(rectangle1_ys[981]), .RECT1_WIDTH(rectangle1_widths[981]), .RECT1_HEIGHT(rectangle1_heights[981]), .RECT1_WEIGHT(rectangle1_weights[981]), .RECT2_X(rectangle2_xs[981]), .RECT2_Y(rectangle2_ys[981]), .RECT2_WIDTH(rectangle2_widths[981]), .RECT2_HEIGHT(rectangle2_heights[981]), .RECT2_WEIGHT(rectangle2_weights[981]), .RECT3_X(rectangle3_xs[981]), .RECT3_Y(rectangle3_ys[981]), .RECT3_WIDTH(rectangle3_widths[981]), .RECT3_HEIGHT(rectangle3_heights[981]), .RECT3_WEIGHT(rectangle3_weights[981]), .FEAT_THRES(feature_thresholds[981]), .FEAT_ABOVE(feature_aboves[981]), .FEAT_BELOW(feature_belows[981])) ac981(.scan_win(scan_win981), .scan_win_std_dev(scan_win_std_dev[981]), .feature_accum(feature_accums[981]));
  accum_calculator #(.RECT1_X(rectangle1_xs[982]), .RECT1_Y(rectangle1_ys[982]), .RECT1_WIDTH(rectangle1_widths[982]), .RECT1_HEIGHT(rectangle1_heights[982]), .RECT1_WEIGHT(rectangle1_weights[982]), .RECT2_X(rectangle2_xs[982]), .RECT2_Y(rectangle2_ys[982]), .RECT2_WIDTH(rectangle2_widths[982]), .RECT2_HEIGHT(rectangle2_heights[982]), .RECT2_WEIGHT(rectangle2_weights[982]), .RECT3_X(rectangle3_xs[982]), .RECT3_Y(rectangle3_ys[982]), .RECT3_WIDTH(rectangle3_widths[982]), .RECT3_HEIGHT(rectangle3_heights[982]), .RECT3_WEIGHT(rectangle3_weights[982]), .FEAT_THRES(feature_thresholds[982]), .FEAT_ABOVE(feature_aboves[982]), .FEAT_BELOW(feature_belows[982])) ac982(.scan_win(scan_win982), .scan_win_std_dev(scan_win_std_dev[982]), .feature_accum(feature_accums[982]));
  accum_calculator #(.RECT1_X(rectangle1_xs[983]), .RECT1_Y(rectangle1_ys[983]), .RECT1_WIDTH(rectangle1_widths[983]), .RECT1_HEIGHT(rectangle1_heights[983]), .RECT1_WEIGHT(rectangle1_weights[983]), .RECT2_X(rectangle2_xs[983]), .RECT2_Y(rectangle2_ys[983]), .RECT2_WIDTH(rectangle2_widths[983]), .RECT2_HEIGHT(rectangle2_heights[983]), .RECT2_WEIGHT(rectangle2_weights[983]), .RECT3_X(rectangle3_xs[983]), .RECT3_Y(rectangle3_ys[983]), .RECT3_WIDTH(rectangle3_widths[983]), .RECT3_HEIGHT(rectangle3_heights[983]), .RECT3_WEIGHT(rectangle3_weights[983]), .FEAT_THRES(feature_thresholds[983]), .FEAT_ABOVE(feature_aboves[983]), .FEAT_BELOW(feature_belows[983])) ac983(.scan_win(scan_win983), .scan_win_std_dev(scan_win_std_dev[983]), .feature_accum(feature_accums[983]));
  accum_calculator #(.RECT1_X(rectangle1_xs[984]), .RECT1_Y(rectangle1_ys[984]), .RECT1_WIDTH(rectangle1_widths[984]), .RECT1_HEIGHT(rectangle1_heights[984]), .RECT1_WEIGHT(rectangle1_weights[984]), .RECT2_X(rectangle2_xs[984]), .RECT2_Y(rectangle2_ys[984]), .RECT2_WIDTH(rectangle2_widths[984]), .RECT2_HEIGHT(rectangle2_heights[984]), .RECT2_WEIGHT(rectangle2_weights[984]), .RECT3_X(rectangle3_xs[984]), .RECT3_Y(rectangle3_ys[984]), .RECT3_WIDTH(rectangle3_widths[984]), .RECT3_HEIGHT(rectangle3_heights[984]), .RECT3_WEIGHT(rectangle3_weights[984]), .FEAT_THRES(feature_thresholds[984]), .FEAT_ABOVE(feature_aboves[984]), .FEAT_BELOW(feature_belows[984])) ac984(.scan_win(scan_win984), .scan_win_std_dev(scan_win_std_dev[984]), .feature_accum(feature_accums[984]));
  accum_calculator #(.RECT1_X(rectangle1_xs[985]), .RECT1_Y(rectangle1_ys[985]), .RECT1_WIDTH(rectangle1_widths[985]), .RECT1_HEIGHT(rectangle1_heights[985]), .RECT1_WEIGHT(rectangle1_weights[985]), .RECT2_X(rectangle2_xs[985]), .RECT2_Y(rectangle2_ys[985]), .RECT2_WIDTH(rectangle2_widths[985]), .RECT2_HEIGHT(rectangle2_heights[985]), .RECT2_WEIGHT(rectangle2_weights[985]), .RECT3_X(rectangle3_xs[985]), .RECT3_Y(rectangle3_ys[985]), .RECT3_WIDTH(rectangle3_widths[985]), .RECT3_HEIGHT(rectangle3_heights[985]), .RECT3_WEIGHT(rectangle3_weights[985]), .FEAT_THRES(feature_thresholds[985]), .FEAT_ABOVE(feature_aboves[985]), .FEAT_BELOW(feature_belows[985])) ac985(.scan_win(scan_win985), .scan_win_std_dev(scan_win_std_dev[985]), .feature_accum(feature_accums[985]));
  accum_calculator #(.RECT1_X(rectangle1_xs[986]), .RECT1_Y(rectangle1_ys[986]), .RECT1_WIDTH(rectangle1_widths[986]), .RECT1_HEIGHT(rectangle1_heights[986]), .RECT1_WEIGHT(rectangle1_weights[986]), .RECT2_X(rectangle2_xs[986]), .RECT2_Y(rectangle2_ys[986]), .RECT2_WIDTH(rectangle2_widths[986]), .RECT2_HEIGHT(rectangle2_heights[986]), .RECT2_WEIGHT(rectangle2_weights[986]), .RECT3_X(rectangle3_xs[986]), .RECT3_Y(rectangle3_ys[986]), .RECT3_WIDTH(rectangle3_widths[986]), .RECT3_HEIGHT(rectangle3_heights[986]), .RECT3_WEIGHT(rectangle3_weights[986]), .FEAT_THRES(feature_thresholds[986]), .FEAT_ABOVE(feature_aboves[986]), .FEAT_BELOW(feature_belows[986])) ac986(.scan_win(scan_win986), .scan_win_std_dev(scan_win_std_dev[986]), .feature_accum(feature_accums[986]));
  accum_calculator #(.RECT1_X(rectangle1_xs[987]), .RECT1_Y(rectangle1_ys[987]), .RECT1_WIDTH(rectangle1_widths[987]), .RECT1_HEIGHT(rectangle1_heights[987]), .RECT1_WEIGHT(rectangle1_weights[987]), .RECT2_X(rectangle2_xs[987]), .RECT2_Y(rectangle2_ys[987]), .RECT2_WIDTH(rectangle2_widths[987]), .RECT2_HEIGHT(rectangle2_heights[987]), .RECT2_WEIGHT(rectangle2_weights[987]), .RECT3_X(rectangle3_xs[987]), .RECT3_Y(rectangle3_ys[987]), .RECT3_WIDTH(rectangle3_widths[987]), .RECT3_HEIGHT(rectangle3_heights[987]), .RECT3_WEIGHT(rectangle3_weights[987]), .FEAT_THRES(feature_thresholds[987]), .FEAT_ABOVE(feature_aboves[987]), .FEAT_BELOW(feature_belows[987])) ac987(.scan_win(scan_win987), .scan_win_std_dev(scan_win_std_dev[987]), .feature_accum(feature_accums[987]));
  accum_calculator #(.RECT1_X(rectangle1_xs[988]), .RECT1_Y(rectangle1_ys[988]), .RECT1_WIDTH(rectangle1_widths[988]), .RECT1_HEIGHT(rectangle1_heights[988]), .RECT1_WEIGHT(rectangle1_weights[988]), .RECT2_X(rectangle2_xs[988]), .RECT2_Y(rectangle2_ys[988]), .RECT2_WIDTH(rectangle2_widths[988]), .RECT2_HEIGHT(rectangle2_heights[988]), .RECT2_WEIGHT(rectangle2_weights[988]), .RECT3_X(rectangle3_xs[988]), .RECT3_Y(rectangle3_ys[988]), .RECT3_WIDTH(rectangle3_widths[988]), .RECT3_HEIGHT(rectangle3_heights[988]), .RECT3_WEIGHT(rectangle3_weights[988]), .FEAT_THRES(feature_thresholds[988]), .FEAT_ABOVE(feature_aboves[988]), .FEAT_BELOW(feature_belows[988])) ac988(.scan_win(scan_win988), .scan_win_std_dev(scan_win_std_dev[988]), .feature_accum(feature_accums[988]));
  accum_calculator #(.RECT1_X(rectangle1_xs[989]), .RECT1_Y(rectangle1_ys[989]), .RECT1_WIDTH(rectangle1_widths[989]), .RECT1_HEIGHT(rectangle1_heights[989]), .RECT1_WEIGHT(rectangle1_weights[989]), .RECT2_X(rectangle2_xs[989]), .RECT2_Y(rectangle2_ys[989]), .RECT2_WIDTH(rectangle2_widths[989]), .RECT2_HEIGHT(rectangle2_heights[989]), .RECT2_WEIGHT(rectangle2_weights[989]), .RECT3_X(rectangle3_xs[989]), .RECT3_Y(rectangle3_ys[989]), .RECT3_WIDTH(rectangle3_widths[989]), .RECT3_HEIGHT(rectangle3_heights[989]), .RECT3_WEIGHT(rectangle3_weights[989]), .FEAT_THRES(feature_thresholds[989]), .FEAT_ABOVE(feature_aboves[989]), .FEAT_BELOW(feature_belows[989])) ac989(.scan_win(scan_win989), .scan_win_std_dev(scan_win_std_dev[989]), .feature_accum(feature_accums[989]));
  accum_calculator #(.RECT1_X(rectangle1_xs[990]), .RECT1_Y(rectangle1_ys[990]), .RECT1_WIDTH(rectangle1_widths[990]), .RECT1_HEIGHT(rectangle1_heights[990]), .RECT1_WEIGHT(rectangle1_weights[990]), .RECT2_X(rectangle2_xs[990]), .RECT2_Y(rectangle2_ys[990]), .RECT2_WIDTH(rectangle2_widths[990]), .RECT2_HEIGHT(rectangle2_heights[990]), .RECT2_WEIGHT(rectangle2_weights[990]), .RECT3_X(rectangle3_xs[990]), .RECT3_Y(rectangle3_ys[990]), .RECT3_WIDTH(rectangle3_widths[990]), .RECT3_HEIGHT(rectangle3_heights[990]), .RECT3_WEIGHT(rectangle3_weights[990]), .FEAT_THRES(feature_thresholds[990]), .FEAT_ABOVE(feature_aboves[990]), .FEAT_BELOW(feature_belows[990])) ac990(.scan_win(scan_win990), .scan_win_std_dev(scan_win_std_dev[990]), .feature_accum(feature_accums[990]));
  accum_calculator #(.RECT1_X(rectangle1_xs[991]), .RECT1_Y(rectangle1_ys[991]), .RECT1_WIDTH(rectangle1_widths[991]), .RECT1_HEIGHT(rectangle1_heights[991]), .RECT1_WEIGHT(rectangle1_weights[991]), .RECT2_X(rectangle2_xs[991]), .RECT2_Y(rectangle2_ys[991]), .RECT2_WIDTH(rectangle2_widths[991]), .RECT2_HEIGHT(rectangle2_heights[991]), .RECT2_WEIGHT(rectangle2_weights[991]), .RECT3_X(rectangle3_xs[991]), .RECT3_Y(rectangle3_ys[991]), .RECT3_WIDTH(rectangle3_widths[991]), .RECT3_HEIGHT(rectangle3_heights[991]), .RECT3_WEIGHT(rectangle3_weights[991]), .FEAT_THRES(feature_thresholds[991]), .FEAT_ABOVE(feature_aboves[991]), .FEAT_BELOW(feature_belows[991])) ac991(.scan_win(scan_win991), .scan_win_std_dev(scan_win_std_dev[991]), .feature_accum(feature_accums[991]));
  accum_calculator #(.RECT1_X(rectangle1_xs[992]), .RECT1_Y(rectangle1_ys[992]), .RECT1_WIDTH(rectangle1_widths[992]), .RECT1_HEIGHT(rectangle1_heights[992]), .RECT1_WEIGHT(rectangle1_weights[992]), .RECT2_X(rectangle2_xs[992]), .RECT2_Y(rectangle2_ys[992]), .RECT2_WIDTH(rectangle2_widths[992]), .RECT2_HEIGHT(rectangle2_heights[992]), .RECT2_WEIGHT(rectangle2_weights[992]), .RECT3_X(rectangle3_xs[992]), .RECT3_Y(rectangle3_ys[992]), .RECT3_WIDTH(rectangle3_widths[992]), .RECT3_HEIGHT(rectangle3_heights[992]), .RECT3_WEIGHT(rectangle3_weights[992]), .FEAT_THRES(feature_thresholds[992]), .FEAT_ABOVE(feature_aboves[992]), .FEAT_BELOW(feature_belows[992])) ac992(.scan_win(scan_win992), .scan_win_std_dev(scan_win_std_dev[992]), .feature_accum(feature_accums[992]));
  accum_calculator #(.RECT1_X(rectangle1_xs[993]), .RECT1_Y(rectangle1_ys[993]), .RECT1_WIDTH(rectangle1_widths[993]), .RECT1_HEIGHT(rectangle1_heights[993]), .RECT1_WEIGHT(rectangle1_weights[993]), .RECT2_X(rectangle2_xs[993]), .RECT2_Y(rectangle2_ys[993]), .RECT2_WIDTH(rectangle2_widths[993]), .RECT2_HEIGHT(rectangle2_heights[993]), .RECT2_WEIGHT(rectangle2_weights[993]), .RECT3_X(rectangle3_xs[993]), .RECT3_Y(rectangle3_ys[993]), .RECT3_WIDTH(rectangle3_widths[993]), .RECT3_HEIGHT(rectangle3_heights[993]), .RECT3_WEIGHT(rectangle3_weights[993]), .FEAT_THRES(feature_thresholds[993]), .FEAT_ABOVE(feature_aboves[993]), .FEAT_BELOW(feature_belows[993])) ac993(.scan_win(scan_win993), .scan_win_std_dev(scan_win_std_dev[993]), .feature_accum(feature_accums[993]));
  accum_calculator #(.RECT1_X(rectangle1_xs[994]), .RECT1_Y(rectangle1_ys[994]), .RECT1_WIDTH(rectangle1_widths[994]), .RECT1_HEIGHT(rectangle1_heights[994]), .RECT1_WEIGHT(rectangle1_weights[994]), .RECT2_X(rectangle2_xs[994]), .RECT2_Y(rectangle2_ys[994]), .RECT2_WIDTH(rectangle2_widths[994]), .RECT2_HEIGHT(rectangle2_heights[994]), .RECT2_WEIGHT(rectangle2_weights[994]), .RECT3_X(rectangle3_xs[994]), .RECT3_Y(rectangle3_ys[994]), .RECT3_WIDTH(rectangle3_widths[994]), .RECT3_HEIGHT(rectangle3_heights[994]), .RECT3_WEIGHT(rectangle3_weights[994]), .FEAT_THRES(feature_thresholds[994]), .FEAT_ABOVE(feature_aboves[994]), .FEAT_BELOW(feature_belows[994])) ac994(.scan_win(scan_win994), .scan_win_std_dev(scan_win_std_dev[994]), .feature_accum(feature_accums[994]));
  accum_calculator #(.RECT1_X(rectangle1_xs[995]), .RECT1_Y(rectangle1_ys[995]), .RECT1_WIDTH(rectangle1_widths[995]), .RECT1_HEIGHT(rectangle1_heights[995]), .RECT1_WEIGHT(rectangle1_weights[995]), .RECT2_X(rectangle2_xs[995]), .RECT2_Y(rectangle2_ys[995]), .RECT2_WIDTH(rectangle2_widths[995]), .RECT2_HEIGHT(rectangle2_heights[995]), .RECT2_WEIGHT(rectangle2_weights[995]), .RECT3_X(rectangle3_xs[995]), .RECT3_Y(rectangle3_ys[995]), .RECT3_WIDTH(rectangle3_widths[995]), .RECT3_HEIGHT(rectangle3_heights[995]), .RECT3_WEIGHT(rectangle3_weights[995]), .FEAT_THRES(feature_thresholds[995]), .FEAT_ABOVE(feature_aboves[995]), .FEAT_BELOW(feature_belows[995])) ac995(.scan_win(scan_win995), .scan_win_std_dev(scan_win_std_dev[995]), .feature_accum(feature_accums[995]));
  accum_calculator #(.RECT1_X(rectangle1_xs[996]), .RECT1_Y(rectangle1_ys[996]), .RECT1_WIDTH(rectangle1_widths[996]), .RECT1_HEIGHT(rectangle1_heights[996]), .RECT1_WEIGHT(rectangle1_weights[996]), .RECT2_X(rectangle2_xs[996]), .RECT2_Y(rectangle2_ys[996]), .RECT2_WIDTH(rectangle2_widths[996]), .RECT2_HEIGHT(rectangle2_heights[996]), .RECT2_WEIGHT(rectangle2_weights[996]), .RECT3_X(rectangle3_xs[996]), .RECT3_Y(rectangle3_ys[996]), .RECT3_WIDTH(rectangle3_widths[996]), .RECT3_HEIGHT(rectangle3_heights[996]), .RECT3_WEIGHT(rectangle3_weights[996]), .FEAT_THRES(feature_thresholds[996]), .FEAT_ABOVE(feature_aboves[996]), .FEAT_BELOW(feature_belows[996])) ac996(.scan_win(scan_win996), .scan_win_std_dev(scan_win_std_dev[996]), .feature_accum(feature_accums[996]));
  accum_calculator #(.RECT1_X(rectangle1_xs[997]), .RECT1_Y(rectangle1_ys[997]), .RECT1_WIDTH(rectangle1_widths[997]), .RECT1_HEIGHT(rectangle1_heights[997]), .RECT1_WEIGHT(rectangle1_weights[997]), .RECT2_X(rectangle2_xs[997]), .RECT2_Y(rectangle2_ys[997]), .RECT2_WIDTH(rectangle2_widths[997]), .RECT2_HEIGHT(rectangle2_heights[997]), .RECT2_WEIGHT(rectangle2_weights[997]), .RECT3_X(rectangle3_xs[997]), .RECT3_Y(rectangle3_ys[997]), .RECT3_WIDTH(rectangle3_widths[997]), .RECT3_HEIGHT(rectangle3_heights[997]), .RECT3_WEIGHT(rectangle3_weights[997]), .FEAT_THRES(feature_thresholds[997]), .FEAT_ABOVE(feature_aboves[997]), .FEAT_BELOW(feature_belows[997])) ac997(.scan_win(scan_win997), .scan_win_std_dev(scan_win_std_dev[997]), .feature_accum(feature_accums[997]));
  accum_calculator #(.RECT1_X(rectangle1_xs[998]), .RECT1_Y(rectangle1_ys[998]), .RECT1_WIDTH(rectangle1_widths[998]), .RECT1_HEIGHT(rectangle1_heights[998]), .RECT1_WEIGHT(rectangle1_weights[998]), .RECT2_X(rectangle2_xs[998]), .RECT2_Y(rectangle2_ys[998]), .RECT2_WIDTH(rectangle2_widths[998]), .RECT2_HEIGHT(rectangle2_heights[998]), .RECT2_WEIGHT(rectangle2_weights[998]), .RECT3_X(rectangle3_xs[998]), .RECT3_Y(rectangle3_ys[998]), .RECT3_WIDTH(rectangle3_widths[998]), .RECT3_HEIGHT(rectangle3_heights[998]), .RECT3_WEIGHT(rectangle3_weights[998]), .FEAT_THRES(feature_thresholds[998]), .FEAT_ABOVE(feature_aboves[998]), .FEAT_BELOW(feature_belows[998])) ac998(.scan_win(scan_win998), .scan_win_std_dev(scan_win_std_dev[998]), .feature_accum(feature_accums[998]));
  accum_calculator #(.RECT1_X(rectangle1_xs[999]), .RECT1_Y(rectangle1_ys[999]), .RECT1_WIDTH(rectangle1_widths[999]), .RECT1_HEIGHT(rectangle1_heights[999]), .RECT1_WEIGHT(rectangle1_weights[999]), .RECT2_X(rectangle2_xs[999]), .RECT2_Y(rectangle2_ys[999]), .RECT2_WIDTH(rectangle2_widths[999]), .RECT2_HEIGHT(rectangle2_heights[999]), .RECT2_WEIGHT(rectangle2_weights[999]), .RECT3_X(rectangle3_xs[999]), .RECT3_Y(rectangle3_ys[999]), .RECT3_WIDTH(rectangle3_widths[999]), .RECT3_HEIGHT(rectangle3_heights[999]), .RECT3_WEIGHT(rectangle3_weights[999]), .FEAT_THRES(feature_thresholds[999]), .FEAT_ABOVE(feature_aboves[999]), .FEAT_BELOW(feature_belows[999])) ac999(.scan_win(scan_win999), .scan_win_std_dev(scan_win_std_dev[999]), .feature_accum(feature_accums[999]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1000]), .RECT1_Y(rectangle1_ys[1000]), .RECT1_WIDTH(rectangle1_widths[1000]), .RECT1_HEIGHT(rectangle1_heights[1000]), .RECT1_WEIGHT(rectangle1_weights[1000]), .RECT2_X(rectangle2_xs[1000]), .RECT2_Y(rectangle2_ys[1000]), .RECT2_WIDTH(rectangle2_widths[1000]), .RECT2_HEIGHT(rectangle2_heights[1000]), .RECT2_WEIGHT(rectangle2_weights[1000]), .RECT3_X(rectangle3_xs[1000]), .RECT3_Y(rectangle3_ys[1000]), .RECT3_WIDTH(rectangle3_widths[1000]), .RECT3_HEIGHT(rectangle3_heights[1000]), .RECT3_WEIGHT(rectangle3_weights[1000]), .FEAT_THRES(feature_thresholds[1000]), .FEAT_ABOVE(feature_aboves[1000]), .FEAT_BELOW(feature_belows[1000])) ac1000(.scan_win(scan_win1000), .scan_win_std_dev(scan_win_std_dev[1000]), .feature_accum(feature_accums[1000]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1001]), .RECT1_Y(rectangle1_ys[1001]), .RECT1_WIDTH(rectangle1_widths[1001]), .RECT1_HEIGHT(rectangle1_heights[1001]), .RECT1_WEIGHT(rectangle1_weights[1001]), .RECT2_X(rectangle2_xs[1001]), .RECT2_Y(rectangle2_ys[1001]), .RECT2_WIDTH(rectangle2_widths[1001]), .RECT2_HEIGHT(rectangle2_heights[1001]), .RECT2_WEIGHT(rectangle2_weights[1001]), .RECT3_X(rectangle3_xs[1001]), .RECT3_Y(rectangle3_ys[1001]), .RECT3_WIDTH(rectangle3_widths[1001]), .RECT3_HEIGHT(rectangle3_heights[1001]), .RECT3_WEIGHT(rectangle3_weights[1001]), .FEAT_THRES(feature_thresholds[1001]), .FEAT_ABOVE(feature_aboves[1001]), .FEAT_BELOW(feature_belows[1001])) ac1001(.scan_win(scan_win1001), .scan_win_std_dev(scan_win_std_dev[1001]), .feature_accum(feature_accums[1001]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1002]), .RECT1_Y(rectangle1_ys[1002]), .RECT1_WIDTH(rectangle1_widths[1002]), .RECT1_HEIGHT(rectangle1_heights[1002]), .RECT1_WEIGHT(rectangle1_weights[1002]), .RECT2_X(rectangle2_xs[1002]), .RECT2_Y(rectangle2_ys[1002]), .RECT2_WIDTH(rectangle2_widths[1002]), .RECT2_HEIGHT(rectangle2_heights[1002]), .RECT2_WEIGHT(rectangle2_weights[1002]), .RECT3_X(rectangle3_xs[1002]), .RECT3_Y(rectangle3_ys[1002]), .RECT3_WIDTH(rectangle3_widths[1002]), .RECT3_HEIGHT(rectangle3_heights[1002]), .RECT3_WEIGHT(rectangle3_weights[1002]), .FEAT_THRES(feature_thresholds[1002]), .FEAT_ABOVE(feature_aboves[1002]), .FEAT_BELOW(feature_belows[1002])) ac1002(.scan_win(scan_win1002), .scan_win_std_dev(scan_win_std_dev[1002]), .feature_accum(feature_accums[1002]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1003]), .RECT1_Y(rectangle1_ys[1003]), .RECT1_WIDTH(rectangle1_widths[1003]), .RECT1_HEIGHT(rectangle1_heights[1003]), .RECT1_WEIGHT(rectangle1_weights[1003]), .RECT2_X(rectangle2_xs[1003]), .RECT2_Y(rectangle2_ys[1003]), .RECT2_WIDTH(rectangle2_widths[1003]), .RECT2_HEIGHT(rectangle2_heights[1003]), .RECT2_WEIGHT(rectangle2_weights[1003]), .RECT3_X(rectangle3_xs[1003]), .RECT3_Y(rectangle3_ys[1003]), .RECT3_WIDTH(rectangle3_widths[1003]), .RECT3_HEIGHT(rectangle3_heights[1003]), .RECT3_WEIGHT(rectangle3_weights[1003]), .FEAT_THRES(feature_thresholds[1003]), .FEAT_ABOVE(feature_aboves[1003]), .FEAT_BELOW(feature_belows[1003])) ac1003(.scan_win(scan_win1003), .scan_win_std_dev(scan_win_std_dev[1003]), .feature_accum(feature_accums[1003]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1004]), .RECT1_Y(rectangle1_ys[1004]), .RECT1_WIDTH(rectangle1_widths[1004]), .RECT1_HEIGHT(rectangle1_heights[1004]), .RECT1_WEIGHT(rectangle1_weights[1004]), .RECT2_X(rectangle2_xs[1004]), .RECT2_Y(rectangle2_ys[1004]), .RECT2_WIDTH(rectangle2_widths[1004]), .RECT2_HEIGHT(rectangle2_heights[1004]), .RECT2_WEIGHT(rectangle2_weights[1004]), .RECT3_X(rectangle3_xs[1004]), .RECT3_Y(rectangle3_ys[1004]), .RECT3_WIDTH(rectangle3_widths[1004]), .RECT3_HEIGHT(rectangle3_heights[1004]), .RECT3_WEIGHT(rectangle3_weights[1004]), .FEAT_THRES(feature_thresholds[1004]), .FEAT_ABOVE(feature_aboves[1004]), .FEAT_BELOW(feature_belows[1004])) ac1004(.scan_win(scan_win1004), .scan_win_std_dev(scan_win_std_dev[1004]), .feature_accum(feature_accums[1004]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1005]), .RECT1_Y(rectangle1_ys[1005]), .RECT1_WIDTH(rectangle1_widths[1005]), .RECT1_HEIGHT(rectangle1_heights[1005]), .RECT1_WEIGHT(rectangle1_weights[1005]), .RECT2_X(rectangle2_xs[1005]), .RECT2_Y(rectangle2_ys[1005]), .RECT2_WIDTH(rectangle2_widths[1005]), .RECT2_HEIGHT(rectangle2_heights[1005]), .RECT2_WEIGHT(rectangle2_weights[1005]), .RECT3_X(rectangle3_xs[1005]), .RECT3_Y(rectangle3_ys[1005]), .RECT3_WIDTH(rectangle3_widths[1005]), .RECT3_HEIGHT(rectangle3_heights[1005]), .RECT3_WEIGHT(rectangle3_weights[1005]), .FEAT_THRES(feature_thresholds[1005]), .FEAT_ABOVE(feature_aboves[1005]), .FEAT_BELOW(feature_belows[1005])) ac1005(.scan_win(scan_win1005), .scan_win_std_dev(scan_win_std_dev[1005]), .feature_accum(feature_accums[1005]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1006]), .RECT1_Y(rectangle1_ys[1006]), .RECT1_WIDTH(rectangle1_widths[1006]), .RECT1_HEIGHT(rectangle1_heights[1006]), .RECT1_WEIGHT(rectangle1_weights[1006]), .RECT2_X(rectangle2_xs[1006]), .RECT2_Y(rectangle2_ys[1006]), .RECT2_WIDTH(rectangle2_widths[1006]), .RECT2_HEIGHT(rectangle2_heights[1006]), .RECT2_WEIGHT(rectangle2_weights[1006]), .RECT3_X(rectangle3_xs[1006]), .RECT3_Y(rectangle3_ys[1006]), .RECT3_WIDTH(rectangle3_widths[1006]), .RECT3_HEIGHT(rectangle3_heights[1006]), .RECT3_WEIGHT(rectangle3_weights[1006]), .FEAT_THRES(feature_thresholds[1006]), .FEAT_ABOVE(feature_aboves[1006]), .FEAT_BELOW(feature_belows[1006])) ac1006(.scan_win(scan_win1006), .scan_win_std_dev(scan_win_std_dev[1006]), .feature_accum(feature_accums[1006]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1007]), .RECT1_Y(rectangle1_ys[1007]), .RECT1_WIDTH(rectangle1_widths[1007]), .RECT1_HEIGHT(rectangle1_heights[1007]), .RECT1_WEIGHT(rectangle1_weights[1007]), .RECT2_X(rectangle2_xs[1007]), .RECT2_Y(rectangle2_ys[1007]), .RECT2_WIDTH(rectangle2_widths[1007]), .RECT2_HEIGHT(rectangle2_heights[1007]), .RECT2_WEIGHT(rectangle2_weights[1007]), .RECT3_X(rectangle3_xs[1007]), .RECT3_Y(rectangle3_ys[1007]), .RECT3_WIDTH(rectangle3_widths[1007]), .RECT3_HEIGHT(rectangle3_heights[1007]), .RECT3_WEIGHT(rectangle3_weights[1007]), .FEAT_THRES(feature_thresholds[1007]), .FEAT_ABOVE(feature_aboves[1007]), .FEAT_BELOW(feature_belows[1007])) ac1007(.scan_win(scan_win1007), .scan_win_std_dev(scan_win_std_dev[1007]), .feature_accum(feature_accums[1007]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1008]), .RECT1_Y(rectangle1_ys[1008]), .RECT1_WIDTH(rectangle1_widths[1008]), .RECT1_HEIGHT(rectangle1_heights[1008]), .RECT1_WEIGHT(rectangle1_weights[1008]), .RECT2_X(rectangle2_xs[1008]), .RECT2_Y(rectangle2_ys[1008]), .RECT2_WIDTH(rectangle2_widths[1008]), .RECT2_HEIGHT(rectangle2_heights[1008]), .RECT2_WEIGHT(rectangle2_weights[1008]), .RECT3_X(rectangle3_xs[1008]), .RECT3_Y(rectangle3_ys[1008]), .RECT3_WIDTH(rectangle3_widths[1008]), .RECT3_HEIGHT(rectangle3_heights[1008]), .RECT3_WEIGHT(rectangle3_weights[1008]), .FEAT_THRES(feature_thresholds[1008]), .FEAT_ABOVE(feature_aboves[1008]), .FEAT_BELOW(feature_belows[1008])) ac1008(.scan_win(scan_win1008), .scan_win_std_dev(scan_win_std_dev[1008]), .feature_accum(feature_accums[1008]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1009]), .RECT1_Y(rectangle1_ys[1009]), .RECT1_WIDTH(rectangle1_widths[1009]), .RECT1_HEIGHT(rectangle1_heights[1009]), .RECT1_WEIGHT(rectangle1_weights[1009]), .RECT2_X(rectangle2_xs[1009]), .RECT2_Y(rectangle2_ys[1009]), .RECT2_WIDTH(rectangle2_widths[1009]), .RECT2_HEIGHT(rectangle2_heights[1009]), .RECT2_WEIGHT(rectangle2_weights[1009]), .RECT3_X(rectangle3_xs[1009]), .RECT3_Y(rectangle3_ys[1009]), .RECT3_WIDTH(rectangle3_widths[1009]), .RECT3_HEIGHT(rectangle3_heights[1009]), .RECT3_WEIGHT(rectangle3_weights[1009]), .FEAT_THRES(feature_thresholds[1009]), .FEAT_ABOVE(feature_aboves[1009]), .FEAT_BELOW(feature_belows[1009])) ac1009(.scan_win(scan_win1009), .scan_win_std_dev(scan_win_std_dev[1009]), .feature_accum(feature_accums[1009]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1010]), .RECT1_Y(rectangle1_ys[1010]), .RECT1_WIDTH(rectangle1_widths[1010]), .RECT1_HEIGHT(rectangle1_heights[1010]), .RECT1_WEIGHT(rectangle1_weights[1010]), .RECT2_X(rectangle2_xs[1010]), .RECT2_Y(rectangle2_ys[1010]), .RECT2_WIDTH(rectangle2_widths[1010]), .RECT2_HEIGHT(rectangle2_heights[1010]), .RECT2_WEIGHT(rectangle2_weights[1010]), .RECT3_X(rectangle3_xs[1010]), .RECT3_Y(rectangle3_ys[1010]), .RECT3_WIDTH(rectangle3_widths[1010]), .RECT3_HEIGHT(rectangle3_heights[1010]), .RECT3_WEIGHT(rectangle3_weights[1010]), .FEAT_THRES(feature_thresholds[1010]), .FEAT_ABOVE(feature_aboves[1010]), .FEAT_BELOW(feature_belows[1010])) ac1010(.scan_win(scan_win1010), .scan_win_std_dev(scan_win_std_dev[1010]), .feature_accum(feature_accums[1010]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1011]), .RECT1_Y(rectangle1_ys[1011]), .RECT1_WIDTH(rectangle1_widths[1011]), .RECT1_HEIGHT(rectangle1_heights[1011]), .RECT1_WEIGHT(rectangle1_weights[1011]), .RECT2_X(rectangle2_xs[1011]), .RECT2_Y(rectangle2_ys[1011]), .RECT2_WIDTH(rectangle2_widths[1011]), .RECT2_HEIGHT(rectangle2_heights[1011]), .RECT2_WEIGHT(rectangle2_weights[1011]), .RECT3_X(rectangle3_xs[1011]), .RECT3_Y(rectangle3_ys[1011]), .RECT3_WIDTH(rectangle3_widths[1011]), .RECT3_HEIGHT(rectangle3_heights[1011]), .RECT3_WEIGHT(rectangle3_weights[1011]), .FEAT_THRES(feature_thresholds[1011]), .FEAT_ABOVE(feature_aboves[1011]), .FEAT_BELOW(feature_belows[1011])) ac1011(.scan_win(scan_win1011), .scan_win_std_dev(scan_win_std_dev[1011]), .feature_accum(feature_accums[1011]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1012]), .RECT1_Y(rectangle1_ys[1012]), .RECT1_WIDTH(rectangle1_widths[1012]), .RECT1_HEIGHT(rectangle1_heights[1012]), .RECT1_WEIGHT(rectangle1_weights[1012]), .RECT2_X(rectangle2_xs[1012]), .RECT2_Y(rectangle2_ys[1012]), .RECT2_WIDTH(rectangle2_widths[1012]), .RECT2_HEIGHT(rectangle2_heights[1012]), .RECT2_WEIGHT(rectangle2_weights[1012]), .RECT3_X(rectangle3_xs[1012]), .RECT3_Y(rectangle3_ys[1012]), .RECT3_WIDTH(rectangle3_widths[1012]), .RECT3_HEIGHT(rectangle3_heights[1012]), .RECT3_WEIGHT(rectangle3_weights[1012]), .FEAT_THRES(feature_thresholds[1012]), .FEAT_ABOVE(feature_aboves[1012]), .FEAT_BELOW(feature_belows[1012])) ac1012(.scan_win(scan_win1012), .scan_win_std_dev(scan_win_std_dev[1012]), .feature_accum(feature_accums[1012]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1013]), .RECT1_Y(rectangle1_ys[1013]), .RECT1_WIDTH(rectangle1_widths[1013]), .RECT1_HEIGHT(rectangle1_heights[1013]), .RECT1_WEIGHT(rectangle1_weights[1013]), .RECT2_X(rectangle2_xs[1013]), .RECT2_Y(rectangle2_ys[1013]), .RECT2_WIDTH(rectangle2_widths[1013]), .RECT2_HEIGHT(rectangle2_heights[1013]), .RECT2_WEIGHT(rectangle2_weights[1013]), .RECT3_X(rectangle3_xs[1013]), .RECT3_Y(rectangle3_ys[1013]), .RECT3_WIDTH(rectangle3_widths[1013]), .RECT3_HEIGHT(rectangle3_heights[1013]), .RECT3_WEIGHT(rectangle3_weights[1013]), .FEAT_THRES(feature_thresholds[1013]), .FEAT_ABOVE(feature_aboves[1013]), .FEAT_BELOW(feature_belows[1013])) ac1013(.scan_win(scan_win1013), .scan_win_std_dev(scan_win_std_dev[1013]), .feature_accum(feature_accums[1013]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1014]), .RECT1_Y(rectangle1_ys[1014]), .RECT1_WIDTH(rectangle1_widths[1014]), .RECT1_HEIGHT(rectangle1_heights[1014]), .RECT1_WEIGHT(rectangle1_weights[1014]), .RECT2_X(rectangle2_xs[1014]), .RECT2_Y(rectangle2_ys[1014]), .RECT2_WIDTH(rectangle2_widths[1014]), .RECT2_HEIGHT(rectangle2_heights[1014]), .RECT2_WEIGHT(rectangle2_weights[1014]), .RECT3_X(rectangle3_xs[1014]), .RECT3_Y(rectangle3_ys[1014]), .RECT3_WIDTH(rectangle3_widths[1014]), .RECT3_HEIGHT(rectangle3_heights[1014]), .RECT3_WEIGHT(rectangle3_weights[1014]), .FEAT_THRES(feature_thresholds[1014]), .FEAT_ABOVE(feature_aboves[1014]), .FEAT_BELOW(feature_belows[1014])) ac1014(.scan_win(scan_win1014), .scan_win_std_dev(scan_win_std_dev[1014]), .feature_accum(feature_accums[1014]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1015]), .RECT1_Y(rectangle1_ys[1015]), .RECT1_WIDTH(rectangle1_widths[1015]), .RECT1_HEIGHT(rectangle1_heights[1015]), .RECT1_WEIGHT(rectangle1_weights[1015]), .RECT2_X(rectangle2_xs[1015]), .RECT2_Y(rectangle2_ys[1015]), .RECT2_WIDTH(rectangle2_widths[1015]), .RECT2_HEIGHT(rectangle2_heights[1015]), .RECT2_WEIGHT(rectangle2_weights[1015]), .RECT3_X(rectangle3_xs[1015]), .RECT3_Y(rectangle3_ys[1015]), .RECT3_WIDTH(rectangle3_widths[1015]), .RECT3_HEIGHT(rectangle3_heights[1015]), .RECT3_WEIGHT(rectangle3_weights[1015]), .FEAT_THRES(feature_thresholds[1015]), .FEAT_ABOVE(feature_aboves[1015]), .FEAT_BELOW(feature_belows[1015])) ac1015(.scan_win(scan_win1015), .scan_win_std_dev(scan_win_std_dev[1015]), .feature_accum(feature_accums[1015]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1016]), .RECT1_Y(rectangle1_ys[1016]), .RECT1_WIDTH(rectangle1_widths[1016]), .RECT1_HEIGHT(rectangle1_heights[1016]), .RECT1_WEIGHT(rectangle1_weights[1016]), .RECT2_X(rectangle2_xs[1016]), .RECT2_Y(rectangle2_ys[1016]), .RECT2_WIDTH(rectangle2_widths[1016]), .RECT2_HEIGHT(rectangle2_heights[1016]), .RECT2_WEIGHT(rectangle2_weights[1016]), .RECT3_X(rectangle3_xs[1016]), .RECT3_Y(rectangle3_ys[1016]), .RECT3_WIDTH(rectangle3_widths[1016]), .RECT3_HEIGHT(rectangle3_heights[1016]), .RECT3_WEIGHT(rectangle3_weights[1016]), .FEAT_THRES(feature_thresholds[1016]), .FEAT_ABOVE(feature_aboves[1016]), .FEAT_BELOW(feature_belows[1016])) ac1016(.scan_win(scan_win1016), .scan_win_std_dev(scan_win_std_dev[1016]), .feature_accum(feature_accums[1016]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1017]), .RECT1_Y(rectangle1_ys[1017]), .RECT1_WIDTH(rectangle1_widths[1017]), .RECT1_HEIGHT(rectangle1_heights[1017]), .RECT1_WEIGHT(rectangle1_weights[1017]), .RECT2_X(rectangle2_xs[1017]), .RECT2_Y(rectangle2_ys[1017]), .RECT2_WIDTH(rectangle2_widths[1017]), .RECT2_HEIGHT(rectangle2_heights[1017]), .RECT2_WEIGHT(rectangle2_weights[1017]), .RECT3_X(rectangle3_xs[1017]), .RECT3_Y(rectangle3_ys[1017]), .RECT3_WIDTH(rectangle3_widths[1017]), .RECT3_HEIGHT(rectangle3_heights[1017]), .RECT3_WEIGHT(rectangle3_weights[1017]), .FEAT_THRES(feature_thresholds[1017]), .FEAT_ABOVE(feature_aboves[1017]), .FEAT_BELOW(feature_belows[1017])) ac1017(.scan_win(scan_win1017), .scan_win_std_dev(scan_win_std_dev[1017]), .feature_accum(feature_accums[1017]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1018]), .RECT1_Y(rectangle1_ys[1018]), .RECT1_WIDTH(rectangle1_widths[1018]), .RECT1_HEIGHT(rectangle1_heights[1018]), .RECT1_WEIGHT(rectangle1_weights[1018]), .RECT2_X(rectangle2_xs[1018]), .RECT2_Y(rectangle2_ys[1018]), .RECT2_WIDTH(rectangle2_widths[1018]), .RECT2_HEIGHT(rectangle2_heights[1018]), .RECT2_WEIGHT(rectangle2_weights[1018]), .RECT3_X(rectangle3_xs[1018]), .RECT3_Y(rectangle3_ys[1018]), .RECT3_WIDTH(rectangle3_widths[1018]), .RECT3_HEIGHT(rectangle3_heights[1018]), .RECT3_WEIGHT(rectangle3_weights[1018]), .FEAT_THRES(feature_thresholds[1018]), .FEAT_ABOVE(feature_aboves[1018]), .FEAT_BELOW(feature_belows[1018])) ac1018(.scan_win(scan_win1018), .scan_win_std_dev(scan_win_std_dev[1018]), .feature_accum(feature_accums[1018]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1019]), .RECT1_Y(rectangle1_ys[1019]), .RECT1_WIDTH(rectangle1_widths[1019]), .RECT1_HEIGHT(rectangle1_heights[1019]), .RECT1_WEIGHT(rectangle1_weights[1019]), .RECT2_X(rectangle2_xs[1019]), .RECT2_Y(rectangle2_ys[1019]), .RECT2_WIDTH(rectangle2_widths[1019]), .RECT2_HEIGHT(rectangle2_heights[1019]), .RECT2_WEIGHT(rectangle2_weights[1019]), .RECT3_X(rectangle3_xs[1019]), .RECT3_Y(rectangle3_ys[1019]), .RECT3_WIDTH(rectangle3_widths[1019]), .RECT3_HEIGHT(rectangle3_heights[1019]), .RECT3_WEIGHT(rectangle3_weights[1019]), .FEAT_THRES(feature_thresholds[1019]), .FEAT_ABOVE(feature_aboves[1019]), .FEAT_BELOW(feature_belows[1019])) ac1019(.scan_win(scan_win1019), .scan_win_std_dev(scan_win_std_dev[1019]), .feature_accum(feature_accums[1019]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1020]), .RECT1_Y(rectangle1_ys[1020]), .RECT1_WIDTH(rectangle1_widths[1020]), .RECT1_HEIGHT(rectangle1_heights[1020]), .RECT1_WEIGHT(rectangle1_weights[1020]), .RECT2_X(rectangle2_xs[1020]), .RECT2_Y(rectangle2_ys[1020]), .RECT2_WIDTH(rectangle2_widths[1020]), .RECT2_HEIGHT(rectangle2_heights[1020]), .RECT2_WEIGHT(rectangle2_weights[1020]), .RECT3_X(rectangle3_xs[1020]), .RECT3_Y(rectangle3_ys[1020]), .RECT3_WIDTH(rectangle3_widths[1020]), .RECT3_HEIGHT(rectangle3_heights[1020]), .RECT3_WEIGHT(rectangle3_weights[1020]), .FEAT_THRES(feature_thresholds[1020]), .FEAT_ABOVE(feature_aboves[1020]), .FEAT_BELOW(feature_belows[1020])) ac1020(.scan_win(scan_win1020), .scan_win_std_dev(scan_win_std_dev[1020]), .feature_accum(feature_accums[1020]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1021]), .RECT1_Y(rectangle1_ys[1021]), .RECT1_WIDTH(rectangle1_widths[1021]), .RECT1_HEIGHT(rectangle1_heights[1021]), .RECT1_WEIGHT(rectangle1_weights[1021]), .RECT2_X(rectangle2_xs[1021]), .RECT2_Y(rectangle2_ys[1021]), .RECT2_WIDTH(rectangle2_widths[1021]), .RECT2_HEIGHT(rectangle2_heights[1021]), .RECT2_WEIGHT(rectangle2_weights[1021]), .RECT3_X(rectangle3_xs[1021]), .RECT3_Y(rectangle3_ys[1021]), .RECT3_WIDTH(rectangle3_widths[1021]), .RECT3_HEIGHT(rectangle3_heights[1021]), .RECT3_WEIGHT(rectangle3_weights[1021]), .FEAT_THRES(feature_thresholds[1021]), .FEAT_ABOVE(feature_aboves[1021]), .FEAT_BELOW(feature_belows[1021])) ac1021(.scan_win(scan_win1021), .scan_win_std_dev(scan_win_std_dev[1021]), .feature_accum(feature_accums[1021]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1022]), .RECT1_Y(rectangle1_ys[1022]), .RECT1_WIDTH(rectangle1_widths[1022]), .RECT1_HEIGHT(rectangle1_heights[1022]), .RECT1_WEIGHT(rectangle1_weights[1022]), .RECT2_X(rectangle2_xs[1022]), .RECT2_Y(rectangle2_ys[1022]), .RECT2_WIDTH(rectangle2_widths[1022]), .RECT2_HEIGHT(rectangle2_heights[1022]), .RECT2_WEIGHT(rectangle2_weights[1022]), .RECT3_X(rectangle3_xs[1022]), .RECT3_Y(rectangle3_ys[1022]), .RECT3_WIDTH(rectangle3_widths[1022]), .RECT3_HEIGHT(rectangle3_heights[1022]), .RECT3_WEIGHT(rectangle3_weights[1022]), .FEAT_THRES(feature_thresholds[1022]), .FEAT_ABOVE(feature_aboves[1022]), .FEAT_BELOW(feature_belows[1022])) ac1022(.scan_win(scan_win1022), .scan_win_std_dev(scan_win_std_dev[1022]), .feature_accum(feature_accums[1022]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1023]), .RECT1_Y(rectangle1_ys[1023]), .RECT1_WIDTH(rectangle1_widths[1023]), .RECT1_HEIGHT(rectangle1_heights[1023]), .RECT1_WEIGHT(rectangle1_weights[1023]), .RECT2_X(rectangle2_xs[1023]), .RECT2_Y(rectangle2_ys[1023]), .RECT2_WIDTH(rectangle2_widths[1023]), .RECT2_HEIGHT(rectangle2_heights[1023]), .RECT2_WEIGHT(rectangle2_weights[1023]), .RECT3_X(rectangle3_xs[1023]), .RECT3_Y(rectangle3_ys[1023]), .RECT3_WIDTH(rectangle3_widths[1023]), .RECT3_HEIGHT(rectangle3_heights[1023]), .RECT3_WEIGHT(rectangle3_weights[1023]), .FEAT_THRES(feature_thresholds[1023]), .FEAT_ABOVE(feature_aboves[1023]), .FEAT_BELOW(feature_belows[1023])) ac1023(.scan_win(scan_win1023), .scan_win_std_dev(scan_win_std_dev[1023]), .feature_accum(feature_accums[1023]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1024]), .RECT1_Y(rectangle1_ys[1024]), .RECT1_WIDTH(rectangle1_widths[1024]), .RECT1_HEIGHT(rectangle1_heights[1024]), .RECT1_WEIGHT(rectangle1_weights[1024]), .RECT2_X(rectangle2_xs[1024]), .RECT2_Y(rectangle2_ys[1024]), .RECT2_WIDTH(rectangle2_widths[1024]), .RECT2_HEIGHT(rectangle2_heights[1024]), .RECT2_WEIGHT(rectangle2_weights[1024]), .RECT3_X(rectangle3_xs[1024]), .RECT3_Y(rectangle3_ys[1024]), .RECT3_WIDTH(rectangle3_widths[1024]), .RECT3_HEIGHT(rectangle3_heights[1024]), .RECT3_WEIGHT(rectangle3_weights[1024]), .FEAT_THRES(feature_thresholds[1024]), .FEAT_ABOVE(feature_aboves[1024]), .FEAT_BELOW(feature_belows[1024])) ac1024(.scan_win(scan_win1024), .scan_win_std_dev(scan_win_std_dev[1024]), .feature_accum(feature_accums[1024]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1025]), .RECT1_Y(rectangle1_ys[1025]), .RECT1_WIDTH(rectangle1_widths[1025]), .RECT1_HEIGHT(rectangle1_heights[1025]), .RECT1_WEIGHT(rectangle1_weights[1025]), .RECT2_X(rectangle2_xs[1025]), .RECT2_Y(rectangle2_ys[1025]), .RECT2_WIDTH(rectangle2_widths[1025]), .RECT2_HEIGHT(rectangle2_heights[1025]), .RECT2_WEIGHT(rectangle2_weights[1025]), .RECT3_X(rectangle3_xs[1025]), .RECT3_Y(rectangle3_ys[1025]), .RECT3_WIDTH(rectangle3_widths[1025]), .RECT3_HEIGHT(rectangle3_heights[1025]), .RECT3_WEIGHT(rectangle3_weights[1025]), .FEAT_THRES(feature_thresholds[1025]), .FEAT_ABOVE(feature_aboves[1025]), .FEAT_BELOW(feature_belows[1025])) ac1025(.scan_win(scan_win1025), .scan_win_std_dev(scan_win_std_dev[1025]), .feature_accum(feature_accums[1025]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1026]), .RECT1_Y(rectangle1_ys[1026]), .RECT1_WIDTH(rectangle1_widths[1026]), .RECT1_HEIGHT(rectangle1_heights[1026]), .RECT1_WEIGHT(rectangle1_weights[1026]), .RECT2_X(rectangle2_xs[1026]), .RECT2_Y(rectangle2_ys[1026]), .RECT2_WIDTH(rectangle2_widths[1026]), .RECT2_HEIGHT(rectangle2_heights[1026]), .RECT2_WEIGHT(rectangle2_weights[1026]), .RECT3_X(rectangle3_xs[1026]), .RECT3_Y(rectangle3_ys[1026]), .RECT3_WIDTH(rectangle3_widths[1026]), .RECT3_HEIGHT(rectangle3_heights[1026]), .RECT3_WEIGHT(rectangle3_weights[1026]), .FEAT_THRES(feature_thresholds[1026]), .FEAT_ABOVE(feature_aboves[1026]), .FEAT_BELOW(feature_belows[1026])) ac1026(.scan_win(scan_win1026), .scan_win_std_dev(scan_win_std_dev[1026]), .feature_accum(feature_accums[1026]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1027]), .RECT1_Y(rectangle1_ys[1027]), .RECT1_WIDTH(rectangle1_widths[1027]), .RECT1_HEIGHT(rectangle1_heights[1027]), .RECT1_WEIGHT(rectangle1_weights[1027]), .RECT2_X(rectangle2_xs[1027]), .RECT2_Y(rectangle2_ys[1027]), .RECT2_WIDTH(rectangle2_widths[1027]), .RECT2_HEIGHT(rectangle2_heights[1027]), .RECT2_WEIGHT(rectangle2_weights[1027]), .RECT3_X(rectangle3_xs[1027]), .RECT3_Y(rectangle3_ys[1027]), .RECT3_WIDTH(rectangle3_widths[1027]), .RECT3_HEIGHT(rectangle3_heights[1027]), .RECT3_WEIGHT(rectangle3_weights[1027]), .FEAT_THRES(feature_thresholds[1027]), .FEAT_ABOVE(feature_aboves[1027]), .FEAT_BELOW(feature_belows[1027])) ac1027(.scan_win(scan_win1027), .scan_win_std_dev(scan_win_std_dev[1027]), .feature_accum(feature_accums[1027]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1028]), .RECT1_Y(rectangle1_ys[1028]), .RECT1_WIDTH(rectangle1_widths[1028]), .RECT1_HEIGHT(rectangle1_heights[1028]), .RECT1_WEIGHT(rectangle1_weights[1028]), .RECT2_X(rectangle2_xs[1028]), .RECT2_Y(rectangle2_ys[1028]), .RECT2_WIDTH(rectangle2_widths[1028]), .RECT2_HEIGHT(rectangle2_heights[1028]), .RECT2_WEIGHT(rectangle2_weights[1028]), .RECT3_X(rectangle3_xs[1028]), .RECT3_Y(rectangle3_ys[1028]), .RECT3_WIDTH(rectangle3_widths[1028]), .RECT3_HEIGHT(rectangle3_heights[1028]), .RECT3_WEIGHT(rectangle3_weights[1028]), .FEAT_THRES(feature_thresholds[1028]), .FEAT_ABOVE(feature_aboves[1028]), .FEAT_BELOW(feature_belows[1028])) ac1028(.scan_win(scan_win1028), .scan_win_std_dev(scan_win_std_dev[1028]), .feature_accum(feature_accums[1028]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1029]), .RECT1_Y(rectangle1_ys[1029]), .RECT1_WIDTH(rectangle1_widths[1029]), .RECT1_HEIGHT(rectangle1_heights[1029]), .RECT1_WEIGHT(rectangle1_weights[1029]), .RECT2_X(rectangle2_xs[1029]), .RECT2_Y(rectangle2_ys[1029]), .RECT2_WIDTH(rectangle2_widths[1029]), .RECT2_HEIGHT(rectangle2_heights[1029]), .RECT2_WEIGHT(rectangle2_weights[1029]), .RECT3_X(rectangle3_xs[1029]), .RECT3_Y(rectangle3_ys[1029]), .RECT3_WIDTH(rectangle3_widths[1029]), .RECT3_HEIGHT(rectangle3_heights[1029]), .RECT3_WEIGHT(rectangle3_weights[1029]), .FEAT_THRES(feature_thresholds[1029]), .FEAT_ABOVE(feature_aboves[1029]), .FEAT_BELOW(feature_belows[1029])) ac1029(.scan_win(scan_win1029), .scan_win_std_dev(scan_win_std_dev[1029]), .feature_accum(feature_accums[1029]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1030]), .RECT1_Y(rectangle1_ys[1030]), .RECT1_WIDTH(rectangle1_widths[1030]), .RECT1_HEIGHT(rectangle1_heights[1030]), .RECT1_WEIGHT(rectangle1_weights[1030]), .RECT2_X(rectangle2_xs[1030]), .RECT2_Y(rectangle2_ys[1030]), .RECT2_WIDTH(rectangle2_widths[1030]), .RECT2_HEIGHT(rectangle2_heights[1030]), .RECT2_WEIGHT(rectangle2_weights[1030]), .RECT3_X(rectangle3_xs[1030]), .RECT3_Y(rectangle3_ys[1030]), .RECT3_WIDTH(rectangle3_widths[1030]), .RECT3_HEIGHT(rectangle3_heights[1030]), .RECT3_WEIGHT(rectangle3_weights[1030]), .FEAT_THRES(feature_thresholds[1030]), .FEAT_ABOVE(feature_aboves[1030]), .FEAT_BELOW(feature_belows[1030])) ac1030(.scan_win(scan_win1030), .scan_win_std_dev(scan_win_std_dev[1030]), .feature_accum(feature_accums[1030]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1031]), .RECT1_Y(rectangle1_ys[1031]), .RECT1_WIDTH(rectangle1_widths[1031]), .RECT1_HEIGHT(rectangle1_heights[1031]), .RECT1_WEIGHT(rectangle1_weights[1031]), .RECT2_X(rectangle2_xs[1031]), .RECT2_Y(rectangle2_ys[1031]), .RECT2_WIDTH(rectangle2_widths[1031]), .RECT2_HEIGHT(rectangle2_heights[1031]), .RECT2_WEIGHT(rectangle2_weights[1031]), .RECT3_X(rectangle3_xs[1031]), .RECT3_Y(rectangle3_ys[1031]), .RECT3_WIDTH(rectangle3_widths[1031]), .RECT3_HEIGHT(rectangle3_heights[1031]), .RECT3_WEIGHT(rectangle3_weights[1031]), .FEAT_THRES(feature_thresholds[1031]), .FEAT_ABOVE(feature_aboves[1031]), .FEAT_BELOW(feature_belows[1031])) ac1031(.scan_win(scan_win1031), .scan_win_std_dev(scan_win_std_dev[1031]), .feature_accum(feature_accums[1031]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1032]), .RECT1_Y(rectangle1_ys[1032]), .RECT1_WIDTH(rectangle1_widths[1032]), .RECT1_HEIGHT(rectangle1_heights[1032]), .RECT1_WEIGHT(rectangle1_weights[1032]), .RECT2_X(rectangle2_xs[1032]), .RECT2_Y(rectangle2_ys[1032]), .RECT2_WIDTH(rectangle2_widths[1032]), .RECT2_HEIGHT(rectangle2_heights[1032]), .RECT2_WEIGHT(rectangle2_weights[1032]), .RECT3_X(rectangle3_xs[1032]), .RECT3_Y(rectangle3_ys[1032]), .RECT3_WIDTH(rectangle3_widths[1032]), .RECT3_HEIGHT(rectangle3_heights[1032]), .RECT3_WEIGHT(rectangle3_weights[1032]), .FEAT_THRES(feature_thresholds[1032]), .FEAT_ABOVE(feature_aboves[1032]), .FEAT_BELOW(feature_belows[1032])) ac1032(.scan_win(scan_win1032), .scan_win_std_dev(scan_win_std_dev[1032]), .feature_accum(feature_accums[1032]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1033]), .RECT1_Y(rectangle1_ys[1033]), .RECT1_WIDTH(rectangle1_widths[1033]), .RECT1_HEIGHT(rectangle1_heights[1033]), .RECT1_WEIGHT(rectangle1_weights[1033]), .RECT2_X(rectangle2_xs[1033]), .RECT2_Y(rectangle2_ys[1033]), .RECT2_WIDTH(rectangle2_widths[1033]), .RECT2_HEIGHT(rectangle2_heights[1033]), .RECT2_WEIGHT(rectangle2_weights[1033]), .RECT3_X(rectangle3_xs[1033]), .RECT3_Y(rectangle3_ys[1033]), .RECT3_WIDTH(rectangle3_widths[1033]), .RECT3_HEIGHT(rectangle3_heights[1033]), .RECT3_WEIGHT(rectangle3_weights[1033]), .FEAT_THRES(feature_thresholds[1033]), .FEAT_ABOVE(feature_aboves[1033]), .FEAT_BELOW(feature_belows[1033])) ac1033(.scan_win(scan_win1033), .scan_win_std_dev(scan_win_std_dev[1033]), .feature_accum(feature_accums[1033]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1034]), .RECT1_Y(rectangle1_ys[1034]), .RECT1_WIDTH(rectangle1_widths[1034]), .RECT1_HEIGHT(rectangle1_heights[1034]), .RECT1_WEIGHT(rectangle1_weights[1034]), .RECT2_X(rectangle2_xs[1034]), .RECT2_Y(rectangle2_ys[1034]), .RECT2_WIDTH(rectangle2_widths[1034]), .RECT2_HEIGHT(rectangle2_heights[1034]), .RECT2_WEIGHT(rectangle2_weights[1034]), .RECT3_X(rectangle3_xs[1034]), .RECT3_Y(rectangle3_ys[1034]), .RECT3_WIDTH(rectangle3_widths[1034]), .RECT3_HEIGHT(rectangle3_heights[1034]), .RECT3_WEIGHT(rectangle3_weights[1034]), .FEAT_THRES(feature_thresholds[1034]), .FEAT_ABOVE(feature_aboves[1034]), .FEAT_BELOW(feature_belows[1034])) ac1034(.scan_win(scan_win1034), .scan_win_std_dev(scan_win_std_dev[1034]), .feature_accum(feature_accums[1034]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1035]), .RECT1_Y(rectangle1_ys[1035]), .RECT1_WIDTH(rectangle1_widths[1035]), .RECT1_HEIGHT(rectangle1_heights[1035]), .RECT1_WEIGHT(rectangle1_weights[1035]), .RECT2_X(rectangle2_xs[1035]), .RECT2_Y(rectangle2_ys[1035]), .RECT2_WIDTH(rectangle2_widths[1035]), .RECT2_HEIGHT(rectangle2_heights[1035]), .RECT2_WEIGHT(rectangle2_weights[1035]), .RECT3_X(rectangle3_xs[1035]), .RECT3_Y(rectangle3_ys[1035]), .RECT3_WIDTH(rectangle3_widths[1035]), .RECT3_HEIGHT(rectangle3_heights[1035]), .RECT3_WEIGHT(rectangle3_weights[1035]), .FEAT_THRES(feature_thresholds[1035]), .FEAT_ABOVE(feature_aboves[1035]), .FEAT_BELOW(feature_belows[1035])) ac1035(.scan_win(scan_win1035), .scan_win_std_dev(scan_win_std_dev[1035]), .feature_accum(feature_accums[1035]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1036]), .RECT1_Y(rectangle1_ys[1036]), .RECT1_WIDTH(rectangle1_widths[1036]), .RECT1_HEIGHT(rectangle1_heights[1036]), .RECT1_WEIGHT(rectangle1_weights[1036]), .RECT2_X(rectangle2_xs[1036]), .RECT2_Y(rectangle2_ys[1036]), .RECT2_WIDTH(rectangle2_widths[1036]), .RECT2_HEIGHT(rectangle2_heights[1036]), .RECT2_WEIGHT(rectangle2_weights[1036]), .RECT3_X(rectangle3_xs[1036]), .RECT3_Y(rectangle3_ys[1036]), .RECT3_WIDTH(rectangle3_widths[1036]), .RECT3_HEIGHT(rectangle3_heights[1036]), .RECT3_WEIGHT(rectangle3_weights[1036]), .FEAT_THRES(feature_thresholds[1036]), .FEAT_ABOVE(feature_aboves[1036]), .FEAT_BELOW(feature_belows[1036])) ac1036(.scan_win(scan_win1036), .scan_win_std_dev(scan_win_std_dev[1036]), .feature_accum(feature_accums[1036]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1037]), .RECT1_Y(rectangle1_ys[1037]), .RECT1_WIDTH(rectangle1_widths[1037]), .RECT1_HEIGHT(rectangle1_heights[1037]), .RECT1_WEIGHT(rectangle1_weights[1037]), .RECT2_X(rectangle2_xs[1037]), .RECT2_Y(rectangle2_ys[1037]), .RECT2_WIDTH(rectangle2_widths[1037]), .RECT2_HEIGHT(rectangle2_heights[1037]), .RECT2_WEIGHT(rectangle2_weights[1037]), .RECT3_X(rectangle3_xs[1037]), .RECT3_Y(rectangle3_ys[1037]), .RECT3_WIDTH(rectangle3_widths[1037]), .RECT3_HEIGHT(rectangle3_heights[1037]), .RECT3_WEIGHT(rectangle3_weights[1037]), .FEAT_THRES(feature_thresholds[1037]), .FEAT_ABOVE(feature_aboves[1037]), .FEAT_BELOW(feature_belows[1037])) ac1037(.scan_win(scan_win1037), .scan_win_std_dev(scan_win_std_dev[1037]), .feature_accum(feature_accums[1037]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1038]), .RECT1_Y(rectangle1_ys[1038]), .RECT1_WIDTH(rectangle1_widths[1038]), .RECT1_HEIGHT(rectangle1_heights[1038]), .RECT1_WEIGHT(rectangle1_weights[1038]), .RECT2_X(rectangle2_xs[1038]), .RECT2_Y(rectangle2_ys[1038]), .RECT2_WIDTH(rectangle2_widths[1038]), .RECT2_HEIGHT(rectangle2_heights[1038]), .RECT2_WEIGHT(rectangle2_weights[1038]), .RECT3_X(rectangle3_xs[1038]), .RECT3_Y(rectangle3_ys[1038]), .RECT3_WIDTH(rectangle3_widths[1038]), .RECT3_HEIGHT(rectangle3_heights[1038]), .RECT3_WEIGHT(rectangle3_weights[1038]), .FEAT_THRES(feature_thresholds[1038]), .FEAT_ABOVE(feature_aboves[1038]), .FEAT_BELOW(feature_belows[1038])) ac1038(.scan_win(scan_win1038), .scan_win_std_dev(scan_win_std_dev[1038]), .feature_accum(feature_accums[1038]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1039]), .RECT1_Y(rectangle1_ys[1039]), .RECT1_WIDTH(rectangle1_widths[1039]), .RECT1_HEIGHT(rectangle1_heights[1039]), .RECT1_WEIGHT(rectangle1_weights[1039]), .RECT2_X(rectangle2_xs[1039]), .RECT2_Y(rectangle2_ys[1039]), .RECT2_WIDTH(rectangle2_widths[1039]), .RECT2_HEIGHT(rectangle2_heights[1039]), .RECT2_WEIGHT(rectangle2_weights[1039]), .RECT3_X(rectangle3_xs[1039]), .RECT3_Y(rectangle3_ys[1039]), .RECT3_WIDTH(rectangle3_widths[1039]), .RECT3_HEIGHT(rectangle3_heights[1039]), .RECT3_WEIGHT(rectangle3_weights[1039]), .FEAT_THRES(feature_thresholds[1039]), .FEAT_ABOVE(feature_aboves[1039]), .FEAT_BELOW(feature_belows[1039])) ac1039(.scan_win(scan_win1039), .scan_win_std_dev(scan_win_std_dev[1039]), .feature_accum(feature_accums[1039]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1040]), .RECT1_Y(rectangle1_ys[1040]), .RECT1_WIDTH(rectangle1_widths[1040]), .RECT1_HEIGHT(rectangle1_heights[1040]), .RECT1_WEIGHT(rectangle1_weights[1040]), .RECT2_X(rectangle2_xs[1040]), .RECT2_Y(rectangle2_ys[1040]), .RECT2_WIDTH(rectangle2_widths[1040]), .RECT2_HEIGHT(rectangle2_heights[1040]), .RECT2_WEIGHT(rectangle2_weights[1040]), .RECT3_X(rectangle3_xs[1040]), .RECT3_Y(rectangle3_ys[1040]), .RECT3_WIDTH(rectangle3_widths[1040]), .RECT3_HEIGHT(rectangle3_heights[1040]), .RECT3_WEIGHT(rectangle3_weights[1040]), .FEAT_THRES(feature_thresholds[1040]), .FEAT_ABOVE(feature_aboves[1040]), .FEAT_BELOW(feature_belows[1040])) ac1040(.scan_win(scan_win1040), .scan_win_std_dev(scan_win_std_dev[1040]), .feature_accum(feature_accums[1040]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1041]), .RECT1_Y(rectangle1_ys[1041]), .RECT1_WIDTH(rectangle1_widths[1041]), .RECT1_HEIGHT(rectangle1_heights[1041]), .RECT1_WEIGHT(rectangle1_weights[1041]), .RECT2_X(rectangle2_xs[1041]), .RECT2_Y(rectangle2_ys[1041]), .RECT2_WIDTH(rectangle2_widths[1041]), .RECT2_HEIGHT(rectangle2_heights[1041]), .RECT2_WEIGHT(rectangle2_weights[1041]), .RECT3_X(rectangle3_xs[1041]), .RECT3_Y(rectangle3_ys[1041]), .RECT3_WIDTH(rectangle3_widths[1041]), .RECT3_HEIGHT(rectangle3_heights[1041]), .RECT3_WEIGHT(rectangle3_weights[1041]), .FEAT_THRES(feature_thresholds[1041]), .FEAT_ABOVE(feature_aboves[1041]), .FEAT_BELOW(feature_belows[1041])) ac1041(.scan_win(scan_win1041), .scan_win_std_dev(scan_win_std_dev[1041]), .feature_accum(feature_accums[1041]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1042]), .RECT1_Y(rectangle1_ys[1042]), .RECT1_WIDTH(rectangle1_widths[1042]), .RECT1_HEIGHT(rectangle1_heights[1042]), .RECT1_WEIGHT(rectangle1_weights[1042]), .RECT2_X(rectangle2_xs[1042]), .RECT2_Y(rectangle2_ys[1042]), .RECT2_WIDTH(rectangle2_widths[1042]), .RECT2_HEIGHT(rectangle2_heights[1042]), .RECT2_WEIGHT(rectangle2_weights[1042]), .RECT3_X(rectangle3_xs[1042]), .RECT3_Y(rectangle3_ys[1042]), .RECT3_WIDTH(rectangle3_widths[1042]), .RECT3_HEIGHT(rectangle3_heights[1042]), .RECT3_WEIGHT(rectangle3_weights[1042]), .FEAT_THRES(feature_thresholds[1042]), .FEAT_ABOVE(feature_aboves[1042]), .FEAT_BELOW(feature_belows[1042])) ac1042(.scan_win(scan_win1042), .scan_win_std_dev(scan_win_std_dev[1042]), .feature_accum(feature_accums[1042]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1043]), .RECT1_Y(rectangle1_ys[1043]), .RECT1_WIDTH(rectangle1_widths[1043]), .RECT1_HEIGHT(rectangle1_heights[1043]), .RECT1_WEIGHT(rectangle1_weights[1043]), .RECT2_X(rectangle2_xs[1043]), .RECT2_Y(rectangle2_ys[1043]), .RECT2_WIDTH(rectangle2_widths[1043]), .RECT2_HEIGHT(rectangle2_heights[1043]), .RECT2_WEIGHT(rectangle2_weights[1043]), .RECT3_X(rectangle3_xs[1043]), .RECT3_Y(rectangle3_ys[1043]), .RECT3_WIDTH(rectangle3_widths[1043]), .RECT3_HEIGHT(rectangle3_heights[1043]), .RECT3_WEIGHT(rectangle3_weights[1043]), .FEAT_THRES(feature_thresholds[1043]), .FEAT_ABOVE(feature_aboves[1043]), .FEAT_BELOW(feature_belows[1043])) ac1043(.scan_win(scan_win1043), .scan_win_std_dev(scan_win_std_dev[1043]), .feature_accum(feature_accums[1043]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1044]), .RECT1_Y(rectangle1_ys[1044]), .RECT1_WIDTH(rectangle1_widths[1044]), .RECT1_HEIGHT(rectangle1_heights[1044]), .RECT1_WEIGHT(rectangle1_weights[1044]), .RECT2_X(rectangle2_xs[1044]), .RECT2_Y(rectangle2_ys[1044]), .RECT2_WIDTH(rectangle2_widths[1044]), .RECT2_HEIGHT(rectangle2_heights[1044]), .RECT2_WEIGHT(rectangle2_weights[1044]), .RECT3_X(rectangle3_xs[1044]), .RECT3_Y(rectangle3_ys[1044]), .RECT3_WIDTH(rectangle3_widths[1044]), .RECT3_HEIGHT(rectangle3_heights[1044]), .RECT3_WEIGHT(rectangle3_weights[1044]), .FEAT_THRES(feature_thresholds[1044]), .FEAT_ABOVE(feature_aboves[1044]), .FEAT_BELOW(feature_belows[1044])) ac1044(.scan_win(scan_win1044), .scan_win_std_dev(scan_win_std_dev[1044]), .feature_accum(feature_accums[1044]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1045]), .RECT1_Y(rectangle1_ys[1045]), .RECT1_WIDTH(rectangle1_widths[1045]), .RECT1_HEIGHT(rectangle1_heights[1045]), .RECT1_WEIGHT(rectangle1_weights[1045]), .RECT2_X(rectangle2_xs[1045]), .RECT2_Y(rectangle2_ys[1045]), .RECT2_WIDTH(rectangle2_widths[1045]), .RECT2_HEIGHT(rectangle2_heights[1045]), .RECT2_WEIGHT(rectangle2_weights[1045]), .RECT3_X(rectangle3_xs[1045]), .RECT3_Y(rectangle3_ys[1045]), .RECT3_WIDTH(rectangle3_widths[1045]), .RECT3_HEIGHT(rectangle3_heights[1045]), .RECT3_WEIGHT(rectangle3_weights[1045]), .FEAT_THRES(feature_thresholds[1045]), .FEAT_ABOVE(feature_aboves[1045]), .FEAT_BELOW(feature_belows[1045])) ac1045(.scan_win(scan_win1045), .scan_win_std_dev(scan_win_std_dev[1045]), .feature_accum(feature_accums[1045]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1046]), .RECT1_Y(rectangle1_ys[1046]), .RECT1_WIDTH(rectangle1_widths[1046]), .RECT1_HEIGHT(rectangle1_heights[1046]), .RECT1_WEIGHT(rectangle1_weights[1046]), .RECT2_X(rectangle2_xs[1046]), .RECT2_Y(rectangle2_ys[1046]), .RECT2_WIDTH(rectangle2_widths[1046]), .RECT2_HEIGHT(rectangle2_heights[1046]), .RECT2_WEIGHT(rectangle2_weights[1046]), .RECT3_X(rectangle3_xs[1046]), .RECT3_Y(rectangle3_ys[1046]), .RECT3_WIDTH(rectangle3_widths[1046]), .RECT3_HEIGHT(rectangle3_heights[1046]), .RECT3_WEIGHT(rectangle3_weights[1046]), .FEAT_THRES(feature_thresholds[1046]), .FEAT_ABOVE(feature_aboves[1046]), .FEAT_BELOW(feature_belows[1046])) ac1046(.scan_win(scan_win1046), .scan_win_std_dev(scan_win_std_dev[1046]), .feature_accum(feature_accums[1046]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1047]), .RECT1_Y(rectangle1_ys[1047]), .RECT1_WIDTH(rectangle1_widths[1047]), .RECT1_HEIGHT(rectangle1_heights[1047]), .RECT1_WEIGHT(rectangle1_weights[1047]), .RECT2_X(rectangle2_xs[1047]), .RECT2_Y(rectangle2_ys[1047]), .RECT2_WIDTH(rectangle2_widths[1047]), .RECT2_HEIGHT(rectangle2_heights[1047]), .RECT2_WEIGHT(rectangle2_weights[1047]), .RECT3_X(rectangle3_xs[1047]), .RECT3_Y(rectangle3_ys[1047]), .RECT3_WIDTH(rectangle3_widths[1047]), .RECT3_HEIGHT(rectangle3_heights[1047]), .RECT3_WEIGHT(rectangle3_weights[1047]), .FEAT_THRES(feature_thresholds[1047]), .FEAT_ABOVE(feature_aboves[1047]), .FEAT_BELOW(feature_belows[1047])) ac1047(.scan_win(scan_win1047), .scan_win_std_dev(scan_win_std_dev[1047]), .feature_accum(feature_accums[1047]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1048]), .RECT1_Y(rectangle1_ys[1048]), .RECT1_WIDTH(rectangle1_widths[1048]), .RECT1_HEIGHT(rectangle1_heights[1048]), .RECT1_WEIGHT(rectangle1_weights[1048]), .RECT2_X(rectangle2_xs[1048]), .RECT2_Y(rectangle2_ys[1048]), .RECT2_WIDTH(rectangle2_widths[1048]), .RECT2_HEIGHT(rectangle2_heights[1048]), .RECT2_WEIGHT(rectangle2_weights[1048]), .RECT3_X(rectangle3_xs[1048]), .RECT3_Y(rectangle3_ys[1048]), .RECT3_WIDTH(rectangle3_widths[1048]), .RECT3_HEIGHT(rectangle3_heights[1048]), .RECT3_WEIGHT(rectangle3_weights[1048]), .FEAT_THRES(feature_thresholds[1048]), .FEAT_ABOVE(feature_aboves[1048]), .FEAT_BELOW(feature_belows[1048])) ac1048(.scan_win(scan_win1048), .scan_win_std_dev(scan_win_std_dev[1048]), .feature_accum(feature_accums[1048]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1049]), .RECT1_Y(rectangle1_ys[1049]), .RECT1_WIDTH(rectangle1_widths[1049]), .RECT1_HEIGHT(rectangle1_heights[1049]), .RECT1_WEIGHT(rectangle1_weights[1049]), .RECT2_X(rectangle2_xs[1049]), .RECT2_Y(rectangle2_ys[1049]), .RECT2_WIDTH(rectangle2_widths[1049]), .RECT2_HEIGHT(rectangle2_heights[1049]), .RECT2_WEIGHT(rectangle2_weights[1049]), .RECT3_X(rectangle3_xs[1049]), .RECT3_Y(rectangle3_ys[1049]), .RECT3_WIDTH(rectangle3_widths[1049]), .RECT3_HEIGHT(rectangle3_heights[1049]), .RECT3_WEIGHT(rectangle3_weights[1049]), .FEAT_THRES(feature_thresholds[1049]), .FEAT_ABOVE(feature_aboves[1049]), .FEAT_BELOW(feature_belows[1049])) ac1049(.scan_win(scan_win1049), .scan_win_std_dev(scan_win_std_dev[1049]), .feature_accum(feature_accums[1049]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1050]), .RECT1_Y(rectangle1_ys[1050]), .RECT1_WIDTH(rectangle1_widths[1050]), .RECT1_HEIGHT(rectangle1_heights[1050]), .RECT1_WEIGHT(rectangle1_weights[1050]), .RECT2_X(rectangle2_xs[1050]), .RECT2_Y(rectangle2_ys[1050]), .RECT2_WIDTH(rectangle2_widths[1050]), .RECT2_HEIGHT(rectangle2_heights[1050]), .RECT2_WEIGHT(rectangle2_weights[1050]), .RECT3_X(rectangle3_xs[1050]), .RECT3_Y(rectangle3_ys[1050]), .RECT3_WIDTH(rectangle3_widths[1050]), .RECT3_HEIGHT(rectangle3_heights[1050]), .RECT3_WEIGHT(rectangle3_weights[1050]), .FEAT_THRES(feature_thresholds[1050]), .FEAT_ABOVE(feature_aboves[1050]), .FEAT_BELOW(feature_belows[1050])) ac1050(.scan_win(scan_win1050), .scan_win_std_dev(scan_win_std_dev[1050]), .feature_accum(feature_accums[1050]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1051]), .RECT1_Y(rectangle1_ys[1051]), .RECT1_WIDTH(rectangle1_widths[1051]), .RECT1_HEIGHT(rectangle1_heights[1051]), .RECT1_WEIGHT(rectangle1_weights[1051]), .RECT2_X(rectangle2_xs[1051]), .RECT2_Y(rectangle2_ys[1051]), .RECT2_WIDTH(rectangle2_widths[1051]), .RECT2_HEIGHT(rectangle2_heights[1051]), .RECT2_WEIGHT(rectangle2_weights[1051]), .RECT3_X(rectangle3_xs[1051]), .RECT3_Y(rectangle3_ys[1051]), .RECT3_WIDTH(rectangle3_widths[1051]), .RECT3_HEIGHT(rectangle3_heights[1051]), .RECT3_WEIGHT(rectangle3_weights[1051]), .FEAT_THRES(feature_thresholds[1051]), .FEAT_ABOVE(feature_aboves[1051]), .FEAT_BELOW(feature_belows[1051])) ac1051(.scan_win(scan_win1051), .scan_win_std_dev(scan_win_std_dev[1051]), .feature_accum(feature_accums[1051]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1052]), .RECT1_Y(rectangle1_ys[1052]), .RECT1_WIDTH(rectangle1_widths[1052]), .RECT1_HEIGHT(rectangle1_heights[1052]), .RECT1_WEIGHT(rectangle1_weights[1052]), .RECT2_X(rectangle2_xs[1052]), .RECT2_Y(rectangle2_ys[1052]), .RECT2_WIDTH(rectangle2_widths[1052]), .RECT2_HEIGHT(rectangle2_heights[1052]), .RECT2_WEIGHT(rectangle2_weights[1052]), .RECT3_X(rectangle3_xs[1052]), .RECT3_Y(rectangle3_ys[1052]), .RECT3_WIDTH(rectangle3_widths[1052]), .RECT3_HEIGHT(rectangle3_heights[1052]), .RECT3_WEIGHT(rectangle3_weights[1052]), .FEAT_THRES(feature_thresholds[1052]), .FEAT_ABOVE(feature_aboves[1052]), .FEAT_BELOW(feature_belows[1052])) ac1052(.scan_win(scan_win1052), .scan_win_std_dev(scan_win_std_dev[1052]), .feature_accum(feature_accums[1052]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1053]), .RECT1_Y(rectangle1_ys[1053]), .RECT1_WIDTH(rectangle1_widths[1053]), .RECT1_HEIGHT(rectangle1_heights[1053]), .RECT1_WEIGHT(rectangle1_weights[1053]), .RECT2_X(rectangle2_xs[1053]), .RECT2_Y(rectangle2_ys[1053]), .RECT2_WIDTH(rectangle2_widths[1053]), .RECT2_HEIGHT(rectangle2_heights[1053]), .RECT2_WEIGHT(rectangle2_weights[1053]), .RECT3_X(rectangle3_xs[1053]), .RECT3_Y(rectangle3_ys[1053]), .RECT3_WIDTH(rectangle3_widths[1053]), .RECT3_HEIGHT(rectangle3_heights[1053]), .RECT3_WEIGHT(rectangle3_weights[1053]), .FEAT_THRES(feature_thresholds[1053]), .FEAT_ABOVE(feature_aboves[1053]), .FEAT_BELOW(feature_belows[1053])) ac1053(.scan_win(scan_win1053), .scan_win_std_dev(scan_win_std_dev[1053]), .feature_accum(feature_accums[1053]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1054]), .RECT1_Y(rectangle1_ys[1054]), .RECT1_WIDTH(rectangle1_widths[1054]), .RECT1_HEIGHT(rectangle1_heights[1054]), .RECT1_WEIGHT(rectangle1_weights[1054]), .RECT2_X(rectangle2_xs[1054]), .RECT2_Y(rectangle2_ys[1054]), .RECT2_WIDTH(rectangle2_widths[1054]), .RECT2_HEIGHT(rectangle2_heights[1054]), .RECT2_WEIGHT(rectangle2_weights[1054]), .RECT3_X(rectangle3_xs[1054]), .RECT3_Y(rectangle3_ys[1054]), .RECT3_WIDTH(rectangle3_widths[1054]), .RECT3_HEIGHT(rectangle3_heights[1054]), .RECT3_WEIGHT(rectangle3_weights[1054]), .FEAT_THRES(feature_thresholds[1054]), .FEAT_ABOVE(feature_aboves[1054]), .FEAT_BELOW(feature_belows[1054])) ac1054(.scan_win(scan_win1054), .scan_win_std_dev(scan_win_std_dev[1054]), .feature_accum(feature_accums[1054]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1055]), .RECT1_Y(rectangle1_ys[1055]), .RECT1_WIDTH(rectangle1_widths[1055]), .RECT1_HEIGHT(rectangle1_heights[1055]), .RECT1_WEIGHT(rectangle1_weights[1055]), .RECT2_X(rectangle2_xs[1055]), .RECT2_Y(rectangle2_ys[1055]), .RECT2_WIDTH(rectangle2_widths[1055]), .RECT2_HEIGHT(rectangle2_heights[1055]), .RECT2_WEIGHT(rectangle2_weights[1055]), .RECT3_X(rectangle3_xs[1055]), .RECT3_Y(rectangle3_ys[1055]), .RECT3_WIDTH(rectangle3_widths[1055]), .RECT3_HEIGHT(rectangle3_heights[1055]), .RECT3_WEIGHT(rectangle3_weights[1055]), .FEAT_THRES(feature_thresholds[1055]), .FEAT_ABOVE(feature_aboves[1055]), .FEAT_BELOW(feature_belows[1055])) ac1055(.scan_win(scan_win1055), .scan_win_std_dev(scan_win_std_dev[1055]), .feature_accum(feature_accums[1055]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1056]), .RECT1_Y(rectangle1_ys[1056]), .RECT1_WIDTH(rectangle1_widths[1056]), .RECT1_HEIGHT(rectangle1_heights[1056]), .RECT1_WEIGHT(rectangle1_weights[1056]), .RECT2_X(rectangle2_xs[1056]), .RECT2_Y(rectangle2_ys[1056]), .RECT2_WIDTH(rectangle2_widths[1056]), .RECT2_HEIGHT(rectangle2_heights[1056]), .RECT2_WEIGHT(rectangle2_weights[1056]), .RECT3_X(rectangle3_xs[1056]), .RECT3_Y(rectangle3_ys[1056]), .RECT3_WIDTH(rectangle3_widths[1056]), .RECT3_HEIGHT(rectangle3_heights[1056]), .RECT3_WEIGHT(rectangle3_weights[1056]), .FEAT_THRES(feature_thresholds[1056]), .FEAT_ABOVE(feature_aboves[1056]), .FEAT_BELOW(feature_belows[1056])) ac1056(.scan_win(scan_win1056), .scan_win_std_dev(scan_win_std_dev[1056]), .feature_accum(feature_accums[1056]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1057]), .RECT1_Y(rectangle1_ys[1057]), .RECT1_WIDTH(rectangle1_widths[1057]), .RECT1_HEIGHT(rectangle1_heights[1057]), .RECT1_WEIGHT(rectangle1_weights[1057]), .RECT2_X(rectangle2_xs[1057]), .RECT2_Y(rectangle2_ys[1057]), .RECT2_WIDTH(rectangle2_widths[1057]), .RECT2_HEIGHT(rectangle2_heights[1057]), .RECT2_WEIGHT(rectangle2_weights[1057]), .RECT3_X(rectangle3_xs[1057]), .RECT3_Y(rectangle3_ys[1057]), .RECT3_WIDTH(rectangle3_widths[1057]), .RECT3_HEIGHT(rectangle3_heights[1057]), .RECT3_WEIGHT(rectangle3_weights[1057]), .FEAT_THRES(feature_thresholds[1057]), .FEAT_ABOVE(feature_aboves[1057]), .FEAT_BELOW(feature_belows[1057])) ac1057(.scan_win(scan_win1057), .scan_win_std_dev(scan_win_std_dev[1057]), .feature_accum(feature_accums[1057]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1058]), .RECT1_Y(rectangle1_ys[1058]), .RECT1_WIDTH(rectangle1_widths[1058]), .RECT1_HEIGHT(rectangle1_heights[1058]), .RECT1_WEIGHT(rectangle1_weights[1058]), .RECT2_X(rectangle2_xs[1058]), .RECT2_Y(rectangle2_ys[1058]), .RECT2_WIDTH(rectangle2_widths[1058]), .RECT2_HEIGHT(rectangle2_heights[1058]), .RECT2_WEIGHT(rectangle2_weights[1058]), .RECT3_X(rectangle3_xs[1058]), .RECT3_Y(rectangle3_ys[1058]), .RECT3_WIDTH(rectangle3_widths[1058]), .RECT3_HEIGHT(rectangle3_heights[1058]), .RECT3_WEIGHT(rectangle3_weights[1058]), .FEAT_THRES(feature_thresholds[1058]), .FEAT_ABOVE(feature_aboves[1058]), .FEAT_BELOW(feature_belows[1058])) ac1058(.scan_win(scan_win1058), .scan_win_std_dev(scan_win_std_dev[1058]), .feature_accum(feature_accums[1058]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1059]), .RECT1_Y(rectangle1_ys[1059]), .RECT1_WIDTH(rectangle1_widths[1059]), .RECT1_HEIGHT(rectangle1_heights[1059]), .RECT1_WEIGHT(rectangle1_weights[1059]), .RECT2_X(rectangle2_xs[1059]), .RECT2_Y(rectangle2_ys[1059]), .RECT2_WIDTH(rectangle2_widths[1059]), .RECT2_HEIGHT(rectangle2_heights[1059]), .RECT2_WEIGHT(rectangle2_weights[1059]), .RECT3_X(rectangle3_xs[1059]), .RECT3_Y(rectangle3_ys[1059]), .RECT3_WIDTH(rectangle3_widths[1059]), .RECT3_HEIGHT(rectangle3_heights[1059]), .RECT3_WEIGHT(rectangle3_weights[1059]), .FEAT_THRES(feature_thresholds[1059]), .FEAT_ABOVE(feature_aboves[1059]), .FEAT_BELOW(feature_belows[1059])) ac1059(.scan_win(scan_win1059), .scan_win_std_dev(scan_win_std_dev[1059]), .feature_accum(feature_accums[1059]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1060]), .RECT1_Y(rectangle1_ys[1060]), .RECT1_WIDTH(rectangle1_widths[1060]), .RECT1_HEIGHT(rectangle1_heights[1060]), .RECT1_WEIGHT(rectangle1_weights[1060]), .RECT2_X(rectangle2_xs[1060]), .RECT2_Y(rectangle2_ys[1060]), .RECT2_WIDTH(rectangle2_widths[1060]), .RECT2_HEIGHT(rectangle2_heights[1060]), .RECT2_WEIGHT(rectangle2_weights[1060]), .RECT3_X(rectangle3_xs[1060]), .RECT3_Y(rectangle3_ys[1060]), .RECT3_WIDTH(rectangle3_widths[1060]), .RECT3_HEIGHT(rectangle3_heights[1060]), .RECT3_WEIGHT(rectangle3_weights[1060]), .FEAT_THRES(feature_thresholds[1060]), .FEAT_ABOVE(feature_aboves[1060]), .FEAT_BELOW(feature_belows[1060])) ac1060(.scan_win(scan_win1060), .scan_win_std_dev(scan_win_std_dev[1060]), .feature_accum(feature_accums[1060]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1061]), .RECT1_Y(rectangle1_ys[1061]), .RECT1_WIDTH(rectangle1_widths[1061]), .RECT1_HEIGHT(rectangle1_heights[1061]), .RECT1_WEIGHT(rectangle1_weights[1061]), .RECT2_X(rectangle2_xs[1061]), .RECT2_Y(rectangle2_ys[1061]), .RECT2_WIDTH(rectangle2_widths[1061]), .RECT2_HEIGHT(rectangle2_heights[1061]), .RECT2_WEIGHT(rectangle2_weights[1061]), .RECT3_X(rectangle3_xs[1061]), .RECT3_Y(rectangle3_ys[1061]), .RECT3_WIDTH(rectangle3_widths[1061]), .RECT3_HEIGHT(rectangle3_heights[1061]), .RECT3_WEIGHT(rectangle3_weights[1061]), .FEAT_THRES(feature_thresholds[1061]), .FEAT_ABOVE(feature_aboves[1061]), .FEAT_BELOW(feature_belows[1061])) ac1061(.scan_win(scan_win1061), .scan_win_std_dev(scan_win_std_dev[1061]), .feature_accum(feature_accums[1061]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1062]), .RECT1_Y(rectangle1_ys[1062]), .RECT1_WIDTH(rectangle1_widths[1062]), .RECT1_HEIGHT(rectangle1_heights[1062]), .RECT1_WEIGHT(rectangle1_weights[1062]), .RECT2_X(rectangle2_xs[1062]), .RECT2_Y(rectangle2_ys[1062]), .RECT2_WIDTH(rectangle2_widths[1062]), .RECT2_HEIGHT(rectangle2_heights[1062]), .RECT2_WEIGHT(rectangle2_weights[1062]), .RECT3_X(rectangle3_xs[1062]), .RECT3_Y(rectangle3_ys[1062]), .RECT3_WIDTH(rectangle3_widths[1062]), .RECT3_HEIGHT(rectangle3_heights[1062]), .RECT3_WEIGHT(rectangle3_weights[1062]), .FEAT_THRES(feature_thresholds[1062]), .FEAT_ABOVE(feature_aboves[1062]), .FEAT_BELOW(feature_belows[1062])) ac1062(.scan_win(scan_win1062), .scan_win_std_dev(scan_win_std_dev[1062]), .feature_accum(feature_accums[1062]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1063]), .RECT1_Y(rectangle1_ys[1063]), .RECT1_WIDTH(rectangle1_widths[1063]), .RECT1_HEIGHT(rectangle1_heights[1063]), .RECT1_WEIGHT(rectangle1_weights[1063]), .RECT2_X(rectangle2_xs[1063]), .RECT2_Y(rectangle2_ys[1063]), .RECT2_WIDTH(rectangle2_widths[1063]), .RECT2_HEIGHT(rectangle2_heights[1063]), .RECT2_WEIGHT(rectangle2_weights[1063]), .RECT3_X(rectangle3_xs[1063]), .RECT3_Y(rectangle3_ys[1063]), .RECT3_WIDTH(rectangle3_widths[1063]), .RECT3_HEIGHT(rectangle3_heights[1063]), .RECT3_WEIGHT(rectangle3_weights[1063]), .FEAT_THRES(feature_thresholds[1063]), .FEAT_ABOVE(feature_aboves[1063]), .FEAT_BELOW(feature_belows[1063])) ac1063(.scan_win(scan_win1063), .scan_win_std_dev(scan_win_std_dev[1063]), .feature_accum(feature_accums[1063]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1064]), .RECT1_Y(rectangle1_ys[1064]), .RECT1_WIDTH(rectangle1_widths[1064]), .RECT1_HEIGHT(rectangle1_heights[1064]), .RECT1_WEIGHT(rectangle1_weights[1064]), .RECT2_X(rectangle2_xs[1064]), .RECT2_Y(rectangle2_ys[1064]), .RECT2_WIDTH(rectangle2_widths[1064]), .RECT2_HEIGHT(rectangle2_heights[1064]), .RECT2_WEIGHT(rectangle2_weights[1064]), .RECT3_X(rectangle3_xs[1064]), .RECT3_Y(rectangle3_ys[1064]), .RECT3_WIDTH(rectangle3_widths[1064]), .RECT3_HEIGHT(rectangle3_heights[1064]), .RECT3_WEIGHT(rectangle3_weights[1064]), .FEAT_THRES(feature_thresholds[1064]), .FEAT_ABOVE(feature_aboves[1064]), .FEAT_BELOW(feature_belows[1064])) ac1064(.scan_win(scan_win1064), .scan_win_std_dev(scan_win_std_dev[1064]), .feature_accum(feature_accums[1064]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1065]), .RECT1_Y(rectangle1_ys[1065]), .RECT1_WIDTH(rectangle1_widths[1065]), .RECT1_HEIGHT(rectangle1_heights[1065]), .RECT1_WEIGHT(rectangle1_weights[1065]), .RECT2_X(rectangle2_xs[1065]), .RECT2_Y(rectangle2_ys[1065]), .RECT2_WIDTH(rectangle2_widths[1065]), .RECT2_HEIGHT(rectangle2_heights[1065]), .RECT2_WEIGHT(rectangle2_weights[1065]), .RECT3_X(rectangle3_xs[1065]), .RECT3_Y(rectangle3_ys[1065]), .RECT3_WIDTH(rectangle3_widths[1065]), .RECT3_HEIGHT(rectangle3_heights[1065]), .RECT3_WEIGHT(rectangle3_weights[1065]), .FEAT_THRES(feature_thresholds[1065]), .FEAT_ABOVE(feature_aboves[1065]), .FEAT_BELOW(feature_belows[1065])) ac1065(.scan_win(scan_win1065), .scan_win_std_dev(scan_win_std_dev[1065]), .feature_accum(feature_accums[1065]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1066]), .RECT1_Y(rectangle1_ys[1066]), .RECT1_WIDTH(rectangle1_widths[1066]), .RECT1_HEIGHT(rectangle1_heights[1066]), .RECT1_WEIGHT(rectangle1_weights[1066]), .RECT2_X(rectangle2_xs[1066]), .RECT2_Y(rectangle2_ys[1066]), .RECT2_WIDTH(rectangle2_widths[1066]), .RECT2_HEIGHT(rectangle2_heights[1066]), .RECT2_WEIGHT(rectangle2_weights[1066]), .RECT3_X(rectangle3_xs[1066]), .RECT3_Y(rectangle3_ys[1066]), .RECT3_WIDTH(rectangle3_widths[1066]), .RECT3_HEIGHT(rectangle3_heights[1066]), .RECT3_WEIGHT(rectangle3_weights[1066]), .FEAT_THRES(feature_thresholds[1066]), .FEAT_ABOVE(feature_aboves[1066]), .FEAT_BELOW(feature_belows[1066])) ac1066(.scan_win(scan_win1066), .scan_win_std_dev(scan_win_std_dev[1066]), .feature_accum(feature_accums[1066]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1067]), .RECT1_Y(rectangle1_ys[1067]), .RECT1_WIDTH(rectangle1_widths[1067]), .RECT1_HEIGHT(rectangle1_heights[1067]), .RECT1_WEIGHT(rectangle1_weights[1067]), .RECT2_X(rectangle2_xs[1067]), .RECT2_Y(rectangle2_ys[1067]), .RECT2_WIDTH(rectangle2_widths[1067]), .RECT2_HEIGHT(rectangle2_heights[1067]), .RECT2_WEIGHT(rectangle2_weights[1067]), .RECT3_X(rectangle3_xs[1067]), .RECT3_Y(rectangle3_ys[1067]), .RECT3_WIDTH(rectangle3_widths[1067]), .RECT3_HEIGHT(rectangle3_heights[1067]), .RECT3_WEIGHT(rectangle3_weights[1067]), .FEAT_THRES(feature_thresholds[1067]), .FEAT_ABOVE(feature_aboves[1067]), .FEAT_BELOW(feature_belows[1067])) ac1067(.scan_win(scan_win1067), .scan_win_std_dev(scan_win_std_dev[1067]), .feature_accum(feature_accums[1067]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1068]), .RECT1_Y(rectangle1_ys[1068]), .RECT1_WIDTH(rectangle1_widths[1068]), .RECT1_HEIGHT(rectangle1_heights[1068]), .RECT1_WEIGHT(rectangle1_weights[1068]), .RECT2_X(rectangle2_xs[1068]), .RECT2_Y(rectangle2_ys[1068]), .RECT2_WIDTH(rectangle2_widths[1068]), .RECT2_HEIGHT(rectangle2_heights[1068]), .RECT2_WEIGHT(rectangle2_weights[1068]), .RECT3_X(rectangle3_xs[1068]), .RECT3_Y(rectangle3_ys[1068]), .RECT3_WIDTH(rectangle3_widths[1068]), .RECT3_HEIGHT(rectangle3_heights[1068]), .RECT3_WEIGHT(rectangle3_weights[1068]), .FEAT_THRES(feature_thresholds[1068]), .FEAT_ABOVE(feature_aboves[1068]), .FEAT_BELOW(feature_belows[1068])) ac1068(.scan_win(scan_win1068), .scan_win_std_dev(scan_win_std_dev[1068]), .feature_accum(feature_accums[1068]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1069]), .RECT1_Y(rectangle1_ys[1069]), .RECT1_WIDTH(rectangle1_widths[1069]), .RECT1_HEIGHT(rectangle1_heights[1069]), .RECT1_WEIGHT(rectangle1_weights[1069]), .RECT2_X(rectangle2_xs[1069]), .RECT2_Y(rectangle2_ys[1069]), .RECT2_WIDTH(rectangle2_widths[1069]), .RECT2_HEIGHT(rectangle2_heights[1069]), .RECT2_WEIGHT(rectangle2_weights[1069]), .RECT3_X(rectangle3_xs[1069]), .RECT3_Y(rectangle3_ys[1069]), .RECT3_WIDTH(rectangle3_widths[1069]), .RECT3_HEIGHT(rectangle3_heights[1069]), .RECT3_WEIGHT(rectangle3_weights[1069]), .FEAT_THRES(feature_thresholds[1069]), .FEAT_ABOVE(feature_aboves[1069]), .FEAT_BELOW(feature_belows[1069])) ac1069(.scan_win(scan_win1069), .scan_win_std_dev(scan_win_std_dev[1069]), .feature_accum(feature_accums[1069]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1070]), .RECT1_Y(rectangle1_ys[1070]), .RECT1_WIDTH(rectangle1_widths[1070]), .RECT1_HEIGHT(rectangle1_heights[1070]), .RECT1_WEIGHT(rectangle1_weights[1070]), .RECT2_X(rectangle2_xs[1070]), .RECT2_Y(rectangle2_ys[1070]), .RECT2_WIDTH(rectangle2_widths[1070]), .RECT2_HEIGHT(rectangle2_heights[1070]), .RECT2_WEIGHT(rectangle2_weights[1070]), .RECT3_X(rectangle3_xs[1070]), .RECT3_Y(rectangle3_ys[1070]), .RECT3_WIDTH(rectangle3_widths[1070]), .RECT3_HEIGHT(rectangle3_heights[1070]), .RECT3_WEIGHT(rectangle3_weights[1070]), .FEAT_THRES(feature_thresholds[1070]), .FEAT_ABOVE(feature_aboves[1070]), .FEAT_BELOW(feature_belows[1070])) ac1070(.scan_win(scan_win1070), .scan_win_std_dev(scan_win_std_dev[1070]), .feature_accum(feature_accums[1070]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1071]), .RECT1_Y(rectangle1_ys[1071]), .RECT1_WIDTH(rectangle1_widths[1071]), .RECT1_HEIGHT(rectangle1_heights[1071]), .RECT1_WEIGHT(rectangle1_weights[1071]), .RECT2_X(rectangle2_xs[1071]), .RECT2_Y(rectangle2_ys[1071]), .RECT2_WIDTH(rectangle2_widths[1071]), .RECT2_HEIGHT(rectangle2_heights[1071]), .RECT2_WEIGHT(rectangle2_weights[1071]), .RECT3_X(rectangle3_xs[1071]), .RECT3_Y(rectangle3_ys[1071]), .RECT3_WIDTH(rectangle3_widths[1071]), .RECT3_HEIGHT(rectangle3_heights[1071]), .RECT3_WEIGHT(rectangle3_weights[1071]), .FEAT_THRES(feature_thresholds[1071]), .FEAT_ABOVE(feature_aboves[1071]), .FEAT_BELOW(feature_belows[1071])) ac1071(.scan_win(scan_win1071), .scan_win_std_dev(scan_win_std_dev[1071]), .feature_accum(feature_accums[1071]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1072]), .RECT1_Y(rectangle1_ys[1072]), .RECT1_WIDTH(rectangle1_widths[1072]), .RECT1_HEIGHT(rectangle1_heights[1072]), .RECT1_WEIGHT(rectangle1_weights[1072]), .RECT2_X(rectangle2_xs[1072]), .RECT2_Y(rectangle2_ys[1072]), .RECT2_WIDTH(rectangle2_widths[1072]), .RECT2_HEIGHT(rectangle2_heights[1072]), .RECT2_WEIGHT(rectangle2_weights[1072]), .RECT3_X(rectangle3_xs[1072]), .RECT3_Y(rectangle3_ys[1072]), .RECT3_WIDTH(rectangle3_widths[1072]), .RECT3_HEIGHT(rectangle3_heights[1072]), .RECT3_WEIGHT(rectangle3_weights[1072]), .FEAT_THRES(feature_thresholds[1072]), .FEAT_ABOVE(feature_aboves[1072]), .FEAT_BELOW(feature_belows[1072])) ac1072(.scan_win(scan_win1072), .scan_win_std_dev(scan_win_std_dev[1072]), .feature_accum(feature_accums[1072]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1073]), .RECT1_Y(rectangle1_ys[1073]), .RECT1_WIDTH(rectangle1_widths[1073]), .RECT1_HEIGHT(rectangle1_heights[1073]), .RECT1_WEIGHT(rectangle1_weights[1073]), .RECT2_X(rectangle2_xs[1073]), .RECT2_Y(rectangle2_ys[1073]), .RECT2_WIDTH(rectangle2_widths[1073]), .RECT2_HEIGHT(rectangle2_heights[1073]), .RECT2_WEIGHT(rectangle2_weights[1073]), .RECT3_X(rectangle3_xs[1073]), .RECT3_Y(rectangle3_ys[1073]), .RECT3_WIDTH(rectangle3_widths[1073]), .RECT3_HEIGHT(rectangle3_heights[1073]), .RECT3_WEIGHT(rectangle3_weights[1073]), .FEAT_THRES(feature_thresholds[1073]), .FEAT_ABOVE(feature_aboves[1073]), .FEAT_BELOW(feature_belows[1073])) ac1073(.scan_win(scan_win1073), .scan_win_std_dev(scan_win_std_dev[1073]), .feature_accum(feature_accums[1073]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1074]), .RECT1_Y(rectangle1_ys[1074]), .RECT1_WIDTH(rectangle1_widths[1074]), .RECT1_HEIGHT(rectangle1_heights[1074]), .RECT1_WEIGHT(rectangle1_weights[1074]), .RECT2_X(rectangle2_xs[1074]), .RECT2_Y(rectangle2_ys[1074]), .RECT2_WIDTH(rectangle2_widths[1074]), .RECT2_HEIGHT(rectangle2_heights[1074]), .RECT2_WEIGHT(rectangle2_weights[1074]), .RECT3_X(rectangle3_xs[1074]), .RECT3_Y(rectangle3_ys[1074]), .RECT3_WIDTH(rectangle3_widths[1074]), .RECT3_HEIGHT(rectangle3_heights[1074]), .RECT3_WEIGHT(rectangle3_weights[1074]), .FEAT_THRES(feature_thresholds[1074]), .FEAT_ABOVE(feature_aboves[1074]), .FEAT_BELOW(feature_belows[1074])) ac1074(.scan_win(scan_win1074), .scan_win_std_dev(scan_win_std_dev[1074]), .feature_accum(feature_accums[1074]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1075]), .RECT1_Y(rectangle1_ys[1075]), .RECT1_WIDTH(rectangle1_widths[1075]), .RECT1_HEIGHT(rectangle1_heights[1075]), .RECT1_WEIGHT(rectangle1_weights[1075]), .RECT2_X(rectangle2_xs[1075]), .RECT2_Y(rectangle2_ys[1075]), .RECT2_WIDTH(rectangle2_widths[1075]), .RECT2_HEIGHT(rectangle2_heights[1075]), .RECT2_WEIGHT(rectangle2_weights[1075]), .RECT3_X(rectangle3_xs[1075]), .RECT3_Y(rectangle3_ys[1075]), .RECT3_WIDTH(rectangle3_widths[1075]), .RECT3_HEIGHT(rectangle3_heights[1075]), .RECT3_WEIGHT(rectangle3_weights[1075]), .FEAT_THRES(feature_thresholds[1075]), .FEAT_ABOVE(feature_aboves[1075]), .FEAT_BELOW(feature_belows[1075])) ac1075(.scan_win(scan_win1075), .scan_win_std_dev(scan_win_std_dev[1075]), .feature_accum(feature_accums[1075]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1076]), .RECT1_Y(rectangle1_ys[1076]), .RECT1_WIDTH(rectangle1_widths[1076]), .RECT1_HEIGHT(rectangle1_heights[1076]), .RECT1_WEIGHT(rectangle1_weights[1076]), .RECT2_X(rectangle2_xs[1076]), .RECT2_Y(rectangle2_ys[1076]), .RECT2_WIDTH(rectangle2_widths[1076]), .RECT2_HEIGHT(rectangle2_heights[1076]), .RECT2_WEIGHT(rectangle2_weights[1076]), .RECT3_X(rectangle3_xs[1076]), .RECT3_Y(rectangle3_ys[1076]), .RECT3_WIDTH(rectangle3_widths[1076]), .RECT3_HEIGHT(rectangle3_heights[1076]), .RECT3_WEIGHT(rectangle3_weights[1076]), .FEAT_THRES(feature_thresholds[1076]), .FEAT_ABOVE(feature_aboves[1076]), .FEAT_BELOW(feature_belows[1076])) ac1076(.scan_win(scan_win1076), .scan_win_std_dev(scan_win_std_dev[1076]), .feature_accum(feature_accums[1076]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1077]), .RECT1_Y(rectangle1_ys[1077]), .RECT1_WIDTH(rectangle1_widths[1077]), .RECT1_HEIGHT(rectangle1_heights[1077]), .RECT1_WEIGHT(rectangle1_weights[1077]), .RECT2_X(rectangle2_xs[1077]), .RECT2_Y(rectangle2_ys[1077]), .RECT2_WIDTH(rectangle2_widths[1077]), .RECT2_HEIGHT(rectangle2_heights[1077]), .RECT2_WEIGHT(rectangle2_weights[1077]), .RECT3_X(rectangle3_xs[1077]), .RECT3_Y(rectangle3_ys[1077]), .RECT3_WIDTH(rectangle3_widths[1077]), .RECT3_HEIGHT(rectangle3_heights[1077]), .RECT3_WEIGHT(rectangle3_weights[1077]), .FEAT_THRES(feature_thresholds[1077]), .FEAT_ABOVE(feature_aboves[1077]), .FEAT_BELOW(feature_belows[1077])) ac1077(.scan_win(scan_win1077), .scan_win_std_dev(scan_win_std_dev[1077]), .feature_accum(feature_accums[1077]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1078]), .RECT1_Y(rectangle1_ys[1078]), .RECT1_WIDTH(rectangle1_widths[1078]), .RECT1_HEIGHT(rectangle1_heights[1078]), .RECT1_WEIGHT(rectangle1_weights[1078]), .RECT2_X(rectangle2_xs[1078]), .RECT2_Y(rectangle2_ys[1078]), .RECT2_WIDTH(rectangle2_widths[1078]), .RECT2_HEIGHT(rectangle2_heights[1078]), .RECT2_WEIGHT(rectangle2_weights[1078]), .RECT3_X(rectangle3_xs[1078]), .RECT3_Y(rectangle3_ys[1078]), .RECT3_WIDTH(rectangle3_widths[1078]), .RECT3_HEIGHT(rectangle3_heights[1078]), .RECT3_WEIGHT(rectangle3_weights[1078]), .FEAT_THRES(feature_thresholds[1078]), .FEAT_ABOVE(feature_aboves[1078]), .FEAT_BELOW(feature_belows[1078])) ac1078(.scan_win(scan_win1078), .scan_win_std_dev(scan_win_std_dev[1078]), .feature_accum(feature_accums[1078]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1079]), .RECT1_Y(rectangle1_ys[1079]), .RECT1_WIDTH(rectangle1_widths[1079]), .RECT1_HEIGHT(rectangle1_heights[1079]), .RECT1_WEIGHT(rectangle1_weights[1079]), .RECT2_X(rectangle2_xs[1079]), .RECT2_Y(rectangle2_ys[1079]), .RECT2_WIDTH(rectangle2_widths[1079]), .RECT2_HEIGHT(rectangle2_heights[1079]), .RECT2_WEIGHT(rectangle2_weights[1079]), .RECT3_X(rectangle3_xs[1079]), .RECT3_Y(rectangle3_ys[1079]), .RECT3_WIDTH(rectangle3_widths[1079]), .RECT3_HEIGHT(rectangle3_heights[1079]), .RECT3_WEIGHT(rectangle3_weights[1079]), .FEAT_THRES(feature_thresholds[1079]), .FEAT_ABOVE(feature_aboves[1079]), .FEAT_BELOW(feature_belows[1079])) ac1079(.scan_win(scan_win1079), .scan_win_std_dev(scan_win_std_dev[1079]), .feature_accum(feature_accums[1079]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1080]), .RECT1_Y(rectangle1_ys[1080]), .RECT1_WIDTH(rectangle1_widths[1080]), .RECT1_HEIGHT(rectangle1_heights[1080]), .RECT1_WEIGHT(rectangle1_weights[1080]), .RECT2_X(rectangle2_xs[1080]), .RECT2_Y(rectangle2_ys[1080]), .RECT2_WIDTH(rectangle2_widths[1080]), .RECT2_HEIGHT(rectangle2_heights[1080]), .RECT2_WEIGHT(rectangle2_weights[1080]), .RECT3_X(rectangle3_xs[1080]), .RECT3_Y(rectangle3_ys[1080]), .RECT3_WIDTH(rectangle3_widths[1080]), .RECT3_HEIGHT(rectangle3_heights[1080]), .RECT3_WEIGHT(rectangle3_weights[1080]), .FEAT_THRES(feature_thresholds[1080]), .FEAT_ABOVE(feature_aboves[1080]), .FEAT_BELOW(feature_belows[1080])) ac1080(.scan_win(scan_win1080), .scan_win_std_dev(scan_win_std_dev[1080]), .feature_accum(feature_accums[1080]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1081]), .RECT1_Y(rectangle1_ys[1081]), .RECT1_WIDTH(rectangle1_widths[1081]), .RECT1_HEIGHT(rectangle1_heights[1081]), .RECT1_WEIGHT(rectangle1_weights[1081]), .RECT2_X(rectangle2_xs[1081]), .RECT2_Y(rectangle2_ys[1081]), .RECT2_WIDTH(rectangle2_widths[1081]), .RECT2_HEIGHT(rectangle2_heights[1081]), .RECT2_WEIGHT(rectangle2_weights[1081]), .RECT3_X(rectangle3_xs[1081]), .RECT3_Y(rectangle3_ys[1081]), .RECT3_WIDTH(rectangle3_widths[1081]), .RECT3_HEIGHT(rectangle3_heights[1081]), .RECT3_WEIGHT(rectangle3_weights[1081]), .FEAT_THRES(feature_thresholds[1081]), .FEAT_ABOVE(feature_aboves[1081]), .FEAT_BELOW(feature_belows[1081])) ac1081(.scan_win(scan_win1081), .scan_win_std_dev(scan_win_std_dev[1081]), .feature_accum(feature_accums[1081]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1082]), .RECT1_Y(rectangle1_ys[1082]), .RECT1_WIDTH(rectangle1_widths[1082]), .RECT1_HEIGHT(rectangle1_heights[1082]), .RECT1_WEIGHT(rectangle1_weights[1082]), .RECT2_X(rectangle2_xs[1082]), .RECT2_Y(rectangle2_ys[1082]), .RECT2_WIDTH(rectangle2_widths[1082]), .RECT2_HEIGHT(rectangle2_heights[1082]), .RECT2_WEIGHT(rectangle2_weights[1082]), .RECT3_X(rectangle3_xs[1082]), .RECT3_Y(rectangle3_ys[1082]), .RECT3_WIDTH(rectangle3_widths[1082]), .RECT3_HEIGHT(rectangle3_heights[1082]), .RECT3_WEIGHT(rectangle3_weights[1082]), .FEAT_THRES(feature_thresholds[1082]), .FEAT_ABOVE(feature_aboves[1082]), .FEAT_BELOW(feature_belows[1082])) ac1082(.scan_win(scan_win1082), .scan_win_std_dev(scan_win_std_dev[1082]), .feature_accum(feature_accums[1082]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1083]), .RECT1_Y(rectangle1_ys[1083]), .RECT1_WIDTH(rectangle1_widths[1083]), .RECT1_HEIGHT(rectangle1_heights[1083]), .RECT1_WEIGHT(rectangle1_weights[1083]), .RECT2_X(rectangle2_xs[1083]), .RECT2_Y(rectangle2_ys[1083]), .RECT2_WIDTH(rectangle2_widths[1083]), .RECT2_HEIGHT(rectangle2_heights[1083]), .RECT2_WEIGHT(rectangle2_weights[1083]), .RECT3_X(rectangle3_xs[1083]), .RECT3_Y(rectangle3_ys[1083]), .RECT3_WIDTH(rectangle3_widths[1083]), .RECT3_HEIGHT(rectangle3_heights[1083]), .RECT3_WEIGHT(rectangle3_weights[1083]), .FEAT_THRES(feature_thresholds[1083]), .FEAT_ABOVE(feature_aboves[1083]), .FEAT_BELOW(feature_belows[1083])) ac1083(.scan_win(scan_win1083), .scan_win_std_dev(scan_win_std_dev[1083]), .feature_accum(feature_accums[1083]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1084]), .RECT1_Y(rectangle1_ys[1084]), .RECT1_WIDTH(rectangle1_widths[1084]), .RECT1_HEIGHT(rectangle1_heights[1084]), .RECT1_WEIGHT(rectangle1_weights[1084]), .RECT2_X(rectangle2_xs[1084]), .RECT2_Y(rectangle2_ys[1084]), .RECT2_WIDTH(rectangle2_widths[1084]), .RECT2_HEIGHT(rectangle2_heights[1084]), .RECT2_WEIGHT(rectangle2_weights[1084]), .RECT3_X(rectangle3_xs[1084]), .RECT3_Y(rectangle3_ys[1084]), .RECT3_WIDTH(rectangle3_widths[1084]), .RECT3_HEIGHT(rectangle3_heights[1084]), .RECT3_WEIGHT(rectangle3_weights[1084]), .FEAT_THRES(feature_thresholds[1084]), .FEAT_ABOVE(feature_aboves[1084]), .FEAT_BELOW(feature_belows[1084])) ac1084(.scan_win(scan_win1084), .scan_win_std_dev(scan_win_std_dev[1084]), .feature_accum(feature_accums[1084]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1085]), .RECT1_Y(rectangle1_ys[1085]), .RECT1_WIDTH(rectangle1_widths[1085]), .RECT1_HEIGHT(rectangle1_heights[1085]), .RECT1_WEIGHT(rectangle1_weights[1085]), .RECT2_X(rectangle2_xs[1085]), .RECT2_Y(rectangle2_ys[1085]), .RECT2_WIDTH(rectangle2_widths[1085]), .RECT2_HEIGHT(rectangle2_heights[1085]), .RECT2_WEIGHT(rectangle2_weights[1085]), .RECT3_X(rectangle3_xs[1085]), .RECT3_Y(rectangle3_ys[1085]), .RECT3_WIDTH(rectangle3_widths[1085]), .RECT3_HEIGHT(rectangle3_heights[1085]), .RECT3_WEIGHT(rectangle3_weights[1085]), .FEAT_THRES(feature_thresholds[1085]), .FEAT_ABOVE(feature_aboves[1085]), .FEAT_BELOW(feature_belows[1085])) ac1085(.scan_win(scan_win1085), .scan_win_std_dev(scan_win_std_dev[1085]), .feature_accum(feature_accums[1085]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1086]), .RECT1_Y(rectangle1_ys[1086]), .RECT1_WIDTH(rectangle1_widths[1086]), .RECT1_HEIGHT(rectangle1_heights[1086]), .RECT1_WEIGHT(rectangle1_weights[1086]), .RECT2_X(rectangle2_xs[1086]), .RECT2_Y(rectangle2_ys[1086]), .RECT2_WIDTH(rectangle2_widths[1086]), .RECT2_HEIGHT(rectangle2_heights[1086]), .RECT2_WEIGHT(rectangle2_weights[1086]), .RECT3_X(rectangle3_xs[1086]), .RECT3_Y(rectangle3_ys[1086]), .RECT3_WIDTH(rectangle3_widths[1086]), .RECT3_HEIGHT(rectangle3_heights[1086]), .RECT3_WEIGHT(rectangle3_weights[1086]), .FEAT_THRES(feature_thresholds[1086]), .FEAT_ABOVE(feature_aboves[1086]), .FEAT_BELOW(feature_belows[1086])) ac1086(.scan_win(scan_win1086), .scan_win_std_dev(scan_win_std_dev[1086]), .feature_accum(feature_accums[1086]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1087]), .RECT1_Y(rectangle1_ys[1087]), .RECT1_WIDTH(rectangle1_widths[1087]), .RECT1_HEIGHT(rectangle1_heights[1087]), .RECT1_WEIGHT(rectangle1_weights[1087]), .RECT2_X(rectangle2_xs[1087]), .RECT2_Y(rectangle2_ys[1087]), .RECT2_WIDTH(rectangle2_widths[1087]), .RECT2_HEIGHT(rectangle2_heights[1087]), .RECT2_WEIGHT(rectangle2_weights[1087]), .RECT3_X(rectangle3_xs[1087]), .RECT3_Y(rectangle3_ys[1087]), .RECT3_WIDTH(rectangle3_widths[1087]), .RECT3_HEIGHT(rectangle3_heights[1087]), .RECT3_WEIGHT(rectangle3_weights[1087]), .FEAT_THRES(feature_thresholds[1087]), .FEAT_ABOVE(feature_aboves[1087]), .FEAT_BELOW(feature_belows[1087])) ac1087(.scan_win(scan_win1087), .scan_win_std_dev(scan_win_std_dev[1087]), .feature_accum(feature_accums[1087]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1088]), .RECT1_Y(rectangle1_ys[1088]), .RECT1_WIDTH(rectangle1_widths[1088]), .RECT1_HEIGHT(rectangle1_heights[1088]), .RECT1_WEIGHT(rectangle1_weights[1088]), .RECT2_X(rectangle2_xs[1088]), .RECT2_Y(rectangle2_ys[1088]), .RECT2_WIDTH(rectangle2_widths[1088]), .RECT2_HEIGHT(rectangle2_heights[1088]), .RECT2_WEIGHT(rectangle2_weights[1088]), .RECT3_X(rectangle3_xs[1088]), .RECT3_Y(rectangle3_ys[1088]), .RECT3_WIDTH(rectangle3_widths[1088]), .RECT3_HEIGHT(rectangle3_heights[1088]), .RECT3_WEIGHT(rectangle3_weights[1088]), .FEAT_THRES(feature_thresholds[1088]), .FEAT_ABOVE(feature_aboves[1088]), .FEAT_BELOW(feature_belows[1088])) ac1088(.scan_win(scan_win1088), .scan_win_std_dev(scan_win_std_dev[1088]), .feature_accum(feature_accums[1088]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1089]), .RECT1_Y(rectangle1_ys[1089]), .RECT1_WIDTH(rectangle1_widths[1089]), .RECT1_HEIGHT(rectangle1_heights[1089]), .RECT1_WEIGHT(rectangle1_weights[1089]), .RECT2_X(rectangle2_xs[1089]), .RECT2_Y(rectangle2_ys[1089]), .RECT2_WIDTH(rectangle2_widths[1089]), .RECT2_HEIGHT(rectangle2_heights[1089]), .RECT2_WEIGHT(rectangle2_weights[1089]), .RECT3_X(rectangle3_xs[1089]), .RECT3_Y(rectangle3_ys[1089]), .RECT3_WIDTH(rectangle3_widths[1089]), .RECT3_HEIGHT(rectangle3_heights[1089]), .RECT3_WEIGHT(rectangle3_weights[1089]), .FEAT_THRES(feature_thresholds[1089]), .FEAT_ABOVE(feature_aboves[1089]), .FEAT_BELOW(feature_belows[1089])) ac1089(.scan_win(scan_win1089), .scan_win_std_dev(scan_win_std_dev[1089]), .feature_accum(feature_accums[1089]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1090]), .RECT1_Y(rectangle1_ys[1090]), .RECT1_WIDTH(rectangle1_widths[1090]), .RECT1_HEIGHT(rectangle1_heights[1090]), .RECT1_WEIGHT(rectangle1_weights[1090]), .RECT2_X(rectangle2_xs[1090]), .RECT2_Y(rectangle2_ys[1090]), .RECT2_WIDTH(rectangle2_widths[1090]), .RECT2_HEIGHT(rectangle2_heights[1090]), .RECT2_WEIGHT(rectangle2_weights[1090]), .RECT3_X(rectangle3_xs[1090]), .RECT3_Y(rectangle3_ys[1090]), .RECT3_WIDTH(rectangle3_widths[1090]), .RECT3_HEIGHT(rectangle3_heights[1090]), .RECT3_WEIGHT(rectangle3_weights[1090]), .FEAT_THRES(feature_thresholds[1090]), .FEAT_ABOVE(feature_aboves[1090]), .FEAT_BELOW(feature_belows[1090])) ac1090(.scan_win(scan_win1090), .scan_win_std_dev(scan_win_std_dev[1090]), .feature_accum(feature_accums[1090]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1091]), .RECT1_Y(rectangle1_ys[1091]), .RECT1_WIDTH(rectangle1_widths[1091]), .RECT1_HEIGHT(rectangle1_heights[1091]), .RECT1_WEIGHT(rectangle1_weights[1091]), .RECT2_X(rectangle2_xs[1091]), .RECT2_Y(rectangle2_ys[1091]), .RECT2_WIDTH(rectangle2_widths[1091]), .RECT2_HEIGHT(rectangle2_heights[1091]), .RECT2_WEIGHT(rectangle2_weights[1091]), .RECT3_X(rectangle3_xs[1091]), .RECT3_Y(rectangle3_ys[1091]), .RECT3_WIDTH(rectangle3_widths[1091]), .RECT3_HEIGHT(rectangle3_heights[1091]), .RECT3_WEIGHT(rectangle3_weights[1091]), .FEAT_THRES(feature_thresholds[1091]), .FEAT_ABOVE(feature_aboves[1091]), .FEAT_BELOW(feature_belows[1091])) ac1091(.scan_win(scan_win1091), .scan_win_std_dev(scan_win_std_dev[1091]), .feature_accum(feature_accums[1091]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1092]), .RECT1_Y(rectangle1_ys[1092]), .RECT1_WIDTH(rectangle1_widths[1092]), .RECT1_HEIGHT(rectangle1_heights[1092]), .RECT1_WEIGHT(rectangle1_weights[1092]), .RECT2_X(rectangle2_xs[1092]), .RECT2_Y(rectangle2_ys[1092]), .RECT2_WIDTH(rectangle2_widths[1092]), .RECT2_HEIGHT(rectangle2_heights[1092]), .RECT2_WEIGHT(rectangle2_weights[1092]), .RECT3_X(rectangle3_xs[1092]), .RECT3_Y(rectangle3_ys[1092]), .RECT3_WIDTH(rectangle3_widths[1092]), .RECT3_HEIGHT(rectangle3_heights[1092]), .RECT3_WEIGHT(rectangle3_weights[1092]), .FEAT_THRES(feature_thresholds[1092]), .FEAT_ABOVE(feature_aboves[1092]), .FEAT_BELOW(feature_belows[1092])) ac1092(.scan_win(scan_win1092), .scan_win_std_dev(scan_win_std_dev[1092]), .feature_accum(feature_accums[1092]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1093]), .RECT1_Y(rectangle1_ys[1093]), .RECT1_WIDTH(rectangle1_widths[1093]), .RECT1_HEIGHT(rectangle1_heights[1093]), .RECT1_WEIGHT(rectangle1_weights[1093]), .RECT2_X(rectangle2_xs[1093]), .RECT2_Y(rectangle2_ys[1093]), .RECT2_WIDTH(rectangle2_widths[1093]), .RECT2_HEIGHT(rectangle2_heights[1093]), .RECT2_WEIGHT(rectangle2_weights[1093]), .RECT3_X(rectangle3_xs[1093]), .RECT3_Y(rectangle3_ys[1093]), .RECT3_WIDTH(rectangle3_widths[1093]), .RECT3_HEIGHT(rectangle3_heights[1093]), .RECT3_WEIGHT(rectangle3_weights[1093]), .FEAT_THRES(feature_thresholds[1093]), .FEAT_ABOVE(feature_aboves[1093]), .FEAT_BELOW(feature_belows[1093])) ac1093(.scan_win(scan_win1093), .scan_win_std_dev(scan_win_std_dev[1093]), .feature_accum(feature_accums[1093]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1094]), .RECT1_Y(rectangle1_ys[1094]), .RECT1_WIDTH(rectangle1_widths[1094]), .RECT1_HEIGHT(rectangle1_heights[1094]), .RECT1_WEIGHT(rectangle1_weights[1094]), .RECT2_X(rectangle2_xs[1094]), .RECT2_Y(rectangle2_ys[1094]), .RECT2_WIDTH(rectangle2_widths[1094]), .RECT2_HEIGHT(rectangle2_heights[1094]), .RECT2_WEIGHT(rectangle2_weights[1094]), .RECT3_X(rectangle3_xs[1094]), .RECT3_Y(rectangle3_ys[1094]), .RECT3_WIDTH(rectangle3_widths[1094]), .RECT3_HEIGHT(rectangle3_heights[1094]), .RECT3_WEIGHT(rectangle3_weights[1094]), .FEAT_THRES(feature_thresholds[1094]), .FEAT_ABOVE(feature_aboves[1094]), .FEAT_BELOW(feature_belows[1094])) ac1094(.scan_win(scan_win1094), .scan_win_std_dev(scan_win_std_dev[1094]), .feature_accum(feature_accums[1094]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1095]), .RECT1_Y(rectangle1_ys[1095]), .RECT1_WIDTH(rectangle1_widths[1095]), .RECT1_HEIGHT(rectangle1_heights[1095]), .RECT1_WEIGHT(rectangle1_weights[1095]), .RECT2_X(rectangle2_xs[1095]), .RECT2_Y(rectangle2_ys[1095]), .RECT2_WIDTH(rectangle2_widths[1095]), .RECT2_HEIGHT(rectangle2_heights[1095]), .RECT2_WEIGHT(rectangle2_weights[1095]), .RECT3_X(rectangle3_xs[1095]), .RECT3_Y(rectangle3_ys[1095]), .RECT3_WIDTH(rectangle3_widths[1095]), .RECT3_HEIGHT(rectangle3_heights[1095]), .RECT3_WEIGHT(rectangle3_weights[1095]), .FEAT_THRES(feature_thresholds[1095]), .FEAT_ABOVE(feature_aboves[1095]), .FEAT_BELOW(feature_belows[1095])) ac1095(.scan_win(scan_win1095), .scan_win_std_dev(scan_win_std_dev[1095]), .feature_accum(feature_accums[1095]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1096]), .RECT1_Y(rectangle1_ys[1096]), .RECT1_WIDTH(rectangle1_widths[1096]), .RECT1_HEIGHT(rectangle1_heights[1096]), .RECT1_WEIGHT(rectangle1_weights[1096]), .RECT2_X(rectangle2_xs[1096]), .RECT2_Y(rectangle2_ys[1096]), .RECT2_WIDTH(rectangle2_widths[1096]), .RECT2_HEIGHT(rectangle2_heights[1096]), .RECT2_WEIGHT(rectangle2_weights[1096]), .RECT3_X(rectangle3_xs[1096]), .RECT3_Y(rectangle3_ys[1096]), .RECT3_WIDTH(rectangle3_widths[1096]), .RECT3_HEIGHT(rectangle3_heights[1096]), .RECT3_WEIGHT(rectangle3_weights[1096]), .FEAT_THRES(feature_thresholds[1096]), .FEAT_ABOVE(feature_aboves[1096]), .FEAT_BELOW(feature_belows[1096])) ac1096(.scan_win(scan_win1096), .scan_win_std_dev(scan_win_std_dev[1096]), .feature_accum(feature_accums[1096]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1097]), .RECT1_Y(rectangle1_ys[1097]), .RECT1_WIDTH(rectangle1_widths[1097]), .RECT1_HEIGHT(rectangle1_heights[1097]), .RECT1_WEIGHT(rectangle1_weights[1097]), .RECT2_X(rectangle2_xs[1097]), .RECT2_Y(rectangle2_ys[1097]), .RECT2_WIDTH(rectangle2_widths[1097]), .RECT2_HEIGHT(rectangle2_heights[1097]), .RECT2_WEIGHT(rectangle2_weights[1097]), .RECT3_X(rectangle3_xs[1097]), .RECT3_Y(rectangle3_ys[1097]), .RECT3_WIDTH(rectangle3_widths[1097]), .RECT3_HEIGHT(rectangle3_heights[1097]), .RECT3_WEIGHT(rectangle3_weights[1097]), .FEAT_THRES(feature_thresholds[1097]), .FEAT_ABOVE(feature_aboves[1097]), .FEAT_BELOW(feature_belows[1097])) ac1097(.scan_win(scan_win1097), .scan_win_std_dev(scan_win_std_dev[1097]), .feature_accum(feature_accums[1097]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1098]), .RECT1_Y(rectangle1_ys[1098]), .RECT1_WIDTH(rectangle1_widths[1098]), .RECT1_HEIGHT(rectangle1_heights[1098]), .RECT1_WEIGHT(rectangle1_weights[1098]), .RECT2_X(rectangle2_xs[1098]), .RECT2_Y(rectangle2_ys[1098]), .RECT2_WIDTH(rectangle2_widths[1098]), .RECT2_HEIGHT(rectangle2_heights[1098]), .RECT2_WEIGHT(rectangle2_weights[1098]), .RECT3_X(rectangle3_xs[1098]), .RECT3_Y(rectangle3_ys[1098]), .RECT3_WIDTH(rectangle3_widths[1098]), .RECT3_HEIGHT(rectangle3_heights[1098]), .RECT3_WEIGHT(rectangle3_weights[1098]), .FEAT_THRES(feature_thresholds[1098]), .FEAT_ABOVE(feature_aboves[1098]), .FEAT_BELOW(feature_belows[1098])) ac1098(.scan_win(scan_win1098), .scan_win_std_dev(scan_win_std_dev[1098]), .feature_accum(feature_accums[1098]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1099]), .RECT1_Y(rectangle1_ys[1099]), .RECT1_WIDTH(rectangle1_widths[1099]), .RECT1_HEIGHT(rectangle1_heights[1099]), .RECT1_WEIGHT(rectangle1_weights[1099]), .RECT2_X(rectangle2_xs[1099]), .RECT2_Y(rectangle2_ys[1099]), .RECT2_WIDTH(rectangle2_widths[1099]), .RECT2_HEIGHT(rectangle2_heights[1099]), .RECT2_WEIGHT(rectangle2_weights[1099]), .RECT3_X(rectangle3_xs[1099]), .RECT3_Y(rectangle3_ys[1099]), .RECT3_WIDTH(rectangle3_widths[1099]), .RECT3_HEIGHT(rectangle3_heights[1099]), .RECT3_WEIGHT(rectangle3_weights[1099]), .FEAT_THRES(feature_thresholds[1099]), .FEAT_ABOVE(feature_aboves[1099]), .FEAT_BELOW(feature_belows[1099])) ac1099(.scan_win(scan_win1099), .scan_win_std_dev(scan_win_std_dev[1099]), .feature_accum(feature_accums[1099]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1100]), .RECT1_Y(rectangle1_ys[1100]), .RECT1_WIDTH(rectangle1_widths[1100]), .RECT1_HEIGHT(rectangle1_heights[1100]), .RECT1_WEIGHT(rectangle1_weights[1100]), .RECT2_X(rectangle2_xs[1100]), .RECT2_Y(rectangle2_ys[1100]), .RECT2_WIDTH(rectangle2_widths[1100]), .RECT2_HEIGHT(rectangle2_heights[1100]), .RECT2_WEIGHT(rectangle2_weights[1100]), .RECT3_X(rectangle3_xs[1100]), .RECT3_Y(rectangle3_ys[1100]), .RECT3_WIDTH(rectangle3_widths[1100]), .RECT3_HEIGHT(rectangle3_heights[1100]), .RECT3_WEIGHT(rectangle3_weights[1100]), .FEAT_THRES(feature_thresholds[1100]), .FEAT_ABOVE(feature_aboves[1100]), .FEAT_BELOW(feature_belows[1100])) ac1100(.scan_win(scan_win1100), .scan_win_std_dev(scan_win_std_dev[1100]), .feature_accum(feature_accums[1100]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1101]), .RECT1_Y(rectangle1_ys[1101]), .RECT1_WIDTH(rectangle1_widths[1101]), .RECT1_HEIGHT(rectangle1_heights[1101]), .RECT1_WEIGHT(rectangle1_weights[1101]), .RECT2_X(rectangle2_xs[1101]), .RECT2_Y(rectangle2_ys[1101]), .RECT2_WIDTH(rectangle2_widths[1101]), .RECT2_HEIGHT(rectangle2_heights[1101]), .RECT2_WEIGHT(rectangle2_weights[1101]), .RECT3_X(rectangle3_xs[1101]), .RECT3_Y(rectangle3_ys[1101]), .RECT3_WIDTH(rectangle3_widths[1101]), .RECT3_HEIGHT(rectangle3_heights[1101]), .RECT3_WEIGHT(rectangle3_weights[1101]), .FEAT_THRES(feature_thresholds[1101]), .FEAT_ABOVE(feature_aboves[1101]), .FEAT_BELOW(feature_belows[1101])) ac1101(.scan_win(scan_win1101), .scan_win_std_dev(scan_win_std_dev[1101]), .feature_accum(feature_accums[1101]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1102]), .RECT1_Y(rectangle1_ys[1102]), .RECT1_WIDTH(rectangle1_widths[1102]), .RECT1_HEIGHT(rectangle1_heights[1102]), .RECT1_WEIGHT(rectangle1_weights[1102]), .RECT2_X(rectangle2_xs[1102]), .RECT2_Y(rectangle2_ys[1102]), .RECT2_WIDTH(rectangle2_widths[1102]), .RECT2_HEIGHT(rectangle2_heights[1102]), .RECT2_WEIGHT(rectangle2_weights[1102]), .RECT3_X(rectangle3_xs[1102]), .RECT3_Y(rectangle3_ys[1102]), .RECT3_WIDTH(rectangle3_widths[1102]), .RECT3_HEIGHT(rectangle3_heights[1102]), .RECT3_WEIGHT(rectangle3_weights[1102]), .FEAT_THRES(feature_thresholds[1102]), .FEAT_ABOVE(feature_aboves[1102]), .FEAT_BELOW(feature_belows[1102])) ac1102(.scan_win(scan_win1102), .scan_win_std_dev(scan_win_std_dev[1102]), .feature_accum(feature_accums[1102]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1103]), .RECT1_Y(rectangle1_ys[1103]), .RECT1_WIDTH(rectangle1_widths[1103]), .RECT1_HEIGHT(rectangle1_heights[1103]), .RECT1_WEIGHT(rectangle1_weights[1103]), .RECT2_X(rectangle2_xs[1103]), .RECT2_Y(rectangle2_ys[1103]), .RECT2_WIDTH(rectangle2_widths[1103]), .RECT2_HEIGHT(rectangle2_heights[1103]), .RECT2_WEIGHT(rectangle2_weights[1103]), .RECT3_X(rectangle3_xs[1103]), .RECT3_Y(rectangle3_ys[1103]), .RECT3_WIDTH(rectangle3_widths[1103]), .RECT3_HEIGHT(rectangle3_heights[1103]), .RECT3_WEIGHT(rectangle3_weights[1103]), .FEAT_THRES(feature_thresholds[1103]), .FEAT_ABOVE(feature_aboves[1103]), .FEAT_BELOW(feature_belows[1103])) ac1103(.scan_win(scan_win1103), .scan_win_std_dev(scan_win_std_dev[1103]), .feature_accum(feature_accums[1103]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1104]), .RECT1_Y(rectangle1_ys[1104]), .RECT1_WIDTH(rectangle1_widths[1104]), .RECT1_HEIGHT(rectangle1_heights[1104]), .RECT1_WEIGHT(rectangle1_weights[1104]), .RECT2_X(rectangle2_xs[1104]), .RECT2_Y(rectangle2_ys[1104]), .RECT2_WIDTH(rectangle2_widths[1104]), .RECT2_HEIGHT(rectangle2_heights[1104]), .RECT2_WEIGHT(rectangle2_weights[1104]), .RECT3_X(rectangle3_xs[1104]), .RECT3_Y(rectangle3_ys[1104]), .RECT3_WIDTH(rectangle3_widths[1104]), .RECT3_HEIGHT(rectangle3_heights[1104]), .RECT3_WEIGHT(rectangle3_weights[1104]), .FEAT_THRES(feature_thresholds[1104]), .FEAT_ABOVE(feature_aboves[1104]), .FEAT_BELOW(feature_belows[1104])) ac1104(.scan_win(scan_win1104), .scan_win_std_dev(scan_win_std_dev[1104]), .feature_accum(feature_accums[1104]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1105]), .RECT1_Y(rectangle1_ys[1105]), .RECT1_WIDTH(rectangle1_widths[1105]), .RECT1_HEIGHT(rectangle1_heights[1105]), .RECT1_WEIGHT(rectangle1_weights[1105]), .RECT2_X(rectangle2_xs[1105]), .RECT2_Y(rectangle2_ys[1105]), .RECT2_WIDTH(rectangle2_widths[1105]), .RECT2_HEIGHT(rectangle2_heights[1105]), .RECT2_WEIGHT(rectangle2_weights[1105]), .RECT3_X(rectangle3_xs[1105]), .RECT3_Y(rectangle3_ys[1105]), .RECT3_WIDTH(rectangle3_widths[1105]), .RECT3_HEIGHT(rectangle3_heights[1105]), .RECT3_WEIGHT(rectangle3_weights[1105]), .FEAT_THRES(feature_thresholds[1105]), .FEAT_ABOVE(feature_aboves[1105]), .FEAT_BELOW(feature_belows[1105])) ac1105(.scan_win(scan_win1105), .scan_win_std_dev(scan_win_std_dev[1105]), .feature_accum(feature_accums[1105]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1106]), .RECT1_Y(rectangle1_ys[1106]), .RECT1_WIDTH(rectangle1_widths[1106]), .RECT1_HEIGHT(rectangle1_heights[1106]), .RECT1_WEIGHT(rectangle1_weights[1106]), .RECT2_X(rectangle2_xs[1106]), .RECT2_Y(rectangle2_ys[1106]), .RECT2_WIDTH(rectangle2_widths[1106]), .RECT2_HEIGHT(rectangle2_heights[1106]), .RECT2_WEIGHT(rectangle2_weights[1106]), .RECT3_X(rectangle3_xs[1106]), .RECT3_Y(rectangle3_ys[1106]), .RECT3_WIDTH(rectangle3_widths[1106]), .RECT3_HEIGHT(rectangle3_heights[1106]), .RECT3_WEIGHT(rectangle3_weights[1106]), .FEAT_THRES(feature_thresholds[1106]), .FEAT_ABOVE(feature_aboves[1106]), .FEAT_BELOW(feature_belows[1106])) ac1106(.scan_win(scan_win1106), .scan_win_std_dev(scan_win_std_dev[1106]), .feature_accum(feature_accums[1106]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1107]), .RECT1_Y(rectangle1_ys[1107]), .RECT1_WIDTH(rectangle1_widths[1107]), .RECT1_HEIGHT(rectangle1_heights[1107]), .RECT1_WEIGHT(rectangle1_weights[1107]), .RECT2_X(rectangle2_xs[1107]), .RECT2_Y(rectangle2_ys[1107]), .RECT2_WIDTH(rectangle2_widths[1107]), .RECT2_HEIGHT(rectangle2_heights[1107]), .RECT2_WEIGHT(rectangle2_weights[1107]), .RECT3_X(rectangle3_xs[1107]), .RECT3_Y(rectangle3_ys[1107]), .RECT3_WIDTH(rectangle3_widths[1107]), .RECT3_HEIGHT(rectangle3_heights[1107]), .RECT3_WEIGHT(rectangle3_weights[1107]), .FEAT_THRES(feature_thresholds[1107]), .FEAT_ABOVE(feature_aboves[1107]), .FEAT_BELOW(feature_belows[1107])) ac1107(.scan_win(scan_win1107), .scan_win_std_dev(scan_win_std_dev[1107]), .feature_accum(feature_accums[1107]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1108]), .RECT1_Y(rectangle1_ys[1108]), .RECT1_WIDTH(rectangle1_widths[1108]), .RECT1_HEIGHT(rectangle1_heights[1108]), .RECT1_WEIGHT(rectangle1_weights[1108]), .RECT2_X(rectangle2_xs[1108]), .RECT2_Y(rectangle2_ys[1108]), .RECT2_WIDTH(rectangle2_widths[1108]), .RECT2_HEIGHT(rectangle2_heights[1108]), .RECT2_WEIGHT(rectangle2_weights[1108]), .RECT3_X(rectangle3_xs[1108]), .RECT3_Y(rectangle3_ys[1108]), .RECT3_WIDTH(rectangle3_widths[1108]), .RECT3_HEIGHT(rectangle3_heights[1108]), .RECT3_WEIGHT(rectangle3_weights[1108]), .FEAT_THRES(feature_thresholds[1108]), .FEAT_ABOVE(feature_aboves[1108]), .FEAT_BELOW(feature_belows[1108])) ac1108(.scan_win(scan_win1108), .scan_win_std_dev(scan_win_std_dev[1108]), .feature_accum(feature_accums[1108]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1109]), .RECT1_Y(rectangle1_ys[1109]), .RECT1_WIDTH(rectangle1_widths[1109]), .RECT1_HEIGHT(rectangle1_heights[1109]), .RECT1_WEIGHT(rectangle1_weights[1109]), .RECT2_X(rectangle2_xs[1109]), .RECT2_Y(rectangle2_ys[1109]), .RECT2_WIDTH(rectangle2_widths[1109]), .RECT2_HEIGHT(rectangle2_heights[1109]), .RECT2_WEIGHT(rectangle2_weights[1109]), .RECT3_X(rectangle3_xs[1109]), .RECT3_Y(rectangle3_ys[1109]), .RECT3_WIDTH(rectangle3_widths[1109]), .RECT3_HEIGHT(rectangle3_heights[1109]), .RECT3_WEIGHT(rectangle3_weights[1109]), .FEAT_THRES(feature_thresholds[1109]), .FEAT_ABOVE(feature_aboves[1109]), .FEAT_BELOW(feature_belows[1109])) ac1109(.scan_win(scan_win1109), .scan_win_std_dev(scan_win_std_dev[1109]), .feature_accum(feature_accums[1109]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1110]), .RECT1_Y(rectangle1_ys[1110]), .RECT1_WIDTH(rectangle1_widths[1110]), .RECT1_HEIGHT(rectangle1_heights[1110]), .RECT1_WEIGHT(rectangle1_weights[1110]), .RECT2_X(rectangle2_xs[1110]), .RECT2_Y(rectangle2_ys[1110]), .RECT2_WIDTH(rectangle2_widths[1110]), .RECT2_HEIGHT(rectangle2_heights[1110]), .RECT2_WEIGHT(rectangle2_weights[1110]), .RECT3_X(rectangle3_xs[1110]), .RECT3_Y(rectangle3_ys[1110]), .RECT3_WIDTH(rectangle3_widths[1110]), .RECT3_HEIGHT(rectangle3_heights[1110]), .RECT3_WEIGHT(rectangle3_weights[1110]), .FEAT_THRES(feature_thresholds[1110]), .FEAT_ABOVE(feature_aboves[1110]), .FEAT_BELOW(feature_belows[1110])) ac1110(.scan_win(scan_win1110), .scan_win_std_dev(scan_win_std_dev[1110]), .feature_accum(feature_accums[1110]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1111]), .RECT1_Y(rectangle1_ys[1111]), .RECT1_WIDTH(rectangle1_widths[1111]), .RECT1_HEIGHT(rectangle1_heights[1111]), .RECT1_WEIGHT(rectangle1_weights[1111]), .RECT2_X(rectangle2_xs[1111]), .RECT2_Y(rectangle2_ys[1111]), .RECT2_WIDTH(rectangle2_widths[1111]), .RECT2_HEIGHT(rectangle2_heights[1111]), .RECT2_WEIGHT(rectangle2_weights[1111]), .RECT3_X(rectangle3_xs[1111]), .RECT3_Y(rectangle3_ys[1111]), .RECT3_WIDTH(rectangle3_widths[1111]), .RECT3_HEIGHT(rectangle3_heights[1111]), .RECT3_WEIGHT(rectangle3_weights[1111]), .FEAT_THRES(feature_thresholds[1111]), .FEAT_ABOVE(feature_aboves[1111]), .FEAT_BELOW(feature_belows[1111])) ac1111(.scan_win(scan_win1111), .scan_win_std_dev(scan_win_std_dev[1111]), .feature_accum(feature_accums[1111]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1112]), .RECT1_Y(rectangle1_ys[1112]), .RECT1_WIDTH(rectangle1_widths[1112]), .RECT1_HEIGHT(rectangle1_heights[1112]), .RECT1_WEIGHT(rectangle1_weights[1112]), .RECT2_X(rectangle2_xs[1112]), .RECT2_Y(rectangle2_ys[1112]), .RECT2_WIDTH(rectangle2_widths[1112]), .RECT2_HEIGHT(rectangle2_heights[1112]), .RECT2_WEIGHT(rectangle2_weights[1112]), .RECT3_X(rectangle3_xs[1112]), .RECT3_Y(rectangle3_ys[1112]), .RECT3_WIDTH(rectangle3_widths[1112]), .RECT3_HEIGHT(rectangle3_heights[1112]), .RECT3_WEIGHT(rectangle3_weights[1112]), .FEAT_THRES(feature_thresholds[1112]), .FEAT_ABOVE(feature_aboves[1112]), .FEAT_BELOW(feature_belows[1112])) ac1112(.scan_win(scan_win1112), .scan_win_std_dev(scan_win_std_dev[1112]), .feature_accum(feature_accums[1112]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1113]), .RECT1_Y(rectangle1_ys[1113]), .RECT1_WIDTH(rectangle1_widths[1113]), .RECT1_HEIGHT(rectangle1_heights[1113]), .RECT1_WEIGHT(rectangle1_weights[1113]), .RECT2_X(rectangle2_xs[1113]), .RECT2_Y(rectangle2_ys[1113]), .RECT2_WIDTH(rectangle2_widths[1113]), .RECT2_HEIGHT(rectangle2_heights[1113]), .RECT2_WEIGHT(rectangle2_weights[1113]), .RECT3_X(rectangle3_xs[1113]), .RECT3_Y(rectangle3_ys[1113]), .RECT3_WIDTH(rectangle3_widths[1113]), .RECT3_HEIGHT(rectangle3_heights[1113]), .RECT3_WEIGHT(rectangle3_weights[1113]), .FEAT_THRES(feature_thresholds[1113]), .FEAT_ABOVE(feature_aboves[1113]), .FEAT_BELOW(feature_belows[1113])) ac1113(.scan_win(scan_win1113), .scan_win_std_dev(scan_win_std_dev[1113]), .feature_accum(feature_accums[1113]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1114]), .RECT1_Y(rectangle1_ys[1114]), .RECT1_WIDTH(rectangle1_widths[1114]), .RECT1_HEIGHT(rectangle1_heights[1114]), .RECT1_WEIGHT(rectangle1_weights[1114]), .RECT2_X(rectangle2_xs[1114]), .RECT2_Y(rectangle2_ys[1114]), .RECT2_WIDTH(rectangle2_widths[1114]), .RECT2_HEIGHT(rectangle2_heights[1114]), .RECT2_WEIGHT(rectangle2_weights[1114]), .RECT3_X(rectangle3_xs[1114]), .RECT3_Y(rectangle3_ys[1114]), .RECT3_WIDTH(rectangle3_widths[1114]), .RECT3_HEIGHT(rectangle3_heights[1114]), .RECT3_WEIGHT(rectangle3_weights[1114]), .FEAT_THRES(feature_thresholds[1114]), .FEAT_ABOVE(feature_aboves[1114]), .FEAT_BELOW(feature_belows[1114])) ac1114(.scan_win(scan_win1114), .scan_win_std_dev(scan_win_std_dev[1114]), .feature_accum(feature_accums[1114]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1115]), .RECT1_Y(rectangle1_ys[1115]), .RECT1_WIDTH(rectangle1_widths[1115]), .RECT1_HEIGHT(rectangle1_heights[1115]), .RECT1_WEIGHT(rectangle1_weights[1115]), .RECT2_X(rectangle2_xs[1115]), .RECT2_Y(rectangle2_ys[1115]), .RECT2_WIDTH(rectangle2_widths[1115]), .RECT2_HEIGHT(rectangle2_heights[1115]), .RECT2_WEIGHT(rectangle2_weights[1115]), .RECT3_X(rectangle3_xs[1115]), .RECT3_Y(rectangle3_ys[1115]), .RECT3_WIDTH(rectangle3_widths[1115]), .RECT3_HEIGHT(rectangle3_heights[1115]), .RECT3_WEIGHT(rectangle3_weights[1115]), .FEAT_THRES(feature_thresholds[1115]), .FEAT_ABOVE(feature_aboves[1115]), .FEAT_BELOW(feature_belows[1115])) ac1115(.scan_win(scan_win1115), .scan_win_std_dev(scan_win_std_dev[1115]), .feature_accum(feature_accums[1115]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1116]), .RECT1_Y(rectangle1_ys[1116]), .RECT1_WIDTH(rectangle1_widths[1116]), .RECT1_HEIGHT(rectangle1_heights[1116]), .RECT1_WEIGHT(rectangle1_weights[1116]), .RECT2_X(rectangle2_xs[1116]), .RECT2_Y(rectangle2_ys[1116]), .RECT2_WIDTH(rectangle2_widths[1116]), .RECT2_HEIGHT(rectangle2_heights[1116]), .RECT2_WEIGHT(rectangle2_weights[1116]), .RECT3_X(rectangle3_xs[1116]), .RECT3_Y(rectangle3_ys[1116]), .RECT3_WIDTH(rectangle3_widths[1116]), .RECT3_HEIGHT(rectangle3_heights[1116]), .RECT3_WEIGHT(rectangle3_weights[1116]), .FEAT_THRES(feature_thresholds[1116]), .FEAT_ABOVE(feature_aboves[1116]), .FEAT_BELOW(feature_belows[1116])) ac1116(.scan_win(scan_win1116), .scan_win_std_dev(scan_win_std_dev[1116]), .feature_accum(feature_accums[1116]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1117]), .RECT1_Y(rectangle1_ys[1117]), .RECT1_WIDTH(rectangle1_widths[1117]), .RECT1_HEIGHT(rectangle1_heights[1117]), .RECT1_WEIGHT(rectangle1_weights[1117]), .RECT2_X(rectangle2_xs[1117]), .RECT2_Y(rectangle2_ys[1117]), .RECT2_WIDTH(rectangle2_widths[1117]), .RECT2_HEIGHT(rectangle2_heights[1117]), .RECT2_WEIGHT(rectangle2_weights[1117]), .RECT3_X(rectangle3_xs[1117]), .RECT3_Y(rectangle3_ys[1117]), .RECT3_WIDTH(rectangle3_widths[1117]), .RECT3_HEIGHT(rectangle3_heights[1117]), .RECT3_WEIGHT(rectangle3_weights[1117]), .FEAT_THRES(feature_thresholds[1117]), .FEAT_ABOVE(feature_aboves[1117]), .FEAT_BELOW(feature_belows[1117])) ac1117(.scan_win(scan_win1117), .scan_win_std_dev(scan_win_std_dev[1117]), .feature_accum(feature_accums[1117]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1118]), .RECT1_Y(rectangle1_ys[1118]), .RECT1_WIDTH(rectangle1_widths[1118]), .RECT1_HEIGHT(rectangle1_heights[1118]), .RECT1_WEIGHT(rectangle1_weights[1118]), .RECT2_X(rectangle2_xs[1118]), .RECT2_Y(rectangle2_ys[1118]), .RECT2_WIDTH(rectangle2_widths[1118]), .RECT2_HEIGHT(rectangle2_heights[1118]), .RECT2_WEIGHT(rectangle2_weights[1118]), .RECT3_X(rectangle3_xs[1118]), .RECT3_Y(rectangle3_ys[1118]), .RECT3_WIDTH(rectangle3_widths[1118]), .RECT3_HEIGHT(rectangle3_heights[1118]), .RECT3_WEIGHT(rectangle3_weights[1118]), .FEAT_THRES(feature_thresholds[1118]), .FEAT_ABOVE(feature_aboves[1118]), .FEAT_BELOW(feature_belows[1118])) ac1118(.scan_win(scan_win1118), .scan_win_std_dev(scan_win_std_dev[1118]), .feature_accum(feature_accums[1118]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1119]), .RECT1_Y(rectangle1_ys[1119]), .RECT1_WIDTH(rectangle1_widths[1119]), .RECT1_HEIGHT(rectangle1_heights[1119]), .RECT1_WEIGHT(rectangle1_weights[1119]), .RECT2_X(rectangle2_xs[1119]), .RECT2_Y(rectangle2_ys[1119]), .RECT2_WIDTH(rectangle2_widths[1119]), .RECT2_HEIGHT(rectangle2_heights[1119]), .RECT2_WEIGHT(rectangle2_weights[1119]), .RECT3_X(rectangle3_xs[1119]), .RECT3_Y(rectangle3_ys[1119]), .RECT3_WIDTH(rectangle3_widths[1119]), .RECT3_HEIGHT(rectangle3_heights[1119]), .RECT3_WEIGHT(rectangle3_weights[1119]), .FEAT_THRES(feature_thresholds[1119]), .FEAT_ABOVE(feature_aboves[1119]), .FEAT_BELOW(feature_belows[1119])) ac1119(.scan_win(scan_win1119), .scan_win_std_dev(scan_win_std_dev[1119]), .feature_accum(feature_accums[1119]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1120]), .RECT1_Y(rectangle1_ys[1120]), .RECT1_WIDTH(rectangle1_widths[1120]), .RECT1_HEIGHT(rectangle1_heights[1120]), .RECT1_WEIGHT(rectangle1_weights[1120]), .RECT2_X(rectangle2_xs[1120]), .RECT2_Y(rectangle2_ys[1120]), .RECT2_WIDTH(rectangle2_widths[1120]), .RECT2_HEIGHT(rectangle2_heights[1120]), .RECT2_WEIGHT(rectangle2_weights[1120]), .RECT3_X(rectangle3_xs[1120]), .RECT3_Y(rectangle3_ys[1120]), .RECT3_WIDTH(rectangle3_widths[1120]), .RECT3_HEIGHT(rectangle3_heights[1120]), .RECT3_WEIGHT(rectangle3_weights[1120]), .FEAT_THRES(feature_thresholds[1120]), .FEAT_ABOVE(feature_aboves[1120]), .FEAT_BELOW(feature_belows[1120])) ac1120(.scan_win(scan_win1120), .scan_win_std_dev(scan_win_std_dev[1120]), .feature_accum(feature_accums[1120]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1121]), .RECT1_Y(rectangle1_ys[1121]), .RECT1_WIDTH(rectangle1_widths[1121]), .RECT1_HEIGHT(rectangle1_heights[1121]), .RECT1_WEIGHT(rectangle1_weights[1121]), .RECT2_X(rectangle2_xs[1121]), .RECT2_Y(rectangle2_ys[1121]), .RECT2_WIDTH(rectangle2_widths[1121]), .RECT2_HEIGHT(rectangle2_heights[1121]), .RECT2_WEIGHT(rectangle2_weights[1121]), .RECT3_X(rectangle3_xs[1121]), .RECT3_Y(rectangle3_ys[1121]), .RECT3_WIDTH(rectangle3_widths[1121]), .RECT3_HEIGHT(rectangle3_heights[1121]), .RECT3_WEIGHT(rectangle3_weights[1121]), .FEAT_THRES(feature_thresholds[1121]), .FEAT_ABOVE(feature_aboves[1121]), .FEAT_BELOW(feature_belows[1121])) ac1121(.scan_win(scan_win1121), .scan_win_std_dev(scan_win_std_dev[1121]), .feature_accum(feature_accums[1121]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1122]), .RECT1_Y(rectangle1_ys[1122]), .RECT1_WIDTH(rectangle1_widths[1122]), .RECT1_HEIGHT(rectangle1_heights[1122]), .RECT1_WEIGHT(rectangle1_weights[1122]), .RECT2_X(rectangle2_xs[1122]), .RECT2_Y(rectangle2_ys[1122]), .RECT2_WIDTH(rectangle2_widths[1122]), .RECT2_HEIGHT(rectangle2_heights[1122]), .RECT2_WEIGHT(rectangle2_weights[1122]), .RECT3_X(rectangle3_xs[1122]), .RECT3_Y(rectangle3_ys[1122]), .RECT3_WIDTH(rectangle3_widths[1122]), .RECT3_HEIGHT(rectangle3_heights[1122]), .RECT3_WEIGHT(rectangle3_weights[1122]), .FEAT_THRES(feature_thresholds[1122]), .FEAT_ABOVE(feature_aboves[1122]), .FEAT_BELOW(feature_belows[1122])) ac1122(.scan_win(scan_win1122), .scan_win_std_dev(scan_win_std_dev[1122]), .feature_accum(feature_accums[1122]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1123]), .RECT1_Y(rectangle1_ys[1123]), .RECT1_WIDTH(rectangle1_widths[1123]), .RECT1_HEIGHT(rectangle1_heights[1123]), .RECT1_WEIGHT(rectangle1_weights[1123]), .RECT2_X(rectangle2_xs[1123]), .RECT2_Y(rectangle2_ys[1123]), .RECT2_WIDTH(rectangle2_widths[1123]), .RECT2_HEIGHT(rectangle2_heights[1123]), .RECT2_WEIGHT(rectangle2_weights[1123]), .RECT3_X(rectangle3_xs[1123]), .RECT3_Y(rectangle3_ys[1123]), .RECT3_WIDTH(rectangle3_widths[1123]), .RECT3_HEIGHT(rectangle3_heights[1123]), .RECT3_WEIGHT(rectangle3_weights[1123]), .FEAT_THRES(feature_thresholds[1123]), .FEAT_ABOVE(feature_aboves[1123]), .FEAT_BELOW(feature_belows[1123])) ac1123(.scan_win(scan_win1123), .scan_win_std_dev(scan_win_std_dev[1123]), .feature_accum(feature_accums[1123]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1124]), .RECT1_Y(rectangle1_ys[1124]), .RECT1_WIDTH(rectangle1_widths[1124]), .RECT1_HEIGHT(rectangle1_heights[1124]), .RECT1_WEIGHT(rectangle1_weights[1124]), .RECT2_X(rectangle2_xs[1124]), .RECT2_Y(rectangle2_ys[1124]), .RECT2_WIDTH(rectangle2_widths[1124]), .RECT2_HEIGHT(rectangle2_heights[1124]), .RECT2_WEIGHT(rectangle2_weights[1124]), .RECT3_X(rectangle3_xs[1124]), .RECT3_Y(rectangle3_ys[1124]), .RECT3_WIDTH(rectangle3_widths[1124]), .RECT3_HEIGHT(rectangle3_heights[1124]), .RECT3_WEIGHT(rectangle3_weights[1124]), .FEAT_THRES(feature_thresholds[1124]), .FEAT_ABOVE(feature_aboves[1124]), .FEAT_BELOW(feature_belows[1124])) ac1124(.scan_win(scan_win1124), .scan_win_std_dev(scan_win_std_dev[1124]), .feature_accum(feature_accums[1124]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1125]), .RECT1_Y(rectangle1_ys[1125]), .RECT1_WIDTH(rectangle1_widths[1125]), .RECT1_HEIGHT(rectangle1_heights[1125]), .RECT1_WEIGHT(rectangle1_weights[1125]), .RECT2_X(rectangle2_xs[1125]), .RECT2_Y(rectangle2_ys[1125]), .RECT2_WIDTH(rectangle2_widths[1125]), .RECT2_HEIGHT(rectangle2_heights[1125]), .RECT2_WEIGHT(rectangle2_weights[1125]), .RECT3_X(rectangle3_xs[1125]), .RECT3_Y(rectangle3_ys[1125]), .RECT3_WIDTH(rectangle3_widths[1125]), .RECT3_HEIGHT(rectangle3_heights[1125]), .RECT3_WEIGHT(rectangle3_weights[1125]), .FEAT_THRES(feature_thresholds[1125]), .FEAT_ABOVE(feature_aboves[1125]), .FEAT_BELOW(feature_belows[1125])) ac1125(.scan_win(scan_win1125), .scan_win_std_dev(scan_win_std_dev[1125]), .feature_accum(feature_accums[1125]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1126]), .RECT1_Y(rectangle1_ys[1126]), .RECT1_WIDTH(rectangle1_widths[1126]), .RECT1_HEIGHT(rectangle1_heights[1126]), .RECT1_WEIGHT(rectangle1_weights[1126]), .RECT2_X(rectangle2_xs[1126]), .RECT2_Y(rectangle2_ys[1126]), .RECT2_WIDTH(rectangle2_widths[1126]), .RECT2_HEIGHT(rectangle2_heights[1126]), .RECT2_WEIGHT(rectangle2_weights[1126]), .RECT3_X(rectangle3_xs[1126]), .RECT3_Y(rectangle3_ys[1126]), .RECT3_WIDTH(rectangle3_widths[1126]), .RECT3_HEIGHT(rectangle3_heights[1126]), .RECT3_WEIGHT(rectangle3_weights[1126]), .FEAT_THRES(feature_thresholds[1126]), .FEAT_ABOVE(feature_aboves[1126]), .FEAT_BELOW(feature_belows[1126])) ac1126(.scan_win(scan_win1126), .scan_win_std_dev(scan_win_std_dev[1126]), .feature_accum(feature_accums[1126]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1127]), .RECT1_Y(rectangle1_ys[1127]), .RECT1_WIDTH(rectangle1_widths[1127]), .RECT1_HEIGHT(rectangle1_heights[1127]), .RECT1_WEIGHT(rectangle1_weights[1127]), .RECT2_X(rectangle2_xs[1127]), .RECT2_Y(rectangle2_ys[1127]), .RECT2_WIDTH(rectangle2_widths[1127]), .RECT2_HEIGHT(rectangle2_heights[1127]), .RECT2_WEIGHT(rectangle2_weights[1127]), .RECT3_X(rectangle3_xs[1127]), .RECT3_Y(rectangle3_ys[1127]), .RECT3_WIDTH(rectangle3_widths[1127]), .RECT3_HEIGHT(rectangle3_heights[1127]), .RECT3_WEIGHT(rectangle3_weights[1127]), .FEAT_THRES(feature_thresholds[1127]), .FEAT_ABOVE(feature_aboves[1127]), .FEAT_BELOW(feature_belows[1127])) ac1127(.scan_win(scan_win1127), .scan_win_std_dev(scan_win_std_dev[1127]), .feature_accum(feature_accums[1127]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1128]), .RECT1_Y(rectangle1_ys[1128]), .RECT1_WIDTH(rectangle1_widths[1128]), .RECT1_HEIGHT(rectangle1_heights[1128]), .RECT1_WEIGHT(rectangle1_weights[1128]), .RECT2_X(rectangle2_xs[1128]), .RECT2_Y(rectangle2_ys[1128]), .RECT2_WIDTH(rectangle2_widths[1128]), .RECT2_HEIGHT(rectangle2_heights[1128]), .RECT2_WEIGHT(rectangle2_weights[1128]), .RECT3_X(rectangle3_xs[1128]), .RECT3_Y(rectangle3_ys[1128]), .RECT3_WIDTH(rectangle3_widths[1128]), .RECT3_HEIGHT(rectangle3_heights[1128]), .RECT3_WEIGHT(rectangle3_weights[1128]), .FEAT_THRES(feature_thresholds[1128]), .FEAT_ABOVE(feature_aboves[1128]), .FEAT_BELOW(feature_belows[1128])) ac1128(.scan_win(scan_win1128), .scan_win_std_dev(scan_win_std_dev[1128]), .feature_accum(feature_accums[1128]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1129]), .RECT1_Y(rectangle1_ys[1129]), .RECT1_WIDTH(rectangle1_widths[1129]), .RECT1_HEIGHT(rectangle1_heights[1129]), .RECT1_WEIGHT(rectangle1_weights[1129]), .RECT2_X(rectangle2_xs[1129]), .RECT2_Y(rectangle2_ys[1129]), .RECT2_WIDTH(rectangle2_widths[1129]), .RECT2_HEIGHT(rectangle2_heights[1129]), .RECT2_WEIGHT(rectangle2_weights[1129]), .RECT3_X(rectangle3_xs[1129]), .RECT3_Y(rectangle3_ys[1129]), .RECT3_WIDTH(rectangle3_widths[1129]), .RECT3_HEIGHT(rectangle3_heights[1129]), .RECT3_WEIGHT(rectangle3_weights[1129]), .FEAT_THRES(feature_thresholds[1129]), .FEAT_ABOVE(feature_aboves[1129]), .FEAT_BELOW(feature_belows[1129])) ac1129(.scan_win(scan_win1129), .scan_win_std_dev(scan_win_std_dev[1129]), .feature_accum(feature_accums[1129]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1130]), .RECT1_Y(rectangle1_ys[1130]), .RECT1_WIDTH(rectangle1_widths[1130]), .RECT1_HEIGHT(rectangle1_heights[1130]), .RECT1_WEIGHT(rectangle1_weights[1130]), .RECT2_X(rectangle2_xs[1130]), .RECT2_Y(rectangle2_ys[1130]), .RECT2_WIDTH(rectangle2_widths[1130]), .RECT2_HEIGHT(rectangle2_heights[1130]), .RECT2_WEIGHT(rectangle2_weights[1130]), .RECT3_X(rectangle3_xs[1130]), .RECT3_Y(rectangle3_ys[1130]), .RECT3_WIDTH(rectangle3_widths[1130]), .RECT3_HEIGHT(rectangle3_heights[1130]), .RECT3_WEIGHT(rectangle3_weights[1130]), .FEAT_THRES(feature_thresholds[1130]), .FEAT_ABOVE(feature_aboves[1130]), .FEAT_BELOW(feature_belows[1130])) ac1130(.scan_win(scan_win1130), .scan_win_std_dev(scan_win_std_dev[1130]), .feature_accum(feature_accums[1130]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1131]), .RECT1_Y(rectangle1_ys[1131]), .RECT1_WIDTH(rectangle1_widths[1131]), .RECT1_HEIGHT(rectangle1_heights[1131]), .RECT1_WEIGHT(rectangle1_weights[1131]), .RECT2_X(rectangle2_xs[1131]), .RECT2_Y(rectangle2_ys[1131]), .RECT2_WIDTH(rectangle2_widths[1131]), .RECT2_HEIGHT(rectangle2_heights[1131]), .RECT2_WEIGHT(rectangle2_weights[1131]), .RECT3_X(rectangle3_xs[1131]), .RECT3_Y(rectangle3_ys[1131]), .RECT3_WIDTH(rectangle3_widths[1131]), .RECT3_HEIGHT(rectangle3_heights[1131]), .RECT3_WEIGHT(rectangle3_weights[1131]), .FEAT_THRES(feature_thresholds[1131]), .FEAT_ABOVE(feature_aboves[1131]), .FEAT_BELOW(feature_belows[1131])) ac1131(.scan_win(scan_win1131), .scan_win_std_dev(scan_win_std_dev[1131]), .feature_accum(feature_accums[1131]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1132]), .RECT1_Y(rectangle1_ys[1132]), .RECT1_WIDTH(rectangle1_widths[1132]), .RECT1_HEIGHT(rectangle1_heights[1132]), .RECT1_WEIGHT(rectangle1_weights[1132]), .RECT2_X(rectangle2_xs[1132]), .RECT2_Y(rectangle2_ys[1132]), .RECT2_WIDTH(rectangle2_widths[1132]), .RECT2_HEIGHT(rectangle2_heights[1132]), .RECT2_WEIGHT(rectangle2_weights[1132]), .RECT3_X(rectangle3_xs[1132]), .RECT3_Y(rectangle3_ys[1132]), .RECT3_WIDTH(rectangle3_widths[1132]), .RECT3_HEIGHT(rectangle3_heights[1132]), .RECT3_WEIGHT(rectangle3_weights[1132]), .FEAT_THRES(feature_thresholds[1132]), .FEAT_ABOVE(feature_aboves[1132]), .FEAT_BELOW(feature_belows[1132])) ac1132(.scan_win(scan_win1132), .scan_win_std_dev(scan_win_std_dev[1132]), .feature_accum(feature_accums[1132]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1133]), .RECT1_Y(rectangle1_ys[1133]), .RECT1_WIDTH(rectangle1_widths[1133]), .RECT1_HEIGHT(rectangle1_heights[1133]), .RECT1_WEIGHT(rectangle1_weights[1133]), .RECT2_X(rectangle2_xs[1133]), .RECT2_Y(rectangle2_ys[1133]), .RECT2_WIDTH(rectangle2_widths[1133]), .RECT2_HEIGHT(rectangle2_heights[1133]), .RECT2_WEIGHT(rectangle2_weights[1133]), .RECT3_X(rectangle3_xs[1133]), .RECT3_Y(rectangle3_ys[1133]), .RECT3_WIDTH(rectangle3_widths[1133]), .RECT3_HEIGHT(rectangle3_heights[1133]), .RECT3_WEIGHT(rectangle3_weights[1133]), .FEAT_THRES(feature_thresholds[1133]), .FEAT_ABOVE(feature_aboves[1133]), .FEAT_BELOW(feature_belows[1133])) ac1133(.scan_win(scan_win1133), .scan_win_std_dev(scan_win_std_dev[1133]), .feature_accum(feature_accums[1133]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1134]), .RECT1_Y(rectangle1_ys[1134]), .RECT1_WIDTH(rectangle1_widths[1134]), .RECT1_HEIGHT(rectangle1_heights[1134]), .RECT1_WEIGHT(rectangle1_weights[1134]), .RECT2_X(rectangle2_xs[1134]), .RECT2_Y(rectangle2_ys[1134]), .RECT2_WIDTH(rectangle2_widths[1134]), .RECT2_HEIGHT(rectangle2_heights[1134]), .RECT2_WEIGHT(rectangle2_weights[1134]), .RECT3_X(rectangle3_xs[1134]), .RECT3_Y(rectangle3_ys[1134]), .RECT3_WIDTH(rectangle3_widths[1134]), .RECT3_HEIGHT(rectangle3_heights[1134]), .RECT3_WEIGHT(rectangle3_weights[1134]), .FEAT_THRES(feature_thresholds[1134]), .FEAT_ABOVE(feature_aboves[1134]), .FEAT_BELOW(feature_belows[1134])) ac1134(.scan_win(scan_win1134), .scan_win_std_dev(scan_win_std_dev[1134]), .feature_accum(feature_accums[1134]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1135]), .RECT1_Y(rectangle1_ys[1135]), .RECT1_WIDTH(rectangle1_widths[1135]), .RECT1_HEIGHT(rectangle1_heights[1135]), .RECT1_WEIGHT(rectangle1_weights[1135]), .RECT2_X(rectangle2_xs[1135]), .RECT2_Y(rectangle2_ys[1135]), .RECT2_WIDTH(rectangle2_widths[1135]), .RECT2_HEIGHT(rectangle2_heights[1135]), .RECT2_WEIGHT(rectangle2_weights[1135]), .RECT3_X(rectangle3_xs[1135]), .RECT3_Y(rectangle3_ys[1135]), .RECT3_WIDTH(rectangle3_widths[1135]), .RECT3_HEIGHT(rectangle3_heights[1135]), .RECT3_WEIGHT(rectangle3_weights[1135]), .FEAT_THRES(feature_thresholds[1135]), .FEAT_ABOVE(feature_aboves[1135]), .FEAT_BELOW(feature_belows[1135])) ac1135(.scan_win(scan_win1135), .scan_win_std_dev(scan_win_std_dev[1135]), .feature_accum(feature_accums[1135]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1136]), .RECT1_Y(rectangle1_ys[1136]), .RECT1_WIDTH(rectangle1_widths[1136]), .RECT1_HEIGHT(rectangle1_heights[1136]), .RECT1_WEIGHT(rectangle1_weights[1136]), .RECT2_X(rectangle2_xs[1136]), .RECT2_Y(rectangle2_ys[1136]), .RECT2_WIDTH(rectangle2_widths[1136]), .RECT2_HEIGHT(rectangle2_heights[1136]), .RECT2_WEIGHT(rectangle2_weights[1136]), .RECT3_X(rectangle3_xs[1136]), .RECT3_Y(rectangle3_ys[1136]), .RECT3_WIDTH(rectangle3_widths[1136]), .RECT3_HEIGHT(rectangle3_heights[1136]), .RECT3_WEIGHT(rectangle3_weights[1136]), .FEAT_THRES(feature_thresholds[1136]), .FEAT_ABOVE(feature_aboves[1136]), .FEAT_BELOW(feature_belows[1136])) ac1136(.scan_win(scan_win1136), .scan_win_std_dev(scan_win_std_dev[1136]), .feature_accum(feature_accums[1136]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1137]), .RECT1_Y(rectangle1_ys[1137]), .RECT1_WIDTH(rectangle1_widths[1137]), .RECT1_HEIGHT(rectangle1_heights[1137]), .RECT1_WEIGHT(rectangle1_weights[1137]), .RECT2_X(rectangle2_xs[1137]), .RECT2_Y(rectangle2_ys[1137]), .RECT2_WIDTH(rectangle2_widths[1137]), .RECT2_HEIGHT(rectangle2_heights[1137]), .RECT2_WEIGHT(rectangle2_weights[1137]), .RECT3_X(rectangle3_xs[1137]), .RECT3_Y(rectangle3_ys[1137]), .RECT3_WIDTH(rectangle3_widths[1137]), .RECT3_HEIGHT(rectangle3_heights[1137]), .RECT3_WEIGHT(rectangle3_weights[1137]), .FEAT_THRES(feature_thresholds[1137]), .FEAT_ABOVE(feature_aboves[1137]), .FEAT_BELOW(feature_belows[1137])) ac1137(.scan_win(scan_win1137), .scan_win_std_dev(scan_win_std_dev[1137]), .feature_accum(feature_accums[1137]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1138]), .RECT1_Y(rectangle1_ys[1138]), .RECT1_WIDTH(rectangle1_widths[1138]), .RECT1_HEIGHT(rectangle1_heights[1138]), .RECT1_WEIGHT(rectangle1_weights[1138]), .RECT2_X(rectangle2_xs[1138]), .RECT2_Y(rectangle2_ys[1138]), .RECT2_WIDTH(rectangle2_widths[1138]), .RECT2_HEIGHT(rectangle2_heights[1138]), .RECT2_WEIGHT(rectangle2_weights[1138]), .RECT3_X(rectangle3_xs[1138]), .RECT3_Y(rectangle3_ys[1138]), .RECT3_WIDTH(rectangle3_widths[1138]), .RECT3_HEIGHT(rectangle3_heights[1138]), .RECT3_WEIGHT(rectangle3_weights[1138]), .FEAT_THRES(feature_thresholds[1138]), .FEAT_ABOVE(feature_aboves[1138]), .FEAT_BELOW(feature_belows[1138])) ac1138(.scan_win(scan_win1138), .scan_win_std_dev(scan_win_std_dev[1138]), .feature_accum(feature_accums[1138]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1139]), .RECT1_Y(rectangle1_ys[1139]), .RECT1_WIDTH(rectangle1_widths[1139]), .RECT1_HEIGHT(rectangle1_heights[1139]), .RECT1_WEIGHT(rectangle1_weights[1139]), .RECT2_X(rectangle2_xs[1139]), .RECT2_Y(rectangle2_ys[1139]), .RECT2_WIDTH(rectangle2_widths[1139]), .RECT2_HEIGHT(rectangle2_heights[1139]), .RECT2_WEIGHT(rectangle2_weights[1139]), .RECT3_X(rectangle3_xs[1139]), .RECT3_Y(rectangle3_ys[1139]), .RECT3_WIDTH(rectangle3_widths[1139]), .RECT3_HEIGHT(rectangle3_heights[1139]), .RECT3_WEIGHT(rectangle3_weights[1139]), .FEAT_THRES(feature_thresholds[1139]), .FEAT_ABOVE(feature_aboves[1139]), .FEAT_BELOW(feature_belows[1139])) ac1139(.scan_win(scan_win1139), .scan_win_std_dev(scan_win_std_dev[1139]), .feature_accum(feature_accums[1139]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1140]), .RECT1_Y(rectangle1_ys[1140]), .RECT1_WIDTH(rectangle1_widths[1140]), .RECT1_HEIGHT(rectangle1_heights[1140]), .RECT1_WEIGHT(rectangle1_weights[1140]), .RECT2_X(rectangle2_xs[1140]), .RECT2_Y(rectangle2_ys[1140]), .RECT2_WIDTH(rectangle2_widths[1140]), .RECT2_HEIGHT(rectangle2_heights[1140]), .RECT2_WEIGHT(rectangle2_weights[1140]), .RECT3_X(rectangle3_xs[1140]), .RECT3_Y(rectangle3_ys[1140]), .RECT3_WIDTH(rectangle3_widths[1140]), .RECT3_HEIGHT(rectangle3_heights[1140]), .RECT3_WEIGHT(rectangle3_weights[1140]), .FEAT_THRES(feature_thresholds[1140]), .FEAT_ABOVE(feature_aboves[1140]), .FEAT_BELOW(feature_belows[1140])) ac1140(.scan_win(scan_win1140), .scan_win_std_dev(scan_win_std_dev[1140]), .feature_accum(feature_accums[1140]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1141]), .RECT1_Y(rectangle1_ys[1141]), .RECT1_WIDTH(rectangle1_widths[1141]), .RECT1_HEIGHT(rectangle1_heights[1141]), .RECT1_WEIGHT(rectangle1_weights[1141]), .RECT2_X(rectangle2_xs[1141]), .RECT2_Y(rectangle2_ys[1141]), .RECT2_WIDTH(rectangle2_widths[1141]), .RECT2_HEIGHT(rectangle2_heights[1141]), .RECT2_WEIGHT(rectangle2_weights[1141]), .RECT3_X(rectangle3_xs[1141]), .RECT3_Y(rectangle3_ys[1141]), .RECT3_WIDTH(rectangle3_widths[1141]), .RECT3_HEIGHT(rectangle3_heights[1141]), .RECT3_WEIGHT(rectangle3_weights[1141]), .FEAT_THRES(feature_thresholds[1141]), .FEAT_ABOVE(feature_aboves[1141]), .FEAT_BELOW(feature_belows[1141])) ac1141(.scan_win(scan_win1141), .scan_win_std_dev(scan_win_std_dev[1141]), .feature_accum(feature_accums[1141]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1142]), .RECT1_Y(rectangle1_ys[1142]), .RECT1_WIDTH(rectangle1_widths[1142]), .RECT1_HEIGHT(rectangle1_heights[1142]), .RECT1_WEIGHT(rectangle1_weights[1142]), .RECT2_X(rectangle2_xs[1142]), .RECT2_Y(rectangle2_ys[1142]), .RECT2_WIDTH(rectangle2_widths[1142]), .RECT2_HEIGHT(rectangle2_heights[1142]), .RECT2_WEIGHT(rectangle2_weights[1142]), .RECT3_X(rectangle3_xs[1142]), .RECT3_Y(rectangle3_ys[1142]), .RECT3_WIDTH(rectangle3_widths[1142]), .RECT3_HEIGHT(rectangle3_heights[1142]), .RECT3_WEIGHT(rectangle3_weights[1142]), .FEAT_THRES(feature_thresholds[1142]), .FEAT_ABOVE(feature_aboves[1142]), .FEAT_BELOW(feature_belows[1142])) ac1142(.scan_win(scan_win1142), .scan_win_std_dev(scan_win_std_dev[1142]), .feature_accum(feature_accums[1142]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1143]), .RECT1_Y(rectangle1_ys[1143]), .RECT1_WIDTH(rectangle1_widths[1143]), .RECT1_HEIGHT(rectangle1_heights[1143]), .RECT1_WEIGHT(rectangle1_weights[1143]), .RECT2_X(rectangle2_xs[1143]), .RECT2_Y(rectangle2_ys[1143]), .RECT2_WIDTH(rectangle2_widths[1143]), .RECT2_HEIGHT(rectangle2_heights[1143]), .RECT2_WEIGHT(rectangle2_weights[1143]), .RECT3_X(rectangle3_xs[1143]), .RECT3_Y(rectangle3_ys[1143]), .RECT3_WIDTH(rectangle3_widths[1143]), .RECT3_HEIGHT(rectangle3_heights[1143]), .RECT3_WEIGHT(rectangle3_weights[1143]), .FEAT_THRES(feature_thresholds[1143]), .FEAT_ABOVE(feature_aboves[1143]), .FEAT_BELOW(feature_belows[1143])) ac1143(.scan_win(scan_win1143), .scan_win_std_dev(scan_win_std_dev[1143]), .feature_accum(feature_accums[1143]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1144]), .RECT1_Y(rectangle1_ys[1144]), .RECT1_WIDTH(rectangle1_widths[1144]), .RECT1_HEIGHT(rectangle1_heights[1144]), .RECT1_WEIGHT(rectangle1_weights[1144]), .RECT2_X(rectangle2_xs[1144]), .RECT2_Y(rectangle2_ys[1144]), .RECT2_WIDTH(rectangle2_widths[1144]), .RECT2_HEIGHT(rectangle2_heights[1144]), .RECT2_WEIGHT(rectangle2_weights[1144]), .RECT3_X(rectangle3_xs[1144]), .RECT3_Y(rectangle3_ys[1144]), .RECT3_WIDTH(rectangle3_widths[1144]), .RECT3_HEIGHT(rectangle3_heights[1144]), .RECT3_WEIGHT(rectangle3_weights[1144]), .FEAT_THRES(feature_thresholds[1144]), .FEAT_ABOVE(feature_aboves[1144]), .FEAT_BELOW(feature_belows[1144])) ac1144(.scan_win(scan_win1144), .scan_win_std_dev(scan_win_std_dev[1144]), .feature_accum(feature_accums[1144]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1145]), .RECT1_Y(rectangle1_ys[1145]), .RECT1_WIDTH(rectangle1_widths[1145]), .RECT1_HEIGHT(rectangle1_heights[1145]), .RECT1_WEIGHT(rectangle1_weights[1145]), .RECT2_X(rectangle2_xs[1145]), .RECT2_Y(rectangle2_ys[1145]), .RECT2_WIDTH(rectangle2_widths[1145]), .RECT2_HEIGHT(rectangle2_heights[1145]), .RECT2_WEIGHT(rectangle2_weights[1145]), .RECT3_X(rectangle3_xs[1145]), .RECT3_Y(rectangle3_ys[1145]), .RECT3_WIDTH(rectangle3_widths[1145]), .RECT3_HEIGHT(rectangle3_heights[1145]), .RECT3_WEIGHT(rectangle3_weights[1145]), .FEAT_THRES(feature_thresholds[1145]), .FEAT_ABOVE(feature_aboves[1145]), .FEAT_BELOW(feature_belows[1145])) ac1145(.scan_win(scan_win1145), .scan_win_std_dev(scan_win_std_dev[1145]), .feature_accum(feature_accums[1145]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1146]), .RECT1_Y(rectangle1_ys[1146]), .RECT1_WIDTH(rectangle1_widths[1146]), .RECT1_HEIGHT(rectangle1_heights[1146]), .RECT1_WEIGHT(rectangle1_weights[1146]), .RECT2_X(rectangle2_xs[1146]), .RECT2_Y(rectangle2_ys[1146]), .RECT2_WIDTH(rectangle2_widths[1146]), .RECT2_HEIGHT(rectangle2_heights[1146]), .RECT2_WEIGHT(rectangle2_weights[1146]), .RECT3_X(rectangle3_xs[1146]), .RECT3_Y(rectangle3_ys[1146]), .RECT3_WIDTH(rectangle3_widths[1146]), .RECT3_HEIGHT(rectangle3_heights[1146]), .RECT3_WEIGHT(rectangle3_weights[1146]), .FEAT_THRES(feature_thresholds[1146]), .FEAT_ABOVE(feature_aboves[1146]), .FEAT_BELOW(feature_belows[1146])) ac1146(.scan_win(scan_win1146), .scan_win_std_dev(scan_win_std_dev[1146]), .feature_accum(feature_accums[1146]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1147]), .RECT1_Y(rectangle1_ys[1147]), .RECT1_WIDTH(rectangle1_widths[1147]), .RECT1_HEIGHT(rectangle1_heights[1147]), .RECT1_WEIGHT(rectangle1_weights[1147]), .RECT2_X(rectangle2_xs[1147]), .RECT2_Y(rectangle2_ys[1147]), .RECT2_WIDTH(rectangle2_widths[1147]), .RECT2_HEIGHT(rectangle2_heights[1147]), .RECT2_WEIGHT(rectangle2_weights[1147]), .RECT3_X(rectangle3_xs[1147]), .RECT3_Y(rectangle3_ys[1147]), .RECT3_WIDTH(rectangle3_widths[1147]), .RECT3_HEIGHT(rectangle3_heights[1147]), .RECT3_WEIGHT(rectangle3_weights[1147]), .FEAT_THRES(feature_thresholds[1147]), .FEAT_ABOVE(feature_aboves[1147]), .FEAT_BELOW(feature_belows[1147])) ac1147(.scan_win(scan_win1147), .scan_win_std_dev(scan_win_std_dev[1147]), .feature_accum(feature_accums[1147]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1148]), .RECT1_Y(rectangle1_ys[1148]), .RECT1_WIDTH(rectangle1_widths[1148]), .RECT1_HEIGHT(rectangle1_heights[1148]), .RECT1_WEIGHT(rectangle1_weights[1148]), .RECT2_X(rectangle2_xs[1148]), .RECT2_Y(rectangle2_ys[1148]), .RECT2_WIDTH(rectangle2_widths[1148]), .RECT2_HEIGHT(rectangle2_heights[1148]), .RECT2_WEIGHT(rectangle2_weights[1148]), .RECT3_X(rectangle3_xs[1148]), .RECT3_Y(rectangle3_ys[1148]), .RECT3_WIDTH(rectangle3_widths[1148]), .RECT3_HEIGHT(rectangle3_heights[1148]), .RECT3_WEIGHT(rectangle3_weights[1148]), .FEAT_THRES(feature_thresholds[1148]), .FEAT_ABOVE(feature_aboves[1148]), .FEAT_BELOW(feature_belows[1148])) ac1148(.scan_win(scan_win1148), .scan_win_std_dev(scan_win_std_dev[1148]), .feature_accum(feature_accums[1148]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1149]), .RECT1_Y(rectangle1_ys[1149]), .RECT1_WIDTH(rectangle1_widths[1149]), .RECT1_HEIGHT(rectangle1_heights[1149]), .RECT1_WEIGHT(rectangle1_weights[1149]), .RECT2_X(rectangle2_xs[1149]), .RECT2_Y(rectangle2_ys[1149]), .RECT2_WIDTH(rectangle2_widths[1149]), .RECT2_HEIGHT(rectangle2_heights[1149]), .RECT2_WEIGHT(rectangle2_weights[1149]), .RECT3_X(rectangle3_xs[1149]), .RECT3_Y(rectangle3_ys[1149]), .RECT3_WIDTH(rectangle3_widths[1149]), .RECT3_HEIGHT(rectangle3_heights[1149]), .RECT3_WEIGHT(rectangle3_weights[1149]), .FEAT_THRES(feature_thresholds[1149]), .FEAT_ABOVE(feature_aboves[1149]), .FEAT_BELOW(feature_belows[1149])) ac1149(.scan_win(scan_win1149), .scan_win_std_dev(scan_win_std_dev[1149]), .feature_accum(feature_accums[1149]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1150]), .RECT1_Y(rectangle1_ys[1150]), .RECT1_WIDTH(rectangle1_widths[1150]), .RECT1_HEIGHT(rectangle1_heights[1150]), .RECT1_WEIGHT(rectangle1_weights[1150]), .RECT2_X(rectangle2_xs[1150]), .RECT2_Y(rectangle2_ys[1150]), .RECT2_WIDTH(rectangle2_widths[1150]), .RECT2_HEIGHT(rectangle2_heights[1150]), .RECT2_WEIGHT(rectangle2_weights[1150]), .RECT3_X(rectangle3_xs[1150]), .RECT3_Y(rectangle3_ys[1150]), .RECT3_WIDTH(rectangle3_widths[1150]), .RECT3_HEIGHT(rectangle3_heights[1150]), .RECT3_WEIGHT(rectangle3_weights[1150]), .FEAT_THRES(feature_thresholds[1150]), .FEAT_ABOVE(feature_aboves[1150]), .FEAT_BELOW(feature_belows[1150])) ac1150(.scan_win(scan_win1150), .scan_win_std_dev(scan_win_std_dev[1150]), .feature_accum(feature_accums[1150]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1151]), .RECT1_Y(rectangle1_ys[1151]), .RECT1_WIDTH(rectangle1_widths[1151]), .RECT1_HEIGHT(rectangle1_heights[1151]), .RECT1_WEIGHT(rectangle1_weights[1151]), .RECT2_X(rectangle2_xs[1151]), .RECT2_Y(rectangle2_ys[1151]), .RECT2_WIDTH(rectangle2_widths[1151]), .RECT2_HEIGHT(rectangle2_heights[1151]), .RECT2_WEIGHT(rectangle2_weights[1151]), .RECT3_X(rectangle3_xs[1151]), .RECT3_Y(rectangle3_ys[1151]), .RECT3_WIDTH(rectangle3_widths[1151]), .RECT3_HEIGHT(rectangle3_heights[1151]), .RECT3_WEIGHT(rectangle3_weights[1151]), .FEAT_THRES(feature_thresholds[1151]), .FEAT_ABOVE(feature_aboves[1151]), .FEAT_BELOW(feature_belows[1151])) ac1151(.scan_win(scan_win1151), .scan_win_std_dev(scan_win_std_dev[1151]), .feature_accum(feature_accums[1151]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1152]), .RECT1_Y(rectangle1_ys[1152]), .RECT1_WIDTH(rectangle1_widths[1152]), .RECT1_HEIGHT(rectangle1_heights[1152]), .RECT1_WEIGHT(rectangle1_weights[1152]), .RECT2_X(rectangle2_xs[1152]), .RECT2_Y(rectangle2_ys[1152]), .RECT2_WIDTH(rectangle2_widths[1152]), .RECT2_HEIGHT(rectangle2_heights[1152]), .RECT2_WEIGHT(rectangle2_weights[1152]), .RECT3_X(rectangle3_xs[1152]), .RECT3_Y(rectangle3_ys[1152]), .RECT3_WIDTH(rectangle3_widths[1152]), .RECT3_HEIGHT(rectangle3_heights[1152]), .RECT3_WEIGHT(rectangle3_weights[1152]), .FEAT_THRES(feature_thresholds[1152]), .FEAT_ABOVE(feature_aboves[1152]), .FEAT_BELOW(feature_belows[1152])) ac1152(.scan_win(scan_win1152), .scan_win_std_dev(scan_win_std_dev[1152]), .feature_accum(feature_accums[1152]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1153]), .RECT1_Y(rectangle1_ys[1153]), .RECT1_WIDTH(rectangle1_widths[1153]), .RECT1_HEIGHT(rectangle1_heights[1153]), .RECT1_WEIGHT(rectangle1_weights[1153]), .RECT2_X(rectangle2_xs[1153]), .RECT2_Y(rectangle2_ys[1153]), .RECT2_WIDTH(rectangle2_widths[1153]), .RECT2_HEIGHT(rectangle2_heights[1153]), .RECT2_WEIGHT(rectangle2_weights[1153]), .RECT3_X(rectangle3_xs[1153]), .RECT3_Y(rectangle3_ys[1153]), .RECT3_WIDTH(rectangle3_widths[1153]), .RECT3_HEIGHT(rectangle3_heights[1153]), .RECT3_WEIGHT(rectangle3_weights[1153]), .FEAT_THRES(feature_thresholds[1153]), .FEAT_ABOVE(feature_aboves[1153]), .FEAT_BELOW(feature_belows[1153])) ac1153(.scan_win(scan_win1153), .scan_win_std_dev(scan_win_std_dev[1153]), .feature_accum(feature_accums[1153]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1154]), .RECT1_Y(rectangle1_ys[1154]), .RECT1_WIDTH(rectangle1_widths[1154]), .RECT1_HEIGHT(rectangle1_heights[1154]), .RECT1_WEIGHT(rectangle1_weights[1154]), .RECT2_X(rectangle2_xs[1154]), .RECT2_Y(rectangle2_ys[1154]), .RECT2_WIDTH(rectangle2_widths[1154]), .RECT2_HEIGHT(rectangle2_heights[1154]), .RECT2_WEIGHT(rectangle2_weights[1154]), .RECT3_X(rectangle3_xs[1154]), .RECT3_Y(rectangle3_ys[1154]), .RECT3_WIDTH(rectangle3_widths[1154]), .RECT3_HEIGHT(rectangle3_heights[1154]), .RECT3_WEIGHT(rectangle3_weights[1154]), .FEAT_THRES(feature_thresholds[1154]), .FEAT_ABOVE(feature_aboves[1154]), .FEAT_BELOW(feature_belows[1154])) ac1154(.scan_win(scan_win1154), .scan_win_std_dev(scan_win_std_dev[1154]), .feature_accum(feature_accums[1154]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1155]), .RECT1_Y(rectangle1_ys[1155]), .RECT1_WIDTH(rectangle1_widths[1155]), .RECT1_HEIGHT(rectangle1_heights[1155]), .RECT1_WEIGHT(rectangle1_weights[1155]), .RECT2_X(rectangle2_xs[1155]), .RECT2_Y(rectangle2_ys[1155]), .RECT2_WIDTH(rectangle2_widths[1155]), .RECT2_HEIGHT(rectangle2_heights[1155]), .RECT2_WEIGHT(rectangle2_weights[1155]), .RECT3_X(rectangle3_xs[1155]), .RECT3_Y(rectangle3_ys[1155]), .RECT3_WIDTH(rectangle3_widths[1155]), .RECT3_HEIGHT(rectangle3_heights[1155]), .RECT3_WEIGHT(rectangle3_weights[1155]), .FEAT_THRES(feature_thresholds[1155]), .FEAT_ABOVE(feature_aboves[1155]), .FEAT_BELOW(feature_belows[1155])) ac1155(.scan_win(scan_win1155), .scan_win_std_dev(scan_win_std_dev[1155]), .feature_accum(feature_accums[1155]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1156]), .RECT1_Y(rectangle1_ys[1156]), .RECT1_WIDTH(rectangle1_widths[1156]), .RECT1_HEIGHT(rectangle1_heights[1156]), .RECT1_WEIGHT(rectangle1_weights[1156]), .RECT2_X(rectangle2_xs[1156]), .RECT2_Y(rectangle2_ys[1156]), .RECT2_WIDTH(rectangle2_widths[1156]), .RECT2_HEIGHT(rectangle2_heights[1156]), .RECT2_WEIGHT(rectangle2_weights[1156]), .RECT3_X(rectangle3_xs[1156]), .RECT3_Y(rectangle3_ys[1156]), .RECT3_WIDTH(rectangle3_widths[1156]), .RECT3_HEIGHT(rectangle3_heights[1156]), .RECT3_WEIGHT(rectangle3_weights[1156]), .FEAT_THRES(feature_thresholds[1156]), .FEAT_ABOVE(feature_aboves[1156]), .FEAT_BELOW(feature_belows[1156])) ac1156(.scan_win(scan_win1156), .scan_win_std_dev(scan_win_std_dev[1156]), .feature_accum(feature_accums[1156]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1157]), .RECT1_Y(rectangle1_ys[1157]), .RECT1_WIDTH(rectangle1_widths[1157]), .RECT1_HEIGHT(rectangle1_heights[1157]), .RECT1_WEIGHT(rectangle1_weights[1157]), .RECT2_X(rectangle2_xs[1157]), .RECT2_Y(rectangle2_ys[1157]), .RECT2_WIDTH(rectangle2_widths[1157]), .RECT2_HEIGHT(rectangle2_heights[1157]), .RECT2_WEIGHT(rectangle2_weights[1157]), .RECT3_X(rectangle3_xs[1157]), .RECT3_Y(rectangle3_ys[1157]), .RECT3_WIDTH(rectangle3_widths[1157]), .RECT3_HEIGHT(rectangle3_heights[1157]), .RECT3_WEIGHT(rectangle3_weights[1157]), .FEAT_THRES(feature_thresholds[1157]), .FEAT_ABOVE(feature_aboves[1157]), .FEAT_BELOW(feature_belows[1157])) ac1157(.scan_win(scan_win1157), .scan_win_std_dev(scan_win_std_dev[1157]), .feature_accum(feature_accums[1157]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1158]), .RECT1_Y(rectangle1_ys[1158]), .RECT1_WIDTH(rectangle1_widths[1158]), .RECT1_HEIGHT(rectangle1_heights[1158]), .RECT1_WEIGHT(rectangle1_weights[1158]), .RECT2_X(rectangle2_xs[1158]), .RECT2_Y(rectangle2_ys[1158]), .RECT2_WIDTH(rectangle2_widths[1158]), .RECT2_HEIGHT(rectangle2_heights[1158]), .RECT2_WEIGHT(rectangle2_weights[1158]), .RECT3_X(rectangle3_xs[1158]), .RECT3_Y(rectangle3_ys[1158]), .RECT3_WIDTH(rectangle3_widths[1158]), .RECT3_HEIGHT(rectangle3_heights[1158]), .RECT3_WEIGHT(rectangle3_weights[1158]), .FEAT_THRES(feature_thresholds[1158]), .FEAT_ABOVE(feature_aboves[1158]), .FEAT_BELOW(feature_belows[1158])) ac1158(.scan_win(scan_win1158), .scan_win_std_dev(scan_win_std_dev[1158]), .feature_accum(feature_accums[1158]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1159]), .RECT1_Y(rectangle1_ys[1159]), .RECT1_WIDTH(rectangle1_widths[1159]), .RECT1_HEIGHT(rectangle1_heights[1159]), .RECT1_WEIGHT(rectangle1_weights[1159]), .RECT2_X(rectangle2_xs[1159]), .RECT2_Y(rectangle2_ys[1159]), .RECT2_WIDTH(rectangle2_widths[1159]), .RECT2_HEIGHT(rectangle2_heights[1159]), .RECT2_WEIGHT(rectangle2_weights[1159]), .RECT3_X(rectangle3_xs[1159]), .RECT3_Y(rectangle3_ys[1159]), .RECT3_WIDTH(rectangle3_widths[1159]), .RECT3_HEIGHT(rectangle3_heights[1159]), .RECT3_WEIGHT(rectangle3_weights[1159]), .FEAT_THRES(feature_thresholds[1159]), .FEAT_ABOVE(feature_aboves[1159]), .FEAT_BELOW(feature_belows[1159])) ac1159(.scan_win(scan_win1159), .scan_win_std_dev(scan_win_std_dev[1159]), .feature_accum(feature_accums[1159]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1160]), .RECT1_Y(rectangle1_ys[1160]), .RECT1_WIDTH(rectangle1_widths[1160]), .RECT1_HEIGHT(rectangle1_heights[1160]), .RECT1_WEIGHT(rectangle1_weights[1160]), .RECT2_X(rectangle2_xs[1160]), .RECT2_Y(rectangle2_ys[1160]), .RECT2_WIDTH(rectangle2_widths[1160]), .RECT2_HEIGHT(rectangle2_heights[1160]), .RECT2_WEIGHT(rectangle2_weights[1160]), .RECT3_X(rectangle3_xs[1160]), .RECT3_Y(rectangle3_ys[1160]), .RECT3_WIDTH(rectangle3_widths[1160]), .RECT3_HEIGHT(rectangle3_heights[1160]), .RECT3_WEIGHT(rectangle3_weights[1160]), .FEAT_THRES(feature_thresholds[1160]), .FEAT_ABOVE(feature_aboves[1160]), .FEAT_BELOW(feature_belows[1160])) ac1160(.scan_win(scan_win1160), .scan_win_std_dev(scan_win_std_dev[1160]), .feature_accum(feature_accums[1160]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1161]), .RECT1_Y(rectangle1_ys[1161]), .RECT1_WIDTH(rectangle1_widths[1161]), .RECT1_HEIGHT(rectangle1_heights[1161]), .RECT1_WEIGHT(rectangle1_weights[1161]), .RECT2_X(rectangle2_xs[1161]), .RECT2_Y(rectangle2_ys[1161]), .RECT2_WIDTH(rectangle2_widths[1161]), .RECT2_HEIGHT(rectangle2_heights[1161]), .RECT2_WEIGHT(rectangle2_weights[1161]), .RECT3_X(rectangle3_xs[1161]), .RECT3_Y(rectangle3_ys[1161]), .RECT3_WIDTH(rectangle3_widths[1161]), .RECT3_HEIGHT(rectangle3_heights[1161]), .RECT3_WEIGHT(rectangle3_weights[1161]), .FEAT_THRES(feature_thresholds[1161]), .FEAT_ABOVE(feature_aboves[1161]), .FEAT_BELOW(feature_belows[1161])) ac1161(.scan_win(scan_win1161), .scan_win_std_dev(scan_win_std_dev[1161]), .feature_accum(feature_accums[1161]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1162]), .RECT1_Y(rectangle1_ys[1162]), .RECT1_WIDTH(rectangle1_widths[1162]), .RECT1_HEIGHT(rectangle1_heights[1162]), .RECT1_WEIGHT(rectangle1_weights[1162]), .RECT2_X(rectangle2_xs[1162]), .RECT2_Y(rectangle2_ys[1162]), .RECT2_WIDTH(rectangle2_widths[1162]), .RECT2_HEIGHT(rectangle2_heights[1162]), .RECT2_WEIGHT(rectangle2_weights[1162]), .RECT3_X(rectangle3_xs[1162]), .RECT3_Y(rectangle3_ys[1162]), .RECT3_WIDTH(rectangle3_widths[1162]), .RECT3_HEIGHT(rectangle3_heights[1162]), .RECT3_WEIGHT(rectangle3_weights[1162]), .FEAT_THRES(feature_thresholds[1162]), .FEAT_ABOVE(feature_aboves[1162]), .FEAT_BELOW(feature_belows[1162])) ac1162(.scan_win(scan_win1162), .scan_win_std_dev(scan_win_std_dev[1162]), .feature_accum(feature_accums[1162]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1163]), .RECT1_Y(rectangle1_ys[1163]), .RECT1_WIDTH(rectangle1_widths[1163]), .RECT1_HEIGHT(rectangle1_heights[1163]), .RECT1_WEIGHT(rectangle1_weights[1163]), .RECT2_X(rectangle2_xs[1163]), .RECT2_Y(rectangle2_ys[1163]), .RECT2_WIDTH(rectangle2_widths[1163]), .RECT2_HEIGHT(rectangle2_heights[1163]), .RECT2_WEIGHT(rectangle2_weights[1163]), .RECT3_X(rectangle3_xs[1163]), .RECT3_Y(rectangle3_ys[1163]), .RECT3_WIDTH(rectangle3_widths[1163]), .RECT3_HEIGHT(rectangle3_heights[1163]), .RECT3_WEIGHT(rectangle3_weights[1163]), .FEAT_THRES(feature_thresholds[1163]), .FEAT_ABOVE(feature_aboves[1163]), .FEAT_BELOW(feature_belows[1163])) ac1163(.scan_win(scan_win1163), .scan_win_std_dev(scan_win_std_dev[1163]), .feature_accum(feature_accums[1163]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1164]), .RECT1_Y(rectangle1_ys[1164]), .RECT1_WIDTH(rectangle1_widths[1164]), .RECT1_HEIGHT(rectangle1_heights[1164]), .RECT1_WEIGHT(rectangle1_weights[1164]), .RECT2_X(rectangle2_xs[1164]), .RECT2_Y(rectangle2_ys[1164]), .RECT2_WIDTH(rectangle2_widths[1164]), .RECT2_HEIGHT(rectangle2_heights[1164]), .RECT2_WEIGHT(rectangle2_weights[1164]), .RECT3_X(rectangle3_xs[1164]), .RECT3_Y(rectangle3_ys[1164]), .RECT3_WIDTH(rectangle3_widths[1164]), .RECT3_HEIGHT(rectangle3_heights[1164]), .RECT3_WEIGHT(rectangle3_weights[1164]), .FEAT_THRES(feature_thresholds[1164]), .FEAT_ABOVE(feature_aboves[1164]), .FEAT_BELOW(feature_belows[1164])) ac1164(.scan_win(scan_win1164), .scan_win_std_dev(scan_win_std_dev[1164]), .feature_accum(feature_accums[1164]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1165]), .RECT1_Y(rectangle1_ys[1165]), .RECT1_WIDTH(rectangle1_widths[1165]), .RECT1_HEIGHT(rectangle1_heights[1165]), .RECT1_WEIGHT(rectangle1_weights[1165]), .RECT2_X(rectangle2_xs[1165]), .RECT2_Y(rectangle2_ys[1165]), .RECT2_WIDTH(rectangle2_widths[1165]), .RECT2_HEIGHT(rectangle2_heights[1165]), .RECT2_WEIGHT(rectangle2_weights[1165]), .RECT3_X(rectangle3_xs[1165]), .RECT3_Y(rectangle3_ys[1165]), .RECT3_WIDTH(rectangle3_widths[1165]), .RECT3_HEIGHT(rectangle3_heights[1165]), .RECT3_WEIGHT(rectangle3_weights[1165]), .FEAT_THRES(feature_thresholds[1165]), .FEAT_ABOVE(feature_aboves[1165]), .FEAT_BELOW(feature_belows[1165])) ac1165(.scan_win(scan_win1165), .scan_win_std_dev(scan_win_std_dev[1165]), .feature_accum(feature_accums[1165]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1166]), .RECT1_Y(rectangle1_ys[1166]), .RECT1_WIDTH(rectangle1_widths[1166]), .RECT1_HEIGHT(rectangle1_heights[1166]), .RECT1_WEIGHT(rectangle1_weights[1166]), .RECT2_X(rectangle2_xs[1166]), .RECT2_Y(rectangle2_ys[1166]), .RECT2_WIDTH(rectangle2_widths[1166]), .RECT2_HEIGHT(rectangle2_heights[1166]), .RECT2_WEIGHT(rectangle2_weights[1166]), .RECT3_X(rectangle3_xs[1166]), .RECT3_Y(rectangle3_ys[1166]), .RECT3_WIDTH(rectangle3_widths[1166]), .RECT3_HEIGHT(rectangle3_heights[1166]), .RECT3_WEIGHT(rectangle3_weights[1166]), .FEAT_THRES(feature_thresholds[1166]), .FEAT_ABOVE(feature_aboves[1166]), .FEAT_BELOW(feature_belows[1166])) ac1166(.scan_win(scan_win1166), .scan_win_std_dev(scan_win_std_dev[1166]), .feature_accum(feature_accums[1166]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1167]), .RECT1_Y(rectangle1_ys[1167]), .RECT1_WIDTH(rectangle1_widths[1167]), .RECT1_HEIGHT(rectangle1_heights[1167]), .RECT1_WEIGHT(rectangle1_weights[1167]), .RECT2_X(rectangle2_xs[1167]), .RECT2_Y(rectangle2_ys[1167]), .RECT2_WIDTH(rectangle2_widths[1167]), .RECT2_HEIGHT(rectangle2_heights[1167]), .RECT2_WEIGHT(rectangle2_weights[1167]), .RECT3_X(rectangle3_xs[1167]), .RECT3_Y(rectangle3_ys[1167]), .RECT3_WIDTH(rectangle3_widths[1167]), .RECT3_HEIGHT(rectangle3_heights[1167]), .RECT3_WEIGHT(rectangle3_weights[1167]), .FEAT_THRES(feature_thresholds[1167]), .FEAT_ABOVE(feature_aboves[1167]), .FEAT_BELOW(feature_belows[1167])) ac1167(.scan_win(scan_win1167), .scan_win_std_dev(scan_win_std_dev[1167]), .feature_accum(feature_accums[1167]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1168]), .RECT1_Y(rectangle1_ys[1168]), .RECT1_WIDTH(rectangle1_widths[1168]), .RECT1_HEIGHT(rectangle1_heights[1168]), .RECT1_WEIGHT(rectangle1_weights[1168]), .RECT2_X(rectangle2_xs[1168]), .RECT2_Y(rectangle2_ys[1168]), .RECT2_WIDTH(rectangle2_widths[1168]), .RECT2_HEIGHT(rectangle2_heights[1168]), .RECT2_WEIGHT(rectangle2_weights[1168]), .RECT3_X(rectangle3_xs[1168]), .RECT3_Y(rectangle3_ys[1168]), .RECT3_WIDTH(rectangle3_widths[1168]), .RECT3_HEIGHT(rectangle3_heights[1168]), .RECT3_WEIGHT(rectangle3_weights[1168]), .FEAT_THRES(feature_thresholds[1168]), .FEAT_ABOVE(feature_aboves[1168]), .FEAT_BELOW(feature_belows[1168])) ac1168(.scan_win(scan_win1168), .scan_win_std_dev(scan_win_std_dev[1168]), .feature_accum(feature_accums[1168]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1169]), .RECT1_Y(rectangle1_ys[1169]), .RECT1_WIDTH(rectangle1_widths[1169]), .RECT1_HEIGHT(rectangle1_heights[1169]), .RECT1_WEIGHT(rectangle1_weights[1169]), .RECT2_X(rectangle2_xs[1169]), .RECT2_Y(rectangle2_ys[1169]), .RECT2_WIDTH(rectangle2_widths[1169]), .RECT2_HEIGHT(rectangle2_heights[1169]), .RECT2_WEIGHT(rectangle2_weights[1169]), .RECT3_X(rectangle3_xs[1169]), .RECT3_Y(rectangle3_ys[1169]), .RECT3_WIDTH(rectangle3_widths[1169]), .RECT3_HEIGHT(rectangle3_heights[1169]), .RECT3_WEIGHT(rectangle3_weights[1169]), .FEAT_THRES(feature_thresholds[1169]), .FEAT_ABOVE(feature_aboves[1169]), .FEAT_BELOW(feature_belows[1169])) ac1169(.scan_win(scan_win1169), .scan_win_std_dev(scan_win_std_dev[1169]), .feature_accum(feature_accums[1169]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1170]), .RECT1_Y(rectangle1_ys[1170]), .RECT1_WIDTH(rectangle1_widths[1170]), .RECT1_HEIGHT(rectangle1_heights[1170]), .RECT1_WEIGHT(rectangle1_weights[1170]), .RECT2_X(rectangle2_xs[1170]), .RECT2_Y(rectangle2_ys[1170]), .RECT2_WIDTH(rectangle2_widths[1170]), .RECT2_HEIGHT(rectangle2_heights[1170]), .RECT2_WEIGHT(rectangle2_weights[1170]), .RECT3_X(rectangle3_xs[1170]), .RECT3_Y(rectangle3_ys[1170]), .RECT3_WIDTH(rectangle3_widths[1170]), .RECT3_HEIGHT(rectangle3_heights[1170]), .RECT3_WEIGHT(rectangle3_weights[1170]), .FEAT_THRES(feature_thresholds[1170]), .FEAT_ABOVE(feature_aboves[1170]), .FEAT_BELOW(feature_belows[1170])) ac1170(.scan_win(scan_win1170), .scan_win_std_dev(scan_win_std_dev[1170]), .feature_accum(feature_accums[1170]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1171]), .RECT1_Y(rectangle1_ys[1171]), .RECT1_WIDTH(rectangle1_widths[1171]), .RECT1_HEIGHT(rectangle1_heights[1171]), .RECT1_WEIGHT(rectangle1_weights[1171]), .RECT2_X(rectangle2_xs[1171]), .RECT2_Y(rectangle2_ys[1171]), .RECT2_WIDTH(rectangle2_widths[1171]), .RECT2_HEIGHT(rectangle2_heights[1171]), .RECT2_WEIGHT(rectangle2_weights[1171]), .RECT3_X(rectangle3_xs[1171]), .RECT3_Y(rectangle3_ys[1171]), .RECT3_WIDTH(rectangle3_widths[1171]), .RECT3_HEIGHT(rectangle3_heights[1171]), .RECT3_WEIGHT(rectangle3_weights[1171]), .FEAT_THRES(feature_thresholds[1171]), .FEAT_ABOVE(feature_aboves[1171]), .FEAT_BELOW(feature_belows[1171])) ac1171(.scan_win(scan_win1171), .scan_win_std_dev(scan_win_std_dev[1171]), .feature_accum(feature_accums[1171]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1172]), .RECT1_Y(rectangle1_ys[1172]), .RECT1_WIDTH(rectangle1_widths[1172]), .RECT1_HEIGHT(rectangle1_heights[1172]), .RECT1_WEIGHT(rectangle1_weights[1172]), .RECT2_X(rectangle2_xs[1172]), .RECT2_Y(rectangle2_ys[1172]), .RECT2_WIDTH(rectangle2_widths[1172]), .RECT2_HEIGHT(rectangle2_heights[1172]), .RECT2_WEIGHT(rectangle2_weights[1172]), .RECT3_X(rectangle3_xs[1172]), .RECT3_Y(rectangle3_ys[1172]), .RECT3_WIDTH(rectangle3_widths[1172]), .RECT3_HEIGHT(rectangle3_heights[1172]), .RECT3_WEIGHT(rectangle3_weights[1172]), .FEAT_THRES(feature_thresholds[1172]), .FEAT_ABOVE(feature_aboves[1172]), .FEAT_BELOW(feature_belows[1172])) ac1172(.scan_win(scan_win1172), .scan_win_std_dev(scan_win_std_dev[1172]), .feature_accum(feature_accums[1172]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1173]), .RECT1_Y(rectangle1_ys[1173]), .RECT1_WIDTH(rectangle1_widths[1173]), .RECT1_HEIGHT(rectangle1_heights[1173]), .RECT1_WEIGHT(rectangle1_weights[1173]), .RECT2_X(rectangle2_xs[1173]), .RECT2_Y(rectangle2_ys[1173]), .RECT2_WIDTH(rectangle2_widths[1173]), .RECT2_HEIGHT(rectangle2_heights[1173]), .RECT2_WEIGHT(rectangle2_weights[1173]), .RECT3_X(rectangle3_xs[1173]), .RECT3_Y(rectangle3_ys[1173]), .RECT3_WIDTH(rectangle3_widths[1173]), .RECT3_HEIGHT(rectangle3_heights[1173]), .RECT3_WEIGHT(rectangle3_weights[1173]), .FEAT_THRES(feature_thresholds[1173]), .FEAT_ABOVE(feature_aboves[1173]), .FEAT_BELOW(feature_belows[1173])) ac1173(.scan_win(scan_win1173), .scan_win_std_dev(scan_win_std_dev[1173]), .feature_accum(feature_accums[1173]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1174]), .RECT1_Y(rectangle1_ys[1174]), .RECT1_WIDTH(rectangle1_widths[1174]), .RECT1_HEIGHT(rectangle1_heights[1174]), .RECT1_WEIGHT(rectangle1_weights[1174]), .RECT2_X(rectangle2_xs[1174]), .RECT2_Y(rectangle2_ys[1174]), .RECT2_WIDTH(rectangle2_widths[1174]), .RECT2_HEIGHT(rectangle2_heights[1174]), .RECT2_WEIGHT(rectangle2_weights[1174]), .RECT3_X(rectangle3_xs[1174]), .RECT3_Y(rectangle3_ys[1174]), .RECT3_WIDTH(rectangle3_widths[1174]), .RECT3_HEIGHT(rectangle3_heights[1174]), .RECT3_WEIGHT(rectangle3_weights[1174]), .FEAT_THRES(feature_thresholds[1174]), .FEAT_ABOVE(feature_aboves[1174]), .FEAT_BELOW(feature_belows[1174])) ac1174(.scan_win(scan_win1174), .scan_win_std_dev(scan_win_std_dev[1174]), .feature_accum(feature_accums[1174]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1175]), .RECT1_Y(rectangle1_ys[1175]), .RECT1_WIDTH(rectangle1_widths[1175]), .RECT1_HEIGHT(rectangle1_heights[1175]), .RECT1_WEIGHT(rectangle1_weights[1175]), .RECT2_X(rectangle2_xs[1175]), .RECT2_Y(rectangle2_ys[1175]), .RECT2_WIDTH(rectangle2_widths[1175]), .RECT2_HEIGHT(rectangle2_heights[1175]), .RECT2_WEIGHT(rectangle2_weights[1175]), .RECT3_X(rectangle3_xs[1175]), .RECT3_Y(rectangle3_ys[1175]), .RECT3_WIDTH(rectangle3_widths[1175]), .RECT3_HEIGHT(rectangle3_heights[1175]), .RECT3_WEIGHT(rectangle3_weights[1175]), .FEAT_THRES(feature_thresholds[1175]), .FEAT_ABOVE(feature_aboves[1175]), .FEAT_BELOW(feature_belows[1175])) ac1175(.scan_win(scan_win1175), .scan_win_std_dev(scan_win_std_dev[1175]), .feature_accum(feature_accums[1175]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1176]), .RECT1_Y(rectangle1_ys[1176]), .RECT1_WIDTH(rectangle1_widths[1176]), .RECT1_HEIGHT(rectangle1_heights[1176]), .RECT1_WEIGHT(rectangle1_weights[1176]), .RECT2_X(rectangle2_xs[1176]), .RECT2_Y(rectangle2_ys[1176]), .RECT2_WIDTH(rectangle2_widths[1176]), .RECT2_HEIGHT(rectangle2_heights[1176]), .RECT2_WEIGHT(rectangle2_weights[1176]), .RECT3_X(rectangle3_xs[1176]), .RECT3_Y(rectangle3_ys[1176]), .RECT3_WIDTH(rectangle3_widths[1176]), .RECT3_HEIGHT(rectangle3_heights[1176]), .RECT3_WEIGHT(rectangle3_weights[1176]), .FEAT_THRES(feature_thresholds[1176]), .FEAT_ABOVE(feature_aboves[1176]), .FEAT_BELOW(feature_belows[1176])) ac1176(.scan_win(scan_win1176), .scan_win_std_dev(scan_win_std_dev[1176]), .feature_accum(feature_accums[1176]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1177]), .RECT1_Y(rectangle1_ys[1177]), .RECT1_WIDTH(rectangle1_widths[1177]), .RECT1_HEIGHT(rectangle1_heights[1177]), .RECT1_WEIGHT(rectangle1_weights[1177]), .RECT2_X(rectangle2_xs[1177]), .RECT2_Y(rectangle2_ys[1177]), .RECT2_WIDTH(rectangle2_widths[1177]), .RECT2_HEIGHT(rectangle2_heights[1177]), .RECT2_WEIGHT(rectangle2_weights[1177]), .RECT3_X(rectangle3_xs[1177]), .RECT3_Y(rectangle3_ys[1177]), .RECT3_WIDTH(rectangle3_widths[1177]), .RECT3_HEIGHT(rectangle3_heights[1177]), .RECT3_WEIGHT(rectangle3_weights[1177]), .FEAT_THRES(feature_thresholds[1177]), .FEAT_ABOVE(feature_aboves[1177]), .FEAT_BELOW(feature_belows[1177])) ac1177(.scan_win(scan_win1177), .scan_win_std_dev(scan_win_std_dev[1177]), .feature_accum(feature_accums[1177]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1178]), .RECT1_Y(rectangle1_ys[1178]), .RECT1_WIDTH(rectangle1_widths[1178]), .RECT1_HEIGHT(rectangle1_heights[1178]), .RECT1_WEIGHT(rectangle1_weights[1178]), .RECT2_X(rectangle2_xs[1178]), .RECT2_Y(rectangle2_ys[1178]), .RECT2_WIDTH(rectangle2_widths[1178]), .RECT2_HEIGHT(rectangle2_heights[1178]), .RECT2_WEIGHT(rectangle2_weights[1178]), .RECT3_X(rectangle3_xs[1178]), .RECT3_Y(rectangle3_ys[1178]), .RECT3_WIDTH(rectangle3_widths[1178]), .RECT3_HEIGHT(rectangle3_heights[1178]), .RECT3_WEIGHT(rectangle3_weights[1178]), .FEAT_THRES(feature_thresholds[1178]), .FEAT_ABOVE(feature_aboves[1178]), .FEAT_BELOW(feature_belows[1178])) ac1178(.scan_win(scan_win1178), .scan_win_std_dev(scan_win_std_dev[1178]), .feature_accum(feature_accums[1178]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1179]), .RECT1_Y(rectangle1_ys[1179]), .RECT1_WIDTH(rectangle1_widths[1179]), .RECT1_HEIGHT(rectangle1_heights[1179]), .RECT1_WEIGHT(rectangle1_weights[1179]), .RECT2_X(rectangle2_xs[1179]), .RECT2_Y(rectangle2_ys[1179]), .RECT2_WIDTH(rectangle2_widths[1179]), .RECT2_HEIGHT(rectangle2_heights[1179]), .RECT2_WEIGHT(rectangle2_weights[1179]), .RECT3_X(rectangle3_xs[1179]), .RECT3_Y(rectangle3_ys[1179]), .RECT3_WIDTH(rectangle3_widths[1179]), .RECT3_HEIGHT(rectangle3_heights[1179]), .RECT3_WEIGHT(rectangle3_weights[1179]), .FEAT_THRES(feature_thresholds[1179]), .FEAT_ABOVE(feature_aboves[1179]), .FEAT_BELOW(feature_belows[1179])) ac1179(.scan_win(scan_win1179), .scan_win_std_dev(scan_win_std_dev[1179]), .feature_accum(feature_accums[1179]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1180]), .RECT1_Y(rectangle1_ys[1180]), .RECT1_WIDTH(rectangle1_widths[1180]), .RECT1_HEIGHT(rectangle1_heights[1180]), .RECT1_WEIGHT(rectangle1_weights[1180]), .RECT2_X(rectangle2_xs[1180]), .RECT2_Y(rectangle2_ys[1180]), .RECT2_WIDTH(rectangle2_widths[1180]), .RECT2_HEIGHT(rectangle2_heights[1180]), .RECT2_WEIGHT(rectangle2_weights[1180]), .RECT3_X(rectangle3_xs[1180]), .RECT3_Y(rectangle3_ys[1180]), .RECT3_WIDTH(rectangle3_widths[1180]), .RECT3_HEIGHT(rectangle3_heights[1180]), .RECT3_WEIGHT(rectangle3_weights[1180]), .FEAT_THRES(feature_thresholds[1180]), .FEAT_ABOVE(feature_aboves[1180]), .FEAT_BELOW(feature_belows[1180])) ac1180(.scan_win(scan_win1180), .scan_win_std_dev(scan_win_std_dev[1180]), .feature_accum(feature_accums[1180]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1181]), .RECT1_Y(rectangle1_ys[1181]), .RECT1_WIDTH(rectangle1_widths[1181]), .RECT1_HEIGHT(rectangle1_heights[1181]), .RECT1_WEIGHT(rectangle1_weights[1181]), .RECT2_X(rectangle2_xs[1181]), .RECT2_Y(rectangle2_ys[1181]), .RECT2_WIDTH(rectangle2_widths[1181]), .RECT2_HEIGHT(rectangle2_heights[1181]), .RECT2_WEIGHT(rectangle2_weights[1181]), .RECT3_X(rectangle3_xs[1181]), .RECT3_Y(rectangle3_ys[1181]), .RECT3_WIDTH(rectangle3_widths[1181]), .RECT3_HEIGHT(rectangle3_heights[1181]), .RECT3_WEIGHT(rectangle3_weights[1181]), .FEAT_THRES(feature_thresholds[1181]), .FEAT_ABOVE(feature_aboves[1181]), .FEAT_BELOW(feature_belows[1181])) ac1181(.scan_win(scan_win1181), .scan_win_std_dev(scan_win_std_dev[1181]), .feature_accum(feature_accums[1181]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1182]), .RECT1_Y(rectangle1_ys[1182]), .RECT1_WIDTH(rectangle1_widths[1182]), .RECT1_HEIGHT(rectangle1_heights[1182]), .RECT1_WEIGHT(rectangle1_weights[1182]), .RECT2_X(rectangle2_xs[1182]), .RECT2_Y(rectangle2_ys[1182]), .RECT2_WIDTH(rectangle2_widths[1182]), .RECT2_HEIGHT(rectangle2_heights[1182]), .RECT2_WEIGHT(rectangle2_weights[1182]), .RECT3_X(rectangle3_xs[1182]), .RECT3_Y(rectangle3_ys[1182]), .RECT3_WIDTH(rectangle3_widths[1182]), .RECT3_HEIGHT(rectangle3_heights[1182]), .RECT3_WEIGHT(rectangle3_weights[1182]), .FEAT_THRES(feature_thresholds[1182]), .FEAT_ABOVE(feature_aboves[1182]), .FEAT_BELOW(feature_belows[1182])) ac1182(.scan_win(scan_win1182), .scan_win_std_dev(scan_win_std_dev[1182]), .feature_accum(feature_accums[1182]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1183]), .RECT1_Y(rectangle1_ys[1183]), .RECT1_WIDTH(rectangle1_widths[1183]), .RECT1_HEIGHT(rectangle1_heights[1183]), .RECT1_WEIGHT(rectangle1_weights[1183]), .RECT2_X(rectangle2_xs[1183]), .RECT2_Y(rectangle2_ys[1183]), .RECT2_WIDTH(rectangle2_widths[1183]), .RECT2_HEIGHT(rectangle2_heights[1183]), .RECT2_WEIGHT(rectangle2_weights[1183]), .RECT3_X(rectangle3_xs[1183]), .RECT3_Y(rectangle3_ys[1183]), .RECT3_WIDTH(rectangle3_widths[1183]), .RECT3_HEIGHT(rectangle3_heights[1183]), .RECT3_WEIGHT(rectangle3_weights[1183]), .FEAT_THRES(feature_thresholds[1183]), .FEAT_ABOVE(feature_aboves[1183]), .FEAT_BELOW(feature_belows[1183])) ac1183(.scan_win(scan_win1183), .scan_win_std_dev(scan_win_std_dev[1183]), .feature_accum(feature_accums[1183]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1184]), .RECT1_Y(rectangle1_ys[1184]), .RECT1_WIDTH(rectangle1_widths[1184]), .RECT1_HEIGHT(rectangle1_heights[1184]), .RECT1_WEIGHT(rectangle1_weights[1184]), .RECT2_X(rectangle2_xs[1184]), .RECT2_Y(rectangle2_ys[1184]), .RECT2_WIDTH(rectangle2_widths[1184]), .RECT2_HEIGHT(rectangle2_heights[1184]), .RECT2_WEIGHT(rectangle2_weights[1184]), .RECT3_X(rectangle3_xs[1184]), .RECT3_Y(rectangle3_ys[1184]), .RECT3_WIDTH(rectangle3_widths[1184]), .RECT3_HEIGHT(rectangle3_heights[1184]), .RECT3_WEIGHT(rectangle3_weights[1184]), .FEAT_THRES(feature_thresholds[1184]), .FEAT_ABOVE(feature_aboves[1184]), .FEAT_BELOW(feature_belows[1184])) ac1184(.scan_win(scan_win1184), .scan_win_std_dev(scan_win_std_dev[1184]), .feature_accum(feature_accums[1184]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1185]), .RECT1_Y(rectangle1_ys[1185]), .RECT1_WIDTH(rectangle1_widths[1185]), .RECT1_HEIGHT(rectangle1_heights[1185]), .RECT1_WEIGHT(rectangle1_weights[1185]), .RECT2_X(rectangle2_xs[1185]), .RECT2_Y(rectangle2_ys[1185]), .RECT2_WIDTH(rectangle2_widths[1185]), .RECT2_HEIGHT(rectangle2_heights[1185]), .RECT2_WEIGHT(rectangle2_weights[1185]), .RECT3_X(rectangle3_xs[1185]), .RECT3_Y(rectangle3_ys[1185]), .RECT3_WIDTH(rectangle3_widths[1185]), .RECT3_HEIGHT(rectangle3_heights[1185]), .RECT3_WEIGHT(rectangle3_weights[1185]), .FEAT_THRES(feature_thresholds[1185]), .FEAT_ABOVE(feature_aboves[1185]), .FEAT_BELOW(feature_belows[1185])) ac1185(.scan_win(scan_win1185), .scan_win_std_dev(scan_win_std_dev[1185]), .feature_accum(feature_accums[1185]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1186]), .RECT1_Y(rectangle1_ys[1186]), .RECT1_WIDTH(rectangle1_widths[1186]), .RECT1_HEIGHT(rectangle1_heights[1186]), .RECT1_WEIGHT(rectangle1_weights[1186]), .RECT2_X(rectangle2_xs[1186]), .RECT2_Y(rectangle2_ys[1186]), .RECT2_WIDTH(rectangle2_widths[1186]), .RECT2_HEIGHT(rectangle2_heights[1186]), .RECT2_WEIGHT(rectangle2_weights[1186]), .RECT3_X(rectangle3_xs[1186]), .RECT3_Y(rectangle3_ys[1186]), .RECT3_WIDTH(rectangle3_widths[1186]), .RECT3_HEIGHT(rectangle3_heights[1186]), .RECT3_WEIGHT(rectangle3_weights[1186]), .FEAT_THRES(feature_thresholds[1186]), .FEAT_ABOVE(feature_aboves[1186]), .FEAT_BELOW(feature_belows[1186])) ac1186(.scan_win(scan_win1186), .scan_win_std_dev(scan_win_std_dev[1186]), .feature_accum(feature_accums[1186]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1187]), .RECT1_Y(rectangle1_ys[1187]), .RECT1_WIDTH(rectangle1_widths[1187]), .RECT1_HEIGHT(rectangle1_heights[1187]), .RECT1_WEIGHT(rectangle1_weights[1187]), .RECT2_X(rectangle2_xs[1187]), .RECT2_Y(rectangle2_ys[1187]), .RECT2_WIDTH(rectangle2_widths[1187]), .RECT2_HEIGHT(rectangle2_heights[1187]), .RECT2_WEIGHT(rectangle2_weights[1187]), .RECT3_X(rectangle3_xs[1187]), .RECT3_Y(rectangle3_ys[1187]), .RECT3_WIDTH(rectangle3_widths[1187]), .RECT3_HEIGHT(rectangle3_heights[1187]), .RECT3_WEIGHT(rectangle3_weights[1187]), .FEAT_THRES(feature_thresholds[1187]), .FEAT_ABOVE(feature_aboves[1187]), .FEAT_BELOW(feature_belows[1187])) ac1187(.scan_win(scan_win1187), .scan_win_std_dev(scan_win_std_dev[1187]), .feature_accum(feature_accums[1187]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1188]), .RECT1_Y(rectangle1_ys[1188]), .RECT1_WIDTH(rectangle1_widths[1188]), .RECT1_HEIGHT(rectangle1_heights[1188]), .RECT1_WEIGHT(rectangle1_weights[1188]), .RECT2_X(rectangle2_xs[1188]), .RECT2_Y(rectangle2_ys[1188]), .RECT2_WIDTH(rectangle2_widths[1188]), .RECT2_HEIGHT(rectangle2_heights[1188]), .RECT2_WEIGHT(rectangle2_weights[1188]), .RECT3_X(rectangle3_xs[1188]), .RECT3_Y(rectangle3_ys[1188]), .RECT3_WIDTH(rectangle3_widths[1188]), .RECT3_HEIGHT(rectangle3_heights[1188]), .RECT3_WEIGHT(rectangle3_weights[1188]), .FEAT_THRES(feature_thresholds[1188]), .FEAT_ABOVE(feature_aboves[1188]), .FEAT_BELOW(feature_belows[1188])) ac1188(.scan_win(scan_win1188), .scan_win_std_dev(scan_win_std_dev[1188]), .feature_accum(feature_accums[1188]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1189]), .RECT1_Y(rectangle1_ys[1189]), .RECT1_WIDTH(rectangle1_widths[1189]), .RECT1_HEIGHT(rectangle1_heights[1189]), .RECT1_WEIGHT(rectangle1_weights[1189]), .RECT2_X(rectangle2_xs[1189]), .RECT2_Y(rectangle2_ys[1189]), .RECT2_WIDTH(rectangle2_widths[1189]), .RECT2_HEIGHT(rectangle2_heights[1189]), .RECT2_WEIGHT(rectangle2_weights[1189]), .RECT3_X(rectangle3_xs[1189]), .RECT3_Y(rectangle3_ys[1189]), .RECT3_WIDTH(rectangle3_widths[1189]), .RECT3_HEIGHT(rectangle3_heights[1189]), .RECT3_WEIGHT(rectangle3_weights[1189]), .FEAT_THRES(feature_thresholds[1189]), .FEAT_ABOVE(feature_aboves[1189]), .FEAT_BELOW(feature_belows[1189])) ac1189(.scan_win(scan_win1189), .scan_win_std_dev(scan_win_std_dev[1189]), .feature_accum(feature_accums[1189]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1190]), .RECT1_Y(rectangle1_ys[1190]), .RECT1_WIDTH(rectangle1_widths[1190]), .RECT1_HEIGHT(rectangle1_heights[1190]), .RECT1_WEIGHT(rectangle1_weights[1190]), .RECT2_X(rectangle2_xs[1190]), .RECT2_Y(rectangle2_ys[1190]), .RECT2_WIDTH(rectangle2_widths[1190]), .RECT2_HEIGHT(rectangle2_heights[1190]), .RECT2_WEIGHT(rectangle2_weights[1190]), .RECT3_X(rectangle3_xs[1190]), .RECT3_Y(rectangle3_ys[1190]), .RECT3_WIDTH(rectangle3_widths[1190]), .RECT3_HEIGHT(rectangle3_heights[1190]), .RECT3_WEIGHT(rectangle3_weights[1190]), .FEAT_THRES(feature_thresholds[1190]), .FEAT_ABOVE(feature_aboves[1190]), .FEAT_BELOW(feature_belows[1190])) ac1190(.scan_win(scan_win1190), .scan_win_std_dev(scan_win_std_dev[1190]), .feature_accum(feature_accums[1190]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1191]), .RECT1_Y(rectangle1_ys[1191]), .RECT1_WIDTH(rectangle1_widths[1191]), .RECT1_HEIGHT(rectangle1_heights[1191]), .RECT1_WEIGHT(rectangle1_weights[1191]), .RECT2_X(rectangle2_xs[1191]), .RECT2_Y(rectangle2_ys[1191]), .RECT2_WIDTH(rectangle2_widths[1191]), .RECT2_HEIGHT(rectangle2_heights[1191]), .RECT2_WEIGHT(rectangle2_weights[1191]), .RECT3_X(rectangle3_xs[1191]), .RECT3_Y(rectangle3_ys[1191]), .RECT3_WIDTH(rectangle3_widths[1191]), .RECT3_HEIGHT(rectangle3_heights[1191]), .RECT3_WEIGHT(rectangle3_weights[1191]), .FEAT_THRES(feature_thresholds[1191]), .FEAT_ABOVE(feature_aboves[1191]), .FEAT_BELOW(feature_belows[1191])) ac1191(.scan_win(scan_win1191), .scan_win_std_dev(scan_win_std_dev[1191]), .feature_accum(feature_accums[1191]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1192]), .RECT1_Y(rectangle1_ys[1192]), .RECT1_WIDTH(rectangle1_widths[1192]), .RECT1_HEIGHT(rectangle1_heights[1192]), .RECT1_WEIGHT(rectangle1_weights[1192]), .RECT2_X(rectangle2_xs[1192]), .RECT2_Y(rectangle2_ys[1192]), .RECT2_WIDTH(rectangle2_widths[1192]), .RECT2_HEIGHT(rectangle2_heights[1192]), .RECT2_WEIGHT(rectangle2_weights[1192]), .RECT3_X(rectangle3_xs[1192]), .RECT3_Y(rectangle3_ys[1192]), .RECT3_WIDTH(rectangle3_widths[1192]), .RECT3_HEIGHT(rectangle3_heights[1192]), .RECT3_WEIGHT(rectangle3_weights[1192]), .FEAT_THRES(feature_thresholds[1192]), .FEAT_ABOVE(feature_aboves[1192]), .FEAT_BELOW(feature_belows[1192])) ac1192(.scan_win(scan_win1192), .scan_win_std_dev(scan_win_std_dev[1192]), .feature_accum(feature_accums[1192]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1193]), .RECT1_Y(rectangle1_ys[1193]), .RECT1_WIDTH(rectangle1_widths[1193]), .RECT1_HEIGHT(rectangle1_heights[1193]), .RECT1_WEIGHT(rectangle1_weights[1193]), .RECT2_X(rectangle2_xs[1193]), .RECT2_Y(rectangle2_ys[1193]), .RECT2_WIDTH(rectangle2_widths[1193]), .RECT2_HEIGHT(rectangle2_heights[1193]), .RECT2_WEIGHT(rectangle2_weights[1193]), .RECT3_X(rectangle3_xs[1193]), .RECT3_Y(rectangle3_ys[1193]), .RECT3_WIDTH(rectangle3_widths[1193]), .RECT3_HEIGHT(rectangle3_heights[1193]), .RECT3_WEIGHT(rectangle3_weights[1193]), .FEAT_THRES(feature_thresholds[1193]), .FEAT_ABOVE(feature_aboves[1193]), .FEAT_BELOW(feature_belows[1193])) ac1193(.scan_win(scan_win1193), .scan_win_std_dev(scan_win_std_dev[1193]), .feature_accum(feature_accums[1193]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1194]), .RECT1_Y(rectangle1_ys[1194]), .RECT1_WIDTH(rectangle1_widths[1194]), .RECT1_HEIGHT(rectangle1_heights[1194]), .RECT1_WEIGHT(rectangle1_weights[1194]), .RECT2_X(rectangle2_xs[1194]), .RECT2_Y(rectangle2_ys[1194]), .RECT2_WIDTH(rectangle2_widths[1194]), .RECT2_HEIGHT(rectangle2_heights[1194]), .RECT2_WEIGHT(rectangle2_weights[1194]), .RECT3_X(rectangle3_xs[1194]), .RECT3_Y(rectangle3_ys[1194]), .RECT3_WIDTH(rectangle3_widths[1194]), .RECT3_HEIGHT(rectangle3_heights[1194]), .RECT3_WEIGHT(rectangle3_weights[1194]), .FEAT_THRES(feature_thresholds[1194]), .FEAT_ABOVE(feature_aboves[1194]), .FEAT_BELOW(feature_belows[1194])) ac1194(.scan_win(scan_win1194), .scan_win_std_dev(scan_win_std_dev[1194]), .feature_accum(feature_accums[1194]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1195]), .RECT1_Y(rectangle1_ys[1195]), .RECT1_WIDTH(rectangle1_widths[1195]), .RECT1_HEIGHT(rectangle1_heights[1195]), .RECT1_WEIGHT(rectangle1_weights[1195]), .RECT2_X(rectangle2_xs[1195]), .RECT2_Y(rectangle2_ys[1195]), .RECT2_WIDTH(rectangle2_widths[1195]), .RECT2_HEIGHT(rectangle2_heights[1195]), .RECT2_WEIGHT(rectangle2_weights[1195]), .RECT3_X(rectangle3_xs[1195]), .RECT3_Y(rectangle3_ys[1195]), .RECT3_WIDTH(rectangle3_widths[1195]), .RECT3_HEIGHT(rectangle3_heights[1195]), .RECT3_WEIGHT(rectangle3_weights[1195]), .FEAT_THRES(feature_thresholds[1195]), .FEAT_ABOVE(feature_aboves[1195]), .FEAT_BELOW(feature_belows[1195])) ac1195(.scan_win(scan_win1195), .scan_win_std_dev(scan_win_std_dev[1195]), .feature_accum(feature_accums[1195]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1196]), .RECT1_Y(rectangle1_ys[1196]), .RECT1_WIDTH(rectangle1_widths[1196]), .RECT1_HEIGHT(rectangle1_heights[1196]), .RECT1_WEIGHT(rectangle1_weights[1196]), .RECT2_X(rectangle2_xs[1196]), .RECT2_Y(rectangle2_ys[1196]), .RECT2_WIDTH(rectangle2_widths[1196]), .RECT2_HEIGHT(rectangle2_heights[1196]), .RECT2_WEIGHT(rectangle2_weights[1196]), .RECT3_X(rectangle3_xs[1196]), .RECT3_Y(rectangle3_ys[1196]), .RECT3_WIDTH(rectangle3_widths[1196]), .RECT3_HEIGHT(rectangle3_heights[1196]), .RECT3_WEIGHT(rectangle3_weights[1196]), .FEAT_THRES(feature_thresholds[1196]), .FEAT_ABOVE(feature_aboves[1196]), .FEAT_BELOW(feature_belows[1196])) ac1196(.scan_win(scan_win1196), .scan_win_std_dev(scan_win_std_dev[1196]), .feature_accum(feature_accums[1196]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1197]), .RECT1_Y(rectangle1_ys[1197]), .RECT1_WIDTH(rectangle1_widths[1197]), .RECT1_HEIGHT(rectangle1_heights[1197]), .RECT1_WEIGHT(rectangle1_weights[1197]), .RECT2_X(rectangle2_xs[1197]), .RECT2_Y(rectangle2_ys[1197]), .RECT2_WIDTH(rectangle2_widths[1197]), .RECT2_HEIGHT(rectangle2_heights[1197]), .RECT2_WEIGHT(rectangle2_weights[1197]), .RECT3_X(rectangle3_xs[1197]), .RECT3_Y(rectangle3_ys[1197]), .RECT3_WIDTH(rectangle3_widths[1197]), .RECT3_HEIGHT(rectangle3_heights[1197]), .RECT3_WEIGHT(rectangle3_weights[1197]), .FEAT_THRES(feature_thresholds[1197]), .FEAT_ABOVE(feature_aboves[1197]), .FEAT_BELOW(feature_belows[1197])) ac1197(.scan_win(scan_win1197), .scan_win_std_dev(scan_win_std_dev[1197]), .feature_accum(feature_accums[1197]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1198]), .RECT1_Y(rectangle1_ys[1198]), .RECT1_WIDTH(rectangle1_widths[1198]), .RECT1_HEIGHT(rectangle1_heights[1198]), .RECT1_WEIGHT(rectangle1_weights[1198]), .RECT2_X(rectangle2_xs[1198]), .RECT2_Y(rectangle2_ys[1198]), .RECT2_WIDTH(rectangle2_widths[1198]), .RECT2_HEIGHT(rectangle2_heights[1198]), .RECT2_WEIGHT(rectangle2_weights[1198]), .RECT3_X(rectangle3_xs[1198]), .RECT3_Y(rectangle3_ys[1198]), .RECT3_WIDTH(rectangle3_widths[1198]), .RECT3_HEIGHT(rectangle3_heights[1198]), .RECT3_WEIGHT(rectangle3_weights[1198]), .FEAT_THRES(feature_thresholds[1198]), .FEAT_ABOVE(feature_aboves[1198]), .FEAT_BELOW(feature_belows[1198])) ac1198(.scan_win(scan_win1198), .scan_win_std_dev(scan_win_std_dev[1198]), .feature_accum(feature_accums[1198]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1199]), .RECT1_Y(rectangle1_ys[1199]), .RECT1_WIDTH(rectangle1_widths[1199]), .RECT1_HEIGHT(rectangle1_heights[1199]), .RECT1_WEIGHT(rectangle1_weights[1199]), .RECT2_X(rectangle2_xs[1199]), .RECT2_Y(rectangle2_ys[1199]), .RECT2_WIDTH(rectangle2_widths[1199]), .RECT2_HEIGHT(rectangle2_heights[1199]), .RECT2_WEIGHT(rectangle2_weights[1199]), .RECT3_X(rectangle3_xs[1199]), .RECT3_Y(rectangle3_ys[1199]), .RECT3_WIDTH(rectangle3_widths[1199]), .RECT3_HEIGHT(rectangle3_heights[1199]), .RECT3_WEIGHT(rectangle3_weights[1199]), .FEAT_THRES(feature_thresholds[1199]), .FEAT_ABOVE(feature_aboves[1199]), .FEAT_BELOW(feature_belows[1199])) ac1199(.scan_win(scan_win1199), .scan_win_std_dev(scan_win_std_dev[1199]), .feature_accum(feature_accums[1199]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1200]), .RECT1_Y(rectangle1_ys[1200]), .RECT1_WIDTH(rectangle1_widths[1200]), .RECT1_HEIGHT(rectangle1_heights[1200]), .RECT1_WEIGHT(rectangle1_weights[1200]), .RECT2_X(rectangle2_xs[1200]), .RECT2_Y(rectangle2_ys[1200]), .RECT2_WIDTH(rectangle2_widths[1200]), .RECT2_HEIGHT(rectangle2_heights[1200]), .RECT2_WEIGHT(rectangle2_weights[1200]), .RECT3_X(rectangle3_xs[1200]), .RECT3_Y(rectangle3_ys[1200]), .RECT3_WIDTH(rectangle3_widths[1200]), .RECT3_HEIGHT(rectangle3_heights[1200]), .RECT3_WEIGHT(rectangle3_weights[1200]), .FEAT_THRES(feature_thresholds[1200]), .FEAT_ABOVE(feature_aboves[1200]), .FEAT_BELOW(feature_belows[1200])) ac1200(.scan_win(scan_win1200), .scan_win_std_dev(scan_win_std_dev[1200]), .feature_accum(feature_accums[1200]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1201]), .RECT1_Y(rectangle1_ys[1201]), .RECT1_WIDTH(rectangle1_widths[1201]), .RECT1_HEIGHT(rectangle1_heights[1201]), .RECT1_WEIGHT(rectangle1_weights[1201]), .RECT2_X(rectangle2_xs[1201]), .RECT2_Y(rectangle2_ys[1201]), .RECT2_WIDTH(rectangle2_widths[1201]), .RECT2_HEIGHT(rectangle2_heights[1201]), .RECT2_WEIGHT(rectangle2_weights[1201]), .RECT3_X(rectangle3_xs[1201]), .RECT3_Y(rectangle3_ys[1201]), .RECT3_WIDTH(rectangle3_widths[1201]), .RECT3_HEIGHT(rectangle3_heights[1201]), .RECT3_WEIGHT(rectangle3_weights[1201]), .FEAT_THRES(feature_thresholds[1201]), .FEAT_ABOVE(feature_aboves[1201]), .FEAT_BELOW(feature_belows[1201])) ac1201(.scan_win(scan_win1201), .scan_win_std_dev(scan_win_std_dev[1201]), .feature_accum(feature_accums[1201]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1202]), .RECT1_Y(rectangle1_ys[1202]), .RECT1_WIDTH(rectangle1_widths[1202]), .RECT1_HEIGHT(rectangle1_heights[1202]), .RECT1_WEIGHT(rectangle1_weights[1202]), .RECT2_X(rectangle2_xs[1202]), .RECT2_Y(rectangle2_ys[1202]), .RECT2_WIDTH(rectangle2_widths[1202]), .RECT2_HEIGHT(rectangle2_heights[1202]), .RECT2_WEIGHT(rectangle2_weights[1202]), .RECT3_X(rectangle3_xs[1202]), .RECT3_Y(rectangle3_ys[1202]), .RECT3_WIDTH(rectangle3_widths[1202]), .RECT3_HEIGHT(rectangle3_heights[1202]), .RECT3_WEIGHT(rectangle3_weights[1202]), .FEAT_THRES(feature_thresholds[1202]), .FEAT_ABOVE(feature_aboves[1202]), .FEAT_BELOW(feature_belows[1202])) ac1202(.scan_win(scan_win1202), .scan_win_std_dev(scan_win_std_dev[1202]), .feature_accum(feature_accums[1202]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1203]), .RECT1_Y(rectangle1_ys[1203]), .RECT1_WIDTH(rectangle1_widths[1203]), .RECT1_HEIGHT(rectangle1_heights[1203]), .RECT1_WEIGHT(rectangle1_weights[1203]), .RECT2_X(rectangle2_xs[1203]), .RECT2_Y(rectangle2_ys[1203]), .RECT2_WIDTH(rectangle2_widths[1203]), .RECT2_HEIGHT(rectangle2_heights[1203]), .RECT2_WEIGHT(rectangle2_weights[1203]), .RECT3_X(rectangle3_xs[1203]), .RECT3_Y(rectangle3_ys[1203]), .RECT3_WIDTH(rectangle3_widths[1203]), .RECT3_HEIGHT(rectangle3_heights[1203]), .RECT3_WEIGHT(rectangle3_weights[1203]), .FEAT_THRES(feature_thresholds[1203]), .FEAT_ABOVE(feature_aboves[1203]), .FEAT_BELOW(feature_belows[1203])) ac1203(.scan_win(scan_win1203), .scan_win_std_dev(scan_win_std_dev[1203]), .feature_accum(feature_accums[1203]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1204]), .RECT1_Y(rectangle1_ys[1204]), .RECT1_WIDTH(rectangle1_widths[1204]), .RECT1_HEIGHT(rectangle1_heights[1204]), .RECT1_WEIGHT(rectangle1_weights[1204]), .RECT2_X(rectangle2_xs[1204]), .RECT2_Y(rectangle2_ys[1204]), .RECT2_WIDTH(rectangle2_widths[1204]), .RECT2_HEIGHT(rectangle2_heights[1204]), .RECT2_WEIGHT(rectangle2_weights[1204]), .RECT3_X(rectangle3_xs[1204]), .RECT3_Y(rectangle3_ys[1204]), .RECT3_WIDTH(rectangle3_widths[1204]), .RECT3_HEIGHT(rectangle3_heights[1204]), .RECT3_WEIGHT(rectangle3_weights[1204]), .FEAT_THRES(feature_thresholds[1204]), .FEAT_ABOVE(feature_aboves[1204]), .FEAT_BELOW(feature_belows[1204])) ac1204(.scan_win(scan_win1204), .scan_win_std_dev(scan_win_std_dev[1204]), .feature_accum(feature_accums[1204]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1205]), .RECT1_Y(rectangle1_ys[1205]), .RECT1_WIDTH(rectangle1_widths[1205]), .RECT1_HEIGHT(rectangle1_heights[1205]), .RECT1_WEIGHT(rectangle1_weights[1205]), .RECT2_X(rectangle2_xs[1205]), .RECT2_Y(rectangle2_ys[1205]), .RECT2_WIDTH(rectangle2_widths[1205]), .RECT2_HEIGHT(rectangle2_heights[1205]), .RECT2_WEIGHT(rectangle2_weights[1205]), .RECT3_X(rectangle3_xs[1205]), .RECT3_Y(rectangle3_ys[1205]), .RECT3_WIDTH(rectangle3_widths[1205]), .RECT3_HEIGHT(rectangle3_heights[1205]), .RECT3_WEIGHT(rectangle3_weights[1205]), .FEAT_THRES(feature_thresholds[1205]), .FEAT_ABOVE(feature_aboves[1205]), .FEAT_BELOW(feature_belows[1205])) ac1205(.scan_win(scan_win1205), .scan_win_std_dev(scan_win_std_dev[1205]), .feature_accum(feature_accums[1205]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1206]), .RECT1_Y(rectangle1_ys[1206]), .RECT1_WIDTH(rectangle1_widths[1206]), .RECT1_HEIGHT(rectangle1_heights[1206]), .RECT1_WEIGHT(rectangle1_weights[1206]), .RECT2_X(rectangle2_xs[1206]), .RECT2_Y(rectangle2_ys[1206]), .RECT2_WIDTH(rectangle2_widths[1206]), .RECT2_HEIGHT(rectangle2_heights[1206]), .RECT2_WEIGHT(rectangle2_weights[1206]), .RECT3_X(rectangle3_xs[1206]), .RECT3_Y(rectangle3_ys[1206]), .RECT3_WIDTH(rectangle3_widths[1206]), .RECT3_HEIGHT(rectangle3_heights[1206]), .RECT3_WEIGHT(rectangle3_weights[1206]), .FEAT_THRES(feature_thresholds[1206]), .FEAT_ABOVE(feature_aboves[1206]), .FEAT_BELOW(feature_belows[1206])) ac1206(.scan_win(scan_win1206), .scan_win_std_dev(scan_win_std_dev[1206]), .feature_accum(feature_accums[1206]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1207]), .RECT1_Y(rectangle1_ys[1207]), .RECT1_WIDTH(rectangle1_widths[1207]), .RECT1_HEIGHT(rectangle1_heights[1207]), .RECT1_WEIGHT(rectangle1_weights[1207]), .RECT2_X(rectangle2_xs[1207]), .RECT2_Y(rectangle2_ys[1207]), .RECT2_WIDTH(rectangle2_widths[1207]), .RECT2_HEIGHT(rectangle2_heights[1207]), .RECT2_WEIGHT(rectangle2_weights[1207]), .RECT3_X(rectangle3_xs[1207]), .RECT3_Y(rectangle3_ys[1207]), .RECT3_WIDTH(rectangle3_widths[1207]), .RECT3_HEIGHT(rectangle3_heights[1207]), .RECT3_WEIGHT(rectangle3_weights[1207]), .FEAT_THRES(feature_thresholds[1207]), .FEAT_ABOVE(feature_aboves[1207]), .FEAT_BELOW(feature_belows[1207])) ac1207(.scan_win(scan_win1207), .scan_win_std_dev(scan_win_std_dev[1207]), .feature_accum(feature_accums[1207]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1208]), .RECT1_Y(rectangle1_ys[1208]), .RECT1_WIDTH(rectangle1_widths[1208]), .RECT1_HEIGHT(rectangle1_heights[1208]), .RECT1_WEIGHT(rectangle1_weights[1208]), .RECT2_X(rectangle2_xs[1208]), .RECT2_Y(rectangle2_ys[1208]), .RECT2_WIDTH(rectangle2_widths[1208]), .RECT2_HEIGHT(rectangle2_heights[1208]), .RECT2_WEIGHT(rectangle2_weights[1208]), .RECT3_X(rectangle3_xs[1208]), .RECT3_Y(rectangle3_ys[1208]), .RECT3_WIDTH(rectangle3_widths[1208]), .RECT3_HEIGHT(rectangle3_heights[1208]), .RECT3_WEIGHT(rectangle3_weights[1208]), .FEAT_THRES(feature_thresholds[1208]), .FEAT_ABOVE(feature_aboves[1208]), .FEAT_BELOW(feature_belows[1208])) ac1208(.scan_win(scan_win1208), .scan_win_std_dev(scan_win_std_dev[1208]), .feature_accum(feature_accums[1208]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1209]), .RECT1_Y(rectangle1_ys[1209]), .RECT1_WIDTH(rectangle1_widths[1209]), .RECT1_HEIGHT(rectangle1_heights[1209]), .RECT1_WEIGHT(rectangle1_weights[1209]), .RECT2_X(rectangle2_xs[1209]), .RECT2_Y(rectangle2_ys[1209]), .RECT2_WIDTH(rectangle2_widths[1209]), .RECT2_HEIGHT(rectangle2_heights[1209]), .RECT2_WEIGHT(rectangle2_weights[1209]), .RECT3_X(rectangle3_xs[1209]), .RECT3_Y(rectangle3_ys[1209]), .RECT3_WIDTH(rectangle3_widths[1209]), .RECT3_HEIGHT(rectangle3_heights[1209]), .RECT3_WEIGHT(rectangle3_weights[1209]), .FEAT_THRES(feature_thresholds[1209]), .FEAT_ABOVE(feature_aboves[1209]), .FEAT_BELOW(feature_belows[1209])) ac1209(.scan_win(scan_win1209), .scan_win_std_dev(scan_win_std_dev[1209]), .feature_accum(feature_accums[1209]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1210]), .RECT1_Y(rectangle1_ys[1210]), .RECT1_WIDTH(rectangle1_widths[1210]), .RECT1_HEIGHT(rectangle1_heights[1210]), .RECT1_WEIGHT(rectangle1_weights[1210]), .RECT2_X(rectangle2_xs[1210]), .RECT2_Y(rectangle2_ys[1210]), .RECT2_WIDTH(rectangle2_widths[1210]), .RECT2_HEIGHT(rectangle2_heights[1210]), .RECT2_WEIGHT(rectangle2_weights[1210]), .RECT3_X(rectangle3_xs[1210]), .RECT3_Y(rectangle3_ys[1210]), .RECT3_WIDTH(rectangle3_widths[1210]), .RECT3_HEIGHT(rectangle3_heights[1210]), .RECT3_WEIGHT(rectangle3_weights[1210]), .FEAT_THRES(feature_thresholds[1210]), .FEAT_ABOVE(feature_aboves[1210]), .FEAT_BELOW(feature_belows[1210])) ac1210(.scan_win(scan_win1210), .scan_win_std_dev(scan_win_std_dev[1210]), .feature_accum(feature_accums[1210]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1211]), .RECT1_Y(rectangle1_ys[1211]), .RECT1_WIDTH(rectangle1_widths[1211]), .RECT1_HEIGHT(rectangle1_heights[1211]), .RECT1_WEIGHT(rectangle1_weights[1211]), .RECT2_X(rectangle2_xs[1211]), .RECT2_Y(rectangle2_ys[1211]), .RECT2_WIDTH(rectangle2_widths[1211]), .RECT2_HEIGHT(rectangle2_heights[1211]), .RECT2_WEIGHT(rectangle2_weights[1211]), .RECT3_X(rectangle3_xs[1211]), .RECT3_Y(rectangle3_ys[1211]), .RECT3_WIDTH(rectangle3_widths[1211]), .RECT3_HEIGHT(rectangle3_heights[1211]), .RECT3_WEIGHT(rectangle3_weights[1211]), .FEAT_THRES(feature_thresholds[1211]), .FEAT_ABOVE(feature_aboves[1211]), .FEAT_BELOW(feature_belows[1211])) ac1211(.scan_win(scan_win1211), .scan_win_std_dev(scan_win_std_dev[1211]), .feature_accum(feature_accums[1211]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1212]), .RECT1_Y(rectangle1_ys[1212]), .RECT1_WIDTH(rectangle1_widths[1212]), .RECT1_HEIGHT(rectangle1_heights[1212]), .RECT1_WEIGHT(rectangle1_weights[1212]), .RECT2_X(rectangle2_xs[1212]), .RECT2_Y(rectangle2_ys[1212]), .RECT2_WIDTH(rectangle2_widths[1212]), .RECT2_HEIGHT(rectangle2_heights[1212]), .RECT2_WEIGHT(rectangle2_weights[1212]), .RECT3_X(rectangle3_xs[1212]), .RECT3_Y(rectangle3_ys[1212]), .RECT3_WIDTH(rectangle3_widths[1212]), .RECT3_HEIGHT(rectangle3_heights[1212]), .RECT3_WEIGHT(rectangle3_weights[1212]), .FEAT_THRES(feature_thresholds[1212]), .FEAT_ABOVE(feature_aboves[1212]), .FEAT_BELOW(feature_belows[1212])) ac1212(.scan_win(scan_win1212), .scan_win_std_dev(scan_win_std_dev[1212]), .feature_accum(feature_accums[1212]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1213]), .RECT1_Y(rectangle1_ys[1213]), .RECT1_WIDTH(rectangle1_widths[1213]), .RECT1_HEIGHT(rectangle1_heights[1213]), .RECT1_WEIGHT(rectangle1_weights[1213]), .RECT2_X(rectangle2_xs[1213]), .RECT2_Y(rectangle2_ys[1213]), .RECT2_WIDTH(rectangle2_widths[1213]), .RECT2_HEIGHT(rectangle2_heights[1213]), .RECT2_WEIGHT(rectangle2_weights[1213]), .RECT3_X(rectangle3_xs[1213]), .RECT3_Y(rectangle3_ys[1213]), .RECT3_WIDTH(rectangle3_widths[1213]), .RECT3_HEIGHT(rectangle3_heights[1213]), .RECT3_WEIGHT(rectangle3_weights[1213]), .FEAT_THRES(feature_thresholds[1213]), .FEAT_ABOVE(feature_aboves[1213]), .FEAT_BELOW(feature_belows[1213])) ac1213(.scan_win(scan_win1213), .scan_win_std_dev(scan_win_std_dev[1213]), .feature_accum(feature_accums[1213]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1214]), .RECT1_Y(rectangle1_ys[1214]), .RECT1_WIDTH(rectangle1_widths[1214]), .RECT1_HEIGHT(rectangle1_heights[1214]), .RECT1_WEIGHT(rectangle1_weights[1214]), .RECT2_X(rectangle2_xs[1214]), .RECT2_Y(rectangle2_ys[1214]), .RECT2_WIDTH(rectangle2_widths[1214]), .RECT2_HEIGHT(rectangle2_heights[1214]), .RECT2_WEIGHT(rectangle2_weights[1214]), .RECT3_X(rectangle3_xs[1214]), .RECT3_Y(rectangle3_ys[1214]), .RECT3_WIDTH(rectangle3_widths[1214]), .RECT3_HEIGHT(rectangle3_heights[1214]), .RECT3_WEIGHT(rectangle3_weights[1214]), .FEAT_THRES(feature_thresholds[1214]), .FEAT_ABOVE(feature_aboves[1214]), .FEAT_BELOW(feature_belows[1214])) ac1214(.scan_win(scan_win1214), .scan_win_std_dev(scan_win_std_dev[1214]), .feature_accum(feature_accums[1214]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1215]), .RECT1_Y(rectangle1_ys[1215]), .RECT1_WIDTH(rectangle1_widths[1215]), .RECT1_HEIGHT(rectangle1_heights[1215]), .RECT1_WEIGHT(rectangle1_weights[1215]), .RECT2_X(rectangle2_xs[1215]), .RECT2_Y(rectangle2_ys[1215]), .RECT2_WIDTH(rectangle2_widths[1215]), .RECT2_HEIGHT(rectangle2_heights[1215]), .RECT2_WEIGHT(rectangle2_weights[1215]), .RECT3_X(rectangle3_xs[1215]), .RECT3_Y(rectangle3_ys[1215]), .RECT3_WIDTH(rectangle3_widths[1215]), .RECT3_HEIGHT(rectangle3_heights[1215]), .RECT3_WEIGHT(rectangle3_weights[1215]), .FEAT_THRES(feature_thresholds[1215]), .FEAT_ABOVE(feature_aboves[1215]), .FEAT_BELOW(feature_belows[1215])) ac1215(.scan_win(scan_win1215), .scan_win_std_dev(scan_win_std_dev[1215]), .feature_accum(feature_accums[1215]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1216]), .RECT1_Y(rectangle1_ys[1216]), .RECT1_WIDTH(rectangle1_widths[1216]), .RECT1_HEIGHT(rectangle1_heights[1216]), .RECT1_WEIGHT(rectangle1_weights[1216]), .RECT2_X(rectangle2_xs[1216]), .RECT2_Y(rectangle2_ys[1216]), .RECT2_WIDTH(rectangle2_widths[1216]), .RECT2_HEIGHT(rectangle2_heights[1216]), .RECT2_WEIGHT(rectangle2_weights[1216]), .RECT3_X(rectangle3_xs[1216]), .RECT3_Y(rectangle3_ys[1216]), .RECT3_WIDTH(rectangle3_widths[1216]), .RECT3_HEIGHT(rectangle3_heights[1216]), .RECT3_WEIGHT(rectangle3_weights[1216]), .FEAT_THRES(feature_thresholds[1216]), .FEAT_ABOVE(feature_aboves[1216]), .FEAT_BELOW(feature_belows[1216])) ac1216(.scan_win(scan_win1216), .scan_win_std_dev(scan_win_std_dev[1216]), .feature_accum(feature_accums[1216]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1217]), .RECT1_Y(rectangle1_ys[1217]), .RECT1_WIDTH(rectangle1_widths[1217]), .RECT1_HEIGHT(rectangle1_heights[1217]), .RECT1_WEIGHT(rectangle1_weights[1217]), .RECT2_X(rectangle2_xs[1217]), .RECT2_Y(rectangle2_ys[1217]), .RECT2_WIDTH(rectangle2_widths[1217]), .RECT2_HEIGHT(rectangle2_heights[1217]), .RECT2_WEIGHT(rectangle2_weights[1217]), .RECT3_X(rectangle3_xs[1217]), .RECT3_Y(rectangle3_ys[1217]), .RECT3_WIDTH(rectangle3_widths[1217]), .RECT3_HEIGHT(rectangle3_heights[1217]), .RECT3_WEIGHT(rectangle3_weights[1217]), .FEAT_THRES(feature_thresholds[1217]), .FEAT_ABOVE(feature_aboves[1217]), .FEAT_BELOW(feature_belows[1217])) ac1217(.scan_win(scan_win1217), .scan_win_std_dev(scan_win_std_dev[1217]), .feature_accum(feature_accums[1217]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1218]), .RECT1_Y(rectangle1_ys[1218]), .RECT1_WIDTH(rectangle1_widths[1218]), .RECT1_HEIGHT(rectangle1_heights[1218]), .RECT1_WEIGHT(rectangle1_weights[1218]), .RECT2_X(rectangle2_xs[1218]), .RECT2_Y(rectangle2_ys[1218]), .RECT2_WIDTH(rectangle2_widths[1218]), .RECT2_HEIGHT(rectangle2_heights[1218]), .RECT2_WEIGHT(rectangle2_weights[1218]), .RECT3_X(rectangle3_xs[1218]), .RECT3_Y(rectangle3_ys[1218]), .RECT3_WIDTH(rectangle3_widths[1218]), .RECT3_HEIGHT(rectangle3_heights[1218]), .RECT3_WEIGHT(rectangle3_weights[1218]), .FEAT_THRES(feature_thresholds[1218]), .FEAT_ABOVE(feature_aboves[1218]), .FEAT_BELOW(feature_belows[1218])) ac1218(.scan_win(scan_win1218), .scan_win_std_dev(scan_win_std_dev[1218]), .feature_accum(feature_accums[1218]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1219]), .RECT1_Y(rectangle1_ys[1219]), .RECT1_WIDTH(rectangle1_widths[1219]), .RECT1_HEIGHT(rectangle1_heights[1219]), .RECT1_WEIGHT(rectangle1_weights[1219]), .RECT2_X(rectangle2_xs[1219]), .RECT2_Y(rectangle2_ys[1219]), .RECT2_WIDTH(rectangle2_widths[1219]), .RECT2_HEIGHT(rectangle2_heights[1219]), .RECT2_WEIGHT(rectangle2_weights[1219]), .RECT3_X(rectangle3_xs[1219]), .RECT3_Y(rectangle3_ys[1219]), .RECT3_WIDTH(rectangle3_widths[1219]), .RECT3_HEIGHT(rectangle3_heights[1219]), .RECT3_WEIGHT(rectangle3_weights[1219]), .FEAT_THRES(feature_thresholds[1219]), .FEAT_ABOVE(feature_aboves[1219]), .FEAT_BELOW(feature_belows[1219])) ac1219(.scan_win(scan_win1219), .scan_win_std_dev(scan_win_std_dev[1219]), .feature_accum(feature_accums[1219]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1220]), .RECT1_Y(rectangle1_ys[1220]), .RECT1_WIDTH(rectangle1_widths[1220]), .RECT1_HEIGHT(rectangle1_heights[1220]), .RECT1_WEIGHT(rectangle1_weights[1220]), .RECT2_X(rectangle2_xs[1220]), .RECT2_Y(rectangle2_ys[1220]), .RECT2_WIDTH(rectangle2_widths[1220]), .RECT2_HEIGHT(rectangle2_heights[1220]), .RECT2_WEIGHT(rectangle2_weights[1220]), .RECT3_X(rectangle3_xs[1220]), .RECT3_Y(rectangle3_ys[1220]), .RECT3_WIDTH(rectangle3_widths[1220]), .RECT3_HEIGHT(rectangle3_heights[1220]), .RECT3_WEIGHT(rectangle3_weights[1220]), .FEAT_THRES(feature_thresholds[1220]), .FEAT_ABOVE(feature_aboves[1220]), .FEAT_BELOW(feature_belows[1220])) ac1220(.scan_win(scan_win1220), .scan_win_std_dev(scan_win_std_dev[1220]), .feature_accum(feature_accums[1220]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1221]), .RECT1_Y(rectangle1_ys[1221]), .RECT1_WIDTH(rectangle1_widths[1221]), .RECT1_HEIGHT(rectangle1_heights[1221]), .RECT1_WEIGHT(rectangle1_weights[1221]), .RECT2_X(rectangle2_xs[1221]), .RECT2_Y(rectangle2_ys[1221]), .RECT2_WIDTH(rectangle2_widths[1221]), .RECT2_HEIGHT(rectangle2_heights[1221]), .RECT2_WEIGHT(rectangle2_weights[1221]), .RECT3_X(rectangle3_xs[1221]), .RECT3_Y(rectangle3_ys[1221]), .RECT3_WIDTH(rectangle3_widths[1221]), .RECT3_HEIGHT(rectangle3_heights[1221]), .RECT3_WEIGHT(rectangle3_weights[1221]), .FEAT_THRES(feature_thresholds[1221]), .FEAT_ABOVE(feature_aboves[1221]), .FEAT_BELOW(feature_belows[1221])) ac1221(.scan_win(scan_win1221), .scan_win_std_dev(scan_win_std_dev[1221]), .feature_accum(feature_accums[1221]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1222]), .RECT1_Y(rectangle1_ys[1222]), .RECT1_WIDTH(rectangle1_widths[1222]), .RECT1_HEIGHT(rectangle1_heights[1222]), .RECT1_WEIGHT(rectangle1_weights[1222]), .RECT2_X(rectangle2_xs[1222]), .RECT2_Y(rectangle2_ys[1222]), .RECT2_WIDTH(rectangle2_widths[1222]), .RECT2_HEIGHT(rectangle2_heights[1222]), .RECT2_WEIGHT(rectangle2_weights[1222]), .RECT3_X(rectangle3_xs[1222]), .RECT3_Y(rectangle3_ys[1222]), .RECT3_WIDTH(rectangle3_widths[1222]), .RECT3_HEIGHT(rectangle3_heights[1222]), .RECT3_WEIGHT(rectangle3_weights[1222]), .FEAT_THRES(feature_thresholds[1222]), .FEAT_ABOVE(feature_aboves[1222]), .FEAT_BELOW(feature_belows[1222])) ac1222(.scan_win(scan_win1222), .scan_win_std_dev(scan_win_std_dev[1222]), .feature_accum(feature_accums[1222]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1223]), .RECT1_Y(rectangle1_ys[1223]), .RECT1_WIDTH(rectangle1_widths[1223]), .RECT1_HEIGHT(rectangle1_heights[1223]), .RECT1_WEIGHT(rectangle1_weights[1223]), .RECT2_X(rectangle2_xs[1223]), .RECT2_Y(rectangle2_ys[1223]), .RECT2_WIDTH(rectangle2_widths[1223]), .RECT2_HEIGHT(rectangle2_heights[1223]), .RECT2_WEIGHT(rectangle2_weights[1223]), .RECT3_X(rectangle3_xs[1223]), .RECT3_Y(rectangle3_ys[1223]), .RECT3_WIDTH(rectangle3_widths[1223]), .RECT3_HEIGHT(rectangle3_heights[1223]), .RECT3_WEIGHT(rectangle3_weights[1223]), .FEAT_THRES(feature_thresholds[1223]), .FEAT_ABOVE(feature_aboves[1223]), .FEAT_BELOW(feature_belows[1223])) ac1223(.scan_win(scan_win1223), .scan_win_std_dev(scan_win_std_dev[1223]), .feature_accum(feature_accums[1223]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1224]), .RECT1_Y(rectangle1_ys[1224]), .RECT1_WIDTH(rectangle1_widths[1224]), .RECT1_HEIGHT(rectangle1_heights[1224]), .RECT1_WEIGHT(rectangle1_weights[1224]), .RECT2_X(rectangle2_xs[1224]), .RECT2_Y(rectangle2_ys[1224]), .RECT2_WIDTH(rectangle2_widths[1224]), .RECT2_HEIGHT(rectangle2_heights[1224]), .RECT2_WEIGHT(rectangle2_weights[1224]), .RECT3_X(rectangle3_xs[1224]), .RECT3_Y(rectangle3_ys[1224]), .RECT3_WIDTH(rectangle3_widths[1224]), .RECT3_HEIGHT(rectangle3_heights[1224]), .RECT3_WEIGHT(rectangle3_weights[1224]), .FEAT_THRES(feature_thresholds[1224]), .FEAT_ABOVE(feature_aboves[1224]), .FEAT_BELOW(feature_belows[1224])) ac1224(.scan_win(scan_win1224), .scan_win_std_dev(scan_win_std_dev[1224]), .feature_accum(feature_accums[1224]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1225]), .RECT1_Y(rectangle1_ys[1225]), .RECT1_WIDTH(rectangle1_widths[1225]), .RECT1_HEIGHT(rectangle1_heights[1225]), .RECT1_WEIGHT(rectangle1_weights[1225]), .RECT2_X(rectangle2_xs[1225]), .RECT2_Y(rectangle2_ys[1225]), .RECT2_WIDTH(rectangle2_widths[1225]), .RECT2_HEIGHT(rectangle2_heights[1225]), .RECT2_WEIGHT(rectangle2_weights[1225]), .RECT3_X(rectangle3_xs[1225]), .RECT3_Y(rectangle3_ys[1225]), .RECT3_WIDTH(rectangle3_widths[1225]), .RECT3_HEIGHT(rectangle3_heights[1225]), .RECT3_WEIGHT(rectangle3_weights[1225]), .FEAT_THRES(feature_thresholds[1225]), .FEAT_ABOVE(feature_aboves[1225]), .FEAT_BELOW(feature_belows[1225])) ac1225(.scan_win(scan_win1225), .scan_win_std_dev(scan_win_std_dev[1225]), .feature_accum(feature_accums[1225]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1226]), .RECT1_Y(rectangle1_ys[1226]), .RECT1_WIDTH(rectangle1_widths[1226]), .RECT1_HEIGHT(rectangle1_heights[1226]), .RECT1_WEIGHT(rectangle1_weights[1226]), .RECT2_X(rectangle2_xs[1226]), .RECT2_Y(rectangle2_ys[1226]), .RECT2_WIDTH(rectangle2_widths[1226]), .RECT2_HEIGHT(rectangle2_heights[1226]), .RECT2_WEIGHT(rectangle2_weights[1226]), .RECT3_X(rectangle3_xs[1226]), .RECT3_Y(rectangle3_ys[1226]), .RECT3_WIDTH(rectangle3_widths[1226]), .RECT3_HEIGHT(rectangle3_heights[1226]), .RECT3_WEIGHT(rectangle3_weights[1226]), .FEAT_THRES(feature_thresholds[1226]), .FEAT_ABOVE(feature_aboves[1226]), .FEAT_BELOW(feature_belows[1226])) ac1226(.scan_win(scan_win1226), .scan_win_std_dev(scan_win_std_dev[1226]), .feature_accum(feature_accums[1226]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1227]), .RECT1_Y(rectangle1_ys[1227]), .RECT1_WIDTH(rectangle1_widths[1227]), .RECT1_HEIGHT(rectangle1_heights[1227]), .RECT1_WEIGHT(rectangle1_weights[1227]), .RECT2_X(rectangle2_xs[1227]), .RECT2_Y(rectangle2_ys[1227]), .RECT2_WIDTH(rectangle2_widths[1227]), .RECT2_HEIGHT(rectangle2_heights[1227]), .RECT2_WEIGHT(rectangle2_weights[1227]), .RECT3_X(rectangle3_xs[1227]), .RECT3_Y(rectangle3_ys[1227]), .RECT3_WIDTH(rectangle3_widths[1227]), .RECT3_HEIGHT(rectangle3_heights[1227]), .RECT3_WEIGHT(rectangle3_weights[1227]), .FEAT_THRES(feature_thresholds[1227]), .FEAT_ABOVE(feature_aboves[1227]), .FEAT_BELOW(feature_belows[1227])) ac1227(.scan_win(scan_win1227), .scan_win_std_dev(scan_win_std_dev[1227]), .feature_accum(feature_accums[1227]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1228]), .RECT1_Y(rectangle1_ys[1228]), .RECT1_WIDTH(rectangle1_widths[1228]), .RECT1_HEIGHT(rectangle1_heights[1228]), .RECT1_WEIGHT(rectangle1_weights[1228]), .RECT2_X(rectangle2_xs[1228]), .RECT2_Y(rectangle2_ys[1228]), .RECT2_WIDTH(rectangle2_widths[1228]), .RECT2_HEIGHT(rectangle2_heights[1228]), .RECT2_WEIGHT(rectangle2_weights[1228]), .RECT3_X(rectangle3_xs[1228]), .RECT3_Y(rectangle3_ys[1228]), .RECT3_WIDTH(rectangle3_widths[1228]), .RECT3_HEIGHT(rectangle3_heights[1228]), .RECT3_WEIGHT(rectangle3_weights[1228]), .FEAT_THRES(feature_thresholds[1228]), .FEAT_ABOVE(feature_aboves[1228]), .FEAT_BELOW(feature_belows[1228])) ac1228(.scan_win(scan_win1228), .scan_win_std_dev(scan_win_std_dev[1228]), .feature_accum(feature_accums[1228]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1229]), .RECT1_Y(rectangle1_ys[1229]), .RECT1_WIDTH(rectangle1_widths[1229]), .RECT1_HEIGHT(rectangle1_heights[1229]), .RECT1_WEIGHT(rectangle1_weights[1229]), .RECT2_X(rectangle2_xs[1229]), .RECT2_Y(rectangle2_ys[1229]), .RECT2_WIDTH(rectangle2_widths[1229]), .RECT2_HEIGHT(rectangle2_heights[1229]), .RECT2_WEIGHT(rectangle2_weights[1229]), .RECT3_X(rectangle3_xs[1229]), .RECT3_Y(rectangle3_ys[1229]), .RECT3_WIDTH(rectangle3_widths[1229]), .RECT3_HEIGHT(rectangle3_heights[1229]), .RECT3_WEIGHT(rectangle3_weights[1229]), .FEAT_THRES(feature_thresholds[1229]), .FEAT_ABOVE(feature_aboves[1229]), .FEAT_BELOW(feature_belows[1229])) ac1229(.scan_win(scan_win1229), .scan_win_std_dev(scan_win_std_dev[1229]), .feature_accum(feature_accums[1229]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1230]), .RECT1_Y(rectangle1_ys[1230]), .RECT1_WIDTH(rectangle1_widths[1230]), .RECT1_HEIGHT(rectangle1_heights[1230]), .RECT1_WEIGHT(rectangle1_weights[1230]), .RECT2_X(rectangle2_xs[1230]), .RECT2_Y(rectangle2_ys[1230]), .RECT2_WIDTH(rectangle2_widths[1230]), .RECT2_HEIGHT(rectangle2_heights[1230]), .RECT2_WEIGHT(rectangle2_weights[1230]), .RECT3_X(rectangle3_xs[1230]), .RECT3_Y(rectangle3_ys[1230]), .RECT3_WIDTH(rectangle3_widths[1230]), .RECT3_HEIGHT(rectangle3_heights[1230]), .RECT3_WEIGHT(rectangle3_weights[1230]), .FEAT_THRES(feature_thresholds[1230]), .FEAT_ABOVE(feature_aboves[1230]), .FEAT_BELOW(feature_belows[1230])) ac1230(.scan_win(scan_win1230), .scan_win_std_dev(scan_win_std_dev[1230]), .feature_accum(feature_accums[1230]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1231]), .RECT1_Y(rectangle1_ys[1231]), .RECT1_WIDTH(rectangle1_widths[1231]), .RECT1_HEIGHT(rectangle1_heights[1231]), .RECT1_WEIGHT(rectangle1_weights[1231]), .RECT2_X(rectangle2_xs[1231]), .RECT2_Y(rectangle2_ys[1231]), .RECT2_WIDTH(rectangle2_widths[1231]), .RECT2_HEIGHT(rectangle2_heights[1231]), .RECT2_WEIGHT(rectangle2_weights[1231]), .RECT3_X(rectangle3_xs[1231]), .RECT3_Y(rectangle3_ys[1231]), .RECT3_WIDTH(rectangle3_widths[1231]), .RECT3_HEIGHT(rectangle3_heights[1231]), .RECT3_WEIGHT(rectangle3_weights[1231]), .FEAT_THRES(feature_thresholds[1231]), .FEAT_ABOVE(feature_aboves[1231]), .FEAT_BELOW(feature_belows[1231])) ac1231(.scan_win(scan_win1231), .scan_win_std_dev(scan_win_std_dev[1231]), .feature_accum(feature_accums[1231]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1232]), .RECT1_Y(rectangle1_ys[1232]), .RECT1_WIDTH(rectangle1_widths[1232]), .RECT1_HEIGHT(rectangle1_heights[1232]), .RECT1_WEIGHT(rectangle1_weights[1232]), .RECT2_X(rectangle2_xs[1232]), .RECT2_Y(rectangle2_ys[1232]), .RECT2_WIDTH(rectangle2_widths[1232]), .RECT2_HEIGHT(rectangle2_heights[1232]), .RECT2_WEIGHT(rectangle2_weights[1232]), .RECT3_X(rectangle3_xs[1232]), .RECT3_Y(rectangle3_ys[1232]), .RECT3_WIDTH(rectangle3_widths[1232]), .RECT3_HEIGHT(rectangle3_heights[1232]), .RECT3_WEIGHT(rectangle3_weights[1232]), .FEAT_THRES(feature_thresholds[1232]), .FEAT_ABOVE(feature_aboves[1232]), .FEAT_BELOW(feature_belows[1232])) ac1232(.scan_win(scan_win1232), .scan_win_std_dev(scan_win_std_dev[1232]), .feature_accum(feature_accums[1232]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1233]), .RECT1_Y(rectangle1_ys[1233]), .RECT1_WIDTH(rectangle1_widths[1233]), .RECT1_HEIGHT(rectangle1_heights[1233]), .RECT1_WEIGHT(rectangle1_weights[1233]), .RECT2_X(rectangle2_xs[1233]), .RECT2_Y(rectangle2_ys[1233]), .RECT2_WIDTH(rectangle2_widths[1233]), .RECT2_HEIGHT(rectangle2_heights[1233]), .RECT2_WEIGHT(rectangle2_weights[1233]), .RECT3_X(rectangle3_xs[1233]), .RECT3_Y(rectangle3_ys[1233]), .RECT3_WIDTH(rectangle3_widths[1233]), .RECT3_HEIGHT(rectangle3_heights[1233]), .RECT3_WEIGHT(rectangle3_weights[1233]), .FEAT_THRES(feature_thresholds[1233]), .FEAT_ABOVE(feature_aboves[1233]), .FEAT_BELOW(feature_belows[1233])) ac1233(.scan_win(scan_win1233), .scan_win_std_dev(scan_win_std_dev[1233]), .feature_accum(feature_accums[1233]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1234]), .RECT1_Y(rectangle1_ys[1234]), .RECT1_WIDTH(rectangle1_widths[1234]), .RECT1_HEIGHT(rectangle1_heights[1234]), .RECT1_WEIGHT(rectangle1_weights[1234]), .RECT2_X(rectangle2_xs[1234]), .RECT2_Y(rectangle2_ys[1234]), .RECT2_WIDTH(rectangle2_widths[1234]), .RECT2_HEIGHT(rectangle2_heights[1234]), .RECT2_WEIGHT(rectangle2_weights[1234]), .RECT3_X(rectangle3_xs[1234]), .RECT3_Y(rectangle3_ys[1234]), .RECT3_WIDTH(rectangle3_widths[1234]), .RECT3_HEIGHT(rectangle3_heights[1234]), .RECT3_WEIGHT(rectangle3_weights[1234]), .FEAT_THRES(feature_thresholds[1234]), .FEAT_ABOVE(feature_aboves[1234]), .FEAT_BELOW(feature_belows[1234])) ac1234(.scan_win(scan_win1234), .scan_win_std_dev(scan_win_std_dev[1234]), .feature_accum(feature_accums[1234]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1235]), .RECT1_Y(rectangle1_ys[1235]), .RECT1_WIDTH(rectangle1_widths[1235]), .RECT1_HEIGHT(rectangle1_heights[1235]), .RECT1_WEIGHT(rectangle1_weights[1235]), .RECT2_X(rectangle2_xs[1235]), .RECT2_Y(rectangle2_ys[1235]), .RECT2_WIDTH(rectangle2_widths[1235]), .RECT2_HEIGHT(rectangle2_heights[1235]), .RECT2_WEIGHT(rectangle2_weights[1235]), .RECT3_X(rectangle3_xs[1235]), .RECT3_Y(rectangle3_ys[1235]), .RECT3_WIDTH(rectangle3_widths[1235]), .RECT3_HEIGHT(rectangle3_heights[1235]), .RECT3_WEIGHT(rectangle3_weights[1235]), .FEAT_THRES(feature_thresholds[1235]), .FEAT_ABOVE(feature_aboves[1235]), .FEAT_BELOW(feature_belows[1235])) ac1235(.scan_win(scan_win1235), .scan_win_std_dev(scan_win_std_dev[1235]), .feature_accum(feature_accums[1235]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1236]), .RECT1_Y(rectangle1_ys[1236]), .RECT1_WIDTH(rectangle1_widths[1236]), .RECT1_HEIGHT(rectangle1_heights[1236]), .RECT1_WEIGHT(rectangle1_weights[1236]), .RECT2_X(rectangle2_xs[1236]), .RECT2_Y(rectangle2_ys[1236]), .RECT2_WIDTH(rectangle2_widths[1236]), .RECT2_HEIGHT(rectangle2_heights[1236]), .RECT2_WEIGHT(rectangle2_weights[1236]), .RECT3_X(rectangle3_xs[1236]), .RECT3_Y(rectangle3_ys[1236]), .RECT3_WIDTH(rectangle3_widths[1236]), .RECT3_HEIGHT(rectangle3_heights[1236]), .RECT3_WEIGHT(rectangle3_weights[1236]), .FEAT_THRES(feature_thresholds[1236]), .FEAT_ABOVE(feature_aboves[1236]), .FEAT_BELOW(feature_belows[1236])) ac1236(.scan_win(scan_win1236), .scan_win_std_dev(scan_win_std_dev[1236]), .feature_accum(feature_accums[1236]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1237]), .RECT1_Y(rectangle1_ys[1237]), .RECT1_WIDTH(rectangle1_widths[1237]), .RECT1_HEIGHT(rectangle1_heights[1237]), .RECT1_WEIGHT(rectangle1_weights[1237]), .RECT2_X(rectangle2_xs[1237]), .RECT2_Y(rectangle2_ys[1237]), .RECT2_WIDTH(rectangle2_widths[1237]), .RECT2_HEIGHT(rectangle2_heights[1237]), .RECT2_WEIGHT(rectangle2_weights[1237]), .RECT3_X(rectangle3_xs[1237]), .RECT3_Y(rectangle3_ys[1237]), .RECT3_WIDTH(rectangle3_widths[1237]), .RECT3_HEIGHT(rectangle3_heights[1237]), .RECT3_WEIGHT(rectangle3_weights[1237]), .FEAT_THRES(feature_thresholds[1237]), .FEAT_ABOVE(feature_aboves[1237]), .FEAT_BELOW(feature_belows[1237])) ac1237(.scan_win(scan_win1237), .scan_win_std_dev(scan_win_std_dev[1237]), .feature_accum(feature_accums[1237]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1238]), .RECT1_Y(rectangle1_ys[1238]), .RECT1_WIDTH(rectangle1_widths[1238]), .RECT1_HEIGHT(rectangle1_heights[1238]), .RECT1_WEIGHT(rectangle1_weights[1238]), .RECT2_X(rectangle2_xs[1238]), .RECT2_Y(rectangle2_ys[1238]), .RECT2_WIDTH(rectangle2_widths[1238]), .RECT2_HEIGHT(rectangle2_heights[1238]), .RECT2_WEIGHT(rectangle2_weights[1238]), .RECT3_X(rectangle3_xs[1238]), .RECT3_Y(rectangle3_ys[1238]), .RECT3_WIDTH(rectangle3_widths[1238]), .RECT3_HEIGHT(rectangle3_heights[1238]), .RECT3_WEIGHT(rectangle3_weights[1238]), .FEAT_THRES(feature_thresholds[1238]), .FEAT_ABOVE(feature_aboves[1238]), .FEAT_BELOW(feature_belows[1238])) ac1238(.scan_win(scan_win1238), .scan_win_std_dev(scan_win_std_dev[1238]), .feature_accum(feature_accums[1238]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1239]), .RECT1_Y(rectangle1_ys[1239]), .RECT1_WIDTH(rectangle1_widths[1239]), .RECT1_HEIGHT(rectangle1_heights[1239]), .RECT1_WEIGHT(rectangle1_weights[1239]), .RECT2_X(rectangle2_xs[1239]), .RECT2_Y(rectangle2_ys[1239]), .RECT2_WIDTH(rectangle2_widths[1239]), .RECT2_HEIGHT(rectangle2_heights[1239]), .RECT2_WEIGHT(rectangle2_weights[1239]), .RECT3_X(rectangle3_xs[1239]), .RECT3_Y(rectangle3_ys[1239]), .RECT3_WIDTH(rectangle3_widths[1239]), .RECT3_HEIGHT(rectangle3_heights[1239]), .RECT3_WEIGHT(rectangle3_weights[1239]), .FEAT_THRES(feature_thresholds[1239]), .FEAT_ABOVE(feature_aboves[1239]), .FEAT_BELOW(feature_belows[1239])) ac1239(.scan_win(scan_win1239), .scan_win_std_dev(scan_win_std_dev[1239]), .feature_accum(feature_accums[1239]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1240]), .RECT1_Y(rectangle1_ys[1240]), .RECT1_WIDTH(rectangle1_widths[1240]), .RECT1_HEIGHT(rectangle1_heights[1240]), .RECT1_WEIGHT(rectangle1_weights[1240]), .RECT2_X(rectangle2_xs[1240]), .RECT2_Y(rectangle2_ys[1240]), .RECT2_WIDTH(rectangle2_widths[1240]), .RECT2_HEIGHT(rectangle2_heights[1240]), .RECT2_WEIGHT(rectangle2_weights[1240]), .RECT3_X(rectangle3_xs[1240]), .RECT3_Y(rectangle3_ys[1240]), .RECT3_WIDTH(rectangle3_widths[1240]), .RECT3_HEIGHT(rectangle3_heights[1240]), .RECT3_WEIGHT(rectangle3_weights[1240]), .FEAT_THRES(feature_thresholds[1240]), .FEAT_ABOVE(feature_aboves[1240]), .FEAT_BELOW(feature_belows[1240])) ac1240(.scan_win(scan_win1240), .scan_win_std_dev(scan_win_std_dev[1240]), .feature_accum(feature_accums[1240]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1241]), .RECT1_Y(rectangle1_ys[1241]), .RECT1_WIDTH(rectangle1_widths[1241]), .RECT1_HEIGHT(rectangle1_heights[1241]), .RECT1_WEIGHT(rectangle1_weights[1241]), .RECT2_X(rectangle2_xs[1241]), .RECT2_Y(rectangle2_ys[1241]), .RECT2_WIDTH(rectangle2_widths[1241]), .RECT2_HEIGHT(rectangle2_heights[1241]), .RECT2_WEIGHT(rectangle2_weights[1241]), .RECT3_X(rectangle3_xs[1241]), .RECT3_Y(rectangle3_ys[1241]), .RECT3_WIDTH(rectangle3_widths[1241]), .RECT3_HEIGHT(rectangle3_heights[1241]), .RECT3_WEIGHT(rectangle3_weights[1241]), .FEAT_THRES(feature_thresholds[1241]), .FEAT_ABOVE(feature_aboves[1241]), .FEAT_BELOW(feature_belows[1241])) ac1241(.scan_win(scan_win1241), .scan_win_std_dev(scan_win_std_dev[1241]), .feature_accum(feature_accums[1241]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1242]), .RECT1_Y(rectangle1_ys[1242]), .RECT1_WIDTH(rectangle1_widths[1242]), .RECT1_HEIGHT(rectangle1_heights[1242]), .RECT1_WEIGHT(rectangle1_weights[1242]), .RECT2_X(rectangle2_xs[1242]), .RECT2_Y(rectangle2_ys[1242]), .RECT2_WIDTH(rectangle2_widths[1242]), .RECT2_HEIGHT(rectangle2_heights[1242]), .RECT2_WEIGHT(rectangle2_weights[1242]), .RECT3_X(rectangle3_xs[1242]), .RECT3_Y(rectangle3_ys[1242]), .RECT3_WIDTH(rectangle3_widths[1242]), .RECT3_HEIGHT(rectangle3_heights[1242]), .RECT3_WEIGHT(rectangle3_weights[1242]), .FEAT_THRES(feature_thresholds[1242]), .FEAT_ABOVE(feature_aboves[1242]), .FEAT_BELOW(feature_belows[1242])) ac1242(.scan_win(scan_win1242), .scan_win_std_dev(scan_win_std_dev[1242]), .feature_accum(feature_accums[1242]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1243]), .RECT1_Y(rectangle1_ys[1243]), .RECT1_WIDTH(rectangle1_widths[1243]), .RECT1_HEIGHT(rectangle1_heights[1243]), .RECT1_WEIGHT(rectangle1_weights[1243]), .RECT2_X(rectangle2_xs[1243]), .RECT2_Y(rectangle2_ys[1243]), .RECT2_WIDTH(rectangle2_widths[1243]), .RECT2_HEIGHT(rectangle2_heights[1243]), .RECT2_WEIGHT(rectangle2_weights[1243]), .RECT3_X(rectangle3_xs[1243]), .RECT3_Y(rectangle3_ys[1243]), .RECT3_WIDTH(rectangle3_widths[1243]), .RECT3_HEIGHT(rectangle3_heights[1243]), .RECT3_WEIGHT(rectangle3_weights[1243]), .FEAT_THRES(feature_thresholds[1243]), .FEAT_ABOVE(feature_aboves[1243]), .FEAT_BELOW(feature_belows[1243])) ac1243(.scan_win(scan_win1243), .scan_win_std_dev(scan_win_std_dev[1243]), .feature_accum(feature_accums[1243]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1244]), .RECT1_Y(rectangle1_ys[1244]), .RECT1_WIDTH(rectangle1_widths[1244]), .RECT1_HEIGHT(rectangle1_heights[1244]), .RECT1_WEIGHT(rectangle1_weights[1244]), .RECT2_X(rectangle2_xs[1244]), .RECT2_Y(rectangle2_ys[1244]), .RECT2_WIDTH(rectangle2_widths[1244]), .RECT2_HEIGHT(rectangle2_heights[1244]), .RECT2_WEIGHT(rectangle2_weights[1244]), .RECT3_X(rectangle3_xs[1244]), .RECT3_Y(rectangle3_ys[1244]), .RECT3_WIDTH(rectangle3_widths[1244]), .RECT3_HEIGHT(rectangle3_heights[1244]), .RECT3_WEIGHT(rectangle3_weights[1244]), .FEAT_THRES(feature_thresholds[1244]), .FEAT_ABOVE(feature_aboves[1244]), .FEAT_BELOW(feature_belows[1244])) ac1244(.scan_win(scan_win1244), .scan_win_std_dev(scan_win_std_dev[1244]), .feature_accum(feature_accums[1244]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1245]), .RECT1_Y(rectangle1_ys[1245]), .RECT1_WIDTH(rectangle1_widths[1245]), .RECT1_HEIGHT(rectangle1_heights[1245]), .RECT1_WEIGHT(rectangle1_weights[1245]), .RECT2_X(rectangle2_xs[1245]), .RECT2_Y(rectangle2_ys[1245]), .RECT2_WIDTH(rectangle2_widths[1245]), .RECT2_HEIGHT(rectangle2_heights[1245]), .RECT2_WEIGHT(rectangle2_weights[1245]), .RECT3_X(rectangle3_xs[1245]), .RECT3_Y(rectangle3_ys[1245]), .RECT3_WIDTH(rectangle3_widths[1245]), .RECT3_HEIGHT(rectangle3_heights[1245]), .RECT3_WEIGHT(rectangle3_weights[1245]), .FEAT_THRES(feature_thresholds[1245]), .FEAT_ABOVE(feature_aboves[1245]), .FEAT_BELOW(feature_belows[1245])) ac1245(.scan_win(scan_win1245), .scan_win_std_dev(scan_win_std_dev[1245]), .feature_accum(feature_accums[1245]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1246]), .RECT1_Y(rectangle1_ys[1246]), .RECT1_WIDTH(rectangle1_widths[1246]), .RECT1_HEIGHT(rectangle1_heights[1246]), .RECT1_WEIGHT(rectangle1_weights[1246]), .RECT2_X(rectangle2_xs[1246]), .RECT2_Y(rectangle2_ys[1246]), .RECT2_WIDTH(rectangle2_widths[1246]), .RECT2_HEIGHT(rectangle2_heights[1246]), .RECT2_WEIGHT(rectangle2_weights[1246]), .RECT3_X(rectangle3_xs[1246]), .RECT3_Y(rectangle3_ys[1246]), .RECT3_WIDTH(rectangle3_widths[1246]), .RECT3_HEIGHT(rectangle3_heights[1246]), .RECT3_WEIGHT(rectangle3_weights[1246]), .FEAT_THRES(feature_thresholds[1246]), .FEAT_ABOVE(feature_aboves[1246]), .FEAT_BELOW(feature_belows[1246])) ac1246(.scan_win(scan_win1246), .scan_win_std_dev(scan_win_std_dev[1246]), .feature_accum(feature_accums[1246]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1247]), .RECT1_Y(rectangle1_ys[1247]), .RECT1_WIDTH(rectangle1_widths[1247]), .RECT1_HEIGHT(rectangle1_heights[1247]), .RECT1_WEIGHT(rectangle1_weights[1247]), .RECT2_X(rectangle2_xs[1247]), .RECT2_Y(rectangle2_ys[1247]), .RECT2_WIDTH(rectangle2_widths[1247]), .RECT2_HEIGHT(rectangle2_heights[1247]), .RECT2_WEIGHT(rectangle2_weights[1247]), .RECT3_X(rectangle3_xs[1247]), .RECT3_Y(rectangle3_ys[1247]), .RECT3_WIDTH(rectangle3_widths[1247]), .RECT3_HEIGHT(rectangle3_heights[1247]), .RECT3_WEIGHT(rectangle3_weights[1247]), .FEAT_THRES(feature_thresholds[1247]), .FEAT_ABOVE(feature_aboves[1247]), .FEAT_BELOW(feature_belows[1247])) ac1247(.scan_win(scan_win1247), .scan_win_std_dev(scan_win_std_dev[1247]), .feature_accum(feature_accums[1247]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1248]), .RECT1_Y(rectangle1_ys[1248]), .RECT1_WIDTH(rectangle1_widths[1248]), .RECT1_HEIGHT(rectangle1_heights[1248]), .RECT1_WEIGHT(rectangle1_weights[1248]), .RECT2_X(rectangle2_xs[1248]), .RECT2_Y(rectangle2_ys[1248]), .RECT2_WIDTH(rectangle2_widths[1248]), .RECT2_HEIGHT(rectangle2_heights[1248]), .RECT2_WEIGHT(rectangle2_weights[1248]), .RECT3_X(rectangle3_xs[1248]), .RECT3_Y(rectangle3_ys[1248]), .RECT3_WIDTH(rectangle3_widths[1248]), .RECT3_HEIGHT(rectangle3_heights[1248]), .RECT3_WEIGHT(rectangle3_weights[1248]), .FEAT_THRES(feature_thresholds[1248]), .FEAT_ABOVE(feature_aboves[1248]), .FEAT_BELOW(feature_belows[1248])) ac1248(.scan_win(scan_win1248), .scan_win_std_dev(scan_win_std_dev[1248]), .feature_accum(feature_accums[1248]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1249]), .RECT1_Y(rectangle1_ys[1249]), .RECT1_WIDTH(rectangle1_widths[1249]), .RECT1_HEIGHT(rectangle1_heights[1249]), .RECT1_WEIGHT(rectangle1_weights[1249]), .RECT2_X(rectangle2_xs[1249]), .RECT2_Y(rectangle2_ys[1249]), .RECT2_WIDTH(rectangle2_widths[1249]), .RECT2_HEIGHT(rectangle2_heights[1249]), .RECT2_WEIGHT(rectangle2_weights[1249]), .RECT3_X(rectangle3_xs[1249]), .RECT3_Y(rectangle3_ys[1249]), .RECT3_WIDTH(rectangle3_widths[1249]), .RECT3_HEIGHT(rectangle3_heights[1249]), .RECT3_WEIGHT(rectangle3_weights[1249]), .FEAT_THRES(feature_thresholds[1249]), .FEAT_ABOVE(feature_aboves[1249]), .FEAT_BELOW(feature_belows[1249])) ac1249(.scan_win(scan_win1249), .scan_win_std_dev(scan_win_std_dev[1249]), .feature_accum(feature_accums[1249]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1250]), .RECT1_Y(rectangle1_ys[1250]), .RECT1_WIDTH(rectangle1_widths[1250]), .RECT1_HEIGHT(rectangle1_heights[1250]), .RECT1_WEIGHT(rectangle1_weights[1250]), .RECT2_X(rectangle2_xs[1250]), .RECT2_Y(rectangle2_ys[1250]), .RECT2_WIDTH(rectangle2_widths[1250]), .RECT2_HEIGHT(rectangle2_heights[1250]), .RECT2_WEIGHT(rectangle2_weights[1250]), .RECT3_X(rectangle3_xs[1250]), .RECT3_Y(rectangle3_ys[1250]), .RECT3_WIDTH(rectangle3_widths[1250]), .RECT3_HEIGHT(rectangle3_heights[1250]), .RECT3_WEIGHT(rectangle3_weights[1250]), .FEAT_THRES(feature_thresholds[1250]), .FEAT_ABOVE(feature_aboves[1250]), .FEAT_BELOW(feature_belows[1250])) ac1250(.scan_win(scan_win1250), .scan_win_std_dev(scan_win_std_dev[1250]), .feature_accum(feature_accums[1250]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1251]), .RECT1_Y(rectangle1_ys[1251]), .RECT1_WIDTH(rectangle1_widths[1251]), .RECT1_HEIGHT(rectangle1_heights[1251]), .RECT1_WEIGHT(rectangle1_weights[1251]), .RECT2_X(rectangle2_xs[1251]), .RECT2_Y(rectangle2_ys[1251]), .RECT2_WIDTH(rectangle2_widths[1251]), .RECT2_HEIGHT(rectangle2_heights[1251]), .RECT2_WEIGHT(rectangle2_weights[1251]), .RECT3_X(rectangle3_xs[1251]), .RECT3_Y(rectangle3_ys[1251]), .RECT3_WIDTH(rectangle3_widths[1251]), .RECT3_HEIGHT(rectangle3_heights[1251]), .RECT3_WEIGHT(rectangle3_weights[1251]), .FEAT_THRES(feature_thresholds[1251]), .FEAT_ABOVE(feature_aboves[1251]), .FEAT_BELOW(feature_belows[1251])) ac1251(.scan_win(scan_win1251), .scan_win_std_dev(scan_win_std_dev[1251]), .feature_accum(feature_accums[1251]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1252]), .RECT1_Y(rectangle1_ys[1252]), .RECT1_WIDTH(rectangle1_widths[1252]), .RECT1_HEIGHT(rectangle1_heights[1252]), .RECT1_WEIGHT(rectangle1_weights[1252]), .RECT2_X(rectangle2_xs[1252]), .RECT2_Y(rectangle2_ys[1252]), .RECT2_WIDTH(rectangle2_widths[1252]), .RECT2_HEIGHT(rectangle2_heights[1252]), .RECT2_WEIGHT(rectangle2_weights[1252]), .RECT3_X(rectangle3_xs[1252]), .RECT3_Y(rectangle3_ys[1252]), .RECT3_WIDTH(rectangle3_widths[1252]), .RECT3_HEIGHT(rectangle3_heights[1252]), .RECT3_WEIGHT(rectangle3_weights[1252]), .FEAT_THRES(feature_thresholds[1252]), .FEAT_ABOVE(feature_aboves[1252]), .FEAT_BELOW(feature_belows[1252])) ac1252(.scan_win(scan_win1252), .scan_win_std_dev(scan_win_std_dev[1252]), .feature_accum(feature_accums[1252]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1253]), .RECT1_Y(rectangle1_ys[1253]), .RECT1_WIDTH(rectangle1_widths[1253]), .RECT1_HEIGHT(rectangle1_heights[1253]), .RECT1_WEIGHT(rectangle1_weights[1253]), .RECT2_X(rectangle2_xs[1253]), .RECT2_Y(rectangle2_ys[1253]), .RECT2_WIDTH(rectangle2_widths[1253]), .RECT2_HEIGHT(rectangle2_heights[1253]), .RECT2_WEIGHT(rectangle2_weights[1253]), .RECT3_X(rectangle3_xs[1253]), .RECT3_Y(rectangle3_ys[1253]), .RECT3_WIDTH(rectangle3_widths[1253]), .RECT3_HEIGHT(rectangle3_heights[1253]), .RECT3_WEIGHT(rectangle3_weights[1253]), .FEAT_THRES(feature_thresholds[1253]), .FEAT_ABOVE(feature_aboves[1253]), .FEAT_BELOW(feature_belows[1253])) ac1253(.scan_win(scan_win1253), .scan_win_std_dev(scan_win_std_dev[1253]), .feature_accum(feature_accums[1253]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1254]), .RECT1_Y(rectangle1_ys[1254]), .RECT1_WIDTH(rectangle1_widths[1254]), .RECT1_HEIGHT(rectangle1_heights[1254]), .RECT1_WEIGHT(rectangle1_weights[1254]), .RECT2_X(rectangle2_xs[1254]), .RECT2_Y(rectangle2_ys[1254]), .RECT2_WIDTH(rectangle2_widths[1254]), .RECT2_HEIGHT(rectangle2_heights[1254]), .RECT2_WEIGHT(rectangle2_weights[1254]), .RECT3_X(rectangle3_xs[1254]), .RECT3_Y(rectangle3_ys[1254]), .RECT3_WIDTH(rectangle3_widths[1254]), .RECT3_HEIGHT(rectangle3_heights[1254]), .RECT3_WEIGHT(rectangle3_weights[1254]), .FEAT_THRES(feature_thresholds[1254]), .FEAT_ABOVE(feature_aboves[1254]), .FEAT_BELOW(feature_belows[1254])) ac1254(.scan_win(scan_win1254), .scan_win_std_dev(scan_win_std_dev[1254]), .feature_accum(feature_accums[1254]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1255]), .RECT1_Y(rectangle1_ys[1255]), .RECT1_WIDTH(rectangle1_widths[1255]), .RECT1_HEIGHT(rectangle1_heights[1255]), .RECT1_WEIGHT(rectangle1_weights[1255]), .RECT2_X(rectangle2_xs[1255]), .RECT2_Y(rectangle2_ys[1255]), .RECT2_WIDTH(rectangle2_widths[1255]), .RECT2_HEIGHT(rectangle2_heights[1255]), .RECT2_WEIGHT(rectangle2_weights[1255]), .RECT3_X(rectangle3_xs[1255]), .RECT3_Y(rectangle3_ys[1255]), .RECT3_WIDTH(rectangle3_widths[1255]), .RECT3_HEIGHT(rectangle3_heights[1255]), .RECT3_WEIGHT(rectangle3_weights[1255]), .FEAT_THRES(feature_thresholds[1255]), .FEAT_ABOVE(feature_aboves[1255]), .FEAT_BELOW(feature_belows[1255])) ac1255(.scan_win(scan_win1255), .scan_win_std_dev(scan_win_std_dev[1255]), .feature_accum(feature_accums[1255]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1256]), .RECT1_Y(rectangle1_ys[1256]), .RECT1_WIDTH(rectangle1_widths[1256]), .RECT1_HEIGHT(rectangle1_heights[1256]), .RECT1_WEIGHT(rectangle1_weights[1256]), .RECT2_X(rectangle2_xs[1256]), .RECT2_Y(rectangle2_ys[1256]), .RECT2_WIDTH(rectangle2_widths[1256]), .RECT2_HEIGHT(rectangle2_heights[1256]), .RECT2_WEIGHT(rectangle2_weights[1256]), .RECT3_X(rectangle3_xs[1256]), .RECT3_Y(rectangle3_ys[1256]), .RECT3_WIDTH(rectangle3_widths[1256]), .RECT3_HEIGHT(rectangle3_heights[1256]), .RECT3_WEIGHT(rectangle3_weights[1256]), .FEAT_THRES(feature_thresholds[1256]), .FEAT_ABOVE(feature_aboves[1256]), .FEAT_BELOW(feature_belows[1256])) ac1256(.scan_win(scan_win1256), .scan_win_std_dev(scan_win_std_dev[1256]), .feature_accum(feature_accums[1256]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1257]), .RECT1_Y(rectangle1_ys[1257]), .RECT1_WIDTH(rectangle1_widths[1257]), .RECT1_HEIGHT(rectangle1_heights[1257]), .RECT1_WEIGHT(rectangle1_weights[1257]), .RECT2_X(rectangle2_xs[1257]), .RECT2_Y(rectangle2_ys[1257]), .RECT2_WIDTH(rectangle2_widths[1257]), .RECT2_HEIGHT(rectangle2_heights[1257]), .RECT2_WEIGHT(rectangle2_weights[1257]), .RECT3_X(rectangle3_xs[1257]), .RECT3_Y(rectangle3_ys[1257]), .RECT3_WIDTH(rectangle3_widths[1257]), .RECT3_HEIGHT(rectangle3_heights[1257]), .RECT3_WEIGHT(rectangle3_weights[1257]), .FEAT_THRES(feature_thresholds[1257]), .FEAT_ABOVE(feature_aboves[1257]), .FEAT_BELOW(feature_belows[1257])) ac1257(.scan_win(scan_win1257), .scan_win_std_dev(scan_win_std_dev[1257]), .feature_accum(feature_accums[1257]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1258]), .RECT1_Y(rectangle1_ys[1258]), .RECT1_WIDTH(rectangle1_widths[1258]), .RECT1_HEIGHT(rectangle1_heights[1258]), .RECT1_WEIGHT(rectangle1_weights[1258]), .RECT2_X(rectangle2_xs[1258]), .RECT2_Y(rectangle2_ys[1258]), .RECT2_WIDTH(rectangle2_widths[1258]), .RECT2_HEIGHT(rectangle2_heights[1258]), .RECT2_WEIGHT(rectangle2_weights[1258]), .RECT3_X(rectangle3_xs[1258]), .RECT3_Y(rectangle3_ys[1258]), .RECT3_WIDTH(rectangle3_widths[1258]), .RECT3_HEIGHT(rectangle3_heights[1258]), .RECT3_WEIGHT(rectangle3_weights[1258]), .FEAT_THRES(feature_thresholds[1258]), .FEAT_ABOVE(feature_aboves[1258]), .FEAT_BELOW(feature_belows[1258])) ac1258(.scan_win(scan_win1258), .scan_win_std_dev(scan_win_std_dev[1258]), .feature_accum(feature_accums[1258]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1259]), .RECT1_Y(rectangle1_ys[1259]), .RECT1_WIDTH(rectangle1_widths[1259]), .RECT1_HEIGHT(rectangle1_heights[1259]), .RECT1_WEIGHT(rectangle1_weights[1259]), .RECT2_X(rectangle2_xs[1259]), .RECT2_Y(rectangle2_ys[1259]), .RECT2_WIDTH(rectangle2_widths[1259]), .RECT2_HEIGHT(rectangle2_heights[1259]), .RECT2_WEIGHT(rectangle2_weights[1259]), .RECT3_X(rectangle3_xs[1259]), .RECT3_Y(rectangle3_ys[1259]), .RECT3_WIDTH(rectangle3_widths[1259]), .RECT3_HEIGHT(rectangle3_heights[1259]), .RECT3_WEIGHT(rectangle3_weights[1259]), .FEAT_THRES(feature_thresholds[1259]), .FEAT_ABOVE(feature_aboves[1259]), .FEAT_BELOW(feature_belows[1259])) ac1259(.scan_win(scan_win1259), .scan_win_std_dev(scan_win_std_dev[1259]), .feature_accum(feature_accums[1259]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1260]), .RECT1_Y(rectangle1_ys[1260]), .RECT1_WIDTH(rectangle1_widths[1260]), .RECT1_HEIGHT(rectangle1_heights[1260]), .RECT1_WEIGHT(rectangle1_weights[1260]), .RECT2_X(rectangle2_xs[1260]), .RECT2_Y(rectangle2_ys[1260]), .RECT2_WIDTH(rectangle2_widths[1260]), .RECT2_HEIGHT(rectangle2_heights[1260]), .RECT2_WEIGHT(rectangle2_weights[1260]), .RECT3_X(rectangle3_xs[1260]), .RECT3_Y(rectangle3_ys[1260]), .RECT3_WIDTH(rectangle3_widths[1260]), .RECT3_HEIGHT(rectangle3_heights[1260]), .RECT3_WEIGHT(rectangle3_weights[1260]), .FEAT_THRES(feature_thresholds[1260]), .FEAT_ABOVE(feature_aboves[1260]), .FEAT_BELOW(feature_belows[1260])) ac1260(.scan_win(scan_win1260), .scan_win_std_dev(scan_win_std_dev[1260]), .feature_accum(feature_accums[1260]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1261]), .RECT1_Y(rectangle1_ys[1261]), .RECT1_WIDTH(rectangle1_widths[1261]), .RECT1_HEIGHT(rectangle1_heights[1261]), .RECT1_WEIGHT(rectangle1_weights[1261]), .RECT2_X(rectangle2_xs[1261]), .RECT2_Y(rectangle2_ys[1261]), .RECT2_WIDTH(rectangle2_widths[1261]), .RECT2_HEIGHT(rectangle2_heights[1261]), .RECT2_WEIGHT(rectangle2_weights[1261]), .RECT3_X(rectangle3_xs[1261]), .RECT3_Y(rectangle3_ys[1261]), .RECT3_WIDTH(rectangle3_widths[1261]), .RECT3_HEIGHT(rectangle3_heights[1261]), .RECT3_WEIGHT(rectangle3_weights[1261]), .FEAT_THRES(feature_thresholds[1261]), .FEAT_ABOVE(feature_aboves[1261]), .FEAT_BELOW(feature_belows[1261])) ac1261(.scan_win(scan_win1261), .scan_win_std_dev(scan_win_std_dev[1261]), .feature_accum(feature_accums[1261]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1262]), .RECT1_Y(rectangle1_ys[1262]), .RECT1_WIDTH(rectangle1_widths[1262]), .RECT1_HEIGHT(rectangle1_heights[1262]), .RECT1_WEIGHT(rectangle1_weights[1262]), .RECT2_X(rectangle2_xs[1262]), .RECT2_Y(rectangle2_ys[1262]), .RECT2_WIDTH(rectangle2_widths[1262]), .RECT2_HEIGHT(rectangle2_heights[1262]), .RECT2_WEIGHT(rectangle2_weights[1262]), .RECT3_X(rectangle3_xs[1262]), .RECT3_Y(rectangle3_ys[1262]), .RECT3_WIDTH(rectangle3_widths[1262]), .RECT3_HEIGHT(rectangle3_heights[1262]), .RECT3_WEIGHT(rectangle3_weights[1262]), .FEAT_THRES(feature_thresholds[1262]), .FEAT_ABOVE(feature_aboves[1262]), .FEAT_BELOW(feature_belows[1262])) ac1262(.scan_win(scan_win1262), .scan_win_std_dev(scan_win_std_dev[1262]), .feature_accum(feature_accums[1262]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1263]), .RECT1_Y(rectangle1_ys[1263]), .RECT1_WIDTH(rectangle1_widths[1263]), .RECT1_HEIGHT(rectangle1_heights[1263]), .RECT1_WEIGHT(rectangle1_weights[1263]), .RECT2_X(rectangle2_xs[1263]), .RECT2_Y(rectangle2_ys[1263]), .RECT2_WIDTH(rectangle2_widths[1263]), .RECT2_HEIGHT(rectangle2_heights[1263]), .RECT2_WEIGHT(rectangle2_weights[1263]), .RECT3_X(rectangle3_xs[1263]), .RECT3_Y(rectangle3_ys[1263]), .RECT3_WIDTH(rectangle3_widths[1263]), .RECT3_HEIGHT(rectangle3_heights[1263]), .RECT3_WEIGHT(rectangle3_weights[1263]), .FEAT_THRES(feature_thresholds[1263]), .FEAT_ABOVE(feature_aboves[1263]), .FEAT_BELOW(feature_belows[1263])) ac1263(.scan_win(scan_win1263), .scan_win_std_dev(scan_win_std_dev[1263]), .feature_accum(feature_accums[1263]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1264]), .RECT1_Y(rectangle1_ys[1264]), .RECT1_WIDTH(rectangle1_widths[1264]), .RECT1_HEIGHT(rectangle1_heights[1264]), .RECT1_WEIGHT(rectangle1_weights[1264]), .RECT2_X(rectangle2_xs[1264]), .RECT2_Y(rectangle2_ys[1264]), .RECT2_WIDTH(rectangle2_widths[1264]), .RECT2_HEIGHT(rectangle2_heights[1264]), .RECT2_WEIGHT(rectangle2_weights[1264]), .RECT3_X(rectangle3_xs[1264]), .RECT3_Y(rectangle3_ys[1264]), .RECT3_WIDTH(rectangle3_widths[1264]), .RECT3_HEIGHT(rectangle3_heights[1264]), .RECT3_WEIGHT(rectangle3_weights[1264]), .FEAT_THRES(feature_thresholds[1264]), .FEAT_ABOVE(feature_aboves[1264]), .FEAT_BELOW(feature_belows[1264])) ac1264(.scan_win(scan_win1264), .scan_win_std_dev(scan_win_std_dev[1264]), .feature_accum(feature_accums[1264]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1265]), .RECT1_Y(rectangle1_ys[1265]), .RECT1_WIDTH(rectangle1_widths[1265]), .RECT1_HEIGHT(rectangle1_heights[1265]), .RECT1_WEIGHT(rectangle1_weights[1265]), .RECT2_X(rectangle2_xs[1265]), .RECT2_Y(rectangle2_ys[1265]), .RECT2_WIDTH(rectangle2_widths[1265]), .RECT2_HEIGHT(rectangle2_heights[1265]), .RECT2_WEIGHT(rectangle2_weights[1265]), .RECT3_X(rectangle3_xs[1265]), .RECT3_Y(rectangle3_ys[1265]), .RECT3_WIDTH(rectangle3_widths[1265]), .RECT3_HEIGHT(rectangle3_heights[1265]), .RECT3_WEIGHT(rectangle3_weights[1265]), .FEAT_THRES(feature_thresholds[1265]), .FEAT_ABOVE(feature_aboves[1265]), .FEAT_BELOW(feature_belows[1265])) ac1265(.scan_win(scan_win1265), .scan_win_std_dev(scan_win_std_dev[1265]), .feature_accum(feature_accums[1265]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1266]), .RECT1_Y(rectangle1_ys[1266]), .RECT1_WIDTH(rectangle1_widths[1266]), .RECT1_HEIGHT(rectangle1_heights[1266]), .RECT1_WEIGHT(rectangle1_weights[1266]), .RECT2_X(rectangle2_xs[1266]), .RECT2_Y(rectangle2_ys[1266]), .RECT2_WIDTH(rectangle2_widths[1266]), .RECT2_HEIGHT(rectangle2_heights[1266]), .RECT2_WEIGHT(rectangle2_weights[1266]), .RECT3_X(rectangle3_xs[1266]), .RECT3_Y(rectangle3_ys[1266]), .RECT3_WIDTH(rectangle3_widths[1266]), .RECT3_HEIGHT(rectangle3_heights[1266]), .RECT3_WEIGHT(rectangle3_weights[1266]), .FEAT_THRES(feature_thresholds[1266]), .FEAT_ABOVE(feature_aboves[1266]), .FEAT_BELOW(feature_belows[1266])) ac1266(.scan_win(scan_win1266), .scan_win_std_dev(scan_win_std_dev[1266]), .feature_accum(feature_accums[1266]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1267]), .RECT1_Y(rectangle1_ys[1267]), .RECT1_WIDTH(rectangle1_widths[1267]), .RECT1_HEIGHT(rectangle1_heights[1267]), .RECT1_WEIGHT(rectangle1_weights[1267]), .RECT2_X(rectangle2_xs[1267]), .RECT2_Y(rectangle2_ys[1267]), .RECT2_WIDTH(rectangle2_widths[1267]), .RECT2_HEIGHT(rectangle2_heights[1267]), .RECT2_WEIGHT(rectangle2_weights[1267]), .RECT3_X(rectangle3_xs[1267]), .RECT3_Y(rectangle3_ys[1267]), .RECT3_WIDTH(rectangle3_widths[1267]), .RECT3_HEIGHT(rectangle3_heights[1267]), .RECT3_WEIGHT(rectangle3_weights[1267]), .FEAT_THRES(feature_thresholds[1267]), .FEAT_ABOVE(feature_aboves[1267]), .FEAT_BELOW(feature_belows[1267])) ac1267(.scan_win(scan_win1267), .scan_win_std_dev(scan_win_std_dev[1267]), .feature_accum(feature_accums[1267]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1268]), .RECT1_Y(rectangle1_ys[1268]), .RECT1_WIDTH(rectangle1_widths[1268]), .RECT1_HEIGHT(rectangle1_heights[1268]), .RECT1_WEIGHT(rectangle1_weights[1268]), .RECT2_X(rectangle2_xs[1268]), .RECT2_Y(rectangle2_ys[1268]), .RECT2_WIDTH(rectangle2_widths[1268]), .RECT2_HEIGHT(rectangle2_heights[1268]), .RECT2_WEIGHT(rectangle2_weights[1268]), .RECT3_X(rectangle3_xs[1268]), .RECT3_Y(rectangle3_ys[1268]), .RECT3_WIDTH(rectangle3_widths[1268]), .RECT3_HEIGHT(rectangle3_heights[1268]), .RECT3_WEIGHT(rectangle3_weights[1268]), .FEAT_THRES(feature_thresholds[1268]), .FEAT_ABOVE(feature_aboves[1268]), .FEAT_BELOW(feature_belows[1268])) ac1268(.scan_win(scan_win1268), .scan_win_std_dev(scan_win_std_dev[1268]), .feature_accum(feature_accums[1268]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1269]), .RECT1_Y(rectangle1_ys[1269]), .RECT1_WIDTH(rectangle1_widths[1269]), .RECT1_HEIGHT(rectangle1_heights[1269]), .RECT1_WEIGHT(rectangle1_weights[1269]), .RECT2_X(rectangle2_xs[1269]), .RECT2_Y(rectangle2_ys[1269]), .RECT2_WIDTH(rectangle2_widths[1269]), .RECT2_HEIGHT(rectangle2_heights[1269]), .RECT2_WEIGHT(rectangle2_weights[1269]), .RECT3_X(rectangle3_xs[1269]), .RECT3_Y(rectangle3_ys[1269]), .RECT3_WIDTH(rectangle3_widths[1269]), .RECT3_HEIGHT(rectangle3_heights[1269]), .RECT3_WEIGHT(rectangle3_weights[1269]), .FEAT_THRES(feature_thresholds[1269]), .FEAT_ABOVE(feature_aboves[1269]), .FEAT_BELOW(feature_belows[1269])) ac1269(.scan_win(scan_win1269), .scan_win_std_dev(scan_win_std_dev[1269]), .feature_accum(feature_accums[1269]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1270]), .RECT1_Y(rectangle1_ys[1270]), .RECT1_WIDTH(rectangle1_widths[1270]), .RECT1_HEIGHT(rectangle1_heights[1270]), .RECT1_WEIGHT(rectangle1_weights[1270]), .RECT2_X(rectangle2_xs[1270]), .RECT2_Y(rectangle2_ys[1270]), .RECT2_WIDTH(rectangle2_widths[1270]), .RECT2_HEIGHT(rectangle2_heights[1270]), .RECT2_WEIGHT(rectangle2_weights[1270]), .RECT3_X(rectangle3_xs[1270]), .RECT3_Y(rectangle3_ys[1270]), .RECT3_WIDTH(rectangle3_widths[1270]), .RECT3_HEIGHT(rectangle3_heights[1270]), .RECT3_WEIGHT(rectangle3_weights[1270]), .FEAT_THRES(feature_thresholds[1270]), .FEAT_ABOVE(feature_aboves[1270]), .FEAT_BELOW(feature_belows[1270])) ac1270(.scan_win(scan_win1270), .scan_win_std_dev(scan_win_std_dev[1270]), .feature_accum(feature_accums[1270]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1271]), .RECT1_Y(rectangle1_ys[1271]), .RECT1_WIDTH(rectangle1_widths[1271]), .RECT1_HEIGHT(rectangle1_heights[1271]), .RECT1_WEIGHT(rectangle1_weights[1271]), .RECT2_X(rectangle2_xs[1271]), .RECT2_Y(rectangle2_ys[1271]), .RECT2_WIDTH(rectangle2_widths[1271]), .RECT2_HEIGHT(rectangle2_heights[1271]), .RECT2_WEIGHT(rectangle2_weights[1271]), .RECT3_X(rectangle3_xs[1271]), .RECT3_Y(rectangle3_ys[1271]), .RECT3_WIDTH(rectangle3_widths[1271]), .RECT3_HEIGHT(rectangle3_heights[1271]), .RECT3_WEIGHT(rectangle3_weights[1271]), .FEAT_THRES(feature_thresholds[1271]), .FEAT_ABOVE(feature_aboves[1271]), .FEAT_BELOW(feature_belows[1271])) ac1271(.scan_win(scan_win1271), .scan_win_std_dev(scan_win_std_dev[1271]), .feature_accum(feature_accums[1271]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1272]), .RECT1_Y(rectangle1_ys[1272]), .RECT1_WIDTH(rectangle1_widths[1272]), .RECT1_HEIGHT(rectangle1_heights[1272]), .RECT1_WEIGHT(rectangle1_weights[1272]), .RECT2_X(rectangle2_xs[1272]), .RECT2_Y(rectangle2_ys[1272]), .RECT2_WIDTH(rectangle2_widths[1272]), .RECT2_HEIGHT(rectangle2_heights[1272]), .RECT2_WEIGHT(rectangle2_weights[1272]), .RECT3_X(rectangle3_xs[1272]), .RECT3_Y(rectangle3_ys[1272]), .RECT3_WIDTH(rectangle3_widths[1272]), .RECT3_HEIGHT(rectangle3_heights[1272]), .RECT3_WEIGHT(rectangle3_weights[1272]), .FEAT_THRES(feature_thresholds[1272]), .FEAT_ABOVE(feature_aboves[1272]), .FEAT_BELOW(feature_belows[1272])) ac1272(.scan_win(scan_win1272), .scan_win_std_dev(scan_win_std_dev[1272]), .feature_accum(feature_accums[1272]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1273]), .RECT1_Y(rectangle1_ys[1273]), .RECT1_WIDTH(rectangle1_widths[1273]), .RECT1_HEIGHT(rectangle1_heights[1273]), .RECT1_WEIGHT(rectangle1_weights[1273]), .RECT2_X(rectangle2_xs[1273]), .RECT2_Y(rectangle2_ys[1273]), .RECT2_WIDTH(rectangle2_widths[1273]), .RECT2_HEIGHT(rectangle2_heights[1273]), .RECT2_WEIGHT(rectangle2_weights[1273]), .RECT3_X(rectangle3_xs[1273]), .RECT3_Y(rectangle3_ys[1273]), .RECT3_WIDTH(rectangle3_widths[1273]), .RECT3_HEIGHT(rectangle3_heights[1273]), .RECT3_WEIGHT(rectangle3_weights[1273]), .FEAT_THRES(feature_thresholds[1273]), .FEAT_ABOVE(feature_aboves[1273]), .FEAT_BELOW(feature_belows[1273])) ac1273(.scan_win(scan_win1273), .scan_win_std_dev(scan_win_std_dev[1273]), .feature_accum(feature_accums[1273]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1274]), .RECT1_Y(rectangle1_ys[1274]), .RECT1_WIDTH(rectangle1_widths[1274]), .RECT1_HEIGHT(rectangle1_heights[1274]), .RECT1_WEIGHT(rectangle1_weights[1274]), .RECT2_X(rectangle2_xs[1274]), .RECT2_Y(rectangle2_ys[1274]), .RECT2_WIDTH(rectangle2_widths[1274]), .RECT2_HEIGHT(rectangle2_heights[1274]), .RECT2_WEIGHT(rectangle2_weights[1274]), .RECT3_X(rectangle3_xs[1274]), .RECT3_Y(rectangle3_ys[1274]), .RECT3_WIDTH(rectangle3_widths[1274]), .RECT3_HEIGHT(rectangle3_heights[1274]), .RECT3_WEIGHT(rectangle3_weights[1274]), .FEAT_THRES(feature_thresholds[1274]), .FEAT_ABOVE(feature_aboves[1274]), .FEAT_BELOW(feature_belows[1274])) ac1274(.scan_win(scan_win1274), .scan_win_std_dev(scan_win_std_dev[1274]), .feature_accum(feature_accums[1274]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1275]), .RECT1_Y(rectangle1_ys[1275]), .RECT1_WIDTH(rectangle1_widths[1275]), .RECT1_HEIGHT(rectangle1_heights[1275]), .RECT1_WEIGHT(rectangle1_weights[1275]), .RECT2_X(rectangle2_xs[1275]), .RECT2_Y(rectangle2_ys[1275]), .RECT2_WIDTH(rectangle2_widths[1275]), .RECT2_HEIGHT(rectangle2_heights[1275]), .RECT2_WEIGHT(rectangle2_weights[1275]), .RECT3_X(rectangle3_xs[1275]), .RECT3_Y(rectangle3_ys[1275]), .RECT3_WIDTH(rectangle3_widths[1275]), .RECT3_HEIGHT(rectangle3_heights[1275]), .RECT3_WEIGHT(rectangle3_weights[1275]), .FEAT_THRES(feature_thresholds[1275]), .FEAT_ABOVE(feature_aboves[1275]), .FEAT_BELOW(feature_belows[1275])) ac1275(.scan_win(scan_win1275), .scan_win_std_dev(scan_win_std_dev[1275]), .feature_accum(feature_accums[1275]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1276]), .RECT1_Y(rectangle1_ys[1276]), .RECT1_WIDTH(rectangle1_widths[1276]), .RECT1_HEIGHT(rectangle1_heights[1276]), .RECT1_WEIGHT(rectangle1_weights[1276]), .RECT2_X(rectangle2_xs[1276]), .RECT2_Y(rectangle2_ys[1276]), .RECT2_WIDTH(rectangle2_widths[1276]), .RECT2_HEIGHT(rectangle2_heights[1276]), .RECT2_WEIGHT(rectangle2_weights[1276]), .RECT3_X(rectangle3_xs[1276]), .RECT3_Y(rectangle3_ys[1276]), .RECT3_WIDTH(rectangle3_widths[1276]), .RECT3_HEIGHT(rectangle3_heights[1276]), .RECT3_WEIGHT(rectangle3_weights[1276]), .FEAT_THRES(feature_thresholds[1276]), .FEAT_ABOVE(feature_aboves[1276]), .FEAT_BELOW(feature_belows[1276])) ac1276(.scan_win(scan_win1276), .scan_win_std_dev(scan_win_std_dev[1276]), .feature_accum(feature_accums[1276]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1277]), .RECT1_Y(rectangle1_ys[1277]), .RECT1_WIDTH(rectangle1_widths[1277]), .RECT1_HEIGHT(rectangle1_heights[1277]), .RECT1_WEIGHT(rectangle1_weights[1277]), .RECT2_X(rectangle2_xs[1277]), .RECT2_Y(rectangle2_ys[1277]), .RECT2_WIDTH(rectangle2_widths[1277]), .RECT2_HEIGHT(rectangle2_heights[1277]), .RECT2_WEIGHT(rectangle2_weights[1277]), .RECT3_X(rectangle3_xs[1277]), .RECT3_Y(rectangle3_ys[1277]), .RECT3_WIDTH(rectangle3_widths[1277]), .RECT3_HEIGHT(rectangle3_heights[1277]), .RECT3_WEIGHT(rectangle3_weights[1277]), .FEAT_THRES(feature_thresholds[1277]), .FEAT_ABOVE(feature_aboves[1277]), .FEAT_BELOW(feature_belows[1277])) ac1277(.scan_win(scan_win1277), .scan_win_std_dev(scan_win_std_dev[1277]), .feature_accum(feature_accums[1277]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1278]), .RECT1_Y(rectangle1_ys[1278]), .RECT1_WIDTH(rectangle1_widths[1278]), .RECT1_HEIGHT(rectangle1_heights[1278]), .RECT1_WEIGHT(rectangle1_weights[1278]), .RECT2_X(rectangle2_xs[1278]), .RECT2_Y(rectangle2_ys[1278]), .RECT2_WIDTH(rectangle2_widths[1278]), .RECT2_HEIGHT(rectangle2_heights[1278]), .RECT2_WEIGHT(rectangle2_weights[1278]), .RECT3_X(rectangle3_xs[1278]), .RECT3_Y(rectangle3_ys[1278]), .RECT3_WIDTH(rectangle3_widths[1278]), .RECT3_HEIGHT(rectangle3_heights[1278]), .RECT3_WEIGHT(rectangle3_weights[1278]), .FEAT_THRES(feature_thresholds[1278]), .FEAT_ABOVE(feature_aboves[1278]), .FEAT_BELOW(feature_belows[1278])) ac1278(.scan_win(scan_win1278), .scan_win_std_dev(scan_win_std_dev[1278]), .feature_accum(feature_accums[1278]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1279]), .RECT1_Y(rectangle1_ys[1279]), .RECT1_WIDTH(rectangle1_widths[1279]), .RECT1_HEIGHT(rectangle1_heights[1279]), .RECT1_WEIGHT(rectangle1_weights[1279]), .RECT2_X(rectangle2_xs[1279]), .RECT2_Y(rectangle2_ys[1279]), .RECT2_WIDTH(rectangle2_widths[1279]), .RECT2_HEIGHT(rectangle2_heights[1279]), .RECT2_WEIGHT(rectangle2_weights[1279]), .RECT3_X(rectangle3_xs[1279]), .RECT3_Y(rectangle3_ys[1279]), .RECT3_WIDTH(rectangle3_widths[1279]), .RECT3_HEIGHT(rectangle3_heights[1279]), .RECT3_WEIGHT(rectangle3_weights[1279]), .FEAT_THRES(feature_thresholds[1279]), .FEAT_ABOVE(feature_aboves[1279]), .FEAT_BELOW(feature_belows[1279])) ac1279(.scan_win(scan_win1279), .scan_win_std_dev(scan_win_std_dev[1279]), .feature_accum(feature_accums[1279]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1280]), .RECT1_Y(rectangle1_ys[1280]), .RECT1_WIDTH(rectangle1_widths[1280]), .RECT1_HEIGHT(rectangle1_heights[1280]), .RECT1_WEIGHT(rectangle1_weights[1280]), .RECT2_X(rectangle2_xs[1280]), .RECT2_Y(rectangle2_ys[1280]), .RECT2_WIDTH(rectangle2_widths[1280]), .RECT2_HEIGHT(rectangle2_heights[1280]), .RECT2_WEIGHT(rectangle2_weights[1280]), .RECT3_X(rectangle3_xs[1280]), .RECT3_Y(rectangle3_ys[1280]), .RECT3_WIDTH(rectangle3_widths[1280]), .RECT3_HEIGHT(rectangle3_heights[1280]), .RECT3_WEIGHT(rectangle3_weights[1280]), .FEAT_THRES(feature_thresholds[1280]), .FEAT_ABOVE(feature_aboves[1280]), .FEAT_BELOW(feature_belows[1280])) ac1280(.scan_win(scan_win1280), .scan_win_std_dev(scan_win_std_dev[1280]), .feature_accum(feature_accums[1280]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1281]), .RECT1_Y(rectangle1_ys[1281]), .RECT1_WIDTH(rectangle1_widths[1281]), .RECT1_HEIGHT(rectangle1_heights[1281]), .RECT1_WEIGHT(rectangle1_weights[1281]), .RECT2_X(rectangle2_xs[1281]), .RECT2_Y(rectangle2_ys[1281]), .RECT2_WIDTH(rectangle2_widths[1281]), .RECT2_HEIGHT(rectangle2_heights[1281]), .RECT2_WEIGHT(rectangle2_weights[1281]), .RECT3_X(rectangle3_xs[1281]), .RECT3_Y(rectangle3_ys[1281]), .RECT3_WIDTH(rectangle3_widths[1281]), .RECT3_HEIGHT(rectangle3_heights[1281]), .RECT3_WEIGHT(rectangle3_weights[1281]), .FEAT_THRES(feature_thresholds[1281]), .FEAT_ABOVE(feature_aboves[1281]), .FEAT_BELOW(feature_belows[1281])) ac1281(.scan_win(scan_win1281), .scan_win_std_dev(scan_win_std_dev[1281]), .feature_accum(feature_accums[1281]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1282]), .RECT1_Y(rectangle1_ys[1282]), .RECT1_WIDTH(rectangle1_widths[1282]), .RECT1_HEIGHT(rectangle1_heights[1282]), .RECT1_WEIGHT(rectangle1_weights[1282]), .RECT2_X(rectangle2_xs[1282]), .RECT2_Y(rectangle2_ys[1282]), .RECT2_WIDTH(rectangle2_widths[1282]), .RECT2_HEIGHT(rectangle2_heights[1282]), .RECT2_WEIGHT(rectangle2_weights[1282]), .RECT3_X(rectangle3_xs[1282]), .RECT3_Y(rectangle3_ys[1282]), .RECT3_WIDTH(rectangle3_widths[1282]), .RECT3_HEIGHT(rectangle3_heights[1282]), .RECT3_WEIGHT(rectangle3_weights[1282]), .FEAT_THRES(feature_thresholds[1282]), .FEAT_ABOVE(feature_aboves[1282]), .FEAT_BELOW(feature_belows[1282])) ac1282(.scan_win(scan_win1282), .scan_win_std_dev(scan_win_std_dev[1282]), .feature_accum(feature_accums[1282]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1283]), .RECT1_Y(rectangle1_ys[1283]), .RECT1_WIDTH(rectangle1_widths[1283]), .RECT1_HEIGHT(rectangle1_heights[1283]), .RECT1_WEIGHT(rectangle1_weights[1283]), .RECT2_X(rectangle2_xs[1283]), .RECT2_Y(rectangle2_ys[1283]), .RECT2_WIDTH(rectangle2_widths[1283]), .RECT2_HEIGHT(rectangle2_heights[1283]), .RECT2_WEIGHT(rectangle2_weights[1283]), .RECT3_X(rectangle3_xs[1283]), .RECT3_Y(rectangle3_ys[1283]), .RECT3_WIDTH(rectangle3_widths[1283]), .RECT3_HEIGHT(rectangle3_heights[1283]), .RECT3_WEIGHT(rectangle3_weights[1283]), .FEAT_THRES(feature_thresholds[1283]), .FEAT_ABOVE(feature_aboves[1283]), .FEAT_BELOW(feature_belows[1283])) ac1283(.scan_win(scan_win1283), .scan_win_std_dev(scan_win_std_dev[1283]), .feature_accum(feature_accums[1283]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1284]), .RECT1_Y(rectangle1_ys[1284]), .RECT1_WIDTH(rectangle1_widths[1284]), .RECT1_HEIGHT(rectangle1_heights[1284]), .RECT1_WEIGHT(rectangle1_weights[1284]), .RECT2_X(rectangle2_xs[1284]), .RECT2_Y(rectangle2_ys[1284]), .RECT2_WIDTH(rectangle2_widths[1284]), .RECT2_HEIGHT(rectangle2_heights[1284]), .RECT2_WEIGHT(rectangle2_weights[1284]), .RECT3_X(rectangle3_xs[1284]), .RECT3_Y(rectangle3_ys[1284]), .RECT3_WIDTH(rectangle3_widths[1284]), .RECT3_HEIGHT(rectangle3_heights[1284]), .RECT3_WEIGHT(rectangle3_weights[1284]), .FEAT_THRES(feature_thresholds[1284]), .FEAT_ABOVE(feature_aboves[1284]), .FEAT_BELOW(feature_belows[1284])) ac1284(.scan_win(scan_win1284), .scan_win_std_dev(scan_win_std_dev[1284]), .feature_accum(feature_accums[1284]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1285]), .RECT1_Y(rectangle1_ys[1285]), .RECT1_WIDTH(rectangle1_widths[1285]), .RECT1_HEIGHT(rectangle1_heights[1285]), .RECT1_WEIGHT(rectangle1_weights[1285]), .RECT2_X(rectangle2_xs[1285]), .RECT2_Y(rectangle2_ys[1285]), .RECT2_WIDTH(rectangle2_widths[1285]), .RECT2_HEIGHT(rectangle2_heights[1285]), .RECT2_WEIGHT(rectangle2_weights[1285]), .RECT3_X(rectangle3_xs[1285]), .RECT3_Y(rectangle3_ys[1285]), .RECT3_WIDTH(rectangle3_widths[1285]), .RECT3_HEIGHT(rectangle3_heights[1285]), .RECT3_WEIGHT(rectangle3_weights[1285]), .FEAT_THRES(feature_thresholds[1285]), .FEAT_ABOVE(feature_aboves[1285]), .FEAT_BELOW(feature_belows[1285])) ac1285(.scan_win(scan_win1285), .scan_win_std_dev(scan_win_std_dev[1285]), .feature_accum(feature_accums[1285]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1286]), .RECT1_Y(rectangle1_ys[1286]), .RECT1_WIDTH(rectangle1_widths[1286]), .RECT1_HEIGHT(rectangle1_heights[1286]), .RECT1_WEIGHT(rectangle1_weights[1286]), .RECT2_X(rectangle2_xs[1286]), .RECT2_Y(rectangle2_ys[1286]), .RECT2_WIDTH(rectangle2_widths[1286]), .RECT2_HEIGHT(rectangle2_heights[1286]), .RECT2_WEIGHT(rectangle2_weights[1286]), .RECT3_X(rectangle3_xs[1286]), .RECT3_Y(rectangle3_ys[1286]), .RECT3_WIDTH(rectangle3_widths[1286]), .RECT3_HEIGHT(rectangle3_heights[1286]), .RECT3_WEIGHT(rectangle3_weights[1286]), .FEAT_THRES(feature_thresholds[1286]), .FEAT_ABOVE(feature_aboves[1286]), .FEAT_BELOW(feature_belows[1286])) ac1286(.scan_win(scan_win1286), .scan_win_std_dev(scan_win_std_dev[1286]), .feature_accum(feature_accums[1286]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1287]), .RECT1_Y(rectangle1_ys[1287]), .RECT1_WIDTH(rectangle1_widths[1287]), .RECT1_HEIGHT(rectangle1_heights[1287]), .RECT1_WEIGHT(rectangle1_weights[1287]), .RECT2_X(rectangle2_xs[1287]), .RECT2_Y(rectangle2_ys[1287]), .RECT2_WIDTH(rectangle2_widths[1287]), .RECT2_HEIGHT(rectangle2_heights[1287]), .RECT2_WEIGHT(rectangle2_weights[1287]), .RECT3_X(rectangle3_xs[1287]), .RECT3_Y(rectangle3_ys[1287]), .RECT3_WIDTH(rectangle3_widths[1287]), .RECT3_HEIGHT(rectangle3_heights[1287]), .RECT3_WEIGHT(rectangle3_weights[1287]), .FEAT_THRES(feature_thresholds[1287]), .FEAT_ABOVE(feature_aboves[1287]), .FEAT_BELOW(feature_belows[1287])) ac1287(.scan_win(scan_win1287), .scan_win_std_dev(scan_win_std_dev[1287]), .feature_accum(feature_accums[1287]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1288]), .RECT1_Y(rectangle1_ys[1288]), .RECT1_WIDTH(rectangle1_widths[1288]), .RECT1_HEIGHT(rectangle1_heights[1288]), .RECT1_WEIGHT(rectangle1_weights[1288]), .RECT2_X(rectangle2_xs[1288]), .RECT2_Y(rectangle2_ys[1288]), .RECT2_WIDTH(rectangle2_widths[1288]), .RECT2_HEIGHT(rectangle2_heights[1288]), .RECT2_WEIGHT(rectangle2_weights[1288]), .RECT3_X(rectangle3_xs[1288]), .RECT3_Y(rectangle3_ys[1288]), .RECT3_WIDTH(rectangle3_widths[1288]), .RECT3_HEIGHT(rectangle3_heights[1288]), .RECT3_WEIGHT(rectangle3_weights[1288]), .FEAT_THRES(feature_thresholds[1288]), .FEAT_ABOVE(feature_aboves[1288]), .FEAT_BELOW(feature_belows[1288])) ac1288(.scan_win(scan_win1288), .scan_win_std_dev(scan_win_std_dev[1288]), .feature_accum(feature_accums[1288]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1289]), .RECT1_Y(rectangle1_ys[1289]), .RECT1_WIDTH(rectangle1_widths[1289]), .RECT1_HEIGHT(rectangle1_heights[1289]), .RECT1_WEIGHT(rectangle1_weights[1289]), .RECT2_X(rectangle2_xs[1289]), .RECT2_Y(rectangle2_ys[1289]), .RECT2_WIDTH(rectangle2_widths[1289]), .RECT2_HEIGHT(rectangle2_heights[1289]), .RECT2_WEIGHT(rectangle2_weights[1289]), .RECT3_X(rectangle3_xs[1289]), .RECT3_Y(rectangle3_ys[1289]), .RECT3_WIDTH(rectangle3_widths[1289]), .RECT3_HEIGHT(rectangle3_heights[1289]), .RECT3_WEIGHT(rectangle3_weights[1289]), .FEAT_THRES(feature_thresholds[1289]), .FEAT_ABOVE(feature_aboves[1289]), .FEAT_BELOW(feature_belows[1289])) ac1289(.scan_win(scan_win1289), .scan_win_std_dev(scan_win_std_dev[1289]), .feature_accum(feature_accums[1289]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1290]), .RECT1_Y(rectangle1_ys[1290]), .RECT1_WIDTH(rectangle1_widths[1290]), .RECT1_HEIGHT(rectangle1_heights[1290]), .RECT1_WEIGHT(rectangle1_weights[1290]), .RECT2_X(rectangle2_xs[1290]), .RECT2_Y(rectangle2_ys[1290]), .RECT2_WIDTH(rectangle2_widths[1290]), .RECT2_HEIGHT(rectangle2_heights[1290]), .RECT2_WEIGHT(rectangle2_weights[1290]), .RECT3_X(rectangle3_xs[1290]), .RECT3_Y(rectangle3_ys[1290]), .RECT3_WIDTH(rectangle3_widths[1290]), .RECT3_HEIGHT(rectangle3_heights[1290]), .RECT3_WEIGHT(rectangle3_weights[1290]), .FEAT_THRES(feature_thresholds[1290]), .FEAT_ABOVE(feature_aboves[1290]), .FEAT_BELOW(feature_belows[1290])) ac1290(.scan_win(scan_win1290), .scan_win_std_dev(scan_win_std_dev[1290]), .feature_accum(feature_accums[1290]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1291]), .RECT1_Y(rectangle1_ys[1291]), .RECT1_WIDTH(rectangle1_widths[1291]), .RECT1_HEIGHT(rectangle1_heights[1291]), .RECT1_WEIGHT(rectangle1_weights[1291]), .RECT2_X(rectangle2_xs[1291]), .RECT2_Y(rectangle2_ys[1291]), .RECT2_WIDTH(rectangle2_widths[1291]), .RECT2_HEIGHT(rectangle2_heights[1291]), .RECT2_WEIGHT(rectangle2_weights[1291]), .RECT3_X(rectangle3_xs[1291]), .RECT3_Y(rectangle3_ys[1291]), .RECT3_WIDTH(rectangle3_widths[1291]), .RECT3_HEIGHT(rectangle3_heights[1291]), .RECT3_WEIGHT(rectangle3_weights[1291]), .FEAT_THRES(feature_thresholds[1291]), .FEAT_ABOVE(feature_aboves[1291]), .FEAT_BELOW(feature_belows[1291])) ac1291(.scan_win(scan_win1291), .scan_win_std_dev(scan_win_std_dev[1291]), .feature_accum(feature_accums[1291]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1292]), .RECT1_Y(rectangle1_ys[1292]), .RECT1_WIDTH(rectangle1_widths[1292]), .RECT1_HEIGHT(rectangle1_heights[1292]), .RECT1_WEIGHT(rectangle1_weights[1292]), .RECT2_X(rectangle2_xs[1292]), .RECT2_Y(rectangle2_ys[1292]), .RECT2_WIDTH(rectangle2_widths[1292]), .RECT2_HEIGHT(rectangle2_heights[1292]), .RECT2_WEIGHT(rectangle2_weights[1292]), .RECT3_X(rectangle3_xs[1292]), .RECT3_Y(rectangle3_ys[1292]), .RECT3_WIDTH(rectangle3_widths[1292]), .RECT3_HEIGHT(rectangle3_heights[1292]), .RECT3_WEIGHT(rectangle3_weights[1292]), .FEAT_THRES(feature_thresholds[1292]), .FEAT_ABOVE(feature_aboves[1292]), .FEAT_BELOW(feature_belows[1292])) ac1292(.scan_win(scan_win1292), .scan_win_std_dev(scan_win_std_dev[1292]), .feature_accum(feature_accums[1292]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1293]), .RECT1_Y(rectangle1_ys[1293]), .RECT1_WIDTH(rectangle1_widths[1293]), .RECT1_HEIGHT(rectangle1_heights[1293]), .RECT1_WEIGHT(rectangle1_weights[1293]), .RECT2_X(rectangle2_xs[1293]), .RECT2_Y(rectangle2_ys[1293]), .RECT2_WIDTH(rectangle2_widths[1293]), .RECT2_HEIGHT(rectangle2_heights[1293]), .RECT2_WEIGHT(rectangle2_weights[1293]), .RECT3_X(rectangle3_xs[1293]), .RECT3_Y(rectangle3_ys[1293]), .RECT3_WIDTH(rectangle3_widths[1293]), .RECT3_HEIGHT(rectangle3_heights[1293]), .RECT3_WEIGHT(rectangle3_weights[1293]), .FEAT_THRES(feature_thresholds[1293]), .FEAT_ABOVE(feature_aboves[1293]), .FEAT_BELOW(feature_belows[1293])) ac1293(.scan_win(scan_win1293), .scan_win_std_dev(scan_win_std_dev[1293]), .feature_accum(feature_accums[1293]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1294]), .RECT1_Y(rectangle1_ys[1294]), .RECT1_WIDTH(rectangle1_widths[1294]), .RECT1_HEIGHT(rectangle1_heights[1294]), .RECT1_WEIGHT(rectangle1_weights[1294]), .RECT2_X(rectangle2_xs[1294]), .RECT2_Y(rectangle2_ys[1294]), .RECT2_WIDTH(rectangle2_widths[1294]), .RECT2_HEIGHT(rectangle2_heights[1294]), .RECT2_WEIGHT(rectangle2_weights[1294]), .RECT3_X(rectangle3_xs[1294]), .RECT3_Y(rectangle3_ys[1294]), .RECT3_WIDTH(rectangle3_widths[1294]), .RECT3_HEIGHT(rectangle3_heights[1294]), .RECT3_WEIGHT(rectangle3_weights[1294]), .FEAT_THRES(feature_thresholds[1294]), .FEAT_ABOVE(feature_aboves[1294]), .FEAT_BELOW(feature_belows[1294])) ac1294(.scan_win(scan_win1294), .scan_win_std_dev(scan_win_std_dev[1294]), .feature_accum(feature_accums[1294]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1295]), .RECT1_Y(rectangle1_ys[1295]), .RECT1_WIDTH(rectangle1_widths[1295]), .RECT1_HEIGHT(rectangle1_heights[1295]), .RECT1_WEIGHT(rectangle1_weights[1295]), .RECT2_X(rectangle2_xs[1295]), .RECT2_Y(rectangle2_ys[1295]), .RECT2_WIDTH(rectangle2_widths[1295]), .RECT2_HEIGHT(rectangle2_heights[1295]), .RECT2_WEIGHT(rectangle2_weights[1295]), .RECT3_X(rectangle3_xs[1295]), .RECT3_Y(rectangle3_ys[1295]), .RECT3_WIDTH(rectangle3_widths[1295]), .RECT3_HEIGHT(rectangle3_heights[1295]), .RECT3_WEIGHT(rectangle3_weights[1295]), .FEAT_THRES(feature_thresholds[1295]), .FEAT_ABOVE(feature_aboves[1295]), .FEAT_BELOW(feature_belows[1295])) ac1295(.scan_win(scan_win1295), .scan_win_std_dev(scan_win_std_dev[1295]), .feature_accum(feature_accums[1295]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1296]), .RECT1_Y(rectangle1_ys[1296]), .RECT1_WIDTH(rectangle1_widths[1296]), .RECT1_HEIGHT(rectangle1_heights[1296]), .RECT1_WEIGHT(rectangle1_weights[1296]), .RECT2_X(rectangle2_xs[1296]), .RECT2_Y(rectangle2_ys[1296]), .RECT2_WIDTH(rectangle2_widths[1296]), .RECT2_HEIGHT(rectangle2_heights[1296]), .RECT2_WEIGHT(rectangle2_weights[1296]), .RECT3_X(rectangle3_xs[1296]), .RECT3_Y(rectangle3_ys[1296]), .RECT3_WIDTH(rectangle3_widths[1296]), .RECT3_HEIGHT(rectangle3_heights[1296]), .RECT3_WEIGHT(rectangle3_weights[1296]), .FEAT_THRES(feature_thresholds[1296]), .FEAT_ABOVE(feature_aboves[1296]), .FEAT_BELOW(feature_belows[1296])) ac1296(.scan_win(scan_win1296), .scan_win_std_dev(scan_win_std_dev[1296]), .feature_accum(feature_accums[1296]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1297]), .RECT1_Y(rectangle1_ys[1297]), .RECT1_WIDTH(rectangle1_widths[1297]), .RECT1_HEIGHT(rectangle1_heights[1297]), .RECT1_WEIGHT(rectangle1_weights[1297]), .RECT2_X(rectangle2_xs[1297]), .RECT2_Y(rectangle2_ys[1297]), .RECT2_WIDTH(rectangle2_widths[1297]), .RECT2_HEIGHT(rectangle2_heights[1297]), .RECT2_WEIGHT(rectangle2_weights[1297]), .RECT3_X(rectangle3_xs[1297]), .RECT3_Y(rectangle3_ys[1297]), .RECT3_WIDTH(rectangle3_widths[1297]), .RECT3_HEIGHT(rectangle3_heights[1297]), .RECT3_WEIGHT(rectangle3_weights[1297]), .FEAT_THRES(feature_thresholds[1297]), .FEAT_ABOVE(feature_aboves[1297]), .FEAT_BELOW(feature_belows[1297])) ac1297(.scan_win(scan_win1297), .scan_win_std_dev(scan_win_std_dev[1297]), .feature_accum(feature_accums[1297]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1298]), .RECT1_Y(rectangle1_ys[1298]), .RECT1_WIDTH(rectangle1_widths[1298]), .RECT1_HEIGHT(rectangle1_heights[1298]), .RECT1_WEIGHT(rectangle1_weights[1298]), .RECT2_X(rectangle2_xs[1298]), .RECT2_Y(rectangle2_ys[1298]), .RECT2_WIDTH(rectangle2_widths[1298]), .RECT2_HEIGHT(rectangle2_heights[1298]), .RECT2_WEIGHT(rectangle2_weights[1298]), .RECT3_X(rectangle3_xs[1298]), .RECT3_Y(rectangle3_ys[1298]), .RECT3_WIDTH(rectangle3_widths[1298]), .RECT3_HEIGHT(rectangle3_heights[1298]), .RECT3_WEIGHT(rectangle3_weights[1298]), .FEAT_THRES(feature_thresholds[1298]), .FEAT_ABOVE(feature_aboves[1298]), .FEAT_BELOW(feature_belows[1298])) ac1298(.scan_win(scan_win1298), .scan_win_std_dev(scan_win_std_dev[1298]), .feature_accum(feature_accums[1298]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1299]), .RECT1_Y(rectangle1_ys[1299]), .RECT1_WIDTH(rectangle1_widths[1299]), .RECT1_HEIGHT(rectangle1_heights[1299]), .RECT1_WEIGHT(rectangle1_weights[1299]), .RECT2_X(rectangle2_xs[1299]), .RECT2_Y(rectangle2_ys[1299]), .RECT2_WIDTH(rectangle2_widths[1299]), .RECT2_HEIGHT(rectangle2_heights[1299]), .RECT2_WEIGHT(rectangle2_weights[1299]), .RECT3_X(rectangle3_xs[1299]), .RECT3_Y(rectangle3_ys[1299]), .RECT3_WIDTH(rectangle3_widths[1299]), .RECT3_HEIGHT(rectangle3_heights[1299]), .RECT3_WEIGHT(rectangle3_weights[1299]), .FEAT_THRES(feature_thresholds[1299]), .FEAT_ABOVE(feature_aboves[1299]), .FEAT_BELOW(feature_belows[1299])) ac1299(.scan_win(scan_win1299), .scan_win_std_dev(scan_win_std_dev[1299]), .feature_accum(feature_accums[1299]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1300]), .RECT1_Y(rectangle1_ys[1300]), .RECT1_WIDTH(rectangle1_widths[1300]), .RECT1_HEIGHT(rectangle1_heights[1300]), .RECT1_WEIGHT(rectangle1_weights[1300]), .RECT2_X(rectangle2_xs[1300]), .RECT2_Y(rectangle2_ys[1300]), .RECT2_WIDTH(rectangle2_widths[1300]), .RECT2_HEIGHT(rectangle2_heights[1300]), .RECT2_WEIGHT(rectangle2_weights[1300]), .RECT3_X(rectangle3_xs[1300]), .RECT3_Y(rectangle3_ys[1300]), .RECT3_WIDTH(rectangle3_widths[1300]), .RECT3_HEIGHT(rectangle3_heights[1300]), .RECT3_WEIGHT(rectangle3_weights[1300]), .FEAT_THRES(feature_thresholds[1300]), .FEAT_ABOVE(feature_aboves[1300]), .FEAT_BELOW(feature_belows[1300])) ac1300(.scan_win(scan_win1300), .scan_win_std_dev(scan_win_std_dev[1300]), .feature_accum(feature_accums[1300]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1301]), .RECT1_Y(rectangle1_ys[1301]), .RECT1_WIDTH(rectangle1_widths[1301]), .RECT1_HEIGHT(rectangle1_heights[1301]), .RECT1_WEIGHT(rectangle1_weights[1301]), .RECT2_X(rectangle2_xs[1301]), .RECT2_Y(rectangle2_ys[1301]), .RECT2_WIDTH(rectangle2_widths[1301]), .RECT2_HEIGHT(rectangle2_heights[1301]), .RECT2_WEIGHT(rectangle2_weights[1301]), .RECT3_X(rectangle3_xs[1301]), .RECT3_Y(rectangle3_ys[1301]), .RECT3_WIDTH(rectangle3_widths[1301]), .RECT3_HEIGHT(rectangle3_heights[1301]), .RECT3_WEIGHT(rectangle3_weights[1301]), .FEAT_THRES(feature_thresholds[1301]), .FEAT_ABOVE(feature_aboves[1301]), .FEAT_BELOW(feature_belows[1301])) ac1301(.scan_win(scan_win1301), .scan_win_std_dev(scan_win_std_dev[1301]), .feature_accum(feature_accums[1301]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1302]), .RECT1_Y(rectangle1_ys[1302]), .RECT1_WIDTH(rectangle1_widths[1302]), .RECT1_HEIGHT(rectangle1_heights[1302]), .RECT1_WEIGHT(rectangle1_weights[1302]), .RECT2_X(rectangle2_xs[1302]), .RECT2_Y(rectangle2_ys[1302]), .RECT2_WIDTH(rectangle2_widths[1302]), .RECT2_HEIGHT(rectangle2_heights[1302]), .RECT2_WEIGHT(rectangle2_weights[1302]), .RECT3_X(rectangle3_xs[1302]), .RECT3_Y(rectangle3_ys[1302]), .RECT3_WIDTH(rectangle3_widths[1302]), .RECT3_HEIGHT(rectangle3_heights[1302]), .RECT3_WEIGHT(rectangle3_weights[1302]), .FEAT_THRES(feature_thresholds[1302]), .FEAT_ABOVE(feature_aboves[1302]), .FEAT_BELOW(feature_belows[1302])) ac1302(.scan_win(scan_win1302), .scan_win_std_dev(scan_win_std_dev[1302]), .feature_accum(feature_accums[1302]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1303]), .RECT1_Y(rectangle1_ys[1303]), .RECT1_WIDTH(rectangle1_widths[1303]), .RECT1_HEIGHT(rectangle1_heights[1303]), .RECT1_WEIGHT(rectangle1_weights[1303]), .RECT2_X(rectangle2_xs[1303]), .RECT2_Y(rectangle2_ys[1303]), .RECT2_WIDTH(rectangle2_widths[1303]), .RECT2_HEIGHT(rectangle2_heights[1303]), .RECT2_WEIGHT(rectangle2_weights[1303]), .RECT3_X(rectangle3_xs[1303]), .RECT3_Y(rectangle3_ys[1303]), .RECT3_WIDTH(rectangle3_widths[1303]), .RECT3_HEIGHT(rectangle3_heights[1303]), .RECT3_WEIGHT(rectangle3_weights[1303]), .FEAT_THRES(feature_thresholds[1303]), .FEAT_ABOVE(feature_aboves[1303]), .FEAT_BELOW(feature_belows[1303])) ac1303(.scan_win(scan_win1303), .scan_win_std_dev(scan_win_std_dev[1303]), .feature_accum(feature_accums[1303]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1304]), .RECT1_Y(rectangle1_ys[1304]), .RECT1_WIDTH(rectangle1_widths[1304]), .RECT1_HEIGHT(rectangle1_heights[1304]), .RECT1_WEIGHT(rectangle1_weights[1304]), .RECT2_X(rectangle2_xs[1304]), .RECT2_Y(rectangle2_ys[1304]), .RECT2_WIDTH(rectangle2_widths[1304]), .RECT2_HEIGHT(rectangle2_heights[1304]), .RECT2_WEIGHT(rectangle2_weights[1304]), .RECT3_X(rectangle3_xs[1304]), .RECT3_Y(rectangle3_ys[1304]), .RECT3_WIDTH(rectangle3_widths[1304]), .RECT3_HEIGHT(rectangle3_heights[1304]), .RECT3_WEIGHT(rectangle3_weights[1304]), .FEAT_THRES(feature_thresholds[1304]), .FEAT_ABOVE(feature_aboves[1304]), .FEAT_BELOW(feature_belows[1304])) ac1304(.scan_win(scan_win1304), .scan_win_std_dev(scan_win_std_dev[1304]), .feature_accum(feature_accums[1304]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1305]), .RECT1_Y(rectangle1_ys[1305]), .RECT1_WIDTH(rectangle1_widths[1305]), .RECT1_HEIGHT(rectangle1_heights[1305]), .RECT1_WEIGHT(rectangle1_weights[1305]), .RECT2_X(rectangle2_xs[1305]), .RECT2_Y(rectangle2_ys[1305]), .RECT2_WIDTH(rectangle2_widths[1305]), .RECT2_HEIGHT(rectangle2_heights[1305]), .RECT2_WEIGHT(rectangle2_weights[1305]), .RECT3_X(rectangle3_xs[1305]), .RECT3_Y(rectangle3_ys[1305]), .RECT3_WIDTH(rectangle3_widths[1305]), .RECT3_HEIGHT(rectangle3_heights[1305]), .RECT3_WEIGHT(rectangle3_weights[1305]), .FEAT_THRES(feature_thresholds[1305]), .FEAT_ABOVE(feature_aboves[1305]), .FEAT_BELOW(feature_belows[1305])) ac1305(.scan_win(scan_win1305), .scan_win_std_dev(scan_win_std_dev[1305]), .feature_accum(feature_accums[1305]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1306]), .RECT1_Y(rectangle1_ys[1306]), .RECT1_WIDTH(rectangle1_widths[1306]), .RECT1_HEIGHT(rectangle1_heights[1306]), .RECT1_WEIGHT(rectangle1_weights[1306]), .RECT2_X(rectangle2_xs[1306]), .RECT2_Y(rectangle2_ys[1306]), .RECT2_WIDTH(rectangle2_widths[1306]), .RECT2_HEIGHT(rectangle2_heights[1306]), .RECT2_WEIGHT(rectangle2_weights[1306]), .RECT3_X(rectangle3_xs[1306]), .RECT3_Y(rectangle3_ys[1306]), .RECT3_WIDTH(rectangle3_widths[1306]), .RECT3_HEIGHT(rectangle3_heights[1306]), .RECT3_WEIGHT(rectangle3_weights[1306]), .FEAT_THRES(feature_thresholds[1306]), .FEAT_ABOVE(feature_aboves[1306]), .FEAT_BELOW(feature_belows[1306])) ac1306(.scan_win(scan_win1306), .scan_win_std_dev(scan_win_std_dev[1306]), .feature_accum(feature_accums[1306]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1307]), .RECT1_Y(rectangle1_ys[1307]), .RECT1_WIDTH(rectangle1_widths[1307]), .RECT1_HEIGHT(rectangle1_heights[1307]), .RECT1_WEIGHT(rectangle1_weights[1307]), .RECT2_X(rectangle2_xs[1307]), .RECT2_Y(rectangle2_ys[1307]), .RECT2_WIDTH(rectangle2_widths[1307]), .RECT2_HEIGHT(rectangle2_heights[1307]), .RECT2_WEIGHT(rectangle2_weights[1307]), .RECT3_X(rectangle3_xs[1307]), .RECT3_Y(rectangle3_ys[1307]), .RECT3_WIDTH(rectangle3_widths[1307]), .RECT3_HEIGHT(rectangle3_heights[1307]), .RECT3_WEIGHT(rectangle3_weights[1307]), .FEAT_THRES(feature_thresholds[1307]), .FEAT_ABOVE(feature_aboves[1307]), .FEAT_BELOW(feature_belows[1307])) ac1307(.scan_win(scan_win1307), .scan_win_std_dev(scan_win_std_dev[1307]), .feature_accum(feature_accums[1307]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1308]), .RECT1_Y(rectangle1_ys[1308]), .RECT1_WIDTH(rectangle1_widths[1308]), .RECT1_HEIGHT(rectangle1_heights[1308]), .RECT1_WEIGHT(rectangle1_weights[1308]), .RECT2_X(rectangle2_xs[1308]), .RECT2_Y(rectangle2_ys[1308]), .RECT2_WIDTH(rectangle2_widths[1308]), .RECT2_HEIGHT(rectangle2_heights[1308]), .RECT2_WEIGHT(rectangle2_weights[1308]), .RECT3_X(rectangle3_xs[1308]), .RECT3_Y(rectangle3_ys[1308]), .RECT3_WIDTH(rectangle3_widths[1308]), .RECT3_HEIGHT(rectangle3_heights[1308]), .RECT3_WEIGHT(rectangle3_weights[1308]), .FEAT_THRES(feature_thresholds[1308]), .FEAT_ABOVE(feature_aboves[1308]), .FEAT_BELOW(feature_belows[1308])) ac1308(.scan_win(scan_win1308), .scan_win_std_dev(scan_win_std_dev[1308]), .feature_accum(feature_accums[1308]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1309]), .RECT1_Y(rectangle1_ys[1309]), .RECT1_WIDTH(rectangle1_widths[1309]), .RECT1_HEIGHT(rectangle1_heights[1309]), .RECT1_WEIGHT(rectangle1_weights[1309]), .RECT2_X(rectangle2_xs[1309]), .RECT2_Y(rectangle2_ys[1309]), .RECT2_WIDTH(rectangle2_widths[1309]), .RECT2_HEIGHT(rectangle2_heights[1309]), .RECT2_WEIGHT(rectangle2_weights[1309]), .RECT3_X(rectangle3_xs[1309]), .RECT3_Y(rectangle3_ys[1309]), .RECT3_WIDTH(rectangle3_widths[1309]), .RECT3_HEIGHT(rectangle3_heights[1309]), .RECT3_WEIGHT(rectangle3_weights[1309]), .FEAT_THRES(feature_thresholds[1309]), .FEAT_ABOVE(feature_aboves[1309]), .FEAT_BELOW(feature_belows[1309])) ac1309(.scan_win(scan_win1309), .scan_win_std_dev(scan_win_std_dev[1309]), .feature_accum(feature_accums[1309]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1310]), .RECT1_Y(rectangle1_ys[1310]), .RECT1_WIDTH(rectangle1_widths[1310]), .RECT1_HEIGHT(rectangle1_heights[1310]), .RECT1_WEIGHT(rectangle1_weights[1310]), .RECT2_X(rectangle2_xs[1310]), .RECT2_Y(rectangle2_ys[1310]), .RECT2_WIDTH(rectangle2_widths[1310]), .RECT2_HEIGHT(rectangle2_heights[1310]), .RECT2_WEIGHT(rectangle2_weights[1310]), .RECT3_X(rectangle3_xs[1310]), .RECT3_Y(rectangle3_ys[1310]), .RECT3_WIDTH(rectangle3_widths[1310]), .RECT3_HEIGHT(rectangle3_heights[1310]), .RECT3_WEIGHT(rectangle3_weights[1310]), .FEAT_THRES(feature_thresholds[1310]), .FEAT_ABOVE(feature_aboves[1310]), .FEAT_BELOW(feature_belows[1310])) ac1310(.scan_win(scan_win1310), .scan_win_std_dev(scan_win_std_dev[1310]), .feature_accum(feature_accums[1310]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1311]), .RECT1_Y(rectangle1_ys[1311]), .RECT1_WIDTH(rectangle1_widths[1311]), .RECT1_HEIGHT(rectangle1_heights[1311]), .RECT1_WEIGHT(rectangle1_weights[1311]), .RECT2_X(rectangle2_xs[1311]), .RECT2_Y(rectangle2_ys[1311]), .RECT2_WIDTH(rectangle2_widths[1311]), .RECT2_HEIGHT(rectangle2_heights[1311]), .RECT2_WEIGHT(rectangle2_weights[1311]), .RECT3_X(rectangle3_xs[1311]), .RECT3_Y(rectangle3_ys[1311]), .RECT3_WIDTH(rectangle3_widths[1311]), .RECT3_HEIGHT(rectangle3_heights[1311]), .RECT3_WEIGHT(rectangle3_weights[1311]), .FEAT_THRES(feature_thresholds[1311]), .FEAT_ABOVE(feature_aboves[1311]), .FEAT_BELOW(feature_belows[1311])) ac1311(.scan_win(scan_win1311), .scan_win_std_dev(scan_win_std_dev[1311]), .feature_accum(feature_accums[1311]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1312]), .RECT1_Y(rectangle1_ys[1312]), .RECT1_WIDTH(rectangle1_widths[1312]), .RECT1_HEIGHT(rectangle1_heights[1312]), .RECT1_WEIGHT(rectangle1_weights[1312]), .RECT2_X(rectangle2_xs[1312]), .RECT2_Y(rectangle2_ys[1312]), .RECT2_WIDTH(rectangle2_widths[1312]), .RECT2_HEIGHT(rectangle2_heights[1312]), .RECT2_WEIGHT(rectangle2_weights[1312]), .RECT3_X(rectangle3_xs[1312]), .RECT3_Y(rectangle3_ys[1312]), .RECT3_WIDTH(rectangle3_widths[1312]), .RECT3_HEIGHT(rectangle3_heights[1312]), .RECT3_WEIGHT(rectangle3_weights[1312]), .FEAT_THRES(feature_thresholds[1312]), .FEAT_ABOVE(feature_aboves[1312]), .FEAT_BELOW(feature_belows[1312])) ac1312(.scan_win(scan_win1312), .scan_win_std_dev(scan_win_std_dev[1312]), .feature_accum(feature_accums[1312]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1313]), .RECT1_Y(rectangle1_ys[1313]), .RECT1_WIDTH(rectangle1_widths[1313]), .RECT1_HEIGHT(rectangle1_heights[1313]), .RECT1_WEIGHT(rectangle1_weights[1313]), .RECT2_X(rectangle2_xs[1313]), .RECT2_Y(rectangle2_ys[1313]), .RECT2_WIDTH(rectangle2_widths[1313]), .RECT2_HEIGHT(rectangle2_heights[1313]), .RECT2_WEIGHT(rectangle2_weights[1313]), .RECT3_X(rectangle3_xs[1313]), .RECT3_Y(rectangle3_ys[1313]), .RECT3_WIDTH(rectangle3_widths[1313]), .RECT3_HEIGHT(rectangle3_heights[1313]), .RECT3_WEIGHT(rectangle3_weights[1313]), .FEAT_THRES(feature_thresholds[1313]), .FEAT_ABOVE(feature_aboves[1313]), .FEAT_BELOW(feature_belows[1313])) ac1313(.scan_win(scan_win1313), .scan_win_std_dev(scan_win_std_dev[1313]), .feature_accum(feature_accums[1313]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1314]), .RECT1_Y(rectangle1_ys[1314]), .RECT1_WIDTH(rectangle1_widths[1314]), .RECT1_HEIGHT(rectangle1_heights[1314]), .RECT1_WEIGHT(rectangle1_weights[1314]), .RECT2_X(rectangle2_xs[1314]), .RECT2_Y(rectangle2_ys[1314]), .RECT2_WIDTH(rectangle2_widths[1314]), .RECT2_HEIGHT(rectangle2_heights[1314]), .RECT2_WEIGHT(rectangle2_weights[1314]), .RECT3_X(rectangle3_xs[1314]), .RECT3_Y(rectangle3_ys[1314]), .RECT3_WIDTH(rectangle3_widths[1314]), .RECT3_HEIGHT(rectangle3_heights[1314]), .RECT3_WEIGHT(rectangle3_weights[1314]), .FEAT_THRES(feature_thresholds[1314]), .FEAT_ABOVE(feature_aboves[1314]), .FEAT_BELOW(feature_belows[1314])) ac1314(.scan_win(scan_win1314), .scan_win_std_dev(scan_win_std_dev[1314]), .feature_accum(feature_accums[1314]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1315]), .RECT1_Y(rectangle1_ys[1315]), .RECT1_WIDTH(rectangle1_widths[1315]), .RECT1_HEIGHT(rectangle1_heights[1315]), .RECT1_WEIGHT(rectangle1_weights[1315]), .RECT2_X(rectangle2_xs[1315]), .RECT2_Y(rectangle2_ys[1315]), .RECT2_WIDTH(rectangle2_widths[1315]), .RECT2_HEIGHT(rectangle2_heights[1315]), .RECT2_WEIGHT(rectangle2_weights[1315]), .RECT3_X(rectangle3_xs[1315]), .RECT3_Y(rectangle3_ys[1315]), .RECT3_WIDTH(rectangle3_widths[1315]), .RECT3_HEIGHT(rectangle3_heights[1315]), .RECT3_WEIGHT(rectangle3_weights[1315]), .FEAT_THRES(feature_thresholds[1315]), .FEAT_ABOVE(feature_aboves[1315]), .FEAT_BELOW(feature_belows[1315])) ac1315(.scan_win(scan_win1315), .scan_win_std_dev(scan_win_std_dev[1315]), .feature_accum(feature_accums[1315]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1316]), .RECT1_Y(rectangle1_ys[1316]), .RECT1_WIDTH(rectangle1_widths[1316]), .RECT1_HEIGHT(rectangle1_heights[1316]), .RECT1_WEIGHT(rectangle1_weights[1316]), .RECT2_X(rectangle2_xs[1316]), .RECT2_Y(rectangle2_ys[1316]), .RECT2_WIDTH(rectangle2_widths[1316]), .RECT2_HEIGHT(rectangle2_heights[1316]), .RECT2_WEIGHT(rectangle2_weights[1316]), .RECT3_X(rectangle3_xs[1316]), .RECT3_Y(rectangle3_ys[1316]), .RECT3_WIDTH(rectangle3_widths[1316]), .RECT3_HEIGHT(rectangle3_heights[1316]), .RECT3_WEIGHT(rectangle3_weights[1316]), .FEAT_THRES(feature_thresholds[1316]), .FEAT_ABOVE(feature_aboves[1316]), .FEAT_BELOW(feature_belows[1316])) ac1316(.scan_win(scan_win1316), .scan_win_std_dev(scan_win_std_dev[1316]), .feature_accum(feature_accums[1316]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1317]), .RECT1_Y(rectangle1_ys[1317]), .RECT1_WIDTH(rectangle1_widths[1317]), .RECT1_HEIGHT(rectangle1_heights[1317]), .RECT1_WEIGHT(rectangle1_weights[1317]), .RECT2_X(rectangle2_xs[1317]), .RECT2_Y(rectangle2_ys[1317]), .RECT2_WIDTH(rectangle2_widths[1317]), .RECT2_HEIGHT(rectangle2_heights[1317]), .RECT2_WEIGHT(rectangle2_weights[1317]), .RECT3_X(rectangle3_xs[1317]), .RECT3_Y(rectangle3_ys[1317]), .RECT3_WIDTH(rectangle3_widths[1317]), .RECT3_HEIGHT(rectangle3_heights[1317]), .RECT3_WEIGHT(rectangle3_weights[1317]), .FEAT_THRES(feature_thresholds[1317]), .FEAT_ABOVE(feature_aboves[1317]), .FEAT_BELOW(feature_belows[1317])) ac1317(.scan_win(scan_win1317), .scan_win_std_dev(scan_win_std_dev[1317]), .feature_accum(feature_accums[1317]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1318]), .RECT1_Y(rectangle1_ys[1318]), .RECT1_WIDTH(rectangle1_widths[1318]), .RECT1_HEIGHT(rectangle1_heights[1318]), .RECT1_WEIGHT(rectangle1_weights[1318]), .RECT2_X(rectangle2_xs[1318]), .RECT2_Y(rectangle2_ys[1318]), .RECT2_WIDTH(rectangle2_widths[1318]), .RECT2_HEIGHT(rectangle2_heights[1318]), .RECT2_WEIGHT(rectangle2_weights[1318]), .RECT3_X(rectangle3_xs[1318]), .RECT3_Y(rectangle3_ys[1318]), .RECT3_WIDTH(rectangle3_widths[1318]), .RECT3_HEIGHT(rectangle3_heights[1318]), .RECT3_WEIGHT(rectangle3_weights[1318]), .FEAT_THRES(feature_thresholds[1318]), .FEAT_ABOVE(feature_aboves[1318]), .FEAT_BELOW(feature_belows[1318])) ac1318(.scan_win(scan_win1318), .scan_win_std_dev(scan_win_std_dev[1318]), .feature_accum(feature_accums[1318]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1319]), .RECT1_Y(rectangle1_ys[1319]), .RECT1_WIDTH(rectangle1_widths[1319]), .RECT1_HEIGHT(rectangle1_heights[1319]), .RECT1_WEIGHT(rectangle1_weights[1319]), .RECT2_X(rectangle2_xs[1319]), .RECT2_Y(rectangle2_ys[1319]), .RECT2_WIDTH(rectangle2_widths[1319]), .RECT2_HEIGHT(rectangle2_heights[1319]), .RECT2_WEIGHT(rectangle2_weights[1319]), .RECT3_X(rectangle3_xs[1319]), .RECT3_Y(rectangle3_ys[1319]), .RECT3_WIDTH(rectangle3_widths[1319]), .RECT3_HEIGHT(rectangle3_heights[1319]), .RECT3_WEIGHT(rectangle3_weights[1319]), .FEAT_THRES(feature_thresholds[1319]), .FEAT_ABOVE(feature_aboves[1319]), .FEAT_BELOW(feature_belows[1319])) ac1319(.scan_win(scan_win1319), .scan_win_std_dev(scan_win_std_dev[1319]), .feature_accum(feature_accums[1319]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1320]), .RECT1_Y(rectangle1_ys[1320]), .RECT1_WIDTH(rectangle1_widths[1320]), .RECT1_HEIGHT(rectangle1_heights[1320]), .RECT1_WEIGHT(rectangle1_weights[1320]), .RECT2_X(rectangle2_xs[1320]), .RECT2_Y(rectangle2_ys[1320]), .RECT2_WIDTH(rectangle2_widths[1320]), .RECT2_HEIGHT(rectangle2_heights[1320]), .RECT2_WEIGHT(rectangle2_weights[1320]), .RECT3_X(rectangle3_xs[1320]), .RECT3_Y(rectangle3_ys[1320]), .RECT3_WIDTH(rectangle3_widths[1320]), .RECT3_HEIGHT(rectangle3_heights[1320]), .RECT3_WEIGHT(rectangle3_weights[1320]), .FEAT_THRES(feature_thresholds[1320]), .FEAT_ABOVE(feature_aboves[1320]), .FEAT_BELOW(feature_belows[1320])) ac1320(.scan_win(scan_win1320), .scan_win_std_dev(scan_win_std_dev[1320]), .feature_accum(feature_accums[1320]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1321]), .RECT1_Y(rectangle1_ys[1321]), .RECT1_WIDTH(rectangle1_widths[1321]), .RECT1_HEIGHT(rectangle1_heights[1321]), .RECT1_WEIGHT(rectangle1_weights[1321]), .RECT2_X(rectangle2_xs[1321]), .RECT2_Y(rectangle2_ys[1321]), .RECT2_WIDTH(rectangle2_widths[1321]), .RECT2_HEIGHT(rectangle2_heights[1321]), .RECT2_WEIGHT(rectangle2_weights[1321]), .RECT3_X(rectangle3_xs[1321]), .RECT3_Y(rectangle3_ys[1321]), .RECT3_WIDTH(rectangle3_widths[1321]), .RECT3_HEIGHT(rectangle3_heights[1321]), .RECT3_WEIGHT(rectangle3_weights[1321]), .FEAT_THRES(feature_thresholds[1321]), .FEAT_ABOVE(feature_aboves[1321]), .FEAT_BELOW(feature_belows[1321])) ac1321(.scan_win(scan_win1321), .scan_win_std_dev(scan_win_std_dev[1321]), .feature_accum(feature_accums[1321]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1322]), .RECT1_Y(rectangle1_ys[1322]), .RECT1_WIDTH(rectangle1_widths[1322]), .RECT1_HEIGHT(rectangle1_heights[1322]), .RECT1_WEIGHT(rectangle1_weights[1322]), .RECT2_X(rectangle2_xs[1322]), .RECT2_Y(rectangle2_ys[1322]), .RECT2_WIDTH(rectangle2_widths[1322]), .RECT2_HEIGHT(rectangle2_heights[1322]), .RECT2_WEIGHT(rectangle2_weights[1322]), .RECT3_X(rectangle3_xs[1322]), .RECT3_Y(rectangle3_ys[1322]), .RECT3_WIDTH(rectangle3_widths[1322]), .RECT3_HEIGHT(rectangle3_heights[1322]), .RECT3_WEIGHT(rectangle3_weights[1322]), .FEAT_THRES(feature_thresholds[1322]), .FEAT_ABOVE(feature_aboves[1322]), .FEAT_BELOW(feature_belows[1322])) ac1322(.scan_win(scan_win1322), .scan_win_std_dev(scan_win_std_dev[1322]), .feature_accum(feature_accums[1322]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1323]), .RECT1_Y(rectangle1_ys[1323]), .RECT1_WIDTH(rectangle1_widths[1323]), .RECT1_HEIGHT(rectangle1_heights[1323]), .RECT1_WEIGHT(rectangle1_weights[1323]), .RECT2_X(rectangle2_xs[1323]), .RECT2_Y(rectangle2_ys[1323]), .RECT2_WIDTH(rectangle2_widths[1323]), .RECT2_HEIGHT(rectangle2_heights[1323]), .RECT2_WEIGHT(rectangle2_weights[1323]), .RECT3_X(rectangle3_xs[1323]), .RECT3_Y(rectangle3_ys[1323]), .RECT3_WIDTH(rectangle3_widths[1323]), .RECT3_HEIGHT(rectangle3_heights[1323]), .RECT3_WEIGHT(rectangle3_weights[1323]), .FEAT_THRES(feature_thresholds[1323]), .FEAT_ABOVE(feature_aboves[1323]), .FEAT_BELOW(feature_belows[1323])) ac1323(.scan_win(scan_win1323), .scan_win_std_dev(scan_win_std_dev[1323]), .feature_accum(feature_accums[1323]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1324]), .RECT1_Y(rectangle1_ys[1324]), .RECT1_WIDTH(rectangle1_widths[1324]), .RECT1_HEIGHT(rectangle1_heights[1324]), .RECT1_WEIGHT(rectangle1_weights[1324]), .RECT2_X(rectangle2_xs[1324]), .RECT2_Y(rectangle2_ys[1324]), .RECT2_WIDTH(rectangle2_widths[1324]), .RECT2_HEIGHT(rectangle2_heights[1324]), .RECT2_WEIGHT(rectangle2_weights[1324]), .RECT3_X(rectangle3_xs[1324]), .RECT3_Y(rectangle3_ys[1324]), .RECT3_WIDTH(rectangle3_widths[1324]), .RECT3_HEIGHT(rectangle3_heights[1324]), .RECT3_WEIGHT(rectangle3_weights[1324]), .FEAT_THRES(feature_thresholds[1324]), .FEAT_ABOVE(feature_aboves[1324]), .FEAT_BELOW(feature_belows[1324])) ac1324(.scan_win(scan_win1324), .scan_win_std_dev(scan_win_std_dev[1324]), .feature_accum(feature_accums[1324]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1325]), .RECT1_Y(rectangle1_ys[1325]), .RECT1_WIDTH(rectangle1_widths[1325]), .RECT1_HEIGHT(rectangle1_heights[1325]), .RECT1_WEIGHT(rectangle1_weights[1325]), .RECT2_X(rectangle2_xs[1325]), .RECT2_Y(rectangle2_ys[1325]), .RECT2_WIDTH(rectangle2_widths[1325]), .RECT2_HEIGHT(rectangle2_heights[1325]), .RECT2_WEIGHT(rectangle2_weights[1325]), .RECT3_X(rectangle3_xs[1325]), .RECT3_Y(rectangle3_ys[1325]), .RECT3_WIDTH(rectangle3_widths[1325]), .RECT3_HEIGHT(rectangle3_heights[1325]), .RECT3_WEIGHT(rectangle3_weights[1325]), .FEAT_THRES(feature_thresholds[1325]), .FEAT_ABOVE(feature_aboves[1325]), .FEAT_BELOW(feature_belows[1325])) ac1325(.scan_win(scan_win1325), .scan_win_std_dev(scan_win_std_dev[1325]), .feature_accum(feature_accums[1325]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1326]), .RECT1_Y(rectangle1_ys[1326]), .RECT1_WIDTH(rectangle1_widths[1326]), .RECT1_HEIGHT(rectangle1_heights[1326]), .RECT1_WEIGHT(rectangle1_weights[1326]), .RECT2_X(rectangle2_xs[1326]), .RECT2_Y(rectangle2_ys[1326]), .RECT2_WIDTH(rectangle2_widths[1326]), .RECT2_HEIGHT(rectangle2_heights[1326]), .RECT2_WEIGHT(rectangle2_weights[1326]), .RECT3_X(rectangle3_xs[1326]), .RECT3_Y(rectangle3_ys[1326]), .RECT3_WIDTH(rectangle3_widths[1326]), .RECT3_HEIGHT(rectangle3_heights[1326]), .RECT3_WEIGHT(rectangle3_weights[1326]), .FEAT_THRES(feature_thresholds[1326]), .FEAT_ABOVE(feature_aboves[1326]), .FEAT_BELOW(feature_belows[1326])) ac1326(.scan_win(scan_win1326), .scan_win_std_dev(scan_win_std_dev[1326]), .feature_accum(feature_accums[1326]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1327]), .RECT1_Y(rectangle1_ys[1327]), .RECT1_WIDTH(rectangle1_widths[1327]), .RECT1_HEIGHT(rectangle1_heights[1327]), .RECT1_WEIGHT(rectangle1_weights[1327]), .RECT2_X(rectangle2_xs[1327]), .RECT2_Y(rectangle2_ys[1327]), .RECT2_WIDTH(rectangle2_widths[1327]), .RECT2_HEIGHT(rectangle2_heights[1327]), .RECT2_WEIGHT(rectangle2_weights[1327]), .RECT3_X(rectangle3_xs[1327]), .RECT3_Y(rectangle3_ys[1327]), .RECT3_WIDTH(rectangle3_widths[1327]), .RECT3_HEIGHT(rectangle3_heights[1327]), .RECT3_WEIGHT(rectangle3_weights[1327]), .FEAT_THRES(feature_thresholds[1327]), .FEAT_ABOVE(feature_aboves[1327]), .FEAT_BELOW(feature_belows[1327])) ac1327(.scan_win(scan_win1327), .scan_win_std_dev(scan_win_std_dev[1327]), .feature_accum(feature_accums[1327]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1328]), .RECT1_Y(rectangle1_ys[1328]), .RECT1_WIDTH(rectangle1_widths[1328]), .RECT1_HEIGHT(rectangle1_heights[1328]), .RECT1_WEIGHT(rectangle1_weights[1328]), .RECT2_X(rectangle2_xs[1328]), .RECT2_Y(rectangle2_ys[1328]), .RECT2_WIDTH(rectangle2_widths[1328]), .RECT2_HEIGHT(rectangle2_heights[1328]), .RECT2_WEIGHT(rectangle2_weights[1328]), .RECT3_X(rectangle3_xs[1328]), .RECT3_Y(rectangle3_ys[1328]), .RECT3_WIDTH(rectangle3_widths[1328]), .RECT3_HEIGHT(rectangle3_heights[1328]), .RECT3_WEIGHT(rectangle3_weights[1328]), .FEAT_THRES(feature_thresholds[1328]), .FEAT_ABOVE(feature_aboves[1328]), .FEAT_BELOW(feature_belows[1328])) ac1328(.scan_win(scan_win1328), .scan_win_std_dev(scan_win_std_dev[1328]), .feature_accum(feature_accums[1328]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1329]), .RECT1_Y(rectangle1_ys[1329]), .RECT1_WIDTH(rectangle1_widths[1329]), .RECT1_HEIGHT(rectangle1_heights[1329]), .RECT1_WEIGHT(rectangle1_weights[1329]), .RECT2_X(rectangle2_xs[1329]), .RECT2_Y(rectangle2_ys[1329]), .RECT2_WIDTH(rectangle2_widths[1329]), .RECT2_HEIGHT(rectangle2_heights[1329]), .RECT2_WEIGHT(rectangle2_weights[1329]), .RECT3_X(rectangle3_xs[1329]), .RECT3_Y(rectangle3_ys[1329]), .RECT3_WIDTH(rectangle3_widths[1329]), .RECT3_HEIGHT(rectangle3_heights[1329]), .RECT3_WEIGHT(rectangle3_weights[1329]), .FEAT_THRES(feature_thresholds[1329]), .FEAT_ABOVE(feature_aboves[1329]), .FEAT_BELOW(feature_belows[1329])) ac1329(.scan_win(scan_win1329), .scan_win_std_dev(scan_win_std_dev[1329]), .feature_accum(feature_accums[1329]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1330]), .RECT1_Y(rectangle1_ys[1330]), .RECT1_WIDTH(rectangle1_widths[1330]), .RECT1_HEIGHT(rectangle1_heights[1330]), .RECT1_WEIGHT(rectangle1_weights[1330]), .RECT2_X(rectangle2_xs[1330]), .RECT2_Y(rectangle2_ys[1330]), .RECT2_WIDTH(rectangle2_widths[1330]), .RECT2_HEIGHT(rectangle2_heights[1330]), .RECT2_WEIGHT(rectangle2_weights[1330]), .RECT3_X(rectangle3_xs[1330]), .RECT3_Y(rectangle3_ys[1330]), .RECT3_WIDTH(rectangle3_widths[1330]), .RECT3_HEIGHT(rectangle3_heights[1330]), .RECT3_WEIGHT(rectangle3_weights[1330]), .FEAT_THRES(feature_thresholds[1330]), .FEAT_ABOVE(feature_aboves[1330]), .FEAT_BELOW(feature_belows[1330])) ac1330(.scan_win(scan_win1330), .scan_win_std_dev(scan_win_std_dev[1330]), .feature_accum(feature_accums[1330]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1331]), .RECT1_Y(rectangle1_ys[1331]), .RECT1_WIDTH(rectangle1_widths[1331]), .RECT1_HEIGHT(rectangle1_heights[1331]), .RECT1_WEIGHT(rectangle1_weights[1331]), .RECT2_X(rectangle2_xs[1331]), .RECT2_Y(rectangle2_ys[1331]), .RECT2_WIDTH(rectangle2_widths[1331]), .RECT2_HEIGHT(rectangle2_heights[1331]), .RECT2_WEIGHT(rectangle2_weights[1331]), .RECT3_X(rectangle3_xs[1331]), .RECT3_Y(rectangle3_ys[1331]), .RECT3_WIDTH(rectangle3_widths[1331]), .RECT3_HEIGHT(rectangle3_heights[1331]), .RECT3_WEIGHT(rectangle3_weights[1331]), .FEAT_THRES(feature_thresholds[1331]), .FEAT_ABOVE(feature_aboves[1331]), .FEAT_BELOW(feature_belows[1331])) ac1331(.scan_win(scan_win1331), .scan_win_std_dev(scan_win_std_dev[1331]), .feature_accum(feature_accums[1331]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1332]), .RECT1_Y(rectangle1_ys[1332]), .RECT1_WIDTH(rectangle1_widths[1332]), .RECT1_HEIGHT(rectangle1_heights[1332]), .RECT1_WEIGHT(rectangle1_weights[1332]), .RECT2_X(rectangle2_xs[1332]), .RECT2_Y(rectangle2_ys[1332]), .RECT2_WIDTH(rectangle2_widths[1332]), .RECT2_HEIGHT(rectangle2_heights[1332]), .RECT2_WEIGHT(rectangle2_weights[1332]), .RECT3_X(rectangle3_xs[1332]), .RECT3_Y(rectangle3_ys[1332]), .RECT3_WIDTH(rectangle3_widths[1332]), .RECT3_HEIGHT(rectangle3_heights[1332]), .RECT3_WEIGHT(rectangle3_weights[1332]), .FEAT_THRES(feature_thresholds[1332]), .FEAT_ABOVE(feature_aboves[1332]), .FEAT_BELOW(feature_belows[1332])) ac1332(.scan_win(scan_win1332), .scan_win_std_dev(scan_win_std_dev[1332]), .feature_accum(feature_accums[1332]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1333]), .RECT1_Y(rectangle1_ys[1333]), .RECT1_WIDTH(rectangle1_widths[1333]), .RECT1_HEIGHT(rectangle1_heights[1333]), .RECT1_WEIGHT(rectangle1_weights[1333]), .RECT2_X(rectangle2_xs[1333]), .RECT2_Y(rectangle2_ys[1333]), .RECT2_WIDTH(rectangle2_widths[1333]), .RECT2_HEIGHT(rectangle2_heights[1333]), .RECT2_WEIGHT(rectangle2_weights[1333]), .RECT3_X(rectangle3_xs[1333]), .RECT3_Y(rectangle3_ys[1333]), .RECT3_WIDTH(rectangle3_widths[1333]), .RECT3_HEIGHT(rectangle3_heights[1333]), .RECT3_WEIGHT(rectangle3_weights[1333]), .FEAT_THRES(feature_thresholds[1333]), .FEAT_ABOVE(feature_aboves[1333]), .FEAT_BELOW(feature_belows[1333])) ac1333(.scan_win(scan_win1333), .scan_win_std_dev(scan_win_std_dev[1333]), .feature_accum(feature_accums[1333]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1334]), .RECT1_Y(rectangle1_ys[1334]), .RECT1_WIDTH(rectangle1_widths[1334]), .RECT1_HEIGHT(rectangle1_heights[1334]), .RECT1_WEIGHT(rectangle1_weights[1334]), .RECT2_X(rectangle2_xs[1334]), .RECT2_Y(rectangle2_ys[1334]), .RECT2_WIDTH(rectangle2_widths[1334]), .RECT2_HEIGHT(rectangle2_heights[1334]), .RECT2_WEIGHT(rectangle2_weights[1334]), .RECT3_X(rectangle3_xs[1334]), .RECT3_Y(rectangle3_ys[1334]), .RECT3_WIDTH(rectangle3_widths[1334]), .RECT3_HEIGHT(rectangle3_heights[1334]), .RECT3_WEIGHT(rectangle3_weights[1334]), .FEAT_THRES(feature_thresholds[1334]), .FEAT_ABOVE(feature_aboves[1334]), .FEAT_BELOW(feature_belows[1334])) ac1334(.scan_win(scan_win1334), .scan_win_std_dev(scan_win_std_dev[1334]), .feature_accum(feature_accums[1334]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1335]), .RECT1_Y(rectangle1_ys[1335]), .RECT1_WIDTH(rectangle1_widths[1335]), .RECT1_HEIGHT(rectangle1_heights[1335]), .RECT1_WEIGHT(rectangle1_weights[1335]), .RECT2_X(rectangle2_xs[1335]), .RECT2_Y(rectangle2_ys[1335]), .RECT2_WIDTH(rectangle2_widths[1335]), .RECT2_HEIGHT(rectangle2_heights[1335]), .RECT2_WEIGHT(rectangle2_weights[1335]), .RECT3_X(rectangle3_xs[1335]), .RECT3_Y(rectangle3_ys[1335]), .RECT3_WIDTH(rectangle3_widths[1335]), .RECT3_HEIGHT(rectangle3_heights[1335]), .RECT3_WEIGHT(rectangle3_weights[1335]), .FEAT_THRES(feature_thresholds[1335]), .FEAT_ABOVE(feature_aboves[1335]), .FEAT_BELOW(feature_belows[1335])) ac1335(.scan_win(scan_win1335), .scan_win_std_dev(scan_win_std_dev[1335]), .feature_accum(feature_accums[1335]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1336]), .RECT1_Y(rectangle1_ys[1336]), .RECT1_WIDTH(rectangle1_widths[1336]), .RECT1_HEIGHT(rectangle1_heights[1336]), .RECT1_WEIGHT(rectangle1_weights[1336]), .RECT2_X(rectangle2_xs[1336]), .RECT2_Y(rectangle2_ys[1336]), .RECT2_WIDTH(rectangle2_widths[1336]), .RECT2_HEIGHT(rectangle2_heights[1336]), .RECT2_WEIGHT(rectangle2_weights[1336]), .RECT3_X(rectangle3_xs[1336]), .RECT3_Y(rectangle3_ys[1336]), .RECT3_WIDTH(rectangle3_widths[1336]), .RECT3_HEIGHT(rectangle3_heights[1336]), .RECT3_WEIGHT(rectangle3_weights[1336]), .FEAT_THRES(feature_thresholds[1336]), .FEAT_ABOVE(feature_aboves[1336]), .FEAT_BELOW(feature_belows[1336])) ac1336(.scan_win(scan_win1336), .scan_win_std_dev(scan_win_std_dev[1336]), .feature_accum(feature_accums[1336]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1337]), .RECT1_Y(rectangle1_ys[1337]), .RECT1_WIDTH(rectangle1_widths[1337]), .RECT1_HEIGHT(rectangle1_heights[1337]), .RECT1_WEIGHT(rectangle1_weights[1337]), .RECT2_X(rectangle2_xs[1337]), .RECT2_Y(rectangle2_ys[1337]), .RECT2_WIDTH(rectangle2_widths[1337]), .RECT2_HEIGHT(rectangle2_heights[1337]), .RECT2_WEIGHT(rectangle2_weights[1337]), .RECT3_X(rectangle3_xs[1337]), .RECT3_Y(rectangle3_ys[1337]), .RECT3_WIDTH(rectangle3_widths[1337]), .RECT3_HEIGHT(rectangle3_heights[1337]), .RECT3_WEIGHT(rectangle3_weights[1337]), .FEAT_THRES(feature_thresholds[1337]), .FEAT_ABOVE(feature_aboves[1337]), .FEAT_BELOW(feature_belows[1337])) ac1337(.scan_win(scan_win1337), .scan_win_std_dev(scan_win_std_dev[1337]), .feature_accum(feature_accums[1337]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1338]), .RECT1_Y(rectangle1_ys[1338]), .RECT1_WIDTH(rectangle1_widths[1338]), .RECT1_HEIGHT(rectangle1_heights[1338]), .RECT1_WEIGHT(rectangle1_weights[1338]), .RECT2_X(rectangle2_xs[1338]), .RECT2_Y(rectangle2_ys[1338]), .RECT2_WIDTH(rectangle2_widths[1338]), .RECT2_HEIGHT(rectangle2_heights[1338]), .RECT2_WEIGHT(rectangle2_weights[1338]), .RECT3_X(rectangle3_xs[1338]), .RECT3_Y(rectangle3_ys[1338]), .RECT3_WIDTH(rectangle3_widths[1338]), .RECT3_HEIGHT(rectangle3_heights[1338]), .RECT3_WEIGHT(rectangle3_weights[1338]), .FEAT_THRES(feature_thresholds[1338]), .FEAT_ABOVE(feature_aboves[1338]), .FEAT_BELOW(feature_belows[1338])) ac1338(.scan_win(scan_win1338), .scan_win_std_dev(scan_win_std_dev[1338]), .feature_accum(feature_accums[1338]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1339]), .RECT1_Y(rectangle1_ys[1339]), .RECT1_WIDTH(rectangle1_widths[1339]), .RECT1_HEIGHT(rectangle1_heights[1339]), .RECT1_WEIGHT(rectangle1_weights[1339]), .RECT2_X(rectangle2_xs[1339]), .RECT2_Y(rectangle2_ys[1339]), .RECT2_WIDTH(rectangle2_widths[1339]), .RECT2_HEIGHT(rectangle2_heights[1339]), .RECT2_WEIGHT(rectangle2_weights[1339]), .RECT3_X(rectangle3_xs[1339]), .RECT3_Y(rectangle3_ys[1339]), .RECT3_WIDTH(rectangle3_widths[1339]), .RECT3_HEIGHT(rectangle3_heights[1339]), .RECT3_WEIGHT(rectangle3_weights[1339]), .FEAT_THRES(feature_thresholds[1339]), .FEAT_ABOVE(feature_aboves[1339]), .FEAT_BELOW(feature_belows[1339])) ac1339(.scan_win(scan_win1339), .scan_win_std_dev(scan_win_std_dev[1339]), .feature_accum(feature_accums[1339]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1340]), .RECT1_Y(rectangle1_ys[1340]), .RECT1_WIDTH(rectangle1_widths[1340]), .RECT1_HEIGHT(rectangle1_heights[1340]), .RECT1_WEIGHT(rectangle1_weights[1340]), .RECT2_X(rectangle2_xs[1340]), .RECT2_Y(rectangle2_ys[1340]), .RECT2_WIDTH(rectangle2_widths[1340]), .RECT2_HEIGHT(rectangle2_heights[1340]), .RECT2_WEIGHT(rectangle2_weights[1340]), .RECT3_X(rectangle3_xs[1340]), .RECT3_Y(rectangle3_ys[1340]), .RECT3_WIDTH(rectangle3_widths[1340]), .RECT3_HEIGHT(rectangle3_heights[1340]), .RECT3_WEIGHT(rectangle3_weights[1340]), .FEAT_THRES(feature_thresholds[1340]), .FEAT_ABOVE(feature_aboves[1340]), .FEAT_BELOW(feature_belows[1340])) ac1340(.scan_win(scan_win1340), .scan_win_std_dev(scan_win_std_dev[1340]), .feature_accum(feature_accums[1340]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1341]), .RECT1_Y(rectangle1_ys[1341]), .RECT1_WIDTH(rectangle1_widths[1341]), .RECT1_HEIGHT(rectangle1_heights[1341]), .RECT1_WEIGHT(rectangle1_weights[1341]), .RECT2_X(rectangle2_xs[1341]), .RECT2_Y(rectangle2_ys[1341]), .RECT2_WIDTH(rectangle2_widths[1341]), .RECT2_HEIGHT(rectangle2_heights[1341]), .RECT2_WEIGHT(rectangle2_weights[1341]), .RECT3_X(rectangle3_xs[1341]), .RECT3_Y(rectangle3_ys[1341]), .RECT3_WIDTH(rectangle3_widths[1341]), .RECT3_HEIGHT(rectangle3_heights[1341]), .RECT3_WEIGHT(rectangle3_weights[1341]), .FEAT_THRES(feature_thresholds[1341]), .FEAT_ABOVE(feature_aboves[1341]), .FEAT_BELOW(feature_belows[1341])) ac1341(.scan_win(scan_win1341), .scan_win_std_dev(scan_win_std_dev[1341]), .feature_accum(feature_accums[1341]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1342]), .RECT1_Y(rectangle1_ys[1342]), .RECT1_WIDTH(rectangle1_widths[1342]), .RECT1_HEIGHT(rectangle1_heights[1342]), .RECT1_WEIGHT(rectangle1_weights[1342]), .RECT2_X(rectangle2_xs[1342]), .RECT2_Y(rectangle2_ys[1342]), .RECT2_WIDTH(rectangle2_widths[1342]), .RECT2_HEIGHT(rectangle2_heights[1342]), .RECT2_WEIGHT(rectangle2_weights[1342]), .RECT3_X(rectangle3_xs[1342]), .RECT3_Y(rectangle3_ys[1342]), .RECT3_WIDTH(rectangle3_widths[1342]), .RECT3_HEIGHT(rectangle3_heights[1342]), .RECT3_WEIGHT(rectangle3_weights[1342]), .FEAT_THRES(feature_thresholds[1342]), .FEAT_ABOVE(feature_aboves[1342]), .FEAT_BELOW(feature_belows[1342])) ac1342(.scan_win(scan_win1342), .scan_win_std_dev(scan_win_std_dev[1342]), .feature_accum(feature_accums[1342]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1343]), .RECT1_Y(rectangle1_ys[1343]), .RECT1_WIDTH(rectangle1_widths[1343]), .RECT1_HEIGHT(rectangle1_heights[1343]), .RECT1_WEIGHT(rectangle1_weights[1343]), .RECT2_X(rectangle2_xs[1343]), .RECT2_Y(rectangle2_ys[1343]), .RECT2_WIDTH(rectangle2_widths[1343]), .RECT2_HEIGHT(rectangle2_heights[1343]), .RECT2_WEIGHT(rectangle2_weights[1343]), .RECT3_X(rectangle3_xs[1343]), .RECT3_Y(rectangle3_ys[1343]), .RECT3_WIDTH(rectangle3_widths[1343]), .RECT3_HEIGHT(rectangle3_heights[1343]), .RECT3_WEIGHT(rectangle3_weights[1343]), .FEAT_THRES(feature_thresholds[1343]), .FEAT_ABOVE(feature_aboves[1343]), .FEAT_BELOW(feature_belows[1343])) ac1343(.scan_win(scan_win1343), .scan_win_std_dev(scan_win_std_dev[1343]), .feature_accum(feature_accums[1343]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1344]), .RECT1_Y(rectangle1_ys[1344]), .RECT1_WIDTH(rectangle1_widths[1344]), .RECT1_HEIGHT(rectangle1_heights[1344]), .RECT1_WEIGHT(rectangle1_weights[1344]), .RECT2_X(rectangle2_xs[1344]), .RECT2_Y(rectangle2_ys[1344]), .RECT2_WIDTH(rectangle2_widths[1344]), .RECT2_HEIGHT(rectangle2_heights[1344]), .RECT2_WEIGHT(rectangle2_weights[1344]), .RECT3_X(rectangle3_xs[1344]), .RECT3_Y(rectangle3_ys[1344]), .RECT3_WIDTH(rectangle3_widths[1344]), .RECT3_HEIGHT(rectangle3_heights[1344]), .RECT3_WEIGHT(rectangle3_weights[1344]), .FEAT_THRES(feature_thresholds[1344]), .FEAT_ABOVE(feature_aboves[1344]), .FEAT_BELOW(feature_belows[1344])) ac1344(.scan_win(scan_win1344), .scan_win_std_dev(scan_win_std_dev[1344]), .feature_accum(feature_accums[1344]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1345]), .RECT1_Y(rectangle1_ys[1345]), .RECT1_WIDTH(rectangle1_widths[1345]), .RECT1_HEIGHT(rectangle1_heights[1345]), .RECT1_WEIGHT(rectangle1_weights[1345]), .RECT2_X(rectangle2_xs[1345]), .RECT2_Y(rectangle2_ys[1345]), .RECT2_WIDTH(rectangle2_widths[1345]), .RECT2_HEIGHT(rectangle2_heights[1345]), .RECT2_WEIGHT(rectangle2_weights[1345]), .RECT3_X(rectangle3_xs[1345]), .RECT3_Y(rectangle3_ys[1345]), .RECT3_WIDTH(rectangle3_widths[1345]), .RECT3_HEIGHT(rectangle3_heights[1345]), .RECT3_WEIGHT(rectangle3_weights[1345]), .FEAT_THRES(feature_thresholds[1345]), .FEAT_ABOVE(feature_aboves[1345]), .FEAT_BELOW(feature_belows[1345])) ac1345(.scan_win(scan_win1345), .scan_win_std_dev(scan_win_std_dev[1345]), .feature_accum(feature_accums[1345]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1346]), .RECT1_Y(rectangle1_ys[1346]), .RECT1_WIDTH(rectangle1_widths[1346]), .RECT1_HEIGHT(rectangle1_heights[1346]), .RECT1_WEIGHT(rectangle1_weights[1346]), .RECT2_X(rectangle2_xs[1346]), .RECT2_Y(rectangle2_ys[1346]), .RECT2_WIDTH(rectangle2_widths[1346]), .RECT2_HEIGHT(rectangle2_heights[1346]), .RECT2_WEIGHT(rectangle2_weights[1346]), .RECT3_X(rectangle3_xs[1346]), .RECT3_Y(rectangle3_ys[1346]), .RECT3_WIDTH(rectangle3_widths[1346]), .RECT3_HEIGHT(rectangle3_heights[1346]), .RECT3_WEIGHT(rectangle3_weights[1346]), .FEAT_THRES(feature_thresholds[1346]), .FEAT_ABOVE(feature_aboves[1346]), .FEAT_BELOW(feature_belows[1346])) ac1346(.scan_win(scan_win1346), .scan_win_std_dev(scan_win_std_dev[1346]), .feature_accum(feature_accums[1346]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1347]), .RECT1_Y(rectangle1_ys[1347]), .RECT1_WIDTH(rectangle1_widths[1347]), .RECT1_HEIGHT(rectangle1_heights[1347]), .RECT1_WEIGHT(rectangle1_weights[1347]), .RECT2_X(rectangle2_xs[1347]), .RECT2_Y(rectangle2_ys[1347]), .RECT2_WIDTH(rectangle2_widths[1347]), .RECT2_HEIGHT(rectangle2_heights[1347]), .RECT2_WEIGHT(rectangle2_weights[1347]), .RECT3_X(rectangle3_xs[1347]), .RECT3_Y(rectangle3_ys[1347]), .RECT3_WIDTH(rectangle3_widths[1347]), .RECT3_HEIGHT(rectangle3_heights[1347]), .RECT3_WEIGHT(rectangle3_weights[1347]), .FEAT_THRES(feature_thresholds[1347]), .FEAT_ABOVE(feature_aboves[1347]), .FEAT_BELOW(feature_belows[1347])) ac1347(.scan_win(scan_win1347), .scan_win_std_dev(scan_win_std_dev[1347]), .feature_accum(feature_accums[1347]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1348]), .RECT1_Y(rectangle1_ys[1348]), .RECT1_WIDTH(rectangle1_widths[1348]), .RECT1_HEIGHT(rectangle1_heights[1348]), .RECT1_WEIGHT(rectangle1_weights[1348]), .RECT2_X(rectangle2_xs[1348]), .RECT2_Y(rectangle2_ys[1348]), .RECT2_WIDTH(rectangle2_widths[1348]), .RECT2_HEIGHT(rectangle2_heights[1348]), .RECT2_WEIGHT(rectangle2_weights[1348]), .RECT3_X(rectangle3_xs[1348]), .RECT3_Y(rectangle3_ys[1348]), .RECT3_WIDTH(rectangle3_widths[1348]), .RECT3_HEIGHT(rectangle3_heights[1348]), .RECT3_WEIGHT(rectangle3_weights[1348]), .FEAT_THRES(feature_thresholds[1348]), .FEAT_ABOVE(feature_aboves[1348]), .FEAT_BELOW(feature_belows[1348])) ac1348(.scan_win(scan_win1348), .scan_win_std_dev(scan_win_std_dev[1348]), .feature_accum(feature_accums[1348]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1349]), .RECT1_Y(rectangle1_ys[1349]), .RECT1_WIDTH(rectangle1_widths[1349]), .RECT1_HEIGHT(rectangle1_heights[1349]), .RECT1_WEIGHT(rectangle1_weights[1349]), .RECT2_X(rectangle2_xs[1349]), .RECT2_Y(rectangle2_ys[1349]), .RECT2_WIDTH(rectangle2_widths[1349]), .RECT2_HEIGHT(rectangle2_heights[1349]), .RECT2_WEIGHT(rectangle2_weights[1349]), .RECT3_X(rectangle3_xs[1349]), .RECT3_Y(rectangle3_ys[1349]), .RECT3_WIDTH(rectangle3_widths[1349]), .RECT3_HEIGHT(rectangle3_heights[1349]), .RECT3_WEIGHT(rectangle3_weights[1349]), .FEAT_THRES(feature_thresholds[1349]), .FEAT_ABOVE(feature_aboves[1349]), .FEAT_BELOW(feature_belows[1349])) ac1349(.scan_win(scan_win1349), .scan_win_std_dev(scan_win_std_dev[1349]), .feature_accum(feature_accums[1349]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1350]), .RECT1_Y(rectangle1_ys[1350]), .RECT1_WIDTH(rectangle1_widths[1350]), .RECT1_HEIGHT(rectangle1_heights[1350]), .RECT1_WEIGHT(rectangle1_weights[1350]), .RECT2_X(rectangle2_xs[1350]), .RECT2_Y(rectangle2_ys[1350]), .RECT2_WIDTH(rectangle2_widths[1350]), .RECT2_HEIGHT(rectangle2_heights[1350]), .RECT2_WEIGHT(rectangle2_weights[1350]), .RECT3_X(rectangle3_xs[1350]), .RECT3_Y(rectangle3_ys[1350]), .RECT3_WIDTH(rectangle3_widths[1350]), .RECT3_HEIGHT(rectangle3_heights[1350]), .RECT3_WEIGHT(rectangle3_weights[1350]), .FEAT_THRES(feature_thresholds[1350]), .FEAT_ABOVE(feature_aboves[1350]), .FEAT_BELOW(feature_belows[1350])) ac1350(.scan_win(scan_win1350), .scan_win_std_dev(scan_win_std_dev[1350]), .feature_accum(feature_accums[1350]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1351]), .RECT1_Y(rectangle1_ys[1351]), .RECT1_WIDTH(rectangle1_widths[1351]), .RECT1_HEIGHT(rectangle1_heights[1351]), .RECT1_WEIGHT(rectangle1_weights[1351]), .RECT2_X(rectangle2_xs[1351]), .RECT2_Y(rectangle2_ys[1351]), .RECT2_WIDTH(rectangle2_widths[1351]), .RECT2_HEIGHT(rectangle2_heights[1351]), .RECT2_WEIGHT(rectangle2_weights[1351]), .RECT3_X(rectangle3_xs[1351]), .RECT3_Y(rectangle3_ys[1351]), .RECT3_WIDTH(rectangle3_widths[1351]), .RECT3_HEIGHT(rectangle3_heights[1351]), .RECT3_WEIGHT(rectangle3_weights[1351]), .FEAT_THRES(feature_thresholds[1351]), .FEAT_ABOVE(feature_aboves[1351]), .FEAT_BELOW(feature_belows[1351])) ac1351(.scan_win(scan_win1351), .scan_win_std_dev(scan_win_std_dev[1351]), .feature_accum(feature_accums[1351]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1352]), .RECT1_Y(rectangle1_ys[1352]), .RECT1_WIDTH(rectangle1_widths[1352]), .RECT1_HEIGHT(rectangle1_heights[1352]), .RECT1_WEIGHT(rectangle1_weights[1352]), .RECT2_X(rectangle2_xs[1352]), .RECT2_Y(rectangle2_ys[1352]), .RECT2_WIDTH(rectangle2_widths[1352]), .RECT2_HEIGHT(rectangle2_heights[1352]), .RECT2_WEIGHT(rectangle2_weights[1352]), .RECT3_X(rectangle3_xs[1352]), .RECT3_Y(rectangle3_ys[1352]), .RECT3_WIDTH(rectangle3_widths[1352]), .RECT3_HEIGHT(rectangle3_heights[1352]), .RECT3_WEIGHT(rectangle3_weights[1352]), .FEAT_THRES(feature_thresholds[1352]), .FEAT_ABOVE(feature_aboves[1352]), .FEAT_BELOW(feature_belows[1352])) ac1352(.scan_win(scan_win1352), .scan_win_std_dev(scan_win_std_dev[1352]), .feature_accum(feature_accums[1352]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1353]), .RECT1_Y(rectangle1_ys[1353]), .RECT1_WIDTH(rectangle1_widths[1353]), .RECT1_HEIGHT(rectangle1_heights[1353]), .RECT1_WEIGHT(rectangle1_weights[1353]), .RECT2_X(rectangle2_xs[1353]), .RECT2_Y(rectangle2_ys[1353]), .RECT2_WIDTH(rectangle2_widths[1353]), .RECT2_HEIGHT(rectangle2_heights[1353]), .RECT2_WEIGHT(rectangle2_weights[1353]), .RECT3_X(rectangle3_xs[1353]), .RECT3_Y(rectangle3_ys[1353]), .RECT3_WIDTH(rectangle3_widths[1353]), .RECT3_HEIGHT(rectangle3_heights[1353]), .RECT3_WEIGHT(rectangle3_weights[1353]), .FEAT_THRES(feature_thresholds[1353]), .FEAT_ABOVE(feature_aboves[1353]), .FEAT_BELOW(feature_belows[1353])) ac1353(.scan_win(scan_win1353), .scan_win_std_dev(scan_win_std_dev[1353]), .feature_accum(feature_accums[1353]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1354]), .RECT1_Y(rectangle1_ys[1354]), .RECT1_WIDTH(rectangle1_widths[1354]), .RECT1_HEIGHT(rectangle1_heights[1354]), .RECT1_WEIGHT(rectangle1_weights[1354]), .RECT2_X(rectangle2_xs[1354]), .RECT2_Y(rectangle2_ys[1354]), .RECT2_WIDTH(rectangle2_widths[1354]), .RECT2_HEIGHT(rectangle2_heights[1354]), .RECT2_WEIGHT(rectangle2_weights[1354]), .RECT3_X(rectangle3_xs[1354]), .RECT3_Y(rectangle3_ys[1354]), .RECT3_WIDTH(rectangle3_widths[1354]), .RECT3_HEIGHT(rectangle3_heights[1354]), .RECT3_WEIGHT(rectangle3_weights[1354]), .FEAT_THRES(feature_thresholds[1354]), .FEAT_ABOVE(feature_aboves[1354]), .FEAT_BELOW(feature_belows[1354])) ac1354(.scan_win(scan_win1354), .scan_win_std_dev(scan_win_std_dev[1354]), .feature_accum(feature_accums[1354]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1355]), .RECT1_Y(rectangle1_ys[1355]), .RECT1_WIDTH(rectangle1_widths[1355]), .RECT1_HEIGHT(rectangle1_heights[1355]), .RECT1_WEIGHT(rectangle1_weights[1355]), .RECT2_X(rectangle2_xs[1355]), .RECT2_Y(rectangle2_ys[1355]), .RECT2_WIDTH(rectangle2_widths[1355]), .RECT2_HEIGHT(rectangle2_heights[1355]), .RECT2_WEIGHT(rectangle2_weights[1355]), .RECT3_X(rectangle3_xs[1355]), .RECT3_Y(rectangle3_ys[1355]), .RECT3_WIDTH(rectangle3_widths[1355]), .RECT3_HEIGHT(rectangle3_heights[1355]), .RECT3_WEIGHT(rectangle3_weights[1355]), .FEAT_THRES(feature_thresholds[1355]), .FEAT_ABOVE(feature_aboves[1355]), .FEAT_BELOW(feature_belows[1355])) ac1355(.scan_win(scan_win1355), .scan_win_std_dev(scan_win_std_dev[1355]), .feature_accum(feature_accums[1355]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1356]), .RECT1_Y(rectangle1_ys[1356]), .RECT1_WIDTH(rectangle1_widths[1356]), .RECT1_HEIGHT(rectangle1_heights[1356]), .RECT1_WEIGHT(rectangle1_weights[1356]), .RECT2_X(rectangle2_xs[1356]), .RECT2_Y(rectangle2_ys[1356]), .RECT2_WIDTH(rectangle2_widths[1356]), .RECT2_HEIGHT(rectangle2_heights[1356]), .RECT2_WEIGHT(rectangle2_weights[1356]), .RECT3_X(rectangle3_xs[1356]), .RECT3_Y(rectangle3_ys[1356]), .RECT3_WIDTH(rectangle3_widths[1356]), .RECT3_HEIGHT(rectangle3_heights[1356]), .RECT3_WEIGHT(rectangle3_weights[1356]), .FEAT_THRES(feature_thresholds[1356]), .FEAT_ABOVE(feature_aboves[1356]), .FEAT_BELOW(feature_belows[1356])) ac1356(.scan_win(scan_win1356), .scan_win_std_dev(scan_win_std_dev[1356]), .feature_accum(feature_accums[1356]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1357]), .RECT1_Y(rectangle1_ys[1357]), .RECT1_WIDTH(rectangle1_widths[1357]), .RECT1_HEIGHT(rectangle1_heights[1357]), .RECT1_WEIGHT(rectangle1_weights[1357]), .RECT2_X(rectangle2_xs[1357]), .RECT2_Y(rectangle2_ys[1357]), .RECT2_WIDTH(rectangle2_widths[1357]), .RECT2_HEIGHT(rectangle2_heights[1357]), .RECT2_WEIGHT(rectangle2_weights[1357]), .RECT3_X(rectangle3_xs[1357]), .RECT3_Y(rectangle3_ys[1357]), .RECT3_WIDTH(rectangle3_widths[1357]), .RECT3_HEIGHT(rectangle3_heights[1357]), .RECT3_WEIGHT(rectangle3_weights[1357]), .FEAT_THRES(feature_thresholds[1357]), .FEAT_ABOVE(feature_aboves[1357]), .FEAT_BELOW(feature_belows[1357])) ac1357(.scan_win(scan_win1357), .scan_win_std_dev(scan_win_std_dev[1357]), .feature_accum(feature_accums[1357]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1358]), .RECT1_Y(rectangle1_ys[1358]), .RECT1_WIDTH(rectangle1_widths[1358]), .RECT1_HEIGHT(rectangle1_heights[1358]), .RECT1_WEIGHT(rectangle1_weights[1358]), .RECT2_X(rectangle2_xs[1358]), .RECT2_Y(rectangle2_ys[1358]), .RECT2_WIDTH(rectangle2_widths[1358]), .RECT2_HEIGHT(rectangle2_heights[1358]), .RECT2_WEIGHT(rectangle2_weights[1358]), .RECT3_X(rectangle3_xs[1358]), .RECT3_Y(rectangle3_ys[1358]), .RECT3_WIDTH(rectangle3_widths[1358]), .RECT3_HEIGHT(rectangle3_heights[1358]), .RECT3_WEIGHT(rectangle3_weights[1358]), .FEAT_THRES(feature_thresholds[1358]), .FEAT_ABOVE(feature_aboves[1358]), .FEAT_BELOW(feature_belows[1358])) ac1358(.scan_win(scan_win1358), .scan_win_std_dev(scan_win_std_dev[1358]), .feature_accum(feature_accums[1358]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1359]), .RECT1_Y(rectangle1_ys[1359]), .RECT1_WIDTH(rectangle1_widths[1359]), .RECT1_HEIGHT(rectangle1_heights[1359]), .RECT1_WEIGHT(rectangle1_weights[1359]), .RECT2_X(rectangle2_xs[1359]), .RECT2_Y(rectangle2_ys[1359]), .RECT2_WIDTH(rectangle2_widths[1359]), .RECT2_HEIGHT(rectangle2_heights[1359]), .RECT2_WEIGHT(rectangle2_weights[1359]), .RECT3_X(rectangle3_xs[1359]), .RECT3_Y(rectangle3_ys[1359]), .RECT3_WIDTH(rectangle3_widths[1359]), .RECT3_HEIGHT(rectangle3_heights[1359]), .RECT3_WEIGHT(rectangle3_weights[1359]), .FEAT_THRES(feature_thresholds[1359]), .FEAT_ABOVE(feature_aboves[1359]), .FEAT_BELOW(feature_belows[1359])) ac1359(.scan_win(scan_win1359), .scan_win_std_dev(scan_win_std_dev[1359]), .feature_accum(feature_accums[1359]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1360]), .RECT1_Y(rectangle1_ys[1360]), .RECT1_WIDTH(rectangle1_widths[1360]), .RECT1_HEIGHT(rectangle1_heights[1360]), .RECT1_WEIGHT(rectangle1_weights[1360]), .RECT2_X(rectangle2_xs[1360]), .RECT2_Y(rectangle2_ys[1360]), .RECT2_WIDTH(rectangle2_widths[1360]), .RECT2_HEIGHT(rectangle2_heights[1360]), .RECT2_WEIGHT(rectangle2_weights[1360]), .RECT3_X(rectangle3_xs[1360]), .RECT3_Y(rectangle3_ys[1360]), .RECT3_WIDTH(rectangle3_widths[1360]), .RECT3_HEIGHT(rectangle3_heights[1360]), .RECT3_WEIGHT(rectangle3_weights[1360]), .FEAT_THRES(feature_thresholds[1360]), .FEAT_ABOVE(feature_aboves[1360]), .FEAT_BELOW(feature_belows[1360])) ac1360(.scan_win(scan_win1360), .scan_win_std_dev(scan_win_std_dev[1360]), .feature_accum(feature_accums[1360]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1361]), .RECT1_Y(rectangle1_ys[1361]), .RECT1_WIDTH(rectangle1_widths[1361]), .RECT1_HEIGHT(rectangle1_heights[1361]), .RECT1_WEIGHT(rectangle1_weights[1361]), .RECT2_X(rectangle2_xs[1361]), .RECT2_Y(rectangle2_ys[1361]), .RECT2_WIDTH(rectangle2_widths[1361]), .RECT2_HEIGHT(rectangle2_heights[1361]), .RECT2_WEIGHT(rectangle2_weights[1361]), .RECT3_X(rectangle3_xs[1361]), .RECT3_Y(rectangle3_ys[1361]), .RECT3_WIDTH(rectangle3_widths[1361]), .RECT3_HEIGHT(rectangle3_heights[1361]), .RECT3_WEIGHT(rectangle3_weights[1361]), .FEAT_THRES(feature_thresholds[1361]), .FEAT_ABOVE(feature_aboves[1361]), .FEAT_BELOW(feature_belows[1361])) ac1361(.scan_win(scan_win1361), .scan_win_std_dev(scan_win_std_dev[1361]), .feature_accum(feature_accums[1361]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1362]), .RECT1_Y(rectangle1_ys[1362]), .RECT1_WIDTH(rectangle1_widths[1362]), .RECT1_HEIGHT(rectangle1_heights[1362]), .RECT1_WEIGHT(rectangle1_weights[1362]), .RECT2_X(rectangle2_xs[1362]), .RECT2_Y(rectangle2_ys[1362]), .RECT2_WIDTH(rectangle2_widths[1362]), .RECT2_HEIGHT(rectangle2_heights[1362]), .RECT2_WEIGHT(rectangle2_weights[1362]), .RECT3_X(rectangle3_xs[1362]), .RECT3_Y(rectangle3_ys[1362]), .RECT3_WIDTH(rectangle3_widths[1362]), .RECT3_HEIGHT(rectangle3_heights[1362]), .RECT3_WEIGHT(rectangle3_weights[1362]), .FEAT_THRES(feature_thresholds[1362]), .FEAT_ABOVE(feature_aboves[1362]), .FEAT_BELOW(feature_belows[1362])) ac1362(.scan_win(scan_win1362), .scan_win_std_dev(scan_win_std_dev[1362]), .feature_accum(feature_accums[1362]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1363]), .RECT1_Y(rectangle1_ys[1363]), .RECT1_WIDTH(rectangle1_widths[1363]), .RECT1_HEIGHT(rectangle1_heights[1363]), .RECT1_WEIGHT(rectangle1_weights[1363]), .RECT2_X(rectangle2_xs[1363]), .RECT2_Y(rectangle2_ys[1363]), .RECT2_WIDTH(rectangle2_widths[1363]), .RECT2_HEIGHT(rectangle2_heights[1363]), .RECT2_WEIGHT(rectangle2_weights[1363]), .RECT3_X(rectangle3_xs[1363]), .RECT3_Y(rectangle3_ys[1363]), .RECT3_WIDTH(rectangle3_widths[1363]), .RECT3_HEIGHT(rectangle3_heights[1363]), .RECT3_WEIGHT(rectangle3_weights[1363]), .FEAT_THRES(feature_thresholds[1363]), .FEAT_ABOVE(feature_aboves[1363]), .FEAT_BELOW(feature_belows[1363])) ac1363(.scan_win(scan_win1363), .scan_win_std_dev(scan_win_std_dev[1363]), .feature_accum(feature_accums[1363]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1364]), .RECT1_Y(rectangle1_ys[1364]), .RECT1_WIDTH(rectangle1_widths[1364]), .RECT1_HEIGHT(rectangle1_heights[1364]), .RECT1_WEIGHT(rectangle1_weights[1364]), .RECT2_X(rectangle2_xs[1364]), .RECT2_Y(rectangle2_ys[1364]), .RECT2_WIDTH(rectangle2_widths[1364]), .RECT2_HEIGHT(rectangle2_heights[1364]), .RECT2_WEIGHT(rectangle2_weights[1364]), .RECT3_X(rectangle3_xs[1364]), .RECT3_Y(rectangle3_ys[1364]), .RECT3_WIDTH(rectangle3_widths[1364]), .RECT3_HEIGHT(rectangle3_heights[1364]), .RECT3_WEIGHT(rectangle3_weights[1364]), .FEAT_THRES(feature_thresholds[1364]), .FEAT_ABOVE(feature_aboves[1364]), .FEAT_BELOW(feature_belows[1364])) ac1364(.scan_win(scan_win1364), .scan_win_std_dev(scan_win_std_dev[1364]), .feature_accum(feature_accums[1364]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1365]), .RECT1_Y(rectangle1_ys[1365]), .RECT1_WIDTH(rectangle1_widths[1365]), .RECT1_HEIGHT(rectangle1_heights[1365]), .RECT1_WEIGHT(rectangle1_weights[1365]), .RECT2_X(rectangle2_xs[1365]), .RECT2_Y(rectangle2_ys[1365]), .RECT2_WIDTH(rectangle2_widths[1365]), .RECT2_HEIGHT(rectangle2_heights[1365]), .RECT2_WEIGHT(rectangle2_weights[1365]), .RECT3_X(rectangle3_xs[1365]), .RECT3_Y(rectangle3_ys[1365]), .RECT3_WIDTH(rectangle3_widths[1365]), .RECT3_HEIGHT(rectangle3_heights[1365]), .RECT3_WEIGHT(rectangle3_weights[1365]), .FEAT_THRES(feature_thresholds[1365]), .FEAT_ABOVE(feature_aboves[1365]), .FEAT_BELOW(feature_belows[1365])) ac1365(.scan_win(scan_win1365), .scan_win_std_dev(scan_win_std_dev[1365]), .feature_accum(feature_accums[1365]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1366]), .RECT1_Y(rectangle1_ys[1366]), .RECT1_WIDTH(rectangle1_widths[1366]), .RECT1_HEIGHT(rectangle1_heights[1366]), .RECT1_WEIGHT(rectangle1_weights[1366]), .RECT2_X(rectangle2_xs[1366]), .RECT2_Y(rectangle2_ys[1366]), .RECT2_WIDTH(rectangle2_widths[1366]), .RECT2_HEIGHT(rectangle2_heights[1366]), .RECT2_WEIGHT(rectangle2_weights[1366]), .RECT3_X(rectangle3_xs[1366]), .RECT3_Y(rectangle3_ys[1366]), .RECT3_WIDTH(rectangle3_widths[1366]), .RECT3_HEIGHT(rectangle3_heights[1366]), .RECT3_WEIGHT(rectangle3_weights[1366]), .FEAT_THRES(feature_thresholds[1366]), .FEAT_ABOVE(feature_aboves[1366]), .FEAT_BELOW(feature_belows[1366])) ac1366(.scan_win(scan_win1366), .scan_win_std_dev(scan_win_std_dev[1366]), .feature_accum(feature_accums[1366]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1367]), .RECT1_Y(rectangle1_ys[1367]), .RECT1_WIDTH(rectangle1_widths[1367]), .RECT1_HEIGHT(rectangle1_heights[1367]), .RECT1_WEIGHT(rectangle1_weights[1367]), .RECT2_X(rectangle2_xs[1367]), .RECT2_Y(rectangle2_ys[1367]), .RECT2_WIDTH(rectangle2_widths[1367]), .RECT2_HEIGHT(rectangle2_heights[1367]), .RECT2_WEIGHT(rectangle2_weights[1367]), .RECT3_X(rectangle3_xs[1367]), .RECT3_Y(rectangle3_ys[1367]), .RECT3_WIDTH(rectangle3_widths[1367]), .RECT3_HEIGHT(rectangle3_heights[1367]), .RECT3_WEIGHT(rectangle3_weights[1367]), .FEAT_THRES(feature_thresholds[1367]), .FEAT_ABOVE(feature_aboves[1367]), .FEAT_BELOW(feature_belows[1367])) ac1367(.scan_win(scan_win1367), .scan_win_std_dev(scan_win_std_dev[1367]), .feature_accum(feature_accums[1367]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1368]), .RECT1_Y(rectangle1_ys[1368]), .RECT1_WIDTH(rectangle1_widths[1368]), .RECT1_HEIGHT(rectangle1_heights[1368]), .RECT1_WEIGHT(rectangle1_weights[1368]), .RECT2_X(rectangle2_xs[1368]), .RECT2_Y(rectangle2_ys[1368]), .RECT2_WIDTH(rectangle2_widths[1368]), .RECT2_HEIGHT(rectangle2_heights[1368]), .RECT2_WEIGHT(rectangle2_weights[1368]), .RECT3_X(rectangle3_xs[1368]), .RECT3_Y(rectangle3_ys[1368]), .RECT3_WIDTH(rectangle3_widths[1368]), .RECT3_HEIGHT(rectangle3_heights[1368]), .RECT3_WEIGHT(rectangle3_weights[1368]), .FEAT_THRES(feature_thresholds[1368]), .FEAT_ABOVE(feature_aboves[1368]), .FEAT_BELOW(feature_belows[1368])) ac1368(.scan_win(scan_win1368), .scan_win_std_dev(scan_win_std_dev[1368]), .feature_accum(feature_accums[1368]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1369]), .RECT1_Y(rectangle1_ys[1369]), .RECT1_WIDTH(rectangle1_widths[1369]), .RECT1_HEIGHT(rectangle1_heights[1369]), .RECT1_WEIGHT(rectangle1_weights[1369]), .RECT2_X(rectangle2_xs[1369]), .RECT2_Y(rectangle2_ys[1369]), .RECT2_WIDTH(rectangle2_widths[1369]), .RECT2_HEIGHT(rectangle2_heights[1369]), .RECT2_WEIGHT(rectangle2_weights[1369]), .RECT3_X(rectangle3_xs[1369]), .RECT3_Y(rectangle3_ys[1369]), .RECT3_WIDTH(rectangle3_widths[1369]), .RECT3_HEIGHT(rectangle3_heights[1369]), .RECT3_WEIGHT(rectangle3_weights[1369]), .FEAT_THRES(feature_thresholds[1369]), .FEAT_ABOVE(feature_aboves[1369]), .FEAT_BELOW(feature_belows[1369])) ac1369(.scan_win(scan_win1369), .scan_win_std_dev(scan_win_std_dev[1369]), .feature_accum(feature_accums[1369]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1370]), .RECT1_Y(rectangle1_ys[1370]), .RECT1_WIDTH(rectangle1_widths[1370]), .RECT1_HEIGHT(rectangle1_heights[1370]), .RECT1_WEIGHT(rectangle1_weights[1370]), .RECT2_X(rectangle2_xs[1370]), .RECT2_Y(rectangle2_ys[1370]), .RECT2_WIDTH(rectangle2_widths[1370]), .RECT2_HEIGHT(rectangle2_heights[1370]), .RECT2_WEIGHT(rectangle2_weights[1370]), .RECT3_X(rectangle3_xs[1370]), .RECT3_Y(rectangle3_ys[1370]), .RECT3_WIDTH(rectangle3_widths[1370]), .RECT3_HEIGHT(rectangle3_heights[1370]), .RECT3_WEIGHT(rectangle3_weights[1370]), .FEAT_THRES(feature_thresholds[1370]), .FEAT_ABOVE(feature_aboves[1370]), .FEAT_BELOW(feature_belows[1370])) ac1370(.scan_win(scan_win1370), .scan_win_std_dev(scan_win_std_dev[1370]), .feature_accum(feature_accums[1370]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1371]), .RECT1_Y(rectangle1_ys[1371]), .RECT1_WIDTH(rectangle1_widths[1371]), .RECT1_HEIGHT(rectangle1_heights[1371]), .RECT1_WEIGHT(rectangle1_weights[1371]), .RECT2_X(rectangle2_xs[1371]), .RECT2_Y(rectangle2_ys[1371]), .RECT2_WIDTH(rectangle2_widths[1371]), .RECT2_HEIGHT(rectangle2_heights[1371]), .RECT2_WEIGHT(rectangle2_weights[1371]), .RECT3_X(rectangle3_xs[1371]), .RECT3_Y(rectangle3_ys[1371]), .RECT3_WIDTH(rectangle3_widths[1371]), .RECT3_HEIGHT(rectangle3_heights[1371]), .RECT3_WEIGHT(rectangle3_weights[1371]), .FEAT_THRES(feature_thresholds[1371]), .FEAT_ABOVE(feature_aboves[1371]), .FEAT_BELOW(feature_belows[1371])) ac1371(.scan_win(scan_win1371), .scan_win_std_dev(scan_win_std_dev[1371]), .feature_accum(feature_accums[1371]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1372]), .RECT1_Y(rectangle1_ys[1372]), .RECT1_WIDTH(rectangle1_widths[1372]), .RECT1_HEIGHT(rectangle1_heights[1372]), .RECT1_WEIGHT(rectangle1_weights[1372]), .RECT2_X(rectangle2_xs[1372]), .RECT2_Y(rectangle2_ys[1372]), .RECT2_WIDTH(rectangle2_widths[1372]), .RECT2_HEIGHT(rectangle2_heights[1372]), .RECT2_WEIGHT(rectangle2_weights[1372]), .RECT3_X(rectangle3_xs[1372]), .RECT3_Y(rectangle3_ys[1372]), .RECT3_WIDTH(rectangle3_widths[1372]), .RECT3_HEIGHT(rectangle3_heights[1372]), .RECT3_WEIGHT(rectangle3_weights[1372]), .FEAT_THRES(feature_thresholds[1372]), .FEAT_ABOVE(feature_aboves[1372]), .FEAT_BELOW(feature_belows[1372])) ac1372(.scan_win(scan_win1372), .scan_win_std_dev(scan_win_std_dev[1372]), .feature_accum(feature_accums[1372]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1373]), .RECT1_Y(rectangle1_ys[1373]), .RECT1_WIDTH(rectangle1_widths[1373]), .RECT1_HEIGHT(rectangle1_heights[1373]), .RECT1_WEIGHT(rectangle1_weights[1373]), .RECT2_X(rectangle2_xs[1373]), .RECT2_Y(rectangle2_ys[1373]), .RECT2_WIDTH(rectangle2_widths[1373]), .RECT2_HEIGHT(rectangle2_heights[1373]), .RECT2_WEIGHT(rectangle2_weights[1373]), .RECT3_X(rectangle3_xs[1373]), .RECT3_Y(rectangle3_ys[1373]), .RECT3_WIDTH(rectangle3_widths[1373]), .RECT3_HEIGHT(rectangle3_heights[1373]), .RECT3_WEIGHT(rectangle3_weights[1373]), .FEAT_THRES(feature_thresholds[1373]), .FEAT_ABOVE(feature_aboves[1373]), .FEAT_BELOW(feature_belows[1373])) ac1373(.scan_win(scan_win1373), .scan_win_std_dev(scan_win_std_dev[1373]), .feature_accum(feature_accums[1373]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1374]), .RECT1_Y(rectangle1_ys[1374]), .RECT1_WIDTH(rectangle1_widths[1374]), .RECT1_HEIGHT(rectangle1_heights[1374]), .RECT1_WEIGHT(rectangle1_weights[1374]), .RECT2_X(rectangle2_xs[1374]), .RECT2_Y(rectangle2_ys[1374]), .RECT2_WIDTH(rectangle2_widths[1374]), .RECT2_HEIGHT(rectangle2_heights[1374]), .RECT2_WEIGHT(rectangle2_weights[1374]), .RECT3_X(rectangle3_xs[1374]), .RECT3_Y(rectangle3_ys[1374]), .RECT3_WIDTH(rectangle3_widths[1374]), .RECT3_HEIGHT(rectangle3_heights[1374]), .RECT3_WEIGHT(rectangle3_weights[1374]), .FEAT_THRES(feature_thresholds[1374]), .FEAT_ABOVE(feature_aboves[1374]), .FEAT_BELOW(feature_belows[1374])) ac1374(.scan_win(scan_win1374), .scan_win_std_dev(scan_win_std_dev[1374]), .feature_accum(feature_accums[1374]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1375]), .RECT1_Y(rectangle1_ys[1375]), .RECT1_WIDTH(rectangle1_widths[1375]), .RECT1_HEIGHT(rectangle1_heights[1375]), .RECT1_WEIGHT(rectangle1_weights[1375]), .RECT2_X(rectangle2_xs[1375]), .RECT2_Y(rectangle2_ys[1375]), .RECT2_WIDTH(rectangle2_widths[1375]), .RECT2_HEIGHT(rectangle2_heights[1375]), .RECT2_WEIGHT(rectangle2_weights[1375]), .RECT3_X(rectangle3_xs[1375]), .RECT3_Y(rectangle3_ys[1375]), .RECT3_WIDTH(rectangle3_widths[1375]), .RECT3_HEIGHT(rectangle3_heights[1375]), .RECT3_WEIGHT(rectangle3_weights[1375]), .FEAT_THRES(feature_thresholds[1375]), .FEAT_ABOVE(feature_aboves[1375]), .FEAT_BELOW(feature_belows[1375])) ac1375(.scan_win(scan_win1375), .scan_win_std_dev(scan_win_std_dev[1375]), .feature_accum(feature_accums[1375]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1376]), .RECT1_Y(rectangle1_ys[1376]), .RECT1_WIDTH(rectangle1_widths[1376]), .RECT1_HEIGHT(rectangle1_heights[1376]), .RECT1_WEIGHT(rectangle1_weights[1376]), .RECT2_X(rectangle2_xs[1376]), .RECT2_Y(rectangle2_ys[1376]), .RECT2_WIDTH(rectangle2_widths[1376]), .RECT2_HEIGHT(rectangle2_heights[1376]), .RECT2_WEIGHT(rectangle2_weights[1376]), .RECT3_X(rectangle3_xs[1376]), .RECT3_Y(rectangle3_ys[1376]), .RECT3_WIDTH(rectangle3_widths[1376]), .RECT3_HEIGHT(rectangle3_heights[1376]), .RECT3_WEIGHT(rectangle3_weights[1376]), .FEAT_THRES(feature_thresholds[1376]), .FEAT_ABOVE(feature_aboves[1376]), .FEAT_BELOW(feature_belows[1376])) ac1376(.scan_win(scan_win1376), .scan_win_std_dev(scan_win_std_dev[1376]), .feature_accum(feature_accums[1376]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1377]), .RECT1_Y(rectangle1_ys[1377]), .RECT1_WIDTH(rectangle1_widths[1377]), .RECT1_HEIGHT(rectangle1_heights[1377]), .RECT1_WEIGHT(rectangle1_weights[1377]), .RECT2_X(rectangle2_xs[1377]), .RECT2_Y(rectangle2_ys[1377]), .RECT2_WIDTH(rectangle2_widths[1377]), .RECT2_HEIGHT(rectangle2_heights[1377]), .RECT2_WEIGHT(rectangle2_weights[1377]), .RECT3_X(rectangle3_xs[1377]), .RECT3_Y(rectangle3_ys[1377]), .RECT3_WIDTH(rectangle3_widths[1377]), .RECT3_HEIGHT(rectangle3_heights[1377]), .RECT3_WEIGHT(rectangle3_weights[1377]), .FEAT_THRES(feature_thresholds[1377]), .FEAT_ABOVE(feature_aboves[1377]), .FEAT_BELOW(feature_belows[1377])) ac1377(.scan_win(scan_win1377), .scan_win_std_dev(scan_win_std_dev[1377]), .feature_accum(feature_accums[1377]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1378]), .RECT1_Y(rectangle1_ys[1378]), .RECT1_WIDTH(rectangle1_widths[1378]), .RECT1_HEIGHT(rectangle1_heights[1378]), .RECT1_WEIGHT(rectangle1_weights[1378]), .RECT2_X(rectangle2_xs[1378]), .RECT2_Y(rectangle2_ys[1378]), .RECT2_WIDTH(rectangle2_widths[1378]), .RECT2_HEIGHT(rectangle2_heights[1378]), .RECT2_WEIGHT(rectangle2_weights[1378]), .RECT3_X(rectangle3_xs[1378]), .RECT3_Y(rectangle3_ys[1378]), .RECT3_WIDTH(rectangle3_widths[1378]), .RECT3_HEIGHT(rectangle3_heights[1378]), .RECT3_WEIGHT(rectangle3_weights[1378]), .FEAT_THRES(feature_thresholds[1378]), .FEAT_ABOVE(feature_aboves[1378]), .FEAT_BELOW(feature_belows[1378])) ac1378(.scan_win(scan_win1378), .scan_win_std_dev(scan_win_std_dev[1378]), .feature_accum(feature_accums[1378]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1379]), .RECT1_Y(rectangle1_ys[1379]), .RECT1_WIDTH(rectangle1_widths[1379]), .RECT1_HEIGHT(rectangle1_heights[1379]), .RECT1_WEIGHT(rectangle1_weights[1379]), .RECT2_X(rectangle2_xs[1379]), .RECT2_Y(rectangle2_ys[1379]), .RECT2_WIDTH(rectangle2_widths[1379]), .RECT2_HEIGHT(rectangle2_heights[1379]), .RECT2_WEIGHT(rectangle2_weights[1379]), .RECT3_X(rectangle3_xs[1379]), .RECT3_Y(rectangle3_ys[1379]), .RECT3_WIDTH(rectangle3_widths[1379]), .RECT3_HEIGHT(rectangle3_heights[1379]), .RECT3_WEIGHT(rectangle3_weights[1379]), .FEAT_THRES(feature_thresholds[1379]), .FEAT_ABOVE(feature_aboves[1379]), .FEAT_BELOW(feature_belows[1379])) ac1379(.scan_win(scan_win1379), .scan_win_std_dev(scan_win_std_dev[1379]), .feature_accum(feature_accums[1379]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1380]), .RECT1_Y(rectangle1_ys[1380]), .RECT1_WIDTH(rectangle1_widths[1380]), .RECT1_HEIGHT(rectangle1_heights[1380]), .RECT1_WEIGHT(rectangle1_weights[1380]), .RECT2_X(rectangle2_xs[1380]), .RECT2_Y(rectangle2_ys[1380]), .RECT2_WIDTH(rectangle2_widths[1380]), .RECT2_HEIGHT(rectangle2_heights[1380]), .RECT2_WEIGHT(rectangle2_weights[1380]), .RECT3_X(rectangle3_xs[1380]), .RECT3_Y(rectangle3_ys[1380]), .RECT3_WIDTH(rectangle3_widths[1380]), .RECT3_HEIGHT(rectangle3_heights[1380]), .RECT3_WEIGHT(rectangle3_weights[1380]), .FEAT_THRES(feature_thresholds[1380]), .FEAT_ABOVE(feature_aboves[1380]), .FEAT_BELOW(feature_belows[1380])) ac1380(.scan_win(scan_win1380), .scan_win_std_dev(scan_win_std_dev[1380]), .feature_accum(feature_accums[1380]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1381]), .RECT1_Y(rectangle1_ys[1381]), .RECT1_WIDTH(rectangle1_widths[1381]), .RECT1_HEIGHT(rectangle1_heights[1381]), .RECT1_WEIGHT(rectangle1_weights[1381]), .RECT2_X(rectangle2_xs[1381]), .RECT2_Y(rectangle2_ys[1381]), .RECT2_WIDTH(rectangle2_widths[1381]), .RECT2_HEIGHT(rectangle2_heights[1381]), .RECT2_WEIGHT(rectangle2_weights[1381]), .RECT3_X(rectangle3_xs[1381]), .RECT3_Y(rectangle3_ys[1381]), .RECT3_WIDTH(rectangle3_widths[1381]), .RECT3_HEIGHT(rectangle3_heights[1381]), .RECT3_WEIGHT(rectangle3_weights[1381]), .FEAT_THRES(feature_thresholds[1381]), .FEAT_ABOVE(feature_aboves[1381]), .FEAT_BELOW(feature_belows[1381])) ac1381(.scan_win(scan_win1381), .scan_win_std_dev(scan_win_std_dev[1381]), .feature_accum(feature_accums[1381]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1382]), .RECT1_Y(rectangle1_ys[1382]), .RECT1_WIDTH(rectangle1_widths[1382]), .RECT1_HEIGHT(rectangle1_heights[1382]), .RECT1_WEIGHT(rectangle1_weights[1382]), .RECT2_X(rectangle2_xs[1382]), .RECT2_Y(rectangle2_ys[1382]), .RECT2_WIDTH(rectangle2_widths[1382]), .RECT2_HEIGHT(rectangle2_heights[1382]), .RECT2_WEIGHT(rectangle2_weights[1382]), .RECT3_X(rectangle3_xs[1382]), .RECT3_Y(rectangle3_ys[1382]), .RECT3_WIDTH(rectangle3_widths[1382]), .RECT3_HEIGHT(rectangle3_heights[1382]), .RECT3_WEIGHT(rectangle3_weights[1382]), .FEAT_THRES(feature_thresholds[1382]), .FEAT_ABOVE(feature_aboves[1382]), .FEAT_BELOW(feature_belows[1382])) ac1382(.scan_win(scan_win1382), .scan_win_std_dev(scan_win_std_dev[1382]), .feature_accum(feature_accums[1382]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1383]), .RECT1_Y(rectangle1_ys[1383]), .RECT1_WIDTH(rectangle1_widths[1383]), .RECT1_HEIGHT(rectangle1_heights[1383]), .RECT1_WEIGHT(rectangle1_weights[1383]), .RECT2_X(rectangle2_xs[1383]), .RECT2_Y(rectangle2_ys[1383]), .RECT2_WIDTH(rectangle2_widths[1383]), .RECT2_HEIGHT(rectangle2_heights[1383]), .RECT2_WEIGHT(rectangle2_weights[1383]), .RECT3_X(rectangle3_xs[1383]), .RECT3_Y(rectangle3_ys[1383]), .RECT3_WIDTH(rectangle3_widths[1383]), .RECT3_HEIGHT(rectangle3_heights[1383]), .RECT3_WEIGHT(rectangle3_weights[1383]), .FEAT_THRES(feature_thresholds[1383]), .FEAT_ABOVE(feature_aboves[1383]), .FEAT_BELOW(feature_belows[1383])) ac1383(.scan_win(scan_win1383), .scan_win_std_dev(scan_win_std_dev[1383]), .feature_accum(feature_accums[1383]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1384]), .RECT1_Y(rectangle1_ys[1384]), .RECT1_WIDTH(rectangle1_widths[1384]), .RECT1_HEIGHT(rectangle1_heights[1384]), .RECT1_WEIGHT(rectangle1_weights[1384]), .RECT2_X(rectangle2_xs[1384]), .RECT2_Y(rectangle2_ys[1384]), .RECT2_WIDTH(rectangle2_widths[1384]), .RECT2_HEIGHT(rectangle2_heights[1384]), .RECT2_WEIGHT(rectangle2_weights[1384]), .RECT3_X(rectangle3_xs[1384]), .RECT3_Y(rectangle3_ys[1384]), .RECT3_WIDTH(rectangle3_widths[1384]), .RECT3_HEIGHT(rectangle3_heights[1384]), .RECT3_WEIGHT(rectangle3_weights[1384]), .FEAT_THRES(feature_thresholds[1384]), .FEAT_ABOVE(feature_aboves[1384]), .FEAT_BELOW(feature_belows[1384])) ac1384(.scan_win(scan_win1384), .scan_win_std_dev(scan_win_std_dev[1384]), .feature_accum(feature_accums[1384]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1385]), .RECT1_Y(rectangle1_ys[1385]), .RECT1_WIDTH(rectangle1_widths[1385]), .RECT1_HEIGHT(rectangle1_heights[1385]), .RECT1_WEIGHT(rectangle1_weights[1385]), .RECT2_X(rectangle2_xs[1385]), .RECT2_Y(rectangle2_ys[1385]), .RECT2_WIDTH(rectangle2_widths[1385]), .RECT2_HEIGHT(rectangle2_heights[1385]), .RECT2_WEIGHT(rectangle2_weights[1385]), .RECT3_X(rectangle3_xs[1385]), .RECT3_Y(rectangle3_ys[1385]), .RECT3_WIDTH(rectangle3_widths[1385]), .RECT3_HEIGHT(rectangle3_heights[1385]), .RECT3_WEIGHT(rectangle3_weights[1385]), .FEAT_THRES(feature_thresholds[1385]), .FEAT_ABOVE(feature_aboves[1385]), .FEAT_BELOW(feature_belows[1385])) ac1385(.scan_win(scan_win1385), .scan_win_std_dev(scan_win_std_dev[1385]), .feature_accum(feature_accums[1385]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1386]), .RECT1_Y(rectangle1_ys[1386]), .RECT1_WIDTH(rectangle1_widths[1386]), .RECT1_HEIGHT(rectangle1_heights[1386]), .RECT1_WEIGHT(rectangle1_weights[1386]), .RECT2_X(rectangle2_xs[1386]), .RECT2_Y(rectangle2_ys[1386]), .RECT2_WIDTH(rectangle2_widths[1386]), .RECT2_HEIGHT(rectangle2_heights[1386]), .RECT2_WEIGHT(rectangle2_weights[1386]), .RECT3_X(rectangle3_xs[1386]), .RECT3_Y(rectangle3_ys[1386]), .RECT3_WIDTH(rectangle3_widths[1386]), .RECT3_HEIGHT(rectangle3_heights[1386]), .RECT3_WEIGHT(rectangle3_weights[1386]), .FEAT_THRES(feature_thresholds[1386]), .FEAT_ABOVE(feature_aboves[1386]), .FEAT_BELOW(feature_belows[1386])) ac1386(.scan_win(scan_win1386), .scan_win_std_dev(scan_win_std_dev[1386]), .feature_accum(feature_accums[1386]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1387]), .RECT1_Y(rectangle1_ys[1387]), .RECT1_WIDTH(rectangle1_widths[1387]), .RECT1_HEIGHT(rectangle1_heights[1387]), .RECT1_WEIGHT(rectangle1_weights[1387]), .RECT2_X(rectangle2_xs[1387]), .RECT2_Y(rectangle2_ys[1387]), .RECT2_WIDTH(rectangle2_widths[1387]), .RECT2_HEIGHT(rectangle2_heights[1387]), .RECT2_WEIGHT(rectangle2_weights[1387]), .RECT3_X(rectangle3_xs[1387]), .RECT3_Y(rectangle3_ys[1387]), .RECT3_WIDTH(rectangle3_widths[1387]), .RECT3_HEIGHT(rectangle3_heights[1387]), .RECT3_WEIGHT(rectangle3_weights[1387]), .FEAT_THRES(feature_thresholds[1387]), .FEAT_ABOVE(feature_aboves[1387]), .FEAT_BELOW(feature_belows[1387])) ac1387(.scan_win(scan_win1387), .scan_win_std_dev(scan_win_std_dev[1387]), .feature_accum(feature_accums[1387]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1388]), .RECT1_Y(rectangle1_ys[1388]), .RECT1_WIDTH(rectangle1_widths[1388]), .RECT1_HEIGHT(rectangle1_heights[1388]), .RECT1_WEIGHT(rectangle1_weights[1388]), .RECT2_X(rectangle2_xs[1388]), .RECT2_Y(rectangle2_ys[1388]), .RECT2_WIDTH(rectangle2_widths[1388]), .RECT2_HEIGHT(rectangle2_heights[1388]), .RECT2_WEIGHT(rectangle2_weights[1388]), .RECT3_X(rectangle3_xs[1388]), .RECT3_Y(rectangle3_ys[1388]), .RECT3_WIDTH(rectangle3_widths[1388]), .RECT3_HEIGHT(rectangle3_heights[1388]), .RECT3_WEIGHT(rectangle3_weights[1388]), .FEAT_THRES(feature_thresholds[1388]), .FEAT_ABOVE(feature_aboves[1388]), .FEAT_BELOW(feature_belows[1388])) ac1388(.scan_win(scan_win1388), .scan_win_std_dev(scan_win_std_dev[1388]), .feature_accum(feature_accums[1388]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1389]), .RECT1_Y(rectangle1_ys[1389]), .RECT1_WIDTH(rectangle1_widths[1389]), .RECT1_HEIGHT(rectangle1_heights[1389]), .RECT1_WEIGHT(rectangle1_weights[1389]), .RECT2_X(rectangle2_xs[1389]), .RECT2_Y(rectangle2_ys[1389]), .RECT2_WIDTH(rectangle2_widths[1389]), .RECT2_HEIGHT(rectangle2_heights[1389]), .RECT2_WEIGHT(rectangle2_weights[1389]), .RECT3_X(rectangle3_xs[1389]), .RECT3_Y(rectangle3_ys[1389]), .RECT3_WIDTH(rectangle3_widths[1389]), .RECT3_HEIGHT(rectangle3_heights[1389]), .RECT3_WEIGHT(rectangle3_weights[1389]), .FEAT_THRES(feature_thresholds[1389]), .FEAT_ABOVE(feature_aboves[1389]), .FEAT_BELOW(feature_belows[1389])) ac1389(.scan_win(scan_win1389), .scan_win_std_dev(scan_win_std_dev[1389]), .feature_accum(feature_accums[1389]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1390]), .RECT1_Y(rectangle1_ys[1390]), .RECT1_WIDTH(rectangle1_widths[1390]), .RECT1_HEIGHT(rectangle1_heights[1390]), .RECT1_WEIGHT(rectangle1_weights[1390]), .RECT2_X(rectangle2_xs[1390]), .RECT2_Y(rectangle2_ys[1390]), .RECT2_WIDTH(rectangle2_widths[1390]), .RECT2_HEIGHT(rectangle2_heights[1390]), .RECT2_WEIGHT(rectangle2_weights[1390]), .RECT3_X(rectangle3_xs[1390]), .RECT3_Y(rectangle3_ys[1390]), .RECT3_WIDTH(rectangle3_widths[1390]), .RECT3_HEIGHT(rectangle3_heights[1390]), .RECT3_WEIGHT(rectangle3_weights[1390]), .FEAT_THRES(feature_thresholds[1390]), .FEAT_ABOVE(feature_aboves[1390]), .FEAT_BELOW(feature_belows[1390])) ac1390(.scan_win(scan_win1390), .scan_win_std_dev(scan_win_std_dev[1390]), .feature_accum(feature_accums[1390]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1391]), .RECT1_Y(rectangle1_ys[1391]), .RECT1_WIDTH(rectangle1_widths[1391]), .RECT1_HEIGHT(rectangle1_heights[1391]), .RECT1_WEIGHT(rectangle1_weights[1391]), .RECT2_X(rectangle2_xs[1391]), .RECT2_Y(rectangle2_ys[1391]), .RECT2_WIDTH(rectangle2_widths[1391]), .RECT2_HEIGHT(rectangle2_heights[1391]), .RECT2_WEIGHT(rectangle2_weights[1391]), .RECT3_X(rectangle3_xs[1391]), .RECT3_Y(rectangle3_ys[1391]), .RECT3_WIDTH(rectangle3_widths[1391]), .RECT3_HEIGHT(rectangle3_heights[1391]), .RECT3_WEIGHT(rectangle3_weights[1391]), .FEAT_THRES(feature_thresholds[1391]), .FEAT_ABOVE(feature_aboves[1391]), .FEAT_BELOW(feature_belows[1391])) ac1391(.scan_win(scan_win1391), .scan_win_std_dev(scan_win_std_dev[1391]), .feature_accum(feature_accums[1391]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1392]), .RECT1_Y(rectangle1_ys[1392]), .RECT1_WIDTH(rectangle1_widths[1392]), .RECT1_HEIGHT(rectangle1_heights[1392]), .RECT1_WEIGHT(rectangle1_weights[1392]), .RECT2_X(rectangle2_xs[1392]), .RECT2_Y(rectangle2_ys[1392]), .RECT2_WIDTH(rectangle2_widths[1392]), .RECT2_HEIGHT(rectangle2_heights[1392]), .RECT2_WEIGHT(rectangle2_weights[1392]), .RECT3_X(rectangle3_xs[1392]), .RECT3_Y(rectangle3_ys[1392]), .RECT3_WIDTH(rectangle3_widths[1392]), .RECT3_HEIGHT(rectangle3_heights[1392]), .RECT3_WEIGHT(rectangle3_weights[1392]), .FEAT_THRES(feature_thresholds[1392]), .FEAT_ABOVE(feature_aboves[1392]), .FEAT_BELOW(feature_belows[1392])) ac1392(.scan_win(scan_win1392), .scan_win_std_dev(scan_win_std_dev[1392]), .feature_accum(feature_accums[1392]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1393]), .RECT1_Y(rectangle1_ys[1393]), .RECT1_WIDTH(rectangle1_widths[1393]), .RECT1_HEIGHT(rectangle1_heights[1393]), .RECT1_WEIGHT(rectangle1_weights[1393]), .RECT2_X(rectangle2_xs[1393]), .RECT2_Y(rectangle2_ys[1393]), .RECT2_WIDTH(rectangle2_widths[1393]), .RECT2_HEIGHT(rectangle2_heights[1393]), .RECT2_WEIGHT(rectangle2_weights[1393]), .RECT3_X(rectangle3_xs[1393]), .RECT3_Y(rectangle3_ys[1393]), .RECT3_WIDTH(rectangle3_widths[1393]), .RECT3_HEIGHT(rectangle3_heights[1393]), .RECT3_WEIGHT(rectangle3_weights[1393]), .FEAT_THRES(feature_thresholds[1393]), .FEAT_ABOVE(feature_aboves[1393]), .FEAT_BELOW(feature_belows[1393])) ac1393(.scan_win(scan_win1393), .scan_win_std_dev(scan_win_std_dev[1393]), .feature_accum(feature_accums[1393]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1394]), .RECT1_Y(rectangle1_ys[1394]), .RECT1_WIDTH(rectangle1_widths[1394]), .RECT1_HEIGHT(rectangle1_heights[1394]), .RECT1_WEIGHT(rectangle1_weights[1394]), .RECT2_X(rectangle2_xs[1394]), .RECT2_Y(rectangle2_ys[1394]), .RECT2_WIDTH(rectangle2_widths[1394]), .RECT2_HEIGHT(rectangle2_heights[1394]), .RECT2_WEIGHT(rectangle2_weights[1394]), .RECT3_X(rectangle3_xs[1394]), .RECT3_Y(rectangle3_ys[1394]), .RECT3_WIDTH(rectangle3_widths[1394]), .RECT3_HEIGHT(rectangle3_heights[1394]), .RECT3_WEIGHT(rectangle3_weights[1394]), .FEAT_THRES(feature_thresholds[1394]), .FEAT_ABOVE(feature_aboves[1394]), .FEAT_BELOW(feature_belows[1394])) ac1394(.scan_win(scan_win1394), .scan_win_std_dev(scan_win_std_dev[1394]), .feature_accum(feature_accums[1394]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1395]), .RECT1_Y(rectangle1_ys[1395]), .RECT1_WIDTH(rectangle1_widths[1395]), .RECT1_HEIGHT(rectangle1_heights[1395]), .RECT1_WEIGHT(rectangle1_weights[1395]), .RECT2_X(rectangle2_xs[1395]), .RECT2_Y(rectangle2_ys[1395]), .RECT2_WIDTH(rectangle2_widths[1395]), .RECT2_HEIGHT(rectangle2_heights[1395]), .RECT2_WEIGHT(rectangle2_weights[1395]), .RECT3_X(rectangle3_xs[1395]), .RECT3_Y(rectangle3_ys[1395]), .RECT3_WIDTH(rectangle3_widths[1395]), .RECT3_HEIGHT(rectangle3_heights[1395]), .RECT3_WEIGHT(rectangle3_weights[1395]), .FEAT_THRES(feature_thresholds[1395]), .FEAT_ABOVE(feature_aboves[1395]), .FEAT_BELOW(feature_belows[1395])) ac1395(.scan_win(scan_win1395), .scan_win_std_dev(scan_win_std_dev[1395]), .feature_accum(feature_accums[1395]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1396]), .RECT1_Y(rectangle1_ys[1396]), .RECT1_WIDTH(rectangle1_widths[1396]), .RECT1_HEIGHT(rectangle1_heights[1396]), .RECT1_WEIGHT(rectangle1_weights[1396]), .RECT2_X(rectangle2_xs[1396]), .RECT2_Y(rectangle2_ys[1396]), .RECT2_WIDTH(rectangle2_widths[1396]), .RECT2_HEIGHT(rectangle2_heights[1396]), .RECT2_WEIGHT(rectangle2_weights[1396]), .RECT3_X(rectangle3_xs[1396]), .RECT3_Y(rectangle3_ys[1396]), .RECT3_WIDTH(rectangle3_widths[1396]), .RECT3_HEIGHT(rectangle3_heights[1396]), .RECT3_WEIGHT(rectangle3_weights[1396]), .FEAT_THRES(feature_thresholds[1396]), .FEAT_ABOVE(feature_aboves[1396]), .FEAT_BELOW(feature_belows[1396])) ac1396(.scan_win(scan_win1396), .scan_win_std_dev(scan_win_std_dev[1396]), .feature_accum(feature_accums[1396]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1397]), .RECT1_Y(rectangle1_ys[1397]), .RECT1_WIDTH(rectangle1_widths[1397]), .RECT1_HEIGHT(rectangle1_heights[1397]), .RECT1_WEIGHT(rectangle1_weights[1397]), .RECT2_X(rectangle2_xs[1397]), .RECT2_Y(rectangle2_ys[1397]), .RECT2_WIDTH(rectangle2_widths[1397]), .RECT2_HEIGHT(rectangle2_heights[1397]), .RECT2_WEIGHT(rectangle2_weights[1397]), .RECT3_X(rectangle3_xs[1397]), .RECT3_Y(rectangle3_ys[1397]), .RECT3_WIDTH(rectangle3_widths[1397]), .RECT3_HEIGHT(rectangle3_heights[1397]), .RECT3_WEIGHT(rectangle3_weights[1397]), .FEAT_THRES(feature_thresholds[1397]), .FEAT_ABOVE(feature_aboves[1397]), .FEAT_BELOW(feature_belows[1397])) ac1397(.scan_win(scan_win1397), .scan_win_std_dev(scan_win_std_dev[1397]), .feature_accum(feature_accums[1397]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1398]), .RECT1_Y(rectangle1_ys[1398]), .RECT1_WIDTH(rectangle1_widths[1398]), .RECT1_HEIGHT(rectangle1_heights[1398]), .RECT1_WEIGHT(rectangle1_weights[1398]), .RECT2_X(rectangle2_xs[1398]), .RECT2_Y(rectangle2_ys[1398]), .RECT2_WIDTH(rectangle2_widths[1398]), .RECT2_HEIGHT(rectangle2_heights[1398]), .RECT2_WEIGHT(rectangle2_weights[1398]), .RECT3_X(rectangle3_xs[1398]), .RECT3_Y(rectangle3_ys[1398]), .RECT3_WIDTH(rectangle3_widths[1398]), .RECT3_HEIGHT(rectangle3_heights[1398]), .RECT3_WEIGHT(rectangle3_weights[1398]), .FEAT_THRES(feature_thresholds[1398]), .FEAT_ABOVE(feature_aboves[1398]), .FEAT_BELOW(feature_belows[1398])) ac1398(.scan_win(scan_win1398), .scan_win_std_dev(scan_win_std_dev[1398]), .feature_accum(feature_accums[1398]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1399]), .RECT1_Y(rectangle1_ys[1399]), .RECT1_WIDTH(rectangle1_widths[1399]), .RECT1_HEIGHT(rectangle1_heights[1399]), .RECT1_WEIGHT(rectangle1_weights[1399]), .RECT2_X(rectangle2_xs[1399]), .RECT2_Y(rectangle2_ys[1399]), .RECT2_WIDTH(rectangle2_widths[1399]), .RECT2_HEIGHT(rectangle2_heights[1399]), .RECT2_WEIGHT(rectangle2_weights[1399]), .RECT3_X(rectangle3_xs[1399]), .RECT3_Y(rectangle3_ys[1399]), .RECT3_WIDTH(rectangle3_widths[1399]), .RECT3_HEIGHT(rectangle3_heights[1399]), .RECT3_WEIGHT(rectangle3_weights[1399]), .FEAT_THRES(feature_thresholds[1399]), .FEAT_ABOVE(feature_aboves[1399]), .FEAT_BELOW(feature_belows[1399])) ac1399(.scan_win(scan_win1399), .scan_win_std_dev(scan_win_std_dev[1399]), .feature_accum(feature_accums[1399]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1400]), .RECT1_Y(rectangle1_ys[1400]), .RECT1_WIDTH(rectangle1_widths[1400]), .RECT1_HEIGHT(rectangle1_heights[1400]), .RECT1_WEIGHT(rectangle1_weights[1400]), .RECT2_X(rectangle2_xs[1400]), .RECT2_Y(rectangle2_ys[1400]), .RECT2_WIDTH(rectangle2_widths[1400]), .RECT2_HEIGHT(rectangle2_heights[1400]), .RECT2_WEIGHT(rectangle2_weights[1400]), .RECT3_X(rectangle3_xs[1400]), .RECT3_Y(rectangle3_ys[1400]), .RECT3_WIDTH(rectangle3_widths[1400]), .RECT3_HEIGHT(rectangle3_heights[1400]), .RECT3_WEIGHT(rectangle3_weights[1400]), .FEAT_THRES(feature_thresholds[1400]), .FEAT_ABOVE(feature_aboves[1400]), .FEAT_BELOW(feature_belows[1400])) ac1400(.scan_win(scan_win1400), .scan_win_std_dev(scan_win_std_dev[1400]), .feature_accum(feature_accums[1400]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1401]), .RECT1_Y(rectangle1_ys[1401]), .RECT1_WIDTH(rectangle1_widths[1401]), .RECT1_HEIGHT(rectangle1_heights[1401]), .RECT1_WEIGHT(rectangle1_weights[1401]), .RECT2_X(rectangle2_xs[1401]), .RECT2_Y(rectangle2_ys[1401]), .RECT2_WIDTH(rectangle2_widths[1401]), .RECT2_HEIGHT(rectangle2_heights[1401]), .RECT2_WEIGHT(rectangle2_weights[1401]), .RECT3_X(rectangle3_xs[1401]), .RECT3_Y(rectangle3_ys[1401]), .RECT3_WIDTH(rectangle3_widths[1401]), .RECT3_HEIGHT(rectangle3_heights[1401]), .RECT3_WEIGHT(rectangle3_weights[1401]), .FEAT_THRES(feature_thresholds[1401]), .FEAT_ABOVE(feature_aboves[1401]), .FEAT_BELOW(feature_belows[1401])) ac1401(.scan_win(scan_win1401), .scan_win_std_dev(scan_win_std_dev[1401]), .feature_accum(feature_accums[1401]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1402]), .RECT1_Y(rectangle1_ys[1402]), .RECT1_WIDTH(rectangle1_widths[1402]), .RECT1_HEIGHT(rectangle1_heights[1402]), .RECT1_WEIGHT(rectangle1_weights[1402]), .RECT2_X(rectangle2_xs[1402]), .RECT2_Y(rectangle2_ys[1402]), .RECT2_WIDTH(rectangle2_widths[1402]), .RECT2_HEIGHT(rectangle2_heights[1402]), .RECT2_WEIGHT(rectangle2_weights[1402]), .RECT3_X(rectangle3_xs[1402]), .RECT3_Y(rectangle3_ys[1402]), .RECT3_WIDTH(rectangle3_widths[1402]), .RECT3_HEIGHT(rectangle3_heights[1402]), .RECT3_WEIGHT(rectangle3_weights[1402]), .FEAT_THRES(feature_thresholds[1402]), .FEAT_ABOVE(feature_aboves[1402]), .FEAT_BELOW(feature_belows[1402])) ac1402(.scan_win(scan_win1402), .scan_win_std_dev(scan_win_std_dev[1402]), .feature_accum(feature_accums[1402]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1403]), .RECT1_Y(rectangle1_ys[1403]), .RECT1_WIDTH(rectangle1_widths[1403]), .RECT1_HEIGHT(rectangle1_heights[1403]), .RECT1_WEIGHT(rectangle1_weights[1403]), .RECT2_X(rectangle2_xs[1403]), .RECT2_Y(rectangle2_ys[1403]), .RECT2_WIDTH(rectangle2_widths[1403]), .RECT2_HEIGHT(rectangle2_heights[1403]), .RECT2_WEIGHT(rectangle2_weights[1403]), .RECT3_X(rectangle3_xs[1403]), .RECT3_Y(rectangle3_ys[1403]), .RECT3_WIDTH(rectangle3_widths[1403]), .RECT3_HEIGHT(rectangle3_heights[1403]), .RECT3_WEIGHT(rectangle3_weights[1403]), .FEAT_THRES(feature_thresholds[1403]), .FEAT_ABOVE(feature_aboves[1403]), .FEAT_BELOW(feature_belows[1403])) ac1403(.scan_win(scan_win1403), .scan_win_std_dev(scan_win_std_dev[1403]), .feature_accum(feature_accums[1403]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1404]), .RECT1_Y(rectangle1_ys[1404]), .RECT1_WIDTH(rectangle1_widths[1404]), .RECT1_HEIGHT(rectangle1_heights[1404]), .RECT1_WEIGHT(rectangle1_weights[1404]), .RECT2_X(rectangle2_xs[1404]), .RECT2_Y(rectangle2_ys[1404]), .RECT2_WIDTH(rectangle2_widths[1404]), .RECT2_HEIGHT(rectangle2_heights[1404]), .RECT2_WEIGHT(rectangle2_weights[1404]), .RECT3_X(rectangle3_xs[1404]), .RECT3_Y(rectangle3_ys[1404]), .RECT3_WIDTH(rectangle3_widths[1404]), .RECT3_HEIGHT(rectangle3_heights[1404]), .RECT3_WEIGHT(rectangle3_weights[1404]), .FEAT_THRES(feature_thresholds[1404]), .FEAT_ABOVE(feature_aboves[1404]), .FEAT_BELOW(feature_belows[1404])) ac1404(.scan_win(scan_win1404), .scan_win_std_dev(scan_win_std_dev[1404]), .feature_accum(feature_accums[1404]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1405]), .RECT1_Y(rectangle1_ys[1405]), .RECT1_WIDTH(rectangle1_widths[1405]), .RECT1_HEIGHT(rectangle1_heights[1405]), .RECT1_WEIGHT(rectangle1_weights[1405]), .RECT2_X(rectangle2_xs[1405]), .RECT2_Y(rectangle2_ys[1405]), .RECT2_WIDTH(rectangle2_widths[1405]), .RECT2_HEIGHT(rectangle2_heights[1405]), .RECT2_WEIGHT(rectangle2_weights[1405]), .RECT3_X(rectangle3_xs[1405]), .RECT3_Y(rectangle3_ys[1405]), .RECT3_WIDTH(rectangle3_widths[1405]), .RECT3_HEIGHT(rectangle3_heights[1405]), .RECT3_WEIGHT(rectangle3_weights[1405]), .FEAT_THRES(feature_thresholds[1405]), .FEAT_ABOVE(feature_aboves[1405]), .FEAT_BELOW(feature_belows[1405])) ac1405(.scan_win(scan_win1405), .scan_win_std_dev(scan_win_std_dev[1405]), .feature_accum(feature_accums[1405]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1406]), .RECT1_Y(rectangle1_ys[1406]), .RECT1_WIDTH(rectangle1_widths[1406]), .RECT1_HEIGHT(rectangle1_heights[1406]), .RECT1_WEIGHT(rectangle1_weights[1406]), .RECT2_X(rectangle2_xs[1406]), .RECT2_Y(rectangle2_ys[1406]), .RECT2_WIDTH(rectangle2_widths[1406]), .RECT2_HEIGHT(rectangle2_heights[1406]), .RECT2_WEIGHT(rectangle2_weights[1406]), .RECT3_X(rectangle3_xs[1406]), .RECT3_Y(rectangle3_ys[1406]), .RECT3_WIDTH(rectangle3_widths[1406]), .RECT3_HEIGHT(rectangle3_heights[1406]), .RECT3_WEIGHT(rectangle3_weights[1406]), .FEAT_THRES(feature_thresholds[1406]), .FEAT_ABOVE(feature_aboves[1406]), .FEAT_BELOW(feature_belows[1406])) ac1406(.scan_win(scan_win1406), .scan_win_std_dev(scan_win_std_dev[1406]), .feature_accum(feature_accums[1406]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1407]), .RECT1_Y(rectangle1_ys[1407]), .RECT1_WIDTH(rectangle1_widths[1407]), .RECT1_HEIGHT(rectangle1_heights[1407]), .RECT1_WEIGHT(rectangle1_weights[1407]), .RECT2_X(rectangle2_xs[1407]), .RECT2_Y(rectangle2_ys[1407]), .RECT2_WIDTH(rectangle2_widths[1407]), .RECT2_HEIGHT(rectangle2_heights[1407]), .RECT2_WEIGHT(rectangle2_weights[1407]), .RECT3_X(rectangle3_xs[1407]), .RECT3_Y(rectangle3_ys[1407]), .RECT3_WIDTH(rectangle3_widths[1407]), .RECT3_HEIGHT(rectangle3_heights[1407]), .RECT3_WEIGHT(rectangle3_weights[1407]), .FEAT_THRES(feature_thresholds[1407]), .FEAT_ABOVE(feature_aboves[1407]), .FEAT_BELOW(feature_belows[1407])) ac1407(.scan_win(scan_win1407), .scan_win_std_dev(scan_win_std_dev[1407]), .feature_accum(feature_accums[1407]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1408]), .RECT1_Y(rectangle1_ys[1408]), .RECT1_WIDTH(rectangle1_widths[1408]), .RECT1_HEIGHT(rectangle1_heights[1408]), .RECT1_WEIGHT(rectangle1_weights[1408]), .RECT2_X(rectangle2_xs[1408]), .RECT2_Y(rectangle2_ys[1408]), .RECT2_WIDTH(rectangle2_widths[1408]), .RECT2_HEIGHT(rectangle2_heights[1408]), .RECT2_WEIGHT(rectangle2_weights[1408]), .RECT3_X(rectangle3_xs[1408]), .RECT3_Y(rectangle3_ys[1408]), .RECT3_WIDTH(rectangle3_widths[1408]), .RECT3_HEIGHT(rectangle3_heights[1408]), .RECT3_WEIGHT(rectangle3_weights[1408]), .FEAT_THRES(feature_thresholds[1408]), .FEAT_ABOVE(feature_aboves[1408]), .FEAT_BELOW(feature_belows[1408])) ac1408(.scan_win(scan_win1408), .scan_win_std_dev(scan_win_std_dev[1408]), .feature_accum(feature_accums[1408]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1409]), .RECT1_Y(rectangle1_ys[1409]), .RECT1_WIDTH(rectangle1_widths[1409]), .RECT1_HEIGHT(rectangle1_heights[1409]), .RECT1_WEIGHT(rectangle1_weights[1409]), .RECT2_X(rectangle2_xs[1409]), .RECT2_Y(rectangle2_ys[1409]), .RECT2_WIDTH(rectangle2_widths[1409]), .RECT2_HEIGHT(rectangle2_heights[1409]), .RECT2_WEIGHT(rectangle2_weights[1409]), .RECT3_X(rectangle3_xs[1409]), .RECT3_Y(rectangle3_ys[1409]), .RECT3_WIDTH(rectangle3_widths[1409]), .RECT3_HEIGHT(rectangle3_heights[1409]), .RECT3_WEIGHT(rectangle3_weights[1409]), .FEAT_THRES(feature_thresholds[1409]), .FEAT_ABOVE(feature_aboves[1409]), .FEAT_BELOW(feature_belows[1409])) ac1409(.scan_win(scan_win1409), .scan_win_std_dev(scan_win_std_dev[1409]), .feature_accum(feature_accums[1409]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1410]), .RECT1_Y(rectangle1_ys[1410]), .RECT1_WIDTH(rectangle1_widths[1410]), .RECT1_HEIGHT(rectangle1_heights[1410]), .RECT1_WEIGHT(rectangle1_weights[1410]), .RECT2_X(rectangle2_xs[1410]), .RECT2_Y(rectangle2_ys[1410]), .RECT2_WIDTH(rectangle2_widths[1410]), .RECT2_HEIGHT(rectangle2_heights[1410]), .RECT2_WEIGHT(rectangle2_weights[1410]), .RECT3_X(rectangle3_xs[1410]), .RECT3_Y(rectangle3_ys[1410]), .RECT3_WIDTH(rectangle3_widths[1410]), .RECT3_HEIGHT(rectangle3_heights[1410]), .RECT3_WEIGHT(rectangle3_weights[1410]), .FEAT_THRES(feature_thresholds[1410]), .FEAT_ABOVE(feature_aboves[1410]), .FEAT_BELOW(feature_belows[1410])) ac1410(.scan_win(scan_win1410), .scan_win_std_dev(scan_win_std_dev[1410]), .feature_accum(feature_accums[1410]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1411]), .RECT1_Y(rectangle1_ys[1411]), .RECT1_WIDTH(rectangle1_widths[1411]), .RECT1_HEIGHT(rectangle1_heights[1411]), .RECT1_WEIGHT(rectangle1_weights[1411]), .RECT2_X(rectangle2_xs[1411]), .RECT2_Y(rectangle2_ys[1411]), .RECT2_WIDTH(rectangle2_widths[1411]), .RECT2_HEIGHT(rectangle2_heights[1411]), .RECT2_WEIGHT(rectangle2_weights[1411]), .RECT3_X(rectangle3_xs[1411]), .RECT3_Y(rectangle3_ys[1411]), .RECT3_WIDTH(rectangle3_widths[1411]), .RECT3_HEIGHT(rectangle3_heights[1411]), .RECT3_WEIGHT(rectangle3_weights[1411]), .FEAT_THRES(feature_thresholds[1411]), .FEAT_ABOVE(feature_aboves[1411]), .FEAT_BELOW(feature_belows[1411])) ac1411(.scan_win(scan_win1411), .scan_win_std_dev(scan_win_std_dev[1411]), .feature_accum(feature_accums[1411]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1412]), .RECT1_Y(rectangle1_ys[1412]), .RECT1_WIDTH(rectangle1_widths[1412]), .RECT1_HEIGHT(rectangle1_heights[1412]), .RECT1_WEIGHT(rectangle1_weights[1412]), .RECT2_X(rectangle2_xs[1412]), .RECT2_Y(rectangle2_ys[1412]), .RECT2_WIDTH(rectangle2_widths[1412]), .RECT2_HEIGHT(rectangle2_heights[1412]), .RECT2_WEIGHT(rectangle2_weights[1412]), .RECT3_X(rectangle3_xs[1412]), .RECT3_Y(rectangle3_ys[1412]), .RECT3_WIDTH(rectangle3_widths[1412]), .RECT3_HEIGHT(rectangle3_heights[1412]), .RECT3_WEIGHT(rectangle3_weights[1412]), .FEAT_THRES(feature_thresholds[1412]), .FEAT_ABOVE(feature_aboves[1412]), .FEAT_BELOW(feature_belows[1412])) ac1412(.scan_win(scan_win1412), .scan_win_std_dev(scan_win_std_dev[1412]), .feature_accum(feature_accums[1412]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1413]), .RECT1_Y(rectangle1_ys[1413]), .RECT1_WIDTH(rectangle1_widths[1413]), .RECT1_HEIGHT(rectangle1_heights[1413]), .RECT1_WEIGHT(rectangle1_weights[1413]), .RECT2_X(rectangle2_xs[1413]), .RECT2_Y(rectangle2_ys[1413]), .RECT2_WIDTH(rectangle2_widths[1413]), .RECT2_HEIGHT(rectangle2_heights[1413]), .RECT2_WEIGHT(rectangle2_weights[1413]), .RECT3_X(rectangle3_xs[1413]), .RECT3_Y(rectangle3_ys[1413]), .RECT3_WIDTH(rectangle3_widths[1413]), .RECT3_HEIGHT(rectangle3_heights[1413]), .RECT3_WEIGHT(rectangle3_weights[1413]), .FEAT_THRES(feature_thresholds[1413]), .FEAT_ABOVE(feature_aboves[1413]), .FEAT_BELOW(feature_belows[1413])) ac1413(.scan_win(scan_win1413), .scan_win_std_dev(scan_win_std_dev[1413]), .feature_accum(feature_accums[1413]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1414]), .RECT1_Y(rectangle1_ys[1414]), .RECT1_WIDTH(rectangle1_widths[1414]), .RECT1_HEIGHT(rectangle1_heights[1414]), .RECT1_WEIGHT(rectangle1_weights[1414]), .RECT2_X(rectangle2_xs[1414]), .RECT2_Y(rectangle2_ys[1414]), .RECT2_WIDTH(rectangle2_widths[1414]), .RECT2_HEIGHT(rectangle2_heights[1414]), .RECT2_WEIGHT(rectangle2_weights[1414]), .RECT3_X(rectangle3_xs[1414]), .RECT3_Y(rectangle3_ys[1414]), .RECT3_WIDTH(rectangle3_widths[1414]), .RECT3_HEIGHT(rectangle3_heights[1414]), .RECT3_WEIGHT(rectangle3_weights[1414]), .FEAT_THRES(feature_thresholds[1414]), .FEAT_ABOVE(feature_aboves[1414]), .FEAT_BELOW(feature_belows[1414])) ac1414(.scan_win(scan_win1414), .scan_win_std_dev(scan_win_std_dev[1414]), .feature_accum(feature_accums[1414]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1415]), .RECT1_Y(rectangle1_ys[1415]), .RECT1_WIDTH(rectangle1_widths[1415]), .RECT1_HEIGHT(rectangle1_heights[1415]), .RECT1_WEIGHT(rectangle1_weights[1415]), .RECT2_X(rectangle2_xs[1415]), .RECT2_Y(rectangle2_ys[1415]), .RECT2_WIDTH(rectangle2_widths[1415]), .RECT2_HEIGHT(rectangle2_heights[1415]), .RECT2_WEIGHT(rectangle2_weights[1415]), .RECT3_X(rectangle3_xs[1415]), .RECT3_Y(rectangle3_ys[1415]), .RECT3_WIDTH(rectangle3_widths[1415]), .RECT3_HEIGHT(rectangle3_heights[1415]), .RECT3_WEIGHT(rectangle3_weights[1415]), .FEAT_THRES(feature_thresholds[1415]), .FEAT_ABOVE(feature_aboves[1415]), .FEAT_BELOW(feature_belows[1415])) ac1415(.scan_win(scan_win1415), .scan_win_std_dev(scan_win_std_dev[1415]), .feature_accum(feature_accums[1415]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1416]), .RECT1_Y(rectangle1_ys[1416]), .RECT1_WIDTH(rectangle1_widths[1416]), .RECT1_HEIGHT(rectangle1_heights[1416]), .RECT1_WEIGHT(rectangle1_weights[1416]), .RECT2_X(rectangle2_xs[1416]), .RECT2_Y(rectangle2_ys[1416]), .RECT2_WIDTH(rectangle2_widths[1416]), .RECT2_HEIGHT(rectangle2_heights[1416]), .RECT2_WEIGHT(rectangle2_weights[1416]), .RECT3_X(rectangle3_xs[1416]), .RECT3_Y(rectangle3_ys[1416]), .RECT3_WIDTH(rectangle3_widths[1416]), .RECT3_HEIGHT(rectangle3_heights[1416]), .RECT3_WEIGHT(rectangle3_weights[1416]), .FEAT_THRES(feature_thresholds[1416]), .FEAT_ABOVE(feature_aboves[1416]), .FEAT_BELOW(feature_belows[1416])) ac1416(.scan_win(scan_win1416), .scan_win_std_dev(scan_win_std_dev[1416]), .feature_accum(feature_accums[1416]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1417]), .RECT1_Y(rectangle1_ys[1417]), .RECT1_WIDTH(rectangle1_widths[1417]), .RECT1_HEIGHT(rectangle1_heights[1417]), .RECT1_WEIGHT(rectangle1_weights[1417]), .RECT2_X(rectangle2_xs[1417]), .RECT2_Y(rectangle2_ys[1417]), .RECT2_WIDTH(rectangle2_widths[1417]), .RECT2_HEIGHT(rectangle2_heights[1417]), .RECT2_WEIGHT(rectangle2_weights[1417]), .RECT3_X(rectangle3_xs[1417]), .RECT3_Y(rectangle3_ys[1417]), .RECT3_WIDTH(rectangle3_widths[1417]), .RECT3_HEIGHT(rectangle3_heights[1417]), .RECT3_WEIGHT(rectangle3_weights[1417]), .FEAT_THRES(feature_thresholds[1417]), .FEAT_ABOVE(feature_aboves[1417]), .FEAT_BELOW(feature_belows[1417])) ac1417(.scan_win(scan_win1417), .scan_win_std_dev(scan_win_std_dev[1417]), .feature_accum(feature_accums[1417]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1418]), .RECT1_Y(rectangle1_ys[1418]), .RECT1_WIDTH(rectangle1_widths[1418]), .RECT1_HEIGHT(rectangle1_heights[1418]), .RECT1_WEIGHT(rectangle1_weights[1418]), .RECT2_X(rectangle2_xs[1418]), .RECT2_Y(rectangle2_ys[1418]), .RECT2_WIDTH(rectangle2_widths[1418]), .RECT2_HEIGHT(rectangle2_heights[1418]), .RECT2_WEIGHT(rectangle2_weights[1418]), .RECT3_X(rectangle3_xs[1418]), .RECT3_Y(rectangle3_ys[1418]), .RECT3_WIDTH(rectangle3_widths[1418]), .RECT3_HEIGHT(rectangle3_heights[1418]), .RECT3_WEIGHT(rectangle3_weights[1418]), .FEAT_THRES(feature_thresholds[1418]), .FEAT_ABOVE(feature_aboves[1418]), .FEAT_BELOW(feature_belows[1418])) ac1418(.scan_win(scan_win1418), .scan_win_std_dev(scan_win_std_dev[1418]), .feature_accum(feature_accums[1418]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1419]), .RECT1_Y(rectangle1_ys[1419]), .RECT1_WIDTH(rectangle1_widths[1419]), .RECT1_HEIGHT(rectangle1_heights[1419]), .RECT1_WEIGHT(rectangle1_weights[1419]), .RECT2_X(rectangle2_xs[1419]), .RECT2_Y(rectangle2_ys[1419]), .RECT2_WIDTH(rectangle2_widths[1419]), .RECT2_HEIGHT(rectangle2_heights[1419]), .RECT2_WEIGHT(rectangle2_weights[1419]), .RECT3_X(rectangle3_xs[1419]), .RECT3_Y(rectangle3_ys[1419]), .RECT3_WIDTH(rectangle3_widths[1419]), .RECT3_HEIGHT(rectangle3_heights[1419]), .RECT3_WEIGHT(rectangle3_weights[1419]), .FEAT_THRES(feature_thresholds[1419]), .FEAT_ABOVE(feature_aboves[1419]), .FEAT_BELOW(feature_belows[1419])) ac1419(.scan_win(scan_win1419), .scan_win_std_dev(scan_win_std_dev[1419]), .feature_accum(feature_accums[1419]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1420]), .RECT1_Y(rectangle1_ys[1420]), .RECT1_WIDTH(rectangle1_widths[1420]), .RECT1_HEIGHT(rectangle1_heights[1420]), .RECT1_WEIGHT(rectangle1_weights[1420]), .RECT2_X(rectangle2_xs[1420]), .RECT2_Y(rectangle2_ys[1420]), .RECT2_WIDTH(rectangle2_widths[1420]), .RECT2_HEIGHT(rectangle2_heights[1420]), .RECT2_WEIGHT(rectangle2_weights[1420]), .RECT3_X(rectangle3_xs[1420]), .RECT3_Y(rectangle3_ys[1420]), .RECT3_WIDTH(rectangle3_widths[1420]), .RECT3_HEIGHT(rectangle3_heights[1420]), .RECT3_WEIGHT(rectangle3_weights[1420]), .FEAT_THRES(feature_thresholds[1420]), .FEAT_ABOVE(feature_aboves[1420]), .FEAT_BELOW(feature_belows[1420])) ac1420(.scan_win(scan_win1420), .scan_win_std_dev(scan_win_std_dev[1420]), .feature_accum(feature_accums[1420]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1421]), .RECT1_Y(rectangle1_ys[1421]), .RECT1_WIDTH(rectangle1_widths[1421]), .RECT1_HEIGHT(rectangle1_heights[1421]), .RECT1_WEIGHT(rectangle1_weights[1421]), .RECT2_X(rectangle2_xs[1421]), .RECT2_Y(rectangle2_ys[1421]), .RECT2_WIDTH(rectangle2_widths[1421]), .RECT2_HEIGHT(rectangle2_heights[1421]), .RECT2_WEIGHT(rectangle2_weights[1421]), .RECT3_X(rectangle3_xs[1421]), .RECT3_Y(rectangle3_ys[1421]), .RECT3_WIDTH(rectangle3_widths[1421]), .RECT3_HEIGHT(rectangle3_heights[1421]), .RECT3_WEIGHT(rectangle3_weights[1421]), .FEAT_THRES(feature_thresholds[1421]), .FEAT_ABOVE(feature_aboves[1421]), .FEAT_BELOW(feature_belows[1421])) ac1421(.scan_win(scan_win1421), .scan_win_std_dev(scan_win_std_dev[1421]), .feature_accum(feature_accums[1421]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1422]), .RECT1_Y(rectangle1_ys[1422]), .RECT1_WIDTH(rectangle1_widths[1422]), .RECT1_HEIGHT(rectangle1_heights[1422]), .RECT1_WEIGHT(rectangle1_weights[1422]), .RECT2_X(rectangle2_xs[1422]), .RECT2_Y(rectangle2_ys[1422]), .RECT2_WIDTH(rectangle2_widths[1422]), .RECT2_HEIGHT(rectangle2_heights[1422]), .RECT2_WEIGHT(rectangle2_weights[1422]), .RECT3_X(rectangle3_xs[1422]), .RECT3_Y(rectangle3_ys[1422]), .RECT3_WIDTH(rectangle3_widths[1422]), .RECT3_HEIGHT(rectangle3_heights[1422]), .RECT3_WEIGHT(rectangle3_weights[1422]), .FEAT_THRES(feature_thresholds[1422]), .FEAT_ABOVE(feature_aboves[1422]), .FEAT_BELOW(feature_belows[1422])) ac1422(.scan_win(scan_win1422), .scan_win_std_dev(scan_win_std_dev[1422]), .feature_accum(feature_accums[1422]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1423]), .RECT1_Y(rectangle1_ys[1423]), .RECT1_WIDTH(rectangle1_widths[1423]), .RECT1_HEIGHT(rectangle1_heights[1423]), .RECT1_WEIGHT(rectangle1_weights[1423]), .RECT2_X(rectangle2_xs[1423]), .RECT2_Y(rectangle2_ys[1423]), .RECT2_WIDTH(rectangle2_widths[1423]), .RECT2_HEIGHT(rectangle2_heights[1423]), .RECT2_WEIGHT(rectangle2_weights[1423]), .RECT3_X(rectangle3_xs[1423]), .RECT3_Y(rectangle3_ys[1423]), .RECT3_WIDTH(rectangle3_widths[1423]), .RECT3_HEIGHT(rectangle3_heights[1423]), .RECT3_WEIGHT(rectangle3_weights[1423]), .FEAT_THRES(feature_thresholds[1423]), .FEAT_ABOVE(feature_aboves[1423]), .FEAT_BELOW(feature_belows[1423])) ac1423(.scan_win(scan_win1423), .scan_win_std_dev(scan_win_std_dev[1423]), .feature_accum(feature_accums[1423]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1424]), .RECT1_Y(rectangle1_ys[1424]), .RECT1_WIDTH(rectangle1_widths[1424]), .RECT1_HEIGHT(rectangle1_heights[1424]), .RECT1_WEIGHT(rectangle1_weights[1424]), .RECT2_X(rectangle2_xs[1424]), .RECT2_Y(rectangle2_ys[1424]), .RECT2_WIDTH(rectangle2_widths[1424]), .RECT2_HEIGHT(rectangle2_heights[1424]), .RECT2_WEIGHT(rectangle2_weights[1424]), .RECT3_X(rectangle3_xs[1424]), .RECT3_Y(rectangle3_ys[1424]), .RECT3_WIDTH(rectangle3_widths[1424]), .RECT3_HEIGHT(rectangle3_heights[1424]), .RECT3_WEIGHT(rectangle3_weights[1424]), .FEAT_THRES(feature_thresholds[1424]), .FEAT_ABOVE(feature_aboves[1424]), .FEAT_BELOW(feature_belows[1424])) ac1424(.scan_win(scan_win1424), .scan_win_std_dev(scan_win_std_dev[1424]), .feature_accum(feature_accums[1424]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1425]), .RECT1_Y(rectangle1_ys[1425]), .RECT1_WIDTH(rectangle1_widths[1425]), .RECT1_HEIGHT(rectangle1_heights[1425]), .RECT1_WEIGHT(rectangle1_weights[1425]), .RECT2_X(rectangle2_xs[1425]), .RECT2_Y(rectangle2_ys[1425]), .RECT2_WIDTH(rectangle2_widths[1425]), .RECT2_HEIGHT(rectangle2_heights[1425]), .RECT2_WEIGHT(rectangle2_weights[1425]), .RECT3_X(rectangle3_xs[1425]), .RECT3_Y(rectangle3_ys[1425]), .RECT3_WIDTH(rectangle3_widths[1425]), .RECT3_HEIGHT(rectangle3_heights[1425]), .RECT3_WEIGHT(rectangle3_weights[1425]), .FEAT_THRES(feature_thresholds[1425]), .FEAT_ABOVE(feature_aboves[1425]), .FEAT_BELOW(feature_belows[1425])) ac1425(.scan_win(scan_win1425), .scan_win_std_dev(scan_win_std_dev[1425]), .feature_accum(feature_accums[1425]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1426]), .RECT1_Y(rectangle1_ys[1426]), .RECT1_WIDTH(rectangle1_widths[1426]), .RECT1_HEIGHT(rectangle1_heights[1426]), .RECT1_WEIGHT(rectangle1_weights[1426]), .RECT2_X(rectangle2_xs[1426]), .RECT2_Y(rectangle2_ys[1426]), .RECT2_WIDTH(rectangle2_widths[1426]), .RECT2_HEIGHT(rectangle2_heights[1426]), .RECT2_WEIGHT(rectangle2_weights[1426]), .RECT3_X(rectangle3_xs[1426]), .RECT3_Y(rectangle3_ys[1426]), .RECT3_WIDTH(rectangle3_widths[1426]), .RECT3_HEIGHT(rectangle3_heights[1426]), .RECT3_WEIGHT(rectangle3_weights[1426]), .FEAT_THRES(feature_thresholds[1426]), .FEAT_ABOVE(feature_aboves[1426]), .FEAT_BELOW(feature_belows[1426])) ac1426(.scan_win(scan_win1426), .scan_win_std_dev(scan_win_std_dev[1426]), .feature_accum(feature_accums[1426]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1427]), .RECT1_Y(rectangle1_ys[1427]), .RECT1_WIDTH(rectangle1_widths[1427]), .RECT1_HEIGHT(rectangle1_heights[1427]), .RECT1_WEIGHT(rectangle1_weights[1427]), .RECT2_X(rectangle2_xs[1427]), .RECT2_Y(rectangle2_ys[1427]), .RECT2_WIDTH(rectangle2_widths[1427]), .RECT2_HEIGHT(rectangle2_heights[1427]), .RECT2_WEIGHT(rectangle2_weights[1427]), .RECT3_X(rectangle3_xs[1427]), .RECT3_Y(rectangle3_ys[1427]), .RECT3_WIDTH(rectangle3_widths[1427]), .RECT3_HEIGHT(rectangle3_heights[1427]), .RECT3_WEIGHT(rectangle3_weights[1427]), .FEAT_THRES(feature_thresholds[1427]), .FEAT_ABOVE(feature_aboves[1427]), .FEAT_BELOW(feature_belows[1427])) ac1427(.scan_win(scan_win1427), .scan_win_std_dev(scan_win_std_dev[1427]), .feature_accum(feature_accums[1427]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1428]), .RECT1_Y(rectangle1_ys[1428]), .RECT1_WIDTH(rectangle1_widths[1428]), .RECT1_HEIGHT(rectangle1_heights[1428]), .RECT1_WEIGHT(rectangle1_weights[1428]), .RECT2_X(rectangle2_xs[1428]), .RECT2_Y(rectangle2_ys[1428]), .RECT2_WIDTH(rectangle2_widths[1428]), .RECT2_HEIGHT(rectangle2_heights[1428]), .RECT2_WEIGHT(rectangle2_weights[1428]), .RECT3_X(rectangle3_xs[1428]), .RECT3_Y(rectangle3_ys[1428]), .RECT3_WIDTH(rectangle3_widths[1428]), .RECT3_HEIGHT(rectangle3_heights[1428]), .RECT3_WEIGHT(rectangle3_weights[1428]), .FEAT_THRES(feature_thresholds[1428]), .FEAT_ABOVE(feature_aboves[1428]), .FEAT_BELOW(feature_belows[1428])) ac1428(.scan_win(scan_win1428), .scan_win_std_dev(scan_win_std_dev[1428]), .feature_accum(feature_accums[1428]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1429]), .RECT1_Y(rectangle1_ys[1429]), .RECT1_WIDTH(rectangle1_widths[1429]), .RECT1_HEIGHT(rectangle1_heights[1429]), .RECT1_WEIGHT(rectangle1_weights[1429]), .RECT2_X(rectangle2_xs[1429]), .RECT2_Y(rectangle2_ys[1429]), .RECT2_WIDTH(rectangle2_widths[1429]), .RECT2_HEIGHT(rectangle2_heights[1429]), .RECT2_WEIGHT(rectangle2_weights[1429]), .RECT3_X(rectangle3_xs[1429]), .RECT3_Y(rectangle3_ys[1429]), .RECT3_WIDTH(rectangle3_widths[1429]), .RECT3_HEIGHT(rectangle3_heights[1429]), .RECT3_WEIGHT(rectangle3_weights[1429]), .FEAT_THRES(feature_thresholds[1429]), .FEAT_ABOVE(feature_aboves[1429]), .FEAT_BELOW(feature_belows[1429])) ac1429(.scan_win(scan_win1429), .scan_win_std_dev(scan_win_std_dev[1429]), .feature_accum(feature_accums[1429]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1430]), .RECT1_Y(rectangle1_ys[1430]), .RECT1_WIDTH(rectangle1_widths[1430]), .RECT1_HEIGHT(rectangle1_heights[1430]), .RECT1_WEIGHT(rectangle1_weights[1430]), .RECT2_X(rectangle2_xs[1430]), .RECT2_Y(rectangle2_ys[1430]), .RECT2_WIDTH(rectangle2_widths[1430]), .RECT2_HEIGHT(rectangle2_heights[1430]), .RECT2_WEIGHT(rectangle2_weights[1430]), .RECT3_X(rectangle3_xs[1430]), .RECT3_Y(rectangle3_ys[1430]), .RECT3_WIDTH(rectangle3_widths[1430]), .RECT3_HEIGHT(rectangle3_heights[1430]), .RECT3_WEIGHT(rectangle3_weights[1430]), .FEAT_THRES(feature_thresholds[1430]), .FEAT_ABOVE(feature_aboves[1430]), .FEAT_BELOW(feature_belows[1430])) ac1430(.scan_win(scan_win1430), .scan_win_std_dev(scan_win_std_dev[1430]), .feature_accum(feature_accums[1430]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1431]), .RECT1_Y(rectangle1_ys[1431]), .RECT1_WIDTH(rectangle1_widths[1431]), .RECT1_HEIGHT(rectangle1_heights[1431]), .RECT1_WEIGHT(rectangle1_weights[1431]), .RECT2_X(rectangle2_xs[1431]), .RECT2_Y(rectangle2_ys[1431]), .RECT2_WIDTH(rectangle2_widths[1431]), .RECT2_HEIGHT(rectangle2_heights[1431]), .RECT2_WEIGHT(rectangle2_weights[1431]), .RECT3_X(rectangle3_xs[1431]), .RECT3_Y(rectangle3_ys[1431]), .RECT3_WIDTH(rectangle3_widths[1431]), .RECT3_HEIGHT(rectangle3_heights[1431]), .RECT3_WEIGHT(rectangle3_weights[1431]), .FEAT_THRES(feature_thresholds[1431]), .FEAT_ABOVE(feature_aboves[1431]), .FEAT_BELOW(feature_belows[1431])) ac1431(.scan_win(scan_win1431), .scan_win_std_dev(scan_win_std_dev[1431]), .feature_accum(feature_accums[1431]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1432]), .RECT1_Y(rectangle1_ys[1432]), .RECT1_WIDTH(rectangle1_widths[1432]), .RECT1_HEIGHT(rectangle1_heights[1432]), .RECT1_WEIGHT(rectangle1_weights[1432]), .RECT2_X(rectangle2_xs[1432]), .RECT2_Y(rectangle2_ys[1432]), .RECT2_WIDTH(rectangle2_widths[1432]), .RECT2_HEIGHT(rectangle2_heights[1432]), .RECT2_WEIGHT(rectangle2_weights[1432]), .RECT3_X(rectangle3_xs[1432]), .RECT3_Y(rectangle3_ys[1432]), .RECT3_WIDTH(rectangle3_widths[1432]), .RECT3_HEIGHT(rectangle3_heights[1432]), .RECT3_WEIGHT(rectangle3_weights[1432]), .FEAT_THRES(feature_thresholds[1432]), .FEAT_ABOVE(feature_aboves[1432]), .FEAT_BELOW(feature_belows[1432])) ac1432(.scan_win(scan_win1432), .scan_win_std_dev(scan_win_std_dev[1432]), .feature_accum(feature_accums[1432]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1433]), .RECT1_Y(rectangle1_ys[1433]), .RECT1_WIDTH(rectangle1_widths[1433]), .RECT1_HEIGHT(rectangle1_heights[1433]), .RECT1_WEIGHT(rectangle1_weights[1433]), .RECT2_X(rectangle2_xs[1433]), .RECT2_Y(rectangle2_ys[1433]), .RECT2_WIDTH(rectangle2_widths[1433]), .RECT2_HEIGHT(rectangle2_heights[1433]), .RECT2_WEIGHT(rectangle2_weights[1433]), .RECT3_X(rectangle3_xs[1433]), .RECT3_Y(rectangle3_ys[1433]), .RECT3_WIDTH(rectangle3_widths[1433]), .RECT3_HEIGHT(rectangle3_heights[1433]), .RECT3_WEIGHT(rectangle3_weights[1433]), .FEAT_THRES(feature_thresholds[1433]), .FEAT_ABOVE(feature_aboves[1433]), .FEAT_BELOW(feature_belows[1433])) ac1433(.scan_win(scan_win1433), .scan_win_std_dev(scan_win_std_dev[1433]), .feature_accum(feature_accums[1433]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1434]), .RECT1_Y(rectangle1_ys[1434]), .RECT1_WIDTH(rectangle1_widths[1434]), .RECT1_HEIGHT(rectangle1_heights[1434]), .RECT1_WEIGHT(rectangle1_weights[1434]), .RECT2_X(rectangle2_xs[1434]), .RECT2_Y(rectangle2_ys[1434]), .RECT2_WIDTH(rectangle2_widths[1434]), .RECT2_HEIGHT(rectangle2_heights[1434]), .RECT2_WEIGHT(rectangle2_weights[1434]), .RECT3_X(rectangle3_xs[1434]), .RECT3_Y(rectangle3_ys[1434]), .RECT3_WIDTH(rectangle3_widths[1434]), .RECT3_HEIGHT(rectangle3_heights[1434]), .RECT3_WEIGHT(rectangle3_weights[1434]), .FEAT_THRES(feature_thresholds[1434]), .FEAT_ABOVE(feature_aboves[1434]), .FEAT_BELOW(feature_belows[1434])) ac1434(.scan_win(scan_win1434), .scan_win_std_dev(scan_win_std_dev[1434]), .feature_accum(feature_accums[1434]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1435]), .RECT1_Y(rectangle1_ys[1435]), .RECT1_WIDTH(rectangle1_widths[1435]), .RECT1_HEIGHT(rectangle1_heights[1435]), .RECT1_WEIGHT(rectangle1_weights[1435]), .RECT2_X(rectangle2_xs[1435]), .RECT2_Y(rectangle2_ys[1435]), .RECT2_WIDTH(rectangle2_widths[1435]), .RECT2_HEIGHT(rectangle2_heights[1435]), .RECT2_WEIGHT(rectangle2_weights[1435]), .RECT3_X(rectangle3_xs[1435]), .RECT3_Y(rectangle3_ys[1435]), .RECT3_WIDTH(rectangle3_widths[1435]), .RECT3_HEIGHT(rectangle3_heights[1435]), .RECT3_WEIGHT(rectangle3_weights[1435]), .FEAT_THRES(feature_thresholds[1435]), .FEAT_ABOVE(feature_aboves[1435]), .FEAT_BELOW(feature_belows[1435])) ac1435(.scan_win(scan_win1435), .scan_win_std_dev(scan_win_std_dev[1435]), .feature_accum(feature_accums[1435]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1436]), .RECT1_Y(rectangle1_ys[1436]), .RECT1_WIDTH(rectangle1_widths[1436]), .RECT1_HEIGHT(rectangle1_heights[1436]), .RECT1_WEIGHT(rectangle1_weights[1436]), .RECT2_X(rectangle2_xs[1436]), .RECT2_Y(rectangle2_ys[1436]), .RECT2_WIDTH(rectangle2_widths[1436]), .RECT2_HEIGHT(rectangle2_heights[1436]), .RECT2_WEIGHT(rectangle2_weights[1436]), .RECT3_X(rectangle3_xs[1436]), .RECT3_Y(rectangle3_ys[1436]), .RECT3_WIDTH(rectangle3_widths[1436]), .RECT3_HEIGHT(rectangle3_heights[1436]), .RECT3_WEIGHT(rectangle3_weights[1436]), .FEAT_THRES(feature_thresholds[1436]), .FEAT_ABOVE(feature_aboves[1436]), .FEAT_BELOW(feature_belows[1436])) ac1436(.scan_win(scan_win1436), .scan_win_std_dev(scan_win_std_dev[1436]), .feature_accum(feature_accums[1436]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1437]), .RECT1_Y(rectangle1_ys[1437]), .RECT1_WIDTH(rectangle1_widths[1437]), .RECT1_HEIGHT(rectangle1_heights[1437]), .RECT1_WEIGHT(rectangle1_weights[1437]), .RECT2_X(rectangle2_xs[1437]), .RECT2_Y(rectangle2_ys[1437]), .RECT2_WIDTH(rectangle2_widths[1437]), .RECT2_HEIGHT(rectangle2_heights[1437]), .RECT2_WEIGHT(rectangle2_weights[1437]), .RECT3_X(rectangle3_xs[1437]), .RECT3_Y(rectangle3_ys[1437]), .RECT3_WIDTH(rectangle3_widths[1437]), .RECT3_HEIGHT(rectangle3_heights[1437]), .RECT3_WEIGHT(rectangle3_weights[1437]), .FEAT_THRES(feature_thresholds[1437]), .FEAT_ABOVE(feature_aboves[1437]), .FEAT_BELOW(feature_belows[1437])) ac1437(.scan_win(scan_win1437), .scan_win_std_dev(scan_win_std_dev[1437]), .feature_accum(feature_accums[1437]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1438]), .RECT1_Y(rectangle1_ys[1438]), .RECT1_WIDTH(rectangle1_widths[1438]), .RECT1_HEIGHT(rectangle1_heights[1438]), .RECT1_WEIGHT(rectangle1_weights[1438]), .RECT2_X(rectangle2_xs[1438]), .RECT2_Y(rectangle2_ys[1438]), .RECT2_WIDTH(rectangle2_widths[1438]), .RECT2_HEIGHT(rectangle2_heights[1438]), .RECT2_WEIGHT(rectangle2_weights[1438]), .RECT3_X(rectangle3_xs[1438]), .RECT3_Y(rectangle3_ys[1438]), .RECT3_WIDTH(rectangle3_widths[1438]), .RECT3_HEIGHT(rectangle3_heights[1438]), .RECT3_WEIGHT(rectangle3_weights[1438]), .FEAT_THRES(feature_thresholds[1438]), .FEAT_ABOVE(feature_aboves[1438]), .FEAT_BELOW(feature_belows[1438])) ac1438(.scan_win(scan_win1438), .scan_win_std_dev(scan_win_std_dev[1438]), .feature_accum(feature_accums[1438]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1439]), .RECT1_Y(rectangle1_ys[1439]), .RECT1_WIDTH(rectangle1_widths[1439]), .RECT1_HEIGHT(rectangle1_heights[1439]), .RECT1_WEIGHT(rectangle1_weights[1439]), .RECT2_X(rectangle2_xs[1439]), .RECT2_Y(rectangle2_ys[1439]), .RECT2_WIDTH(rectangle2_widths[1439]), .RECT2_HEIGHT(rectangle2_heights[1439]), .RECT2_WEIGHT(rectangle2_weights[1439]), .RECT3_X(rectangle3_xs[1439]), .RECT3_Y(rectangle3_ys[1439]), .RECT3_WIDTH(rectangle3_widths[1439]), .RECT3_HEIGHT(rectangle3_heights[1439]), .RECT3_WEIGHT(rectangle3_weights[1439]), .FEAT_THRES(feature_thresholds[1439]), .FEAT_ABOVE(feature_aboves[1439]), .FEAT_BELOW(feature_belows[1439])) ac1439(.scan_win(scan_win1439), .scan_win_std_dev(scan_win_std_dev[1439]), .feature_accum(feature_accums[1439]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1440]), .RECT1_Y(rectangle1_ys[1440]), .RECT1_WIDTH(rectangle1_widths[1440]), .RECT1_HEIGHT(rectangle1_heights[1440]), .RECT1_WEIGHT(rectangle1_weights[1440]), .RECT2_X(rectangle2_xs[1440]), .RECT2_Y(rectangle2_ys[1440]), .RECT2_WIDTH(rectangle2_widths[1440]), .RECT2_HEIGHT(rectangle2_heights[1440]), .RECT2_WEIGHT(rectangle2_weights[1440]), .RECT3_X(rectangle3_xs[1440]), .RECT3_Y(rectangle3_ys[1440]), .RECT3_WIDTH(rectangle3_widths[1440]), .RECT3_HEIGHT(rectangle3_heights[1440]), .RECT3_WEIGHT(rectangle3_weights[1440]), .FEAT_THRES(feature_thresholds[1440]), .FEAT_ABOVE(feature_aboves[1440]), .FEAT_BELOW(feature_belows[1440])) ac1440(.scan_win(scan_win1440), .scan_win_std_dev(scan_win_std_dev[1440]), .feature_accum(feature_accums[1440]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1441]), .RECT1_Y(rectangle1_ys[1441]), .RECT1_WIDTH(rectangle1_widths[1441]), .RECT1_HEIGHT(rectangle1_heights[1441]), .RECT1_WEIGHT(rectangle1_weights[1441]), .RECT2_X(rectangle2_xs[1441]), .RECT2_Y(rectangle2_ys[1441]), .RECT2_WIDTH(rectangle2_widths[1441]), .RECT2_HEIGHT(rectangle2_heights[1441]), .RECT2_WEIGHT(rectangle2_weights[1441]), .RECT3_X(rectangle3_xs[1441]), .RECT3_Y(rectangle3_ys[1441]), .RECT3_WIDTH(rectangle3_widths[1441]), .RECT3_HEIGHT(rectangle3_heights[1441]), .RECT3_WEIGHT(rectangle3_weights[1441]), .FEAT_THRES(feature_thresholds[1441]), .FEAT_ABOVE(feature_aboves[1441]), .FEAT_BELOW(feature_belows[1441])) ac1441(.scan_win(scan_win1441), .scan_win_std_dev(scan_win_std_dev[1441]), .feature_accum(feature_accums[1441]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1442]), .RECT1_Y(rectangle1_ys[1442]), .RECT1_WIDTH(rectangle1_widths[1442]), .RECT1_HEIGHT(rectangle1_heights[1442]), .RECT1_WEIGHT(rectangle1_weights[1442]), .RECT2_X(rectangle2_xs[1442]), .RECT2_Y(rectangle2_ys[1442]), .RECT2_WIDTH(rectangle2_widths[1442]), .RECT2_HEIGHT(rectangle2_heights[1442]), .RECT2_WEIGHT(rectangle2_weights[1442]), .RECT3_X(rectangle3_xs[1442]), .RECT3_Y(rectangle3_ys[1442]), .RECT3_WIDTH(rectangle3_widths[1442]), .RECT3_HEIGHT(rectangle3_heights[1442]), .RECT3_WEIGHT(rectangle3_weights[1442]), .FEAT_THRES(feature_thresholds[1442]), .FEAT_ABOVE(feature_aboves[1442]), .FEAT_BELOW(feature_belows[1442])) ac1442(.scan_win(scan_win1442), .scan_win_std_dev(scan_win_std_dev[1442]), .feature_accum(feature_accums[1442]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1443]), .RECT1_Y(rectangle1_ys[1443]), .RECT1_WIDTH(rectangle1_widths[1443]), .RECT1_HEIGHT(rectangle1_heights[1443]), .RECT1_WEIGHT(rectangle1_weights[1443]), .RECT2_X(rectangle2_xs[1443]), .RECT2_Y(rectangle2_ys[1443]), .RECT2_WIDTH(rectangle2_widths[1443]), .RECT2_HEIGHT(rectangle2_heights[1443]), .RECT2_WEIGHT(rectangle2_weights[1443]), .RECT3_X(rectangle3_xs[1443]), .RECT3_Y(rectangle3_ys[1443]), .RECT3_WIDTH(rectangle3_widths[1443]), .RECT3_HEIGHT(rectangle3_heights[1443]), .RECT3_WEIGHT(rectangle3_weights[1443]), .FEAT_THRES(feature_thresholds[1443]), .FEAT_ABOVE(feature_aboves[1443]), .FEAT_BELOW(feature_belows[1443])) ac1443(.scan_win(scan_win1443), .scan_win_std_dev(scan_win_std_dev[1443]), .feature_accum(feature_accums[1443]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1444]), .RECT1_Y(rectangle1_ys[1444]), .RECT1_WIDTH(rectangle1_widths[1444]), .RECT1_HEIGHT(rectangle1_heights[1444]), .RECT1_WEIGHT(rectangle1_weights[1444]), .RECT2_X(rectangle2_xs[1444]), .RECT2_Y(rectangle2_ys[1444]), .RECT2_WIDTH(rectangle2_widths[1444]), .RECT2_HEIGHT(rectangle2_heights[1444]), .RECT2_WEIGHT(rectangle2_weights[1444]), .RECT3_X(rectangle3_xs[1444]), .RECT3_Y(rectangle3_ys[1444]), .RECT3_WIDTH(rectangle3_widths[1444]), .RECT3_HEIGHT(rectangle3_heights[1444]), .RECT3_WEIGHT(rectangle3_weights[1444]), .FEAT_THRES(feature_thresholds[1444]), .FEAT_ABOVE(feature_aboves[1444]), .FEAT_BELOW(feature_belows[1444])) ac1444(.scan_win(scan_win1444), .scan_win_std_dev(scan_win_std_dev[1444]), .feature_accum(feature_accums[1444]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1445]), .RECT1_Y(rectangle1_ys[1445]), .RECT1_WIDTH(rectangle1_widths[1445]), .RECT1_HEIGHT(rectangle1_heights[1445]), .RECT1_WEIGHT(rectangle1_weights[1445]), .RECT2_X(rectangle2_xs[1445]), .RECT2_Y(rectangle2_ys[1445]), .RECT2_WIDTH(rectangle2_widths[1445]), .RECT2_HEIGHT(rectangle2_heights[1445]), .RECT2_WEIGHT(rectangle2_weights[1445]), .RECT3_X(rectangle3_xs[1445]), .RECT3_Y(rectangle3_ys[1445]), .RECT3_WIDTH(rectangle3_widths[1445]), .RECT3_HEIGHT(rectangle3_heights[1445]), .RECT3_WEIGHT(rectangle3_weights[1445]), .FEAT_THRES(feature_thresholds[1445]), .FEAT_ABOVE(feature_aboves[1445]), .FEAT_BELOW(feature_belows[1445])) ac1445(.scan_win(scan_win1445), .scan_win_std_dev(scan_win_std_dev[1445]), .feature_accum(feature_accums[1445]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1446]), .RECT1_Y(rectangle1_ys[1446]), .RECT1_WIDTH(rectangle1_widths[1446]), .RECT1_HEIGHT(rectangle1_heights[1446]), .RECT1_WEIGHT(rectangle1_weights[1446]), .RECT2_X(rectangle2_xs[1446]), .RECT2_Y(rectangle2_ys[1446]), .RECT2_WIDTH(rectangle2_widths[1446]), .RECT2_HEIGHT(rectangle2_heights[1446]), .RECT2_WEIGHT(rectangle2_weights[1446]), .RECT3_X(rectangle3_xs[1446]), .RECT3_Y(rectangle3_ys[1446]), .RECT3_WIDTH(rectangle3_widths[1446]), .RECT3_HEIGHT(rectangle3_heights[1446]), .RECT3_WEIGHT(rectangle3_weights[1446]), .FEAT_THRES(feature_thresholds[1446]), .FEAT_ABOVE(feature_aboves[1446]), .FEAT_BELOW(feature_belows[1446])) ac1446(.scan_win(scan_win1446), .scan_win_std_dev(scan_win_std_dev[1446]), .feature_accum(feature_accums[1446]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1447]), .RECT1_Y(rectangle1_ys[1447]), .RECT1_WIDTH(rectangle1_widths[1447]), .RECT1_HEIGHT(rectangle1_heights[1447]), .RECT1_WEIGHT(rectangle1_weights[1447]), .RECT2_X(rectangle2_xs[1447]), .RECT2_Y(rectangle2_ys[1447]), .RECT2_WIDTH(rectangle2_widths[1447]), .RECT2_HEIGHT(rectangle2_heights[1447]), .RECT2_WEIGHT(rectangle2_weights[1447]), .RECT3_X(rectangle3_xs[1447]), .RECT3_Y(rectangle3_ys[1447]), .RECT3_WIDTH(rectangle3_widths[1447]), .RECT3_HEIGHT(rectangle3_heights[1447]), .RECT3_WEIGHT(rectangle3_weights[1447]), .FEAT_THRES(feature_thresholds[1447]), .FEAT_ABOVE(feature_aboves[1447]), .FEAT_BELOW(feature_belows[1447])) ac1447(.scan_win(scan_win1447), .scan_win_std_dev(scan_win_std_dev[1447]), .feature_accum(feature_accums[1447]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1448]), .RECT1_Y(rectangle1_ys[1448]), .RECT1_WIDTH(rectangle1_widths[1448]), .RECT1_HEIGHT(rectangle1_heights[1448]), .RECT1_WEIGHT(rectangle1_weights[1448]), .RECT2_X(rectangle2_xs[1448]), .RECT2_Y(rectangle2_ys[1448]), .RECT2_WIDTH(rectangle2_widths[1448]), .RECT2_HEIGHT(rectangle2_heights[1448]), .RECT2_WEIGHT(rectangle2_weights[1448]), .RECT3_X(rectangle3_xs[1448]), .RECT3_Y(rectangle3_ys[1448]), .RECT3_WIDTH(rectangle3_widths[1448]), .RECT3_HEIGHT(rectangle3_heights[1448]), .RECT3_WEIGHT(rectangle3_weights[1448]), .FEAT_THRES(feature_thresholds[1448]), .FEAT_ABOVE(feature_aboves[1448]), .FEAT_BELOW(feature_belows[1448])) ac1448(.scan_win(scan_win1448), .scan_win_std_dev(scan_win_std_dev[1448]), .feature_accum(feature_accums[1448]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1449]), .RECT1_Y(rectangle1_ys[1449]), .RECT1_WIDTH(rectangle1_widths[1449]), .RECT1_HEIGHT(rectangle1_heights[1449]), .RECT1_WEIGHT(rectangle1_weights[1449]), .RECT2_X(rectangle2_xs[1449]), .RECT2_Y(rectangle2_ys[1449]), .RECT2_WIDTH(rectangle2_widths[1449]), .RECT2_HEIGHT(rectangle2_heights[1449]), .RECT2_WEIGHT(rectangle2_weights[1449]), .RECT3_X(rectangle3_xs[1449]), .RECT3_Y(rectangle3_ys[1449]), .RECT3_WIDTH(rectangle3_widths[1449]), .RECT3_HEIGHT(rectangle3_heights[1449]), .RECT3_WEIGHT(rectangle3_weights[1449]), .FEAT_THRES(feature_thresholds[1449]), .FEAT_ABOVE(feature_aboves[1449]), .FEAT_BELOW(feature_belows[1449])) ac1449(.scan_win(scan_win1449), .scan_win_std_dev(scan_win_std_dev[1449]), .feature_accum(feature_accums[1449]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1450]), .RECT1_Y(rectangle1_ys[1450]), .RECT1_WIDTH(rectangle1_widths[1450]), .RECT1_HEIGHT(rectangle1_heights[1450]), .RECT1_WEIGHT(rectangle1_weights[1450]), .RECT2_X(rectangle2_xs[1450]), .RECT2_Y(rectangle2_ys[1450]), .RECT2_WIDTH(rectangle2_widths[1450]), .RECT2_HEIGHT(rectangle2_heights[1450]), .RECT2_WEIGHT(rectangle2_weights[1450]), .RECT3_X(rectangle3_xs[1450]), .RECT3_Y(rectangle3_ys[1450]), .RECT3_WIDTH(rectangle3_widths[1450]), .RECT3_HEIGHT(rectangle3_heights[1450]), .RECT3_WEIGHT(rectangle3_weights[1450]), .FEAT_THRES(feature_thresholds[1450]), .FEAT_ABOVE(feature_aboves[1450]), .FEAT_BELOW(feature_belows[1450])) ac1450(.scan_win(scan_win1450), .scan_win_std_dev(scan_win_std_dev[1450]), .feature_accum(feature_accums[1450]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1451]), .RECT1_Y(rectangle1_ys[1451]), .RECT1_WIDTH(rectangle1_widths[1451]), .RECT1_HEIGHT(rectangle1_heights[1451]), .RECT1_WEIGHT(rectangle1_weights[1451]), .RECT2_X(rectangle2_xs[1451]), .RECT2_Y(rectangle2_ys[1451]), .RECT2_WIDTH(rectangle2_widths[1451]), .RECT2_HEIGHT(rectangle2_heights[1451]), .RECT2_WEIGHT(rectangle2_weights[1451]), .RECT3_X(rectangle3_xs[1451]), .RECT3_Y(rectangle3_ys[1451]), .RECT3_WIDTH(rectangle3_widths[1451]), .RECT3_HEIGHT(rectangle3_heights[1451]), .RECT3_WEIGHT(rectangle3_weights[1451]), .FEAT_THRES(feature_thresholds[1451]), .FEAT_ABOVE(feature_aboves[1451]), .FEAT_BELOW(feature_belows[1451])) ac1451(.scan_win(scan_win1451), .scan_win_std_dev(scan_win_std_dev[1451]), .feature_accum(feature_accums[1451]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1452]), .RECT1_Y(rectangle1_ys[1452]), .RECT1_WIDTH(rectangle1_widths[1452]), .RECT1_HEIGHT(rectangle1_heights[1452]), .RECT1_WEIGHT(rectangle1_weights[1452]), .RECT2_X(rectangle2_xs[1452]), .RECT2_Y(rectangle2_ys[1452]), .RECT2_WIDTH(rectangle2_widths[1452]), .RECT2_HEIGHT(rectangle2_heights[1452]), .RECT2_WEIGHT(rectangle2_weights[1452]), .RECT3_X(rectangle3_xs[1452]), .RECT3_Y(rectangle3_ys[1452]), .RECT3_WIDTH(rectangle3_widths[1452]), .RECT3_HEIGHT(rectangle3_heights[1452]), .RECT3_WEIGHT(rectangle3_weights[1452]), .FEAT_THRES(feature_thresholds[1452]), .FEAT_ABOVE(feature_aboves[1452]), .FEAT_BELOW(feature_belows[1452])) ac1452(.scan_win(scan_win1452), .scan_win_std_dev(scan_win_std_dev[1452]), .feature_accum(feature_accums[1452]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1453]), .RECT1_Y(rectangle1_ys[1453]), .RECT1_WIDTH(rectangle1_widths[1453]), .RECT1_HEIGHT(rectangle1_heights[1453]), .RECT1_WEIGHT(rectangle1_weights[1453]), .RECT2_X(rectangle2_xs[1453]), .RECT2_Y(rectangle2_ys[1453]), .RECT2_WIDTH(rectangle2_widths[1453]), .RECT2_HEIGHT(rectangle2_heights[1453]), .RECT2_WEIGHT(rectangle2_weights[1453]), .RECT3_X(rectangle3_xs[1453]), .RECT3_Y(rectangle3_ys[1453]), .RECT3_WIDTH(rectangle3_widths[1453]), .RECT3_HEIGHT(rectangle3_heights[1453]), .RECT3_WEIGHT(rectangle3_weights[1453]), .FEAT_THRES(feature_thresholds[1453]), .FEAT_ABOVE(feature_aboves[1453]), .FEAT_BELOW(feature_belows[1453])) ac1453(.scan_win(scan_win1453), .scan_win_std_dev(scan_win_std_dev[1453]), .feature_accum(feature_accums[1453]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1454]), .RECT1_Y(rectangle1_ys[1454]), .RECT1_WIDTH(rectangle1_widths[1454]), .RECT1_HEIGHT(rectangle1_heights[1454]), .RECT1_WEIGHT(rectangle1_weights[1454]), .RECT2_X(rectangle2_xs[1454]), .RECT2_Y(rectangle2_ys[1454]), .RECT2_WIDTH(rectangle2_widths[1454]), .RECT2_HEIGHT(rectangle2_heights[1454]), .RECT2_WEIGHT(rectangle2_weights[1454]), .RECT3_X(rectangle3_xs[1454]), .RECT3_Y(rectangle3_ys[1454]), .RECT3_WIDTH(rectangle3_widths[1454]), .RECT3_HEIGHT(rectangle3_heights[1454]), .RECT3_WEIGHT(rectangle3_weights[1454]), .FEAT_THRES(feature_thresholds[1454]), .FEAT_ABOVE(feature_aboves[1454]), .FEAT_BELOW(feature_belows[1454])) ac1454(.scan_win(scan_win1454), .scan_win_std_dev(scan_win_std_dev[1454]), .feature_accum(feature_accums[1454]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1455]), .RECT1_Y(rectangle1_ys[1455]), .RECT1_WIDTH(rectangle1_widths[1455]), .RECT1_HEIGHT(rectangle1_heights[1455]), .RECT1_WEIGHT(rectangle1_weights[1455]), .RECT2_X(rectangle2_xs[1455]), .RECT2_Y(rectangle2_ys[1455]), .RECT2_WIDTH(rectangle2_widths[1455]), .RECT2_HEIGHT(rectangle2_heights[1455]), .RECT2_WEIGHT(rectangle2_weights[1455]), .RECT3_X(rectangle3_xs[1455]), .RECT3_Y(rectangle3_ys[1455]), .RECT3_WIDTH(rectangle3_widths[1455]), .RECT3_HEIGHT(rectangle3_heights[1455]), .RECT3_WEIGHT(rectangle3_weights[1455]), .FEAT_THRES(feature_thresholds[1455]), .FEAT_ABOVE(feature_aboves[1455]), .FEAT_BELOW(feature_belows[1455])) ac1455(.scan_win(scan_win1455), .scan_win_std_dev(scan_win_std_dev[1455]), .feature_accum(feature_accums[1455]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1456]), .RECT1_Y(rectangle1_ys[1456]), .RECT1_WIDTH(rectangle1_widths[1456]), .RECT1_HEIGHT(rectangle1_heights[1456]), .RECT1_WEIGHT(rectangle1_weights[1456]), .RECT2_X(rectangle2_xs[1456]), .RECT2_Y(rectangle2_ys[1456]), .RECT2_WIDTH(rectangle2_widths[1456]), .RECT2_HEIGHT(rectangle2_heights[1456]), .RECT2_WEIGHT(rectangle2_weights[1456]), .RECT3_X(rectangle3_xs[1456]), .RECT3_Y(rectangle3_ys[1456]), .RECT3_WIDTH(rectangle3_widths[1456]), .RECT3_HEIGHT(rectangle3_heights[1456]), .RECT3_WEIGHT(rectangle3_weights[1456]), .FEAT_THRES(feature_thresholds[1456]), .FEAT_ABOVE(feature_aboves[1456]), .FEAT_BELOW(feature_belows[1456])) ac1456(.scan_win(scan_win1456), .scan_win_std_dev(scan_win_std_dev[1456]), .feature_accum(feature_accums[1456]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1457]), .RECT1_Y(rectangle1_ys[1457]), .RECT1_WIDTH(rectangle1_widths[1457]), .RECT1_HEIGHT(rectangle1_heights[1457]), .RECT1_WEIGHT(rectangle1_weights[1457]), .RECT2_X(rectangle2_xs[1457]), .RECT2_Y(rectangle2_ys[1457]), .RECT2_WIDTH(rectangle2_widths[1457]), .RECT2_HEIGHT(rectangle2_heights[1457]), .RECT2_WEIGHT(rectangle2_weights[1457]), .RECT3_X(rectangle3_xs[1457]), .RECT3_Y(rectangle3_ys[1457]), .RECT3_WIDTH(rectangle3_widths[1457]), .RECT3_HEIGHT(rectangle3_heights[1457]), .RECT3_WEIGHT(rectangle3_weights[1457]), .FEAT_THRES(feature_thresholds[1457]), .FEAT_ABOVE(feature_aboves[1457]), .FEAT_BELOW(feature_belows[1457])) ac1457(.scan_win(scan_win1457), .scan_win_std_dev(scan_win_std_dev[1457]), .feature_accum(feature_accums[1457]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1458]), .RECT1_Y(rectangle1_ys[1458]), .RECT1_WIDTH(rectangle1_widths[1458]), .RECT1_HEIGHT(rectangle1_heights[1458]), .RECT1_WEIGHT(rectangle1_weights[1458]), .RECT2_X(rectangle2_xs[1458]), .RECT2_Y(rectangle2_ys[1458]), .RECT2_WIDTH(rectangle2_widths[1458]), .RECT2_HEIGHT(rectangle2_heights[1458]), .RECT2_WEIGHT(rectangle2_weights[1458]), .RECT3_X(rectangle3_xs[1458]), .RECT3_Y(rectangle3_ys[1458]), .RECT3_WIDTH(rectangle3_widths[1458]), .RECT3_HEIGHT(rectangle3_heights[1458]), .RECT3_WEIGHT(rectangle3_weights[1458]), .FEAT_THRES(feature_thresholds[1458]), .FEAT_ABOVE(feature_aboves[1458]), .FEAT_BELOW(feature_belows[1458])) ac1458(.scan_win(scan_win1458), .scan_win_std_dev(scan_win_std_dev[1458]), .feature_accum(feature_accums[1458]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1459]), .RECT1_Y(rectangle1_ys[1459]), .RECT1_WIDTH(rectangle1_widths[1459]), .RECT1_HEIGHT(rectangle1_heights[1459]), .RECT1_WEIGHT(rectangle1_weights[1459]), .RECT2_X(rectangle2_xs[1459]), .RECT2_Y(rectangle2_ys[1459]), .RECT2_WIDTH(rectangle2_widths[1459]), .RECT2_HEIGHT(rectangle2_heights[1459]), .RECT2_WEIGHT(rectangle2_weights[1459]), .RECT3_X(rectangle3_xs[1459]), .RECT3_Y(rectangle3_ys[1459]), .RECT3_WIDTH(rectangle3_widths[1459]), .RECT3_HEIGHT(rectangle3_heights[1459]), .RECT3_WEIGHT(rectangle3_weights[1459]), .FEAT_THRES(feature_thresholds[1459]), .FEAT_ABOVE(feature_aboves[1459]), .FEAT_BELOW(feature_belows[1459])) ac1459(.scan_win(scan_win1459), .scan_win_std_dev(scan_win_std_dev[1459]), .feature_accum(feature_accums[1459]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1460]), .RECT1_Y(rectangle1_ys[1460]), .RECT1_WIDTH(rectangle1_widths[1460]), .RECT1_HEIGHT(rectangle1_heights[1460]), .RECT1_WEIGHT(rectangle1_weights[1460]), .RECT2_X(rectangle2_xs[1460]), .RECT2_Y(rectangle2_ys[1460]), .RECT2_WIDTH(rectangle2_widths[1460]), .RECT2_HEIGHT(rectangle2_heights[1460]), .RECT2_WEIGHT(rectangle2_weights[1460]), .RECT3_X(rectangle3_xs[1460]), .RECT3_Y(rectangle3_ys[1460]), .RECT3_WIDTH(rectangle3_widths[1460]), .RECT3_HEIGHT(rectangle3_heights[1460]), .RECT3_WEIGHT(rectangle3_weights[1460]), .FEAT_THRES(feature_thresholds[1460]), .FEAT_ABOVE(feature_aboves[1460]), .FEAT_BELOW(feature_belows[1460])) ac1460(.scan_win(scan_win1460), .scan_win_std_dev(scan_win_std_dev[1460]), .feature_accum(feature_accums[1460]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1461]), .RECT1_Y(rectangle1_ys[1461]), .RECT1_WIDTH(rectangle1_widths[1461]), .RECT1_HEIGHT(rectangle1_heights[1461]), .RECT1_WEIGHT(rectangle1_weights[1461]), .RECT2_X(rectangle2_xs[1461]), .RECT2_Y(rectangle2_ys[1461]), .RECT2_WIDTH(rectangle2_widths[1461]), .RECT2_HEIGHT(rectangle2_heights[1461]), .RECT2_WEIGHT(rectangle2_weights[1461]), .RECT3_X(rectangle3_xs[1461]), .RECT3_Y(rectangle3_ys[1461]), .RECT3_WIDTH(rectangle3_widths[1461]), .RECT3_HEIGHT(rectangle3_heights[1461]), .RECT3_WEIGHT(rectangle3_weights[1461]), .FEAT_THRES(feature_thresholds[1461]), .FEAT_ABOVE(feature_aboves[1461]), .FEAT_BELOW(feature_belows[1461])) ac1461(.scan_win(scan_win1461), .scan_win_std_dev(scan_win_std_dev[1461]), .feature_accum(feature_accums[1461]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1462]), .RECT1_Y(rectangle1_ys[1462]), .RECT1_WIDTH(rectangle1_widths[1462]), .RECT1_HEIGHT(rectangle1_heights[1462]), .RECT1_WEIGHT(rectangle1_weights[1462]), .RECT2_X(rectangle2_xs[1462]), .RECT2_Y(rectangle2_ys[1462]), .RECT2_WIDTH(rectangle2_widths[1462]), .RECT2_HEIGHT(rectangle2_heights[1462]), .RECT2_WEIGHT(rectangle2_weights[1462]), .RECT3_X(rectangle3_xs[1462]), .RECT3_Y(rectangle3_ys[1462]), .RECT3_WIDTH(rectangle3_widths[1462]), .RECT3_HEIGHT(rectangle3_heights[1462]), .RECT3_WEIGHT(rectangle3_weights[1462]), .FEAT_THRES(feature_thresholds[1462]), .FEAT_ABOVE(feature_aboves[1462]), .FEAT_BELOW(feature_belows[1462])) ac1462(.scan_win(scan_win1462), .scan_win_std_dev(scan_win_std_dev[1462]), .feature_accum(feature_accums[1462]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1463]), .RECT1_Y(rectangle1_ys[1463]), .RECT1_WIDTH(rectangle1_widths[1463]), .RECT1_HEIGHT(rectangle1_heights[1463]), .RECT1_WEIGHT(rectangle1_weights[1463]), .RECT2_X(rectangle2_xs[1463]), .RECT2_Y(rectangle2_ys[1463]), .RECT2_WIDTH(rectangle2_widths[1463]), .RECT2_HEIGHT(rectangle2_heights[1463]), .RECT2_WEIGHT(rectangle2_weights[1463]), .RECT3_X(rectangle3_xs[1463]), .RECT3_Y(rectangle3_ys[1463]), .RECT3_WIDTH(rectangle3_widths[1463]), .RECT3_HEIGHT(rectangle3_heights[1463]), .RECT3_WEIGHT(rectangle3_weights[1463]), .FEAT_THRES(feature_thresholds[1463]), .FEAT_ABOVE(feature_aboves[1463]), .FEAT_BELOW(feature_belows[1463])) ac1463(.scan_win(scan_win1463), .scan_win_std_dev(scan_win_std_dev[1463]), .feature_accum(feature_accums[1463]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1464]), .RECT1_Y(rectangle1_ys[1464]), .RECT1_WIDTH(rectangle1_widths[1464]), .RECT1_HEIGHT(rectangle1_heights[1464]), .RECT1_WEIGHT(rectangle1_weights[1464]), .RECT2_X(rectangle2_xs[1464]), .RECT2_Y(rectangle2_ys[1464]), .RECT2_WIDTH(rectangle2_widths[1464]), .RECT2_HEIGHT(rectangle2_heights[1464]), .RECT2_WEIGHT(rectangle2_weights[1464]), .RECT3_X(rectangle3_xs[1464]), .RECT3_Y(rectangle3_ys[1464]), .RECT3_WIDTH(rectangle3_widths[1464]), .RECT3_HEIGHT(rectangle3_heights[1464]), .RECT3_WEIGHT(rectangle3_weights[1464]), .FEAT_THRES(feature_thresholds[1464]), .FEAT_ABOVE(feature_aboves[1464]), .FEAT_BELOW(feature_belows[1464])) ac1464(.scan_win(scan_win1464), .scan_win_std_dev(scan_win_std_dev[1464]), .feature_accum(feature_accums[1464]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1465]), .RECT1_Y(rectangle1_ys[1465]), .RECT1_WIDTH(rectangle1_widths[1465]), .RECT1_HEIGHT(rectangle1_heights[1465]), .RECT1_WEIGHT(rectangle1_weights[1465]), .RECT2_X(rectangle2_xs[1465]), .RECT2_Y(rectangle2_ys[1465]), .RECT2_WIDTH(rectangle2_widths[1465]), .RECT2_HEIGHT(rectangle2_heights[1465]), .RECT2_WEIGHT(rectangle2_weights[1465]), .RECT3_X(rectangle3_xs[1465]), .RECT3_Y(rectangle3_ys[1465]), .RECT3_WIDTH(rectangle3_widths[1465]), .RECT3_HEIGHT(rectangle3_heights[1465]), .RECT3_WEIGHT(rectangle3_weights[1465]), .FEAT_THRES(feature_thresholds[1465]), .FEAT_ABOVE(feature_aboves[1465]), .FEAT_BELOW(feature_belows[1465])) ac1465(.scan_win(scan_win1465), .scan_win_std_dev(scan_win_std_dev[1465]), .feature_accum(feature_accums[1465]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1466]), .RECT1_Y(rectangle1_ys[1466]), .RECT1_WIDTH(rectangle1_widths[1466]), .RECT1_HEIGHT(rectangle1_heights[1466]), .RECT1_WEIGHT(rectangle1_weights[1466]), .RECT2_X(rectangle2_xs[1466]), .RECT2_Y(rectangle2_ys[1466]), .RECT2_WIDTH(rectangle2_widths[1466]), .RECT2_HEIGHT(rectangle2_heights[1466]), .RECT2_WEIGHT(rectangle2_weights[1466]), .RECT3_X(rectangle3_xs[1466]), .RECT3_Y(rectangle3_ys[1466]), .RECT3_WIDTH(rectangle3_widths[1466]), .RECT3_HEIGHT(rectangle3_heights[1466]), .RECT3_WEIGHT(rectangle3_weights[1466]), .FEAT_THRES(feature_thresholds[1466]), .FEAT_ABOVE(feature_aboves[1466]), .FEAT_BELOW(feature_belows[1466])) ac1466(.scan_win(scan_win1466), .scan_win_std_dev(scan_win_std_dev[1466]), .feature_accum(feature_accums[1466]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1467]), .RECT1_Y(rectangle1_ys[1467]), .RECT1_WIDTH(rectangle1_widths[1467]), .RECT1_HEIGHT(rectangle1_heights[1467]), .RECT1_WEIGHT(rectangle1_weights[1467]), .RECT2_X(rectangle2_xs[1467]), .RECT2_Y(rectangle2_ys[1467]), .RECT2_WIDTH(rectangle2_widths[1467]), .RECT2_HEIGHT(rectangle2_heights[1467]), .RECT2_WEIGHT(rectangle2_weights[1467]), .RECT3_X(rectangle3_xs[1467]), .RECT3_Y(rectangle3_ys[1467]), .RECT3_WIDTH(rectangle3_widths[1467]), .RECT3_HEIGHT(rectangle3_heights[1467]), .RECT3_WEIGHT(rectangle3_weights[1467]), .FEAT_THRES(feature_thresholds[1467]), .FEAT_ABOVE(feature_aboves[1467]), .FEAT_BELOW(feature_belows[1467])) ac1467(.scan_win(scan_win1467), .scan_win_std_dev(scan_win_std_dev[1467]), .feature_accum(feature_accums[1467]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1468]), .RECT1_Y(rectangle1_ys[1468]), .RECT1_WIDTH(rectangle1_widths[1468]), .RECT1_HEIGHT(rectangle1_heights[1468]), .RECT1_WEIGHT(rectangle1_weights[1468]), .RECT2_X(rectangle2_xs[1468]), .RECT2_Y(rectangle2_ys[1468]), .RECT2_WIDTH(rectangle2_widths[1468]), .RECT2_HEIGHT(rectangle2_heights[1468]), .RECT2_WEIGHT(rectangle2_weights[1468]), .RECT3_X(rectangle3_xs[1468]), .RECT3_Y(rectangle3_ys[1468]), .RECT3_WIDTH(rectangle3_widths[1468]), .RECT3_HEIGHT(rectangle3_heights[1468]), .RECT3_WEIGHT(rectangle3_weights[1468]), .FEAT_THRES(feature_thresholds[1468]), .FEAT_ABOVE(feature_aboves[1468]), .FEAT_BELOW(feature_belows[1468])) ac1468(.scan_win(scan_win1468), .scan_win_std_dev(scan_win_std_dev[1468]), .feature_accum(feature_accums[1468]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1469]), .RECT1_Y(rectangle1_ys[1469]), .RECT1_WIDTH(rectangle1_widths[1469]), .RECT1_HEIGHT(rectangle1_heights[1469]), .RECT1_WEIGHT(rectangle1_weights[1469]), .RECT2_X(rectangle2_xs[1469]), .RECT2_Y(rectangle2_ys[1469]), .RECT2_WIDTH(rectangle2_widths[1469]), .RECT2_HEIGHT(rectangle2_heights[1469]), .RECT2_WEIGHT(rectangle2_weights[1469]), .RECT3_X(rectangle3_xs[1469]), .RECT3_Y(rectangle3_ys[1469]), .RECT3_WIDTH(rectangle3_widths[1469]), .RECT3_HEIGHT(rectangle3_heights[1469]), .RECT3_WEIGHT(rectangle3_weights[1469]), .FEAT_THRES(feature_thresholds[1469]), .FEAT_ABOVE(feature_aboves[1469]), .FEAT_BELOW(feature_belows[1469])) ac1469(.scan_win(scan_win1469), .scan_win_std_dev(scan_win_std_dev[1469]), .feature_accum(feature_accums[1469]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1470]), .RECT1_Y(rectangle1_ys[1470]), .RECT1_WIDTH(rectangle1_widths[1470]), .RECT1_HEIGHT(rectangle1_heights[1470]), .RECT1_WEIGHT(rectangle1_weights[1470]), .RECT2_X(rectangle2_xs[1470]), .RECT2_Y(rectangle2_ys[1470]), .RECT2_WIDTH(rectangle2_widths[1470]), .RECT2_HEIGHT(rectangle2_heights[1470]), .RECT2_WEIGHT(rectangle2_weights[1470]), .RECT3_X(rectangle3_xs[1470]), .RECT3_Y(rectangle3_ys[1470]), .RECT3_WIDTH(rectangle3_widths[1470]), .RECT3_HEIGHT(rectangle3_heights[1470]), .RECT3_WEIGHT(rectangle3_weights[1470]), .FEAT_THRES(feature_thresholds[1470]), .FEAT_ABOVE(feature_aboves[1470]), .FEAT_BELOW(feature_belows[1470])) ac1470(.scan_win(scan_win1470), .scan_win_std_dev(scan_win_std_dev[1470]), .feature_accum(feature_accums[1470]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1471]), .RECT1_Y(rectangle1_ys[1471]), .RECT1_WIDTH(rectangle1_widths[1471]), .RECT1_HEIGHT(rectangle1_heights[1471]), .RECT1_WEIGHT(rectangle1_weights[1471]), .RECT2_X(rectangle2_xs[1471]), .RECT2_Y(rectangle2_ys[1471]), .RECT2_WIDTH(rectangle2_widths[1471]), .RECT2_HEIGHT(rectangle2_heights[1471]), .RECT2_WEIGHT(rectangle2_weights[1471]), .RECT3_X(rectangle3_xs[1471]), .RECT3_Y(rectangle3_ys[1471]), .RECT3_WIDTH(rectangle3_widths[1471]), .RECT3_HEIGHT(rectangle3_heights[1471]), .RECT3_WEIGHT(rectangle3_weights[1471]), .FEAT_THRES(feature_thresholds[1471]), .FEAT_ABOVE(feature_aboves[1471]), .FEAT_BELOW(feature_belows[1471])) ac1471(.scan_win(scan_win1471), .scan_win_std_dev(scan_win_std_dev[1471]), .feature_accum(feature_accums[1471]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1472]), .RECT1_Y(rectangle1_ys[1472]), .RECT1_WIDTH(rectangle1_widths[1472]), .RECT1_HEIGHT(rectangle1_heights[1472]), .RECT1_WEIGHT(rectangle1_weights[1472]), .RECT2_X(rectangle2_xs[1472]), .RECT2_Y(rectangle2_ys[1472]), .RECT2_WIDTH(rectangle2_widths[1472]), .RECT2_HEIGHT(rectangle2_heights[1472]), .RECT2_WEIGHT(rectangle2_weights[1472]), .RECT3_X(rectangle3_xs[1472]), .RECT3_Y(rectangle3_ys[1472]), .RECT3_WIDTH(rectangle3_widths[1472]), .RECT3_HEIGHT(rectangle3_heights[1472]), .RECT3_WEIGHT(rectangle3_weights[1472]), .FEAT_THRES(feature_thresholds[1472]), .FEAT_ABOVE(feature_aboves[1472]), .FEAT_BELOW(feature_belows[1472])) ac1472(.scan_win(scan_win1472), .scan_win_std_dev(scan_win_std_dev[1472]), .feature_accum(feature_accums[1472]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1473]), .RECT1_Y(rectangle1_ys[1473]), .RECT1_WIDTH(rectangle1_widths[1473]), .RECT1_HEIGHT(rectangle1_heights[1473]), .RECT1_WEIGHT(rectangle1_weights[1473]), .RECT2_X(rectangle2_xs[1473]), .RECT2_Y(rectangle2_ys[1473]), .RECT2_WIDTH(rectangle2_widths[1473]), .RECT2_HEIGHT(rectangle2_heights[1473]), .RECT2_WEIGHT(rectangle2_weights[1473]), .RECT3_X(rectangle3_xs[1473]), .RECT3_Y(rectangle3_ys[1473]), .RECT3_WIDTH(rectangle3_widths[1473]), .RECT3_HEIGHT(rectangle3_heights[1473]), .RECT3_WEIGHT(rectangle3_weights[1473]), .FEAT_THRES(feature_thresholds[1473]), .FEAT_ABOVE(feature_aboves[1473]), .FEAT_BELOW(feature_belows[1473])) ac1473(.scan_win(scan_win1473), .scan_win_std_dev(scan_win_std_dev[1473]), .feature_accum(feature_accums[1473]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1474]), .RECT1_Y(rectangle1_ys[1474]), .RECT1_WIDTH(rectangle1_widths[1474]), .RECT1_HEIGHT(rectangle1_heights[1474]), .RECT1_WEIGHT(rectangle1_weights[1474]), .RECT2_X(rectangle2_xs[1474]), .RECT2_Y(rectangle2_ys[1474]), .RECT2_WIDTH(rectangle2_widths[1474]), .RECT2_HEIGHT(rectangle2_heights[1474]), .RECT2_WEIGHT(rectangle2_weights[1474]), .RECT3_X(rectangle3_xs[1474]), .RECT3_Y(rectangle3_ys[1474]), .RECT3_WIDTH(rectangle3_widths[1474]), .RECT3_HEIGHT(rectangle3_heights[1474]), .RECT3_WEIGHT(rectangle3_weights[1474]), .FEAT_THRES(feature_thresholds[1474]), .FEAT_ABOVE(feature_aboves[1474]), .FEAT_BELOW(feature_belows[1474])) ac1474(.scan_win(scan_win1474), .scan_win_std_dev(scan_win_std_dev[1474]), .feature_accum(feature_accums[1474]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1475]), .RECT1_Y(rectangle1_ys[1475]), .RECT1_WIDTH(rectangle1_widths[1475]), .RECT1_HEIGHT(rectangle1_heights[1475]), .RECT1_WEIGHT(rectangle1_weights[1475]), .RECT2_X(rectangle2_xs[1475]), .RECT2_Y(rectangle2_ys[1475]), .RECT2_WIDTH(rectangle2_widths[1475]), .RECT2_HEIGHT(rectangle2_heights[1475]), .RECT2_WEIGHT(rectangle2_weights[1475]), .RECT3_X(rectangle3_xs[1475]), .RECT3_Y(rectangle3_ys[1475]), .RECT3_WIDTH(rectangle3_widths[1475]), .RECT3_HEIGHT(rectangle3_heights[1475]), .RECT3_WEIGHT(rectangle3_weights[1475]), .FEAT_THRES(feature_thresholds[1475]), .FEAT_ABOVE(feature_aboves[1475]), .FEAT_BELOW(feature_belows[1475])) ac1475(.scan_win(scan_win1475), .scan_win_std_dev(scan_win_std_dev[1475]), .feature_accum(feature_accums[1475]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1476]), .RECT1_Y(rectangle1_ys[1476]), .RECT1_WIDTH(rectangle1_widths[1476]), .RECT1_HEIGHT(rectangle1_heights[1476]), .RECT1_WEIGHT(rectangle1_weights[1476]), .RECT2_X(rectangle2_xs[1476]), .RECT2_Y(rectangle2_ys[1476]), .RECT2_WIDTH(rectangle2_widths[1476]), .RECT2_HEIGHT(rectangle2_heights[1476]), .RECT2_WEIGHT(rectangle2_weights[1476]), .RECT3_X(rectangle3_xs[1476]), .RECT3_Y(rectangle3_ys[1476]), .RECT3_WIDTH(rectangle3_widths[1476]), .RECT3_HEIGHT(rectangle3_heights[1476]), .RECT3_WEIGHT(rectangle3_weights[1476]), .FEAT_THRES(feature_thresholds[1476]), .FEAT_ABOVE(feature_aboves[1476]), .FEAT_BELOW(feature_belows[1476])) ac1476(.scan_win(scan_win1476), .scan_win_std_dev(scan_win_std_dev[1476]), .feature_accum(feature_accums[1476]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1477]), .RECT1_Y(rectangle1_ys[1477]), .RECT1_WIDTH(rectangle1_widths[1477]), .RECT1_HEIGHT(rectangle1_heights[1477]), .RECT1_WEIGHT(rectangle1_weights[1477]), .RECT2_X(rectangle2_xs[1477]), .RECT2_Y(rectangle2_ys[1477]), .RECT2_WIDTH(rectangle2_widths[1477]), .RECT2_HEIGHT(rectangle2_heights[1477]), .RECT2_WEIGHT(rectangle2_weights[1477]), .RECT3_X(rectangle3_xs[1477]), .RECT3_Y(rectangle3_ys[1477]), .RECT3_WIDTH(rectangle3_widths[1477]), .RECT3_HEIGHT(rectangle3_heights[1477]), .RECT3_WEIGHT(rectangle3_weights[1477]), .FEAT_THRES(feature_thresholds[1477]), .FEAT_ABOVE(feature_aboves[1477]), .FEAT_BELOW(feature_belows[1477])) ac1477(.scan_win(scan_win1477), .scan_win_std_dev(scan_win_std_dev[1477]), .feature_accum(feature_accums[1477]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1478]), .RECT1_Y(rectangle1_ys[1478]), .RECT1_WIDTH(rectangle1_widths[1478]), .RECT1_HEIGHT(rectangle1_heights[1478]), .RECT1_WEIGHT(rectangle1_weights[1478]), .RECT2_X(rectangle2_xs[1478]), .RECT2_Y(rectangle2_ys[1478]), .RECT2_WIDTH(rectangle2_widths[1478]), .RECT2_HEIGHT(rectangle2_heights[1478]), .RECT2_WEIGHT(rectangle2_weights[1478]), .RECT3_X(rectangle3_xs[1478]), .RECT3_Y(rectangle3_ys[1478]), .RECT3_WIDTH(rectangle3_widths[1478]), .RECT3_HEIGHT(rectangle3_heights[1478]), .RECT3_WEIGHT(rectangle3_weights[1478]), .FEAT_THRES(feature_thresholds[1478]), .FEAT_ABOVE(feature_aboves[1478]), .FEAT_BELOW(feature_belows[1478])) ac1478(.scan_win(scan_win1478), .scan_win_std_dev(scan_win_std_dev[1478]), .feature_accum(feature_accums[1478]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1479]), .RECT1_Y(rectangle1_ys[1479]), .RECT1_WIDTH(rectangle1_widths[1479]), .RECT1_HEIGHT(rectangle1_heights[1479]), .RECT1_WEIGHT(rectangle1_weights[1479]), .RECT2_X(rectangle2_xs[1479]), .RECT2_Y(rectangle2_ys[1479]), .RECT2_WIDTH(rectangle2_widths[1479]), .RECT2_HEIGHT(rectangle2_heights[1479]), .RECT2_WEIGHT(rectangle2_weights[1479]), .RECT3_X(rectangle3_xs[1479]), .RECT3_Y(rectangle3_ys[1479]), .RECT3_WIDTH(rectangle3_widths[1479]), .RECT3_HEIGHT(rectangle3_heights[1479]), .RECT3_WEIGHT(rectangle3_weights[1479]), .FEAT_THRES(feature_thresholds[1479]), .FEAT_ABOVE(feature_aboves[1479]), .FEAT_BELOW(feature_belows[1479])) ac1479(.scan_win(scan_win1479), .scan_win_std_dev(scan_win_std_dev[1479]), .feature_accum(feature_accums[1479]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1480]), .RECT1_Y(rectangle1_ys[1480]), .RECT1_WIDTH(rectangle1_widths[1480]), .RECT1_HEIGHT(rectangle1_heights[1480]), .RECT1_WEIGHT(rectangle1_weights[1480]), .RECT2_X(rectangle2_xs[1480]), .RECT2_Y(rectangle2_ys[1480]), .RECT2_WIDTH(rectangle2_widths[1480]), .RECT2_HEIGHT(rectangle2_heights[1480]), .RECT2_WEIGHT(rectangle2_weights[1480]), .RECT3_X(rectangle3_xs[1480]), .RECT3_Y(rectangle3_ys[1480]), .RECT3_WIDTH(rectangle3_widths[1480]), .RECT3_HEIGHT(rectangle3_heights[1480]), .RECT3_WEIGHT(rectangle3_weights[1480]), .FEAT_THRES(feature_thresholds[1480]), .FEAT_ABOVE(feature_aboves[1480]), .FEAT_BELOW(feature_belows[1480])) ac1480(.scan_win(scan_win1480), .scan_win_std_dev(scan_win_std_dev[1480]), .feature_accum(feature_accums[1480]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1481]), .RECT1_Y(rectangle1_ys[1481]), .RECT1_WIDTH(rectangle1_widths[1481]), .RECT1_HEIGHT(rectangle1_heights[1481]), .RECT1_WEIGHT(rectangle1_weights[1481]), .RECT2_X(rectangle2_xs[1481]), .RECT2_Y(rectangle2_ys[1481]), .RECT2_WIDTH(rectangle2_widths[1481]), .RECT2_HEIGHT(rectangle2_heights[1481]), .RECT2_WEIGHT(rectangle2_weights[1481]), .RECT3_X(rectangle3_xs[1481]), .RECT3_Y(rectangle3_ys[1481]), .RECT3_WIDTH(rectangle3_widths[1481]), .RECT3_HEIGHT(rectangle3_heights[1481]), .RECT3_WEIGHT(rectangle3_weights[1481]), .FEAT_THRES(feature_thresholds[1481]), .FEAT_ABOVE(feature_aboves[1481]), .FEAT_BELOW(feature_belows[1481])) ac1481(.scan_win(scan_win1481), .scan_win_std_dev(scan_win_std_dev[1481]), .feature_accum(feature_accums[1481]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1482]), .RECT1_Y(rectangle1_ys[1482]), .RECT1_WIDTH(rectangle1_widths[1482]), .RECT1_HEIGHT(rectangle1_heights[1482]), .RECT1_WEIGHT(rectangle1_weights[1482]), .RECT2_X(rectangle2_xs[1482]), .RECT2_Y(rectangle2_ys[1482]), .RECT2_WIDTH(rectangle2_widths[1482]), .RECT2_HEIGHT(rectangle2_heights[1482]), .RECT2_WEIGHT(rectangle2_weights[1482]), .RECT3_X(rectangle3_xs[1482]), .RECT3_Y(rectangle3_ys[1482]), .RECT3_WIDTH(rectangle3_widths[1482]), .RECT3_HEIGHT(rectangle3_heights[1482]), .RECT3_WEIGHT(rectangle3_weights[1482]), .FEAT_THRES(feature_thresholds[1482]), .FEAT_ABOVE(feature_aboves[1482]), .FEAT_BELOW(feature_belows[1482])) ac1482(.scan_win(scan_win1482), .scan_win_std_dev(scan_win_std_dev[1482]), .feature_accum(feature_accums[1482]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1483]), .RECT1_Y(rectangle1_ys[1483]), .RECT1_WIDTH(rectangle1_widths[1483]), .RECT1_HEIGHT(rectangle1_heights[1483]), .RECT1_WEIGHT(rectangle1_weights[1483]), .RECT2_X(rectangle2_xs[1483]), .RECT2_Y(rectangle2_ys[1483]), .RECT2_WIDTH(rectangle2_widths[1483]), .RECT2_HEIGHT(rectangle2_heights[1483]), .RECT2_WEIGHT(rectangle2_weights[1483]), .RECT3_X(rectangle3_xs[1483]), .RECT3_Y(rectangle3_ys[1483]), .RECT3_WIDTH(rectangle3_widths[1483]), .RECT3_HEIGHT(rectangle3_heights[1483]), .RECT3_WEIGHT(rectangle3_weights[1483]), .FEAT_THRES(feature_thresholds[1483]), .FEAT_ABOVE(feature_aboves[1483]), .FEAT_BELOW(feature_belows[1483])) ac1483(.scan_win(scan_win1483), .scan_win_std_dev(scan_win_std_dev[1483]), .feature_accum(feature_accums[1483]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1484]), .RECT1_Y(rectangle1_ys[1484]), .RECT1_WIDTH(rectangle1_widths[1484]), .RECT1_HEIGHT(rectangle1_heights[1484]), .RECT1_WEIGHT(rectangle1_weights[1484]), .RECT2_X(rectangle2_xs[1484]), .RECT2_Y(rectangle2_ys[1484]), .RECT2_WIDTH(rectangle2_widths[1484]), .RECT2_HEIGHT(rectangle2_heights[1484]), .RECT2_WEIGHT(rectangle2_weights[1484]), .RECT3_X(rectangle3_xs[1484]), .RECT3_Y(rectangle3_ys[1484]), .RECT3_WIDTH(rectangle3_widths[1484]), .RECT3_HEIGHT(rectangle3_heights[1484]), .RECT3_WEIGHT(rectangle3_weights[1484]), .FEAT_THRES(feature_thresholds[1484]), .FEAT_ABOVE(feature_aboves[1484]), .FEAT_BELOW(feature_belows[1484])) ac1484(.scan_win(scan_win1484), .scan_win_std_dev(scan_win_std_dev[1484]), .feature_accum(feature_accums[1484]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1485]), .RECT1_Y(rectangle1_ys[1485]), .RECT1_WIDTH(rectangle1_widths[1485]), .RECT1_HEIGHT(rectangle1_heights[1485]), .RECT1_WEIGHT(rectangle1_weights[1485]), .RECT2_X(rectangle2_xs[1485]), .RECT2_Y(rectangle2_ys[1485]), .RECT2_WIDTH(rectangle2_widths[1485]), .RECT2_HEIGHT(rectangle2_heights[1485]), .RECT2_WEIGHT(rectangle2_weights[1485]), .RECT3_X(rectangle3_xs[1485]), .RECT3_Y(rectangle3_ys[1485]), .RECT3_WIDTH(rectangle3_widths[1485]), .RECT3_HEIGHT(rectangle3_heights[1485]), .RECT3_WEIGHT(rectangle3_weights[1485]), .FEAT_THRES(feature_thresholds[1485]), .FEAT_ABOVE(feature_aboves[1485]), .FEAT_BELOW(feature_belows[1485])) ac1485(.scan_win(scan_win1485), .scan_win_std_dev(scan_win_std_dev[1485]), .feature_accum(feature_accums[1485]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1486]), .RECT1_Y(rectangle1_ys[1486]), .RECT1_WIDTH(rectangle1_widths[1486]), .RECT1_HEIGHT(rectangle1_heights[1486]), .RECT1_WEIGHT(rectangle1_weights[1486]), .RECT2_X(rectangle2_xs[1486]), .RECT2_Y(rectangle2_ys[1486]), .RECT2_WIDTH(rectangle2_widths[1486]), .RECT2_HEIGHT(rectangle2_heights[1486]), .RECT2_WEIGHT(rectangle2_weights[1486]), .RECT3_X(rectangle3_xs[1486]), .RECT3_Y(rectangle3_ys[1486]), .RECT3_WIDTH(rectangle3_widths[1486]), .RECT3_HEIGHT(rectangle3_heights[1486]), .RECT3_WEIGHT(rectangle3_weights[1486]), .FEAT_THRES(feature_thresholds[1486]), .FEAT_ABOVE(feature_aboves[1486]), .FEAT_BELOW(feature_belows[1486])) ac1486(.scan_win(scan_win1486), .scan_win_std_dev(scan_win_std_dev[1486]), .feature_accum(feature_accums[1486]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1487]), .RECT1_Y(rectangle1_ys[1487]), .RECT1_WIDTH(rectangle1_widths[1487]), .RECT1_HEIGHT(rectangle1_heights[1487]), .RECT1_WEIGHT(rectangle1_weights[1487]), .RECT2_X(rectangle2_xs[1487]), .RECT2_Y(rectangle2_ys[1487]), .RECT2_WIDTH(rectangle2_widths[1487]), .RECT2_HEIGHT(rectangle2_heights[1487]), .RECT2_WEIGHT(rectangle2_weights[1487]), .RECT3_X(rectangle3_xs[1487]), .RECT3_Y(rectangle3_ys[1487]), .RECT3_WIDTH(rectangle3_widths[1487]), .RECT3_HEIGHT(rectangle3_heights[1487]), .RECT3_WEIGHT(rectangle3_weights[1487]), .FEAT_THRES(feature_thresholds[1487]), .FEAT_ABOVE(feature_aboves[1487]), .FEAT_BELOW(feature_belows[1487])) ac1487(.scan_win(scan_win1487), .scan_win_std_dev(scan_win_std_dev[1487]), .feature_accum(feature_accums[1487]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1488]), .RECT1_Y(rectangle1_ys[1488]), .RECT1_WIDTH(rectangle1_widths[1488]), .RECT1_HEIGHT(rectangle1_heights[1488]), .RECT1_WEIGHT(rectangle1_weights[1488]), .RECT2_X(rectangle2_xs[1488]), .RECT2_Y(rectangle2_ys[1488]), .RECT2_WIDTH(rectangle2_widths[1488]), .RECT2_HEIGHT(rectangle2_heights[1488]), .RECT2_WEIGHT(rectangle2_weights[1488]), .RECT3_X(rectangle3_xs[1488]), .RECT3_Y(rectangle3_ys[1488]), .RECT3_WIDTH(rectangle3_widths[1488]), .RECT3_HEIGHT(rectangle3_heights[1488]), .RECT3_WEIGHT(rectangle3_weights[1488]), .FEAT_THRES(feature_thresholds[1488]), .FEAT_ABOVE(feature_aboves[1488]), .FEAT_BELOW(feature_belows[1488])) ac1488(.scan_win(scan_win1488), .scan_win_std_dev(scan_win_std_dev[1488]), .feature_accum(feature_accums[1488]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1489]), .RECT1_Y(rectangle1_ys[1489]), .RECT1_WIDTH(rectangle1_widths[1489]), .RECT1_HEIGHT(rectangle1_heights[1489]), .RECT1_WEIGHT(rectangle1_weights[1489]), .RECT2_X(rectangle2_xs[1489]), .RECT2_Y(rectangle2_ys[1489]), .RECT2_WIDTH(rectangle2_widths[1489]), .RECT2_HEIGHT(rectangle2_heights[1489]), .RECT2_WEIGHT(rectangle2_weights[1489]), .RECT3_X(rectangle3_xs[1489]), .RECT3_Y(rectangle3_ys[1489]), .RECT3_WIDTH(rectangle3_widths[1489]), .RECT3_HEIGHT(rectangle3_heights[1489]), .RECT3_WEIGHT(rectangle3_weights[1489]), .FEAT_THRES(feature_thresholds[1489]), .FEAT_ABOVE(feature_aboves[1489]), .FEAT_BELOW(feature_belows[1489])) ac1489(.scan_win(scan_win1489), .scan_win_std_dev(scan_win_std_dev[1489]), .feature_accum(feature_accums[1489]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1490]), .RECT1_Y(rectangle1_ys[1490]), .RECT1_WIDTH(rectangle1_widths[1490]), .RECT1_HEIGHT(rectangle1_heights[1490]), .RECT1_WEIGHT(rectangle1_weights[1490]), .RECT2_X(rectangle2_xs[1490]), .RECT2_Y(rectangle2_ys[1490]), .RECT2_WIDTH(rectangle2_widths[1490]), .RECT2_HEIGHT(rectangle2_heights[1490]), .RECT2_WEIGHT(rectangle2_weights[1490]), .RECT3_X(rectangle3_xs[1490]), .RECT3_Y(rectangle3_ys[1490]), .RECT3_WIDTH(rectangle3_widths[1490]), .RECT3_HEIGHT(rectangle3_heights[1490]), .RECT3_WEIGHT(rectangle3_weights[1490]), .FEAT_THRES(feature_thresholds[1490]), .FEAT_ABOVE(feature_aboves[1490]), .FEAT_BELOW(feature_belows[1490])) ac1490(.scan_win(scan_win1490), .scan_win_std_dev(scan_win_std_dev[1490]), .feature_accum(feature_accums[1490]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1491]), .RECT1_Y(rectangle1_ys[1491]), .RECT1_WIDTH(rectangle1_widths[1491]), .RECT1_HEIGHT(rectangle1_heights[1491]), .RECT1_WEIGHT(rectangle1_weights[1491]), .RECT2_X(rectangle2_xs[1491]), .RECT2_Y(rectangle2_ys[1491]), .RECT2_WIDTH(rectangle2_widths[1491]), .RECT2_HEIGHT(rectangle2_heights[1491]), .RECT2_WEIGHT(rectangle2_weights[1491]), .RECT3_X(rectangle3_xs[1491]), .RECT3_Y(rectangle3_ys[1491]), .RECT3_WIDTH(rectangle3_widths[1491]), .RECT3_HEIGHT(rectangle3_heights[1491]), .RECT3_WEIGHT(rectangle3_weights[1491]), .FEAT_THRES(feature_thresholds[1491]), .FEAT_ABOVE(feature_aboves[1491]), .FEAT_BELOW(feature_belows[1491])) ac1491(.scan_win(scan_win1491), .scan_win_std_dev(scan_win_std_dev[1491]), .feature_accum(feature_accums[1491]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1492]), .RECT1_Y(rectangle1_ys[1492]), .RECT1_WIDTH(rectangle1_widths[1492]), .RECT1_HEIGHT(rectangle1_heights[1492]), .RECT1_WEIGHT(rectangle1_weights[1492]), .RECT2_X(rectangle2_xs[1492]), .RECT2_Y(rectangle2_ys[1492]), .RECT2_WIDTH(rectangle2_widths[1492]), .RECT2_HEIGHT(rectangle2_heights[1492]), .RECT2_WEIGHT(rectangle2_weights[1492]), .RECT3_X(rectangle3_xs[1492]), .RECT3_Y(rectangle3_ys[1492]), .RECT3_WIDTH(rectangle3_widths[1492]), .RECT3_HEIGHT(rectangle3_heights[1492]), .RECT3_WEIGHT(rectangle3_weights[1492]), .FEAT_THRES(feature_thresholds[1492]), .FEAT_ABOVE(feature_aboves[1492]), .FEAT_BELOW(feature_belows[1492])) ac1492(.scan_win(scan_win1492), .scan_win_std_dev(scan_win_std_dev[1492]), .feature_accum(feature_accums[1492]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1493]), .RECT1_Y(rectangle1_ys[1493]), .RECT1_WIDTH(rectangle1_widths[1493]), .RECT1_HEIGHT(rectangle1_heights[1493]), .RECT1_WEIGHT(rectangle1_weights[1493]), .RECT2_X(rectangle2_xs[1493]), .RECT2_Y(rectangle2_ys[1493]), .RECT2_WIDTH(rectangle2_widths[1493]), .RECT2_HEIGHT(rectangle2_heights[1493]), .RECT2_WEIGHT(rectangle2_weights[1493]), .RECT3_X(rectangle3_xs[1493]), .RECT3_Y(rectangle3_ys[1493]), .RECT3_WIDTH(rectangle3_widths[1493]), .RECT3_HEIGHT(rectangle3_heights[1493]), .RECT3_WEIGHT(rectangle3_weights[1493]), .FEAT_THRES(feature_thresholds[1493]), .FEAT_ABOVE(feature_aboves[1493]), .FEAT_BELOW(feature_belows[1493])) ac1493(.scan_win(scan_win1493), .scan_win_std_dev(scan_win_std_dev[1493]), .feature_accum(feature_accums[1493]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1494]), .RECT1_Y(rectangle1_ys[1494]), .RECT1_WIDTH(rectangle1_widths[1494]), .RECT1_HEIGHT(rectangle1_heights[1494]), .RECT1_WEIGHT(rectangle1_weights[1494]), .RECT2_X(rectangle2_xs[1494]), .RECT2_Y(rectangle2_ys[1494]), .RECT2_WIDTH(rectangle2_widths[1494]), .RECT2_HEIGHT(rectangle2_heights[1494]), .RECT2_WEIGHT(rectangle2_weights[1494]), .RECT3_X(rectangle3_xs[1494]), .RECT3_Y(rectangle3_ys[1494]), .RECT3_WIDTH(rectangle3_widths[1494]), .RECT3_HEIGHT(rectangle3_heights[1494]), .RECT3_WEIGHT(rectangle3_weights[1494]), .FEAT_THRES(feature_thresholds[1494]), .FEAT_ABOVE(feature_aboves[1494]), .FEAT_BELOW(feature_belows[1494])) ac1494(.scan_win(scan_win1494), .scan_win_std_dev(scan_win_std_dev[1494]), .feature_accum(feature_accums[1494]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1495]), .RECT1_Y(rectangle1_ys[1495]), .RECT1_WIDTH(rectangle1_widths[1495]), .RECT1_HEIGHT(rectangle1_heights[1495]), .RECT1_WEIGHT(rectangle1_weights[1495]), .RECT2_X(rectangle2_xs[1495]), .RECT2_Y(rectangle2_ys[1495]), .RECT2_WIDTH(rectangle2_widths[1495]), .RECT2_HEIGHT(rectangle2_heights[1495]), .RECT2_WEIGHT(rectangle2_weights[1495]), .RECT3_X(rectangle3_xs[1495]), .RECT3_Y(rectangle3_ys[1495]), .RECT3_WIDTH(rectangle3_widths[1495]), .RECT3_HEIGHT(rectangle3_heights[1495]), .RECT3_WEIGHT(rectangle3_weights[1495]), .FEAT_THRES(feature_thresholds[1495]), .FEAT_ABOVE(feature_aboves[1495]), .FEAT_BELOW(feature_belows[1495])) ac1495(.scan_win(scan_win1495), .scan_win_std_dev(scan_win_std_dev[1495]), .feature_accum(feature_accums[1495]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1496]), .RECT1_Y(rectangle1_ys[1496]), .RECT1_WIDTH(rectangle1_widths[1496]), .RECT1_HEIGHT(rectangle1_heights[1496]), .RECT1_WEIGHT(rectangle1_weights[1496]), .RECT2_X(rectangle2_xs[1496]), .RECT2_Y(rectangle2_ys[1496]), .RECT2_WIDTH(rectangle2_widths[1496]), .RECT2_HEIGHT(rectangle2_heights[1496]), .RECT2_WEIGHT(rectangle2_weights[1496]), .RECT3_X(rectangle3_xs[1496]), .RECT3_Y(rectangle3_ys[1496]), .RECT3_WIDTH(rectangle3_widths[1496]), .RECT3_HEIGHT(rectangle3_heights[1496]), .RECT3_WEIGHT(rectangle3_weights[1496]), .FEAT_THRES(feature_thresholds[1496]), .FEAT_ABOVE(feature_aboves[1496]), .FEAT_BELOW(feature_belows[1496])) ac1496(.scan_win(scan_win1496), .scan_win_std_dev(scan_win_std_dev[1496]), .feature_accum(feature_accums[1496]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1497]), .RECT1_Y(rectangle1_ys[1497]), .RECT1_WIDTH(rectangle1_widths[1497]), .RECT1_HEIGHT(rectangle1_heights[1497]), .RECT1_WEIGHT(rectangle1_weights[1497]), .RECT2_X(rectangle2_xs[1497]), .RECT2_Y(rectangle2_ys[1497]), .RECT2_WIDTH(rectangle2_widths[1497]), .RECT2_HEIGHT(rectangle2_heights[1497]), .RECT2_WEIGHT(rectangle2_weights[1497]), .RECT3_X(rectangle3_xs[1497]), .RECT3_Y(rectangle3_ys[1497]), .RECT3_WIDTH(rectangle3_widths[1497]), .RECT3_HEIGHT(rectangle3_heights[1497]), .RECT3_WEIGHT(rectangle3_weights[1497]), .FEAT_THRES(feature_thresholds[1497]), .FEAT_ABOVE(feature_aboves[1497]), .FEAT_BELOW(feature_belows[1497])) ac1497(.scan_win(scan_win1497), .scan_win_std_dev(scan_win_std_dev[1497]), .feature_accum(feature_accums[1497]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1498]), .RECT1_Y(rectangle1_ys[1498]), .RECT1_WIDTH(rectangle1_widths[1498]), .RECT1_HEIGHT(rectangle1_heights[1498]), .RECT1_WEIGHT(rectangle1_weights[1498]), .RECT2_X(rectangle2_xs[1498]), .RECT2_Y(rectangle2_ys[1498]), .RECT2_WIDTH(rectangle2_widths[1498]), .RECT2_HEIGHT(rectangle2_heights[1498]), .RECT2_WEIGHT(rectangle2_weights[1498]), .RECT3_X(rectangle3_xs[1498]), .RECT3_Y(rectangle3_ys[1498]), .RECT3_WIDTH(rectangle3_widths[1498]), .RECT3_HEIGHT(rectangle3_heights[1498]), .RECT3_WEIGHT(rectangle3_weights[1498]), .FEAT_THRES(feature_thresholds[1498]), .FEAT_ABOVE(feature_aboves[1498]), .FEAT_BELOW(feature_belows[1498])) ac1498(.scan_win(scan_win1498), .scan_win_std_dev(scan_win_std_dev[1498]), .feature_accum(feature_accums[1498]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1499]), .RECT1_Y(rectangle1_ys[1499]), .RECT1_WIDTH(rectangle1_widths[1499]), .RECT1_HEIGHT(rectangle1_heights[1499]), .RECT1_WEIGHT(rectangle1_weights[1499]), .RECT2_X(rectangle2_xs[1499]), .RECT2_Y(rectangle2_ys[1499]), .RECT2_WIDTH(rectangle2_widths[1499]), .RECT2_HEIGHT(rectangle2_heights[1499]), .RECT2_WEIGHT(rectangle2_weights[1499]), .RECT3_X(rectangle3_xs[1499]), .RECT3_Y(rectangle3_ys[1499]), .RECT3_WIDTH(rectangle3_widths[1499]), .RECT3_HEIGHT(rectangle3_heights[1499]), .RECT3_WEIGHT(rectangle3_weights[1499]), .FEAT_THRES(feature_thresholds[1499]), .FEAT_ABOVE(feature_aboves[1499]), .FEAT_BELOW(feature_belows[1499])) ac1499(.scan_win(scan_win1499), .scan_win_std_dev(scan_win_std_dev[1499]), .feature_accum(feature_accums[1499]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1500]), .RECT1_Y(rectangle1_ys[1500]), .RECT1_WIDTH(rectangle1_widths[1500]), .RECT1_HEIGHT(rectangle1_heights[1500]), .RECT1_WEIGHT(rectangle1_weights[1500]), .RECT2_X(rectangle2_xs[1500]), .RECT2_Y(rectangle2_ys[1500]), .RECT2_WIDTH(rectangle2_widths[1500]), .RECT2_HEIGHT(rectangle2_heights[1500]), .RECT2_WEIGHT(rectangle2_weights[1500]), .RECT3_X(rectangle3_xs[1500]), .RECT3_Y(rectangle3_ys[1500]), .RECT3_WIDTH(rectangle3_widths[1500]), .RECT3_HEIGHT(rectangle3_heights[1500]), .RECT3_WEIGHT(rectangle3_weights[1500]), .FEAT_THRES(feature_thresholds[1500]), .FEAT_ABOVE(feature_aboves[1500]), .FEAT_BELOW(feature_belows[1500])) ac1500(.scan_win(scan_win1500), .scan_win_std_dev(scan_win_std_dev[1500]), .feature_accum(feature_accums[1500]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1501]), .RECT1_Y(rectangle1_ys[1501]), .RECT1_WIDTH(rectangle1_widths[1501]), .RECT1_HEIGHT(rectangle1_heights[1501]), .RECT1_WEIGHT(rectangle1_weights[1501]), .RECT2_X(rectangle2_xs[1501]), .RECT2_Y(rectangle2_ys[1501]), .RECT2_WIDTH(rectangle2_widths[1501]), .RECT2_HEIGHT(rectangle2_heights[1501]), .RECT2_WEIGHT(rectangle2_weights[1501]), .RECT3_X(rectangle3_xs[1501]), .RECT3_Y(rectangle3_ys[1501]), .RECT3_WIDTH(rectangle3_widths[1501]), .RECT3_HEIGHT(rectangle3_heights[1501]), .RECT3_WEIGHT(rectangle3_weights[1501]), .FEAT_THRES(feature_thresholds[1501]), .FEAT_ABOVE(feature_aboves[1501]), .FEAT_BELOW(feature_belows[1501])) ac1501(.scan_win(scan_win1501), .scan_win_std_dev(scan_win_std_dev[1501]), .feature_accum(feature_accums[1501]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1502]), .RECT1_Y(rectangle1_ys[1502]), .RECT1_WIDTH(rectangle1_widths[1502]), .RECT1_HEIGHT(rectangle1_heights[1502]), .RECT1_WEIGHT(rectangle1_weights[1502]), .RECT2_X(rectangle2_xs[1502]), .RECT2_Y(rectangle2_ys[1502]), .RECT2_WIDTH(rectangle2_widths[1502]), .RECT2_HEIGHT(rectangle2_heights[1502]), .RECT2_WEIGHT(rectangle2_weights[1502]), .RECT3_X(rectangle3_xs[1502]), .RECT3_Y(rectangle3_ys[1502]), .RECT3_WIDTH(rectangle3_widths[1502]), .RECT3_HEIGHT(rectangle3_heights[1502]), .RECT3_WEIGHT(rectangle3_weights[1502]), .FEAT_THRES(feature_thresholds[1502]), .FEAT_ABOVE(feature_aboves[1502]), .FEAT_BELOW(feature_belows[1502])) ac1502(.scan_win(scan_win1502), .scan_win_std_dev(scan_win_std_dev[1502]), .feature_accum(feature_accums[1502]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1503]), .RECT1_Y(rectangle1_ys[1503]), .RECT1_WIDTH(rectangle1_widths[1503]), .RECT1_HEIGHT(rectangle1_heights[1503]), .RECT1_WEIGHT(rectangle1_weights[1503]), .RECT2_X(rectangle2_xs[1503]), .RECT2_Y(rectangle2_ys[1503]), .RECT2_WIDTH(rectangle2_widths[1503]), .RECT2_HEIGHT(rectangle2_heights[1503]), .RECT2_WEIGHT(rectangle2_weights[1503]), .RECT3_X(rectangle3_xs[1503]), .RECT3_Y(rectangle3_ys[1503]), .RECT3_WIDTH(rectangle3_widths[1503]), .RECT3_HEIGHT(rectangle3_heights[1503]), .RECT3_WEIGHT(rectangle3_weights[1503]), .FEAT_THRES(feature_thresholds[1503]), .FEAT_ABOVE(feature_aboves[1503]), .FEAT_BELOW(feature_belows[1503])) ac1503(.scan_win(scan_win1503), .scan_win_std_dev(scan_win_std_dev[1503]), .feature_accum(feature_accums[1503]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1504]), .RECT1_Y(rectangle1_ys[1504]), .RECT1_WIDTH(rectangle1_widths[1504]), .RECT1_HEIGHT(rectangle1_heights[1504]), .RECT1_WEIGHT(rectangle1_weights[1504]), .RECT2_X(rectangle2_xs[1504]), .RECT2_Y(rectangle2_ys[1504]), .RECT2_WIDTH(rectangle2_widths[1504]), .RECT2_HEIGHT(rectangle2_heights[1504]), .RECT2_WEIGHT(rectangle2_weights[1504]), .RECT3_X(rectangle3_xs[1504]), .RECT3_Y(rectangle3_ys[1504]), .RECT3_WIDTH(rectangle3_widths[1504]), .RECT3_HEIGHT(rectangle3_heights[1504]), .RECT3_WEIGHT(rectangle3_weights[1504]), .FEAT_THRES(feature_thresholds[1504]), .FEAT_ABOVE(feature_aboves[1504]), .FEAT_BELOW(feature_belows[1504])) ac1504(.scan_win(scan_win1504), .scan_win_std_dev(scan_win_std_dev[1504]), .feature_accum(feature_accums[1504]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1505]), .RECT1_Y(rectangle1_ys[1505]), .RECT1_WIDTH(rectangle1_widths[1505]), .RECT1_HEIGHT(rectangle1_heights[1505]), .RECT1_WEIGHT(rectangle1_weights[1505]), .RECT2_X(rectangle2_xs[1505]), .RECT2_Y(rectangle2_ys[1505]), .RECT2_WIDTH(rectangle2_widths[1505]), .RECT2_HEIGHT(rectangle2_heights[1505]), .RECT2_WEIGHT(rectangle2_weights[1505]), .RECT3_X(rectangle3_xs[1505]), .RECT3_Y(rectangle3_ys[1505]), .RECT3_WIDTH(rectangle3_widths[1505]), .RECT3_HEIGHT(rectangle3_heights[1505]), .RECT3_WEIGHT(rectangle3_weights[1505]), .FEAT_THRES(feature_thresholds[1505]), .FEAT_ABOVE(feature_aboves[1505]), .FEAT_BELOW(feature_belows[1505])) ac1505(.scan_win(scan_win1505), .scan_win_std_dev(scan_win_std_dev[1505]), .feature_accum(feature_accums[1505]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1506]), .RECT1_Y(rectangle1_ys[1506]), .RECT1_WIDTH(rectangle1_widths[1506]), .RECT1_HEIGHT(rectangle1_heights[1506]), .RECT1_WEIGHT(rectangle1_weights[1506]), .RECT2_X(rectangle2_xs[1506]), .RECT2_Y(rectangle2_ys[1506]), .RECT2_WIDTH(rectangle2_widths[1506]), .RECT2_HEIGHT(rectangle2_heights[1506]), .RECT2_WEIGHT(rectangle2_weights[1506]), .RECT3_X(rectangle3_xs[1506]), .RECT3_Y(rectangle3_ys[1506]), .RECT3_WIDTH(rectangle3_widths[1506]), .RECT3_HEIGHT(rectangle3_heights[1506]), .RECT3_WEIGHT(rectangle3_weights[1506]), .FEAT_THRES(feature_thresholds[1506]), .FEAT_ABOVE(feature_aboves[1506]), .FEAT_BELOW(feature_belows[1506])) ac1506(.scan_win(scan_win1506), .scan_win_std_dev(scan_win_std_dev[1506]), .feature_accum(feature_accums[1506]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1507]), .RECT1_Y(rectangle1_ys[1507]), .RECT1_WIDTH(rectangle1_widths[1507]), .RECT1_HEIGHT(rectangle1_heights[1507]), .RECT1_WEIGHT(rectangle1_weights[1507]), .RECT2_X(rectangle2_xs[1507]), .RECT2_Y(rectangle2_ys[1507]), .RECT2_WIDTH(rectangle2_widths[1507]), .RECT2_HEIGHT(rectangle2_heights[1507]), .RECT2_WEIGHT(rectangle2_weights[1507]), .RECT3_X(rectangle3_xs[1507]), .RECT3_Y(rectangle3_ys[1507]), .RECT3_WIDTH(rectangle3_widths[1507]), .RECT3_HEIGHT(rectangle3_heights[1507]), .RECT3_WEIGHT(rectangle3_weights[1507]), .FEAT_THRES(feature_thresholds[1507]), .FEAT_ABOVE(feature_aboves[1507]), .FEAT_BELOW(feature_belows[1507])) ac1507(.scan_win(scan_win1507), .scan_win_std_dev(scan_win_std_dev[1507]), .feature_accum(feature_accums[1507]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1508]), .RECT1_Y(rectangle1_ys[1508]), .RECT1_WIDTH(rectangle1_widths[1508]), .RECT1_HEIGHT(rectangle1_heights[1508]), .RECT1_WEIGHT(rectangle1_weights[1508]), .RECT2_X(rectangle2_xs[1508]), .RECT2_Y(rectangle2_ys[1508]), .RECT2_WIDTH(rectangle2_widths[1508]), .RECT2_HEIGHT(rectangle2_heights[1508]), .RECT2_WEIGHT(rectangle2_weights[1508]), .RECT3_X(rectangle3_xs[1508]), .RECT3_Y(rectangle3_ys[1508]), .RECT3_WIDTH(rectangle3_widths[1508]), .RECT3_HEIGHT(rectangle3_heights[1508]), .RECT3_WEIGHT(rectangle3_weights[1508]), .FEAT_THRES(feature_thresholds[1508]), .FEAT_ABOVE(feature_aboves[1508]), .FEAT_BELOW(feature_belows[1508])) ac1508(.scan_win(scan_win1508), .scan_win_std_dev(scan_win_std_dev[1508]), .feature_accum(feature_accums[1508]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1509]), .RECT1_Y(rectangle1_ys[1509]), .RECT1_WIDTH(rectangle1_widths[1509]), .RECT1_HEIGHT(rectangle1_heights[1509]), .RECT1_WEIGHT(rectangle1_weights[1509]), .RECT2_X(rectangle2_xs[1509]), .RECT2_Y(rectangle2_ys[1509]), .RECT2_WIDTH(rectangle2_widths[1509]), .RECT2_HEIGHT(rectangle2_heights[1509]), .RECT2_WEIGHT(rectangle2_weights[1509]), .RECT3_X(rectangle3_xs[1509]), .RECT3_Y(rectangle3_ys[1509]), .RECT3_WIDTH(rectangle3_widths[1509]), .RECT3_HEIGHT(rectangle3_heights[1509]), .RECT3_WEIGHT(rectangle3_weights[1509]), .FEAT_THRES(feature_thresholds[1509]), .FEAT_ABOVE(feature_aboves[1509]), .FEAT_BELOW(feature_belows[1509])) ac1509(.scan_win(scan_win1509), .scan_win_std_dev(scan_win_std_dev[1509]), .feature_accum(feature_accums[1509]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1510]), .RECT1_Y(rectangle1_ys[1510]), .RECT1_WIDTH(rectangle1_widths[1510]), .RECT1_HEIGHT(rectangle1_heights[1510]), .RECT1_WEIGHT(rectangle1_weights[1510]), .RECT2_X(rectangle2_xs[1510]), .RECT2_Y(rectangle2_ys[1510]), .RECT2_WIDTH(rectangle2_widths[1510]), .RECT2_HEIGHT(rectangle2_heights[1510]), .RECT2_WEIGHT(rectangle2_weights[1510]), .RECT3_X(rectangle3_xs[1510]), .RECT3_Y(rectangle3_ys[1510]), .RECT3_WIDTH(rectangle3_widths[1510]), .RECT3_HEIGHT(rectangle3_heights[1510]), .RECT3_WEIGHT(rectangle3_weights[1510]), .FEAT_THRES(feature_thresholds[1510]), .FEAT_ABOVE(feature_aboves[1510]), .FEAT_BELOW(feature_belows[1510])) ac1510(.scan_win(scan_win1510), .scan_win_std_dev(scan_win_std_dev[1510]), .feature_accum(feature_accums[1510]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1511]), .RECT1_Y(rectangle1_ys[1511]), .RECT1_WIDTH(rectangle1_widths[1511]), .RECT1_HEIGHT(rectangle1_heights[1511]), .RECT1_WEIGHT(rectangle1_weights[1511]), .RECT2_X(rectangle2_xs[1511]), .RECT2_Y(rectangle2_ys[1511]), .RECT2_WIDTH(rectangle2_widths[1511]), .RECT2_HEIGHT(rectangle2_heights[1511]), .RECT2_WEIGHT(rectangle2_weights[1511]), .RECT3_X(rectangle3_xs[1511]), .RECT3_Y(rectangle3_ys[1511]), .RECT3_WIDTH(rectangle3_widths[1511]), .RECT3_HEIGHT(rectangle3_heights[1511]), .RECT3_WEIGHT(rectangle3_weights[1511]), .FEAT_THRES(feature_thresholds[1511]), .FEAT_ABOVE(feature_aboves[1511]), .FEAT_BELOW(feature_belows[1511])) ac1511(.scan_win(scan_win1511), .scan_win_std_dev(scan_win_std_dev[1511]), .feature_accum(feature_accums[1511]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1512]), .RECT1_Y(rectangle1_ys[1512]), .RECT1_WIDTH(rectangle1_widths[1512]), .RECT1_HEIGHT(rectangle1_heights[1512]), .RECT1_WEIGHT(rectangle1_weights[1512]), .RECT2_X(rectangle2_xs[1512]), .RECT2_Y(rectangle2_ys[1512]), .RECT2_WIDTH(rectangle2_widths[1512]), .RECT2_HEIGHT(rectangle2_heights[1512]), .RECT2_WEIGHT(rectangle2_weights[1512]), .RECT3_X(rectangle3_xs[1512]), .RECT3_Y(rectangle3_ys[1512]), .RECT3_WIDTH(rectangle3_widths[1512]), .RECT3_HEIGHT(rectangle3_heights[1512]), .RECT3_WEIGHT(rectangle3_weights[1512]), .FEAT_THRES(feature_thresholds[1512]), .FEAT_ABOVE(feature_aboves[1512]), .FEAT_BELOW(feature_belows[1512])) ac1512(.scan_win(scan_win1512), .scan_win_std_dev(scan_win_std_dev[1512]), .feature_accum(feature_accums[1512]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1513]), .RECT1_Y(rectangle1_ys[1513]), .RECT1_WIDTH(rectangle1_widths[1513]), .RECT1_HEIGHT(rectangle1_heights[1513]), .RECT1_WEIGHT(rectangle1_weights[1513]), .RECT2_X(rectangle2_xs[1513]), .RECT2_Y(rectangle2_ys[1513]), .RECT2_WIDTH(rectangle2_widths[1513]), .RECT2_HEIGHT(rectangle2_heights[1513]), .RECT2_WEIGHT(rectangle2_weights[1513]), .RECT3_X(rectangle3_xs[1513]), .RECT3_Y(rectangle3_ys[1513]), .RECT3_WIDTH(rectangle3_widths[1513]), .RECT3_HEIGHT(rectangle3_heights[1513]), .RECT3_WEIGHT(rectangle3_weights[1513]), .FEAT_THRES(feature_thresholds[1513]), .FEAT_ABOVE(feature_aboves[1513]), .FEAT_BELOW(feature_belows[1513])) ac1513(.scan_win(scan_win1513), .scan_win_std_dev(scan_win_std_dev[1513]), .feature_accum(feature_accums[1513]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1514]), .RECT1_Y(rectangle1_ys[1514]), .RECT1_WIDTH(rectangle1_widths[1514]), .RECT1_HEIGHT(rectangle1_heights[1514]), .RECT1_WEIGHT(rectangle1_weights[1514]), .RECT2_X(rectangle2_xs[1514]), .RECT2_Y(rectangle2_ys[1514]), .RECT2_WIDTH(rectangle2_widths[1514]), .RECT2_HEIGHT(rectangle2_heights[1514]), .RECT2_WEIGHT(rectangle2_weights[1514]), .RECT3_X(rectangle3_xs[1514]), .RECT3_Y(rectangle3_ys[1514]), .RECT3_WIDTH(rectangle3_widths[1514]), .RECT3_HEIGHT(rectangle3_heights[1514]), .RECT3_WEIGHT(rectangle3_weights[1514]), .FEAT_THRES(feature_thresholds[1514]), .FEAT_ABOVE(feature_aboves[1514]), .FEAT_BELOW(feature_belows[1514])) ac1514(.scan_win(scan_win1514), .scan_win_std_dev(scan_win_std_dev[1514]), .feature_accum(feature_accums[1514]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1515]), .RECT1_Y(rectangle1_ys[1515]), .RECT1_WIDTH(rectangle1_widths[1515]), .RECT1_HEIGHT(rectangle1_heights[1515]), .RECT1_WEIGHT(rectangle1_weights[1515]), .RECT2_X(rectangle2_xs[1515]), .RECT2_Y(rectangle2_ys[1515]), .RECT2_WIDTH(rectangle2_widths[1515]), .RECT2_HEIGHT(rectangle2_heights[1515]), .RECT2_WEIGHT(rectangle2_weights[1515]), .RECT3_X(rectangle3_xs[1515]), .RECT3_Y(rectangle3_ys[1515]), .RECT3_WIDTH(rectangle3_widths[1515]), .RECT3_HEIGHT(rectangle3_heights[1515]), .RECT3_WEIGHT(rectangle3_weights[1515]), .FEAT_THRES(feature_thresholds[1515]), .FEAT_ABOVE(feature_aboves[1515]), .FEAT_BELOW(feature_belows[1515])) ac1515(.scan_win(scan_win1515), .scan_win_std_dev(scan_win_std_dev[1515]), .feature_accum(feature_accums[1515]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1516]), .RECT1_Y(rectangle1_ys[1516]), .RECT1_WIDTH(rectangle1_widths[1516]), .RECT1_HEIGHT(rectangle1_heights[1516]), .RECT1_WEIGHT(rectangle1_weights[1516]), .RECT2_X(rectangle2_xs[1516]), .RECT2_Y(rectangle2_ys[1516]), .RECT2_WIDTH(rectangle2_widths[1516]), .RECT2_HEIGHT(rectangle2_heights[1516]), .RECT2_WEIGHT(rectangle2_weights[1516]), .RECT3_X(rectangle3_xs[1516]), .RECT3_Y(rectangle3_ys[1516]), .RECT3_WIDTH(rectangle3_widths[1516]), .RECT3_HEIGHT(rectangle3_heights[1516]), .RECT3_WEIGHT(rectangle3_weights[1516]), .FEAT_THRES(feature_thresholds[1516]), .FEAT_ABOVE(feature_aboves[1516]), .FEAT_BELOW(feature_belows[1516])) ac1516(.scan_win(scan_win1516), .scan_win_std_dev(scan_win_std_dev[1516]), .feature_accum(feature_accums[1516]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1517]), .RECT1_Y(rectangle1_ys[1517]), .RECT1_WIDTH(rectangle1_widths[1517]), .RECT1_HEIGHT(rectangle1_heights[1517]), .RECT1_WEIGHT(rectangle1_weights[1517]), .RECT2_X(rectangle2_xs[1517]), .RECT2_Y(rectangle2_ys[1517]), .RECT2_WIDTH(rectangle2_widths[1517]), .RECT2_HEIGHT(rectangle2_heights[1517]), .RECT2_WEIGHT(rectangle2_weights[1517]), .RECT3_X(rectangle3_xs[1517]), .RECT3_Y(rectangle3_ys[1517]), .RECT3_WIDTH(rectangle3_widths[1517]), .RECT3_HEIGHT(rectangle3_heights[1517]), .RECT3_WEIGHT(rectangle3_weights[1517]), .FEAT_THRES(feature_thresholds[1517]), .FEAT_ABOVE(feature_aboves[1517]), .FEAT_BELOW(feature_belows[1517])) ac1517(.scan_win(scan_win1517), .scan_win_std_dev(scan_win_std_dev[1517]), .feature_accum(feature_accums[1517]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1518]), .RECT1_Y(rectangle1_ys[1518]), .RECT1_WIDTH(rectangle1_widths[1518]), .RECT1_HEIGHT(rectangle1_heights[1518]), .RECT1_WEIGHT(rectangle1_weights[1518]), .RECT2_X(rectangle2_xs[1518]), .RECT2_Y(rectangle2_ys[1518]), .RECT2_WIDTH(rectangle2_widths[1518]), .RECT2_HEIGHT(rectangle2_heights[1518]), .RECT2_WEIGHT(rectangle2_weights[1518]), .RECT3_X(rectangle3_xs[1518]), .RECT3_Y(rectangle3_ys[1518]), .RECT3_WIDTH(rectangle3_widths[1518]), .RECT3_HEIGHT(rectangle3_heights[1518]), .RECT3_WEIGHT(rectangle3_weights[1518]), .FEAT_THRES(feature_thresholds[1518]), .FEAT_ABOVE(feature_aboves[1518]), .FEAT_BELOW(feature_belows[1518])) ac1518(.scan_win(scan_win1518), .scan_win_std_dev(scan_win_std_dev[1518]), .feature_accum(feature_accums[1518]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1519]), .RECT1_Y(rectangle1_ys[1519]), .RECT1_WIDTH(rectangle1_widths[1519]), .RECT1_HEIGHT(rectangle1_heights[1519]), .RECT1_WEIGHT(rectangle1_weights[1519]), .RECT2_X(rectangle2_xs[1519]), .RECT2_Y(rectangle2_ys[1519]), .RECT2_WIDTH(rectangle2_widths[1519]), .RECT2_HEIGHT(rectangle2_heights[1519]), .RECT2_WEIGHT(rectangle2_weights[1519]), .RECT3_X(rectangle3_xs[1519]), .RECT3_Y(rectangle3_ys[1519]), .RECT3_WIDTH(rectangle3_widths[1519]), .RECT3_HEIGHT(rectangle3_heights[1519]), .RECT3_WEIGHT(rectangle3_weights[1519]), .FEAT_THRES(feature_thresholds[1519]), .FEAT_ABOVE(feature_aboves[1519]), .FEAT_BELOW(feature_belows[1519])) ac1519(.scan_win(scan_win1519), .scan_win_std_dev(scan_win_std_dev[1519]), .feature_accum(feature_accums[1519]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1520]), .RECT1_Y(rectangle1_ys[1520]), .RECT1_WIDTH(rectangle1_widths[1520]), .RECT1_HEIGHT(rectangle1_heights[1520]), .RECT1_WEIGHT(rectangle1_weights[1520]), .RECT2_X(rectangle2_xs[1520]), .RECT2_Y(rectangle2_ys[1520]), .RECT2_WIDTH(rectangle2_widths[1520]), .RECT2_HEIGHT(rectangle2_heights[1520]), .RECT2_WEIGHT(rectangle2_weights[1520]), .RECT3_X(rectangle3_xs[1520]), .RECT3_Y(rectangle3_ys[1520]), .RECT3_WIDTH(rectangle3_widths[1520]), .RECT3_HEIGHT(rectangle3_heights[1520]), .RECT3_WEIGHT(rectangle3_weights[1520]), .FEAT_THRES(feature_thresholds[1520]), .FEAT_ABOVE(feature_aboves[1520]), .FEAT_BELOW(feature_belows[1520])) ac1520(.scan_win(scan_win1520), .scan_win_std_dev(scan_win_std_dev[1520]), .feature_accum(feature_accums[1520]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1521]), .RECT1_Y(rectangle1_ys[1521]), .RECT1_WIDTH(rectangle1_widths[1521]), .RECT1_HEIGHT(rectangle1_heights[1521]), .RECT1_WEIGHT(rectangle1_weights[1521]), .RECT2_X(rectangle2_xs[1521]), .RECT2_Y(rectangle2_ys[1521]), .RECT2_WIDTH(rectangle2_widths[1521]), .RECT2_HEIGHT(rectangle2_heights[1521]), .RECT2_WEIGHT(rectangle2_weights[1521]), .RECT3_X(rectangle3_xs[1521]), .RECT3_Y(rectangle3_ys[1521]), .RECT3_WIDTH(rectangle3_widths[1521]), .RECT3_HEIGHT(rectangle3_heights[1521]), .RECT3_WEIGHT(rectangle3_weights[1521]), .FEAT_THRES(feature_thresholds[1521]), .FEAT_ABOVE(feature_aboves[1521]), .FEAT_BELOW(feature_belows[1521])) ac1521(.scan_win(scan_win1521), .scan_win_std_dev(scan_win_std_dev[1521]), .feature_accum(feature_accums[1521]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1522]), .RECT1_Y(rectangle1_ys[1522]), .RECT1_WIDTH(rectangle1_widths[1522]), .RECT1_HEIGHT(rectangle1_heights[1522]), .RECT1_WEIGHT(rectangle1_weights[1522]), .RECT2_X(rectangle2_xs[1522]), .RECT2_Y(rectangle2_ys[1522]), .RECT2_WIDTH(rectangle2_widths[1522]), .RECT2_HEIGHT(rectangle2_heights[1522]), .RECT2_WEIGHT(rectangle2_weights[1522]), .RECT3_X(rectangle3_xs[1522]), .RECT3_Y(rectangle3_ys[1522]), .RECT3_WIDTH(rectangle3_widths[1522]), .RECT3_HEIGHT(rectangle3_heights[1522]), .RECT3_WEIGHT(rectangle3_weights[1522]), .FEAT_THRES(feature_thresholds[1522]), .FEAT_ABOVE(feature_aboves[1522]), .FEAT_BELOW(feature_belows[1522])) ac1522(.scan_win(scan_win1522), .scan_win_std_dev(scan_win_std_dev[1522]), .feature_accum(feature_accums[1522]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1523]), .RECT1_Y(rectangle1_ys[1523]), .RECT1_WIDTH(rectangle1_widths[1523]), .RECT1_HEIGHT(rectangle1_heights[1523]), .RECT1_WEIGHT(rectangle1_weights[1523]), .RECT2_X(rectangle2_xs[1523]), .RECT2_Y(rectangle2_ys[1523]), .RECT2_WIDTH(rectangle2_widths[1523]), .RECT2_HEIGHT(rectangle2_heights[1523]), .RECT2_WEIGHT(rectangle2_weights[1523]), .RECT3_X(rectangle3_xs[1523]), .RECT3_Y(rectangle3_ys[1523]), .RECT3_WIDTH(rectangle3_widths[1523]), .RECT3_HEIGHT(rectangle3_heights[1523]), .RECT3_WEIGHT(rectangle3_weights[1523]), .FEAT_THRES(feature_thresholds[1523]), .FEAT_ABOVE(feature_aboves[1523]), .FEAT_BELOW(feature_belows[1523])) ac1523(.scan_win(scan_win1523), .scan_win_std_dev(scan_win_std_dev[1523]), .feature_accum(feature_accums[1523]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1524]), .RECT1_Y(rectangle1_ys[1524]), .RECT1_WIDTH(rectangle1_widths[1524]), .RECT1_HEIGHT(rectangle1_heights[1524]), .RECT1_WEIGHT(rectangle1_weights[1524]), .RECT2_X(rectangle2_xs[1524]), .RECT2_Y(rectangle2_ys[1524]), .RECT2_WIDTH(rectangle2_widths[1524]), .RECT2_HEIGHT(rectangle2_heights[1524]), .RECT2_WEIGHT(rectangle2_weights[1524]), .RECT3_X(rectangle3_xs[1524]), .RECT3_Y(rectangle3_ys[1524]), .RECT3_WIDTH(rectangle3_widths[1524]), .RECT3_HEIGHT(rectangle3_heights[1524]), .RECT3_WEIGHT(rectangle3_weights[1524]), .FEAT_THRES(feature_thresholds[1524]), .FEAT_ABOVE(feature_aboves[1524]), .FEAT_BELOW(feature_belows[1524])) ac1524(.scan_win(scan_win1524), .scan_win_std_dev(scan_win_std_dev[1524]), .feature_accum(feature_accums[1524]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1525]), .RECT1_Y(rectangle1_ys[1525]), .RECT1_WIDTH(rectangle1_widths[1525]), .RECT1_HEIGHT(rectangle1_heights[1525]), .RECT1_WEIGHT(rectangle1_weights[1525]), .RECT2_X(rectangle2_xs[1525]), .RECT2_Y(rectangle2_ys[1525]), .RECT2_WIDTH(rectangle2_widths[1525]), .RECT2_HEIGHT(rectangle2_heights[1525]), .RECT2_WEIGHT(rectangle2_weights[1525]), .RECT3_X(rectangle3_xs[1525]), .RECT3_Y(rectangle3_ys[1525]), .RECT3_WIDTH(rectangle3_widths[1525]), .RECT3_HEIGHT(rectangle3_heights[1525]), .RECT3_WEIGHT(rectangle3_weights[1525]), .FEAT_THRES(feature_thresholds[1525]), .FEAT_ABOVE(feature_aboves[1525]), .FEAT_BELOW(feature_belows[1525])) ac1525(.scan_win(scan_win1525), .scan_win_std_dev(scan_win_std_dev[1525]), .feature_accum(feature_accums[1525]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1526]), .RECT1_Y(rectangle1_ys[1526]), .RECT1_WIDTH(rectangle1_widths[1526]), .RECT1_HEIGHT(rectangle1_heights[1526]), .RECT1_WEIGHT(rectangle1_weights[1526]), .RECT2_X(rectangle2_xs[1526]), .RECT2_Y(rectangle2_ys[1526]), .RECT2_WIDTH(rectangle2_widths[1526]), .RECT2_HEIGHT(rectangle2_heights[1526]), .RECT2_WEIGHT(rectangle2_weights[1526]), .RECT3_X(rectangle3_xs[1526]), .RECT3_Y(rectangle3_ys[1526]), .RECT3_WIDTH(rectangle3_widths[1526]), .RECT3_HEIGHT(rectangle3_heights[1526]), .RECT3_WEIGHT(rectangle3_weights[1526]), .FEAT_THRES(feature_thresholds[1526]), .FEAT_ABOVE(feature_aboves[1526]), .FEAT_BELOW(feature_belows[1526])) ac1526(.scan_win(scan_win1526), .scan_win_std_dev(scan_win_std_dev[1526]), .feature_accum(feature_accums[1526]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1527]), .RECT1_Y(rectangle1_ys[1527]), .RECT1_WIDTH(rectangle1_widths[1527]), .RECT1_HEIGHT(rectangle1_heights[1527]), .RECT1_WEIGHT(rectangle1_weights[1527]), .RECT2_X(rectangle2_xs[1527]), .RECT2_Y(rectangle2_ys[1527]), .RECT2_WIDTH(rectangle2_widths[1527]), .RECT2_HEIGHT(rectangle2_heights[1527]), .RECT2_WEIGHT(rectangle2_weights[1527]), .RECT3_X(rectangle3_xs[1527]), .RECT3_Y(rectangle3_ys[1527]), .RECT3_WIDTH(rectangle3_widths[1527]), .RECT3_HEIGHT(rectangle3_heights[1527]), .RECT3_WEIGHT(rectangle3_weights[1527]), .FEAT_THRES(feature_thresholds[1527]), .FEAT_ABOVE(feature_aboves[1527]), .FEAT_BELOW(feature_belows[1527])) ac1527(.scan_win(scan_win1527), .scan_win_std_dev(scan_win_std_dev[1527]), .feature_accum(feature_accums[1527]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1528]), .RECT1_Y(rectangle1_ys[1528]), .RECT1_WIDTH(rectangle1_widths[1528]), .RECT1_HEIGHT(rectangle1_heights[1528]), .RECT1_WEIGHT(rectangle1_weights[1528]), .RECT2_X(rectangle2_xs[1528]), .RECT2_Y(rectangle2_ys[1528]), .RECT2_WIDTH(rectangle2_widths[1528]), .RECT2_HEIGHT(rectangle2_heights[1528]), .RECT2_WEIGHT(rectangle2_weights[1528]), .RECT3_X(rectangle3_xs[1528]), .RECT3_Y(rectangle3_ys[1528]), .RECT3_WIDTH(rectangle3_widths[1528]), .RECT3_HEIGHT(rectangle3_heights[1528]), .RECT3_WEIGHT(rectangle3_weights[1528]), .FEAT_THRES(feature_thresholds[1528]), .FEAT_ABOVE(feature_aboves[1528]), .FEAT_BELOW(feature_belows[1528])) ac1528(.scan_win(scan_win1528), .scan_win_std_dev(scan_win_std_dev[1528]), .feature_accum(feature_accums[1528]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1529]), .RECT1_Y(rectangle1_ys[1529]), .RECT1_WIDTH(rectangle1_widths[1529]), .RECT1_HEIGHT(rectangle1_heights[1529]), .RECT1_WEIGHT(rectangle1_weights[1529]), .RECT2_X(rectangle2_xs[1529]), .RECT2_Y(rectangle2_ys[1529]), .RECT2_WIDTH(rectangle2_widths[1529]), .RECT2_HEIGHT(rectangle2_heights[1529]), .RECT2_WEIGHT(rectangle2_weights[1529]), .RECT3_X(rectangle3_xs[1529]), .RECT3_Y(rectangle3_ys[1529]), .RECT3_WIDTH(rectangle3_widths[1529]), .RECT3_HEIGHT(rectangle3_heights[1529]), .RECT3_WEIGHT(rectangle3_weights[1529]), .FEAT_THRES(feature_thresholds[1529]), .FEAT_ABOVE(feature_aboves[1529]), .FEAT_BELOW(feature_belows[1529])) ac1529(.scan_win(scan_win1529), .scan_win_std_dev(scan_win_std_dev[1529]), .feature_accum(feature_accums[1529]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1530]), .RECT1_Y(rectangle1_ys[1530]), .RECT1_WIDTH(rectangle1_widths[1530]), .RECT1_HEIGHT(rectangle1_heights[1530]), .RECT1_WEIGHT(rectangle1_weights[1530]), .RECT2_X(rectangle2_xs[1530]), .RECT2_Y(rectangle2_ys[1530]), .RECT2_WIDTH(rectangle2_widths[1530]), .RECT2_HEIGHT(rectangle2_heights[1530]), .RECT2_WEIGHT(rectangle2_weights[1530]), .RECT3_X(rectangle3_xs[1530]), .RECT3_Y(rectangle3_ys[1530]), .RECT3_WIDTH(rectangle3_widths[1530]), .RECT3_HEIGHT(rectangle3_heights[1530]), .RECT3_WEIGHT(rectangle3_weights[1530]), .FEAT_THRES(feature_thresholds[1530]), .FEAT_ABOVE(feature_aboves[1530]), .FEAT_BELOW(feature_belows[1530])) ac1530(.scan_win(scan_win1530), .scan_win_std_dev(scan_win_std_dev[1530]), .feature_accum(feature_accums[1530]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1531]), .RECT1_Y(rectangle1_ys[1531]), .RECT1_WIDTH(rectangle1_widths[1531]), .RECT1_HEIGHT(rectangle1_heights[1531]), .RECT1_WEIGHT(rectangle1_weights[1531]), .RECT2_X(rectangle2_xs[1531]), .RECT2_Y(rectangle2_ys[1531]), .RECT2_WIDTH(rectangle2_widths[1531]), .RECT2_HEIGHT(rectangle2_heights[1531]), .RECT2_WEIGHT(rectangle2_weights[1531]), .RECT3_X(rectangle3_xs[1531]), .RECT3_Y(rectangle3_ys[1531]), .RECT3_WIDTH(rectangle3_widths[1531]), .RECT3_HEIGHT(rectangle3_heights[1531]), .RECT3_WEIGHT(rectangle3_weights[1531]), .FEAT_THRES(feature_thresholds[1531]), .FEAT_ABOVE(feature_aboves[1531]), .FEAT_BELOW(feature_belows[1531])) ac1531(.scan_win(scan_win1531), .scan_win_std_dev(scan_win_std_dev[1531]), .feature_accum(feature_accums[1531]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1532]), .RECT1_Y(rectangle1_ys[1532]), .RECT1_WIDTH(rectangle1_widths[1532]), .RECT1_HEIGHT(rectangle1_heights[1532]), .RECT1_WEIGHT(rectangle1_weights[1532]), .RECT2_X(rectangle2_xs[1532]), .RECT2_Y(rectangle2_ys[1532]), .RECT2_WIDTH(rectangle2_widths[1532]), .RECT2_HEIGHT(rectangle2_heights[1532]), .RECT2_WEIGHT(rectangle2_weights[1532]), .RECT3_X(rectangle3_xs[1532]), .RECT3_Y(rectangle3_ys[1532]), .RECT3_WIDTH(rectangle3_widths[1532]), .RECT3_HEIGHT(rectangle3_heights[1532]), .RECT3_WEIGHT(rectangle3_weights[1532]), .FEAT_THRES(feature_thresholds[1532]), .FEAT_ABOVE(feature_aboves[1532]), .FEAT_BELOW(feature_belows[1532])) ac1532(.scan_win(scan_win1532), .scan_win_std_dev(scan_win_std_dev[1532]), .feature_accum(feature_accums[1532]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1533]), .RECT1_Y(rectangle1_ys[1533]), .RECT1_WIDTH(rectangle1_widths[1533]), .RECT1_HEIGHT(rectangle1_heights[1533]), .RECT1_WEIGHT(rectangle1_weights[1533]), .RECT2_X(rectangle2_xs[1533]), .RECT2_Y(rectangle2_ys[1533]), .RECT2_WIDTH(rectangle2_widths[1533]), .RECT2_HEIGHT(rectangle2_heights[1533]), .RECT2_WEIGHT(rectangle2_weights[1533]), .RECT3_X(rectangle3_xs[1533]), .RECT3_Y(rectangle3_ys[1533]), .RECT3_WIDTH(rectangle3_widths[1533]), .RECT3_HEIGHT(rectangle3_heights[1533]), .RECT3_WEIGHT(rectangle3_weights[1533]), .FEAT_THRES(feature_thresholds[1533]), .FEAT_ABOVE(feature_aboves[1533]), .FEAT_BELOW(feature_belows[1533])) ac1533(.scan_win(scan_win1533), .scan_win_std_dev(scan_win_std_dev[1533]), .feature_accum(feature_accums[1533]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1534]), .RECT1_Y(rectangle1_ys[1534]), .RECT1_WIDTH(rectangle1_widths[1534]), .RECT1_HEIGHT(rectangle1_heights[1534]), .RECT1_WEIGHT(rectangle1_weights[1534]), .RECT2_X(rectangle2_xs[1534]), .RECT2_Y(rectangle2_ys[1534]), .RECT2_WIDTH(rectangle2_widths[1534]), .RECT2_HEIGHT(rectangle2_heights[1534]), .RECT2_WEIGHT(rectangle2_weights[1534]), .RECT3_X(rectangle3_xs[1534]), .RECT3_Y(rectangle3_ys[1534]), .RECT3_WIDTH(rectangle3_widths[1534]), .RECT3_HEIGHT(rectangle3_heights[1534]), .RECT3_WEIGHT(rectangle3_weights[1534]), .FEAT_THRES(feature_thresholds[1534]), .FEAT_ABOVE(feature_aboves[1534]), .FEAT_BELOW(feature_belows[1534])) ac1534(.scan_win(scan_win1534), .scan_win_std_dev(scan_win_std_dev[1534]), .feature_accum(feature_accums[1534]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1535]), .RECT1_Y(rectangle1_ys[1535]), .RECT1_WIDTH(rectangle1_widths[1535]), .RECT1_HEIGHT(rectangle1_heights[1535]), .RECT1_WEIGHT(rectangle1_weights[1535]), .RECT2_X(rectangle2_xs[1535]), .RECT2_Y(rectangle2_ys[1535]), .RECT2_WIDTH(rectangle2_widths[1535]), .RECT2_HEIGHT(rectangle2_heights[1535]), .RECT2_WEIGHT(rectangle2_weights[1535]), .RECT3_X(rectangle3_xs[1535]), .RECT3_Y(rectangle3_ys[1535]), .RECT3_WIDTH(rectangle3_widths[1535]), .RECT3_HEIGHT(rectangle3_heights[1535]), .RECT3_WEIGHT(rectangle3_weights[1535]), .FEAT_THRES(feature_thresholds[1535]), .FEAT_ABOVE(feature_aboves[1535]), .FEAT_BELOW(feature_belows[1535])) ac1535(.scan_win(scan_win1535), .scan_win_std_dev(scan_win_std_dev[1535]), .feature_accum(feature_accums[1535]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1536]), .RECT1_Y(rectangle1_ys[1536]), .RECT1_WIDTH(rectangle1_widths[1536]), .RECT1_HEIGHT(rectangle1_heights[1536]), .RECT1_WEIGHT(rectangle1_weights[1536]), .RECT2_X(rectangle2_xs[1536]), .RECT2_Y(rectangle2_ys[1536]), .RECT2_WIDTH(rectangle2_widths[1536]), .RECT2_HEIGHT(rectangle2_heights[1536]), .RECT2_WEIGHT(rectangle2_weights[1536]), .RECT3_X(rectangle3_xs[1536]), .RECT3_Y(rectangle3_ys[1536]), .RECT3_WIDTH(rectangle3_widths[1536]), .RECT3_HEIGHT(rectangle3_heights[1536]), .RECT3_WEIGHT(rectangle3_weights[1536]), .FEAT_THRES(feature_thresholds[1536]), .FEAT_ABOVE(feature_aboves[1536]), .FEAT_BELOW(feature_belows[1536])) ac1536(.scan_win(scan_win1536), .scan_win_std_dev(scan_win_std_dev[1536]), .feature_accum(feature_accums[1536]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1537]), .RECT1_Y(rectangle1_ys[1537]), .RECT1_WIDTH(rectangle1_widths[1537]), .RECT1_HEIGHT(rectangle1_heights[1537]), .RECT1_WEIGHT(rectangle1_weights[1537]), .RECT2_X(rectangle2_xs[1537]), .RECT2_Y(rectangle2_ys[1537]), .RECT2_WIDTH(rectangle2_widths[1537]), .RECT2_HEIGHT(rectangle2_heights[1537]), .RECT2_WEIGHT(rectangle2_weights[1537]), .RECT3_X(rectangle3_xs[1537]), .RECT3_Y(rectangle3_ys[1537]), .RECT3_WIDTH(rectangle3_widths[1537]), .RECT3_HEIGHT(rectangle3_heights[1537]), .RECT3_WEIGHT(rectangle3_weights[1537]), .FEAT_THRES(feature_thresholds[1537]), .FEAT_ABOVE(feature_aboves[1537]), .FEAT_BELOW(feature_belows[1537])) ac1537(.scan_win(scan_win1537), .scan_win_std_dev(scan_win_std_dev[1537]), .feature_accum(feature_accums[1537]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1538]), .RECT1_Y(rectangle1_ys[1538]), .RECT1_WIDTH(rectangle1_widths[1538]), .RECT1_HEIGHT(rectangle1_heights[1538]), .RECT1_WEIGHT(rectangle1_weights[1538]), .RECT2_X(rectangle2_xs[1538]), .RECT2_Y(rectangle2_ys[1538]), .RECT2_WIDTH(rectangle2_widths[1538]), .RECT2_HEIGHT(rectangle2_heights[1538]), .RECT2_WEIGHT(rectangle2_weights[1538]), .RECT3_X(rectangle3_xs[1538]), .RECT3_Y(rectangle3_ys[1538]), .RECT3_WIDTH(rectangle3_widths[1538]), .RECT3_HEIGHT(rectangle3_heights[1538]), .RECT3_WEIGHT(rectangle3_weights[1538]), .FEAT_THRES(feature_thresholds[1538]), .FEAT_ABOVE(feature_aboves[1538]), .FEAT_BELOW(feature_belows[1538])) ac1538(.scan_win(scan_win1538), .scan_win_std_dev(scan_win_std_dev[1538]), .feature_accum(feature_accums[1538]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1539]), .RECT1_Y(rectangle1_ys[1539]), .RECT1_WIDTH(rectangle1_widths[1539]), .RECT1_HEIGHT(rectangle1_heights[1539]), .RECT1_WEIGHT(rectangle1_weights[1539]), .RECT2_X(rectangle2_xs[1539]), .RECT2_Y(rectangle2_ys[1539]), .RECT2_WIDTH(rectangle2_widths[1539]), .RECT2_HEIGHT(rectangle2_heights[1539]), .RECT2_WEIGHT(rectangle2_weights[1539]), .RECT3_X(rectangle3_xs[1539]), .RECT3_Y(rectangle3_ys[1539]), .RECT3_WIDTH(rectangle3_widths[1539]), .RECT3_HEIGHT(rectangle3_heights[1539]), .RECT3_WEIGHT(rectangle3_weights[1539]), .FEAT_THRES(feature_thresholds[1539]), .FEAT_ABOVE(feature_aboves[1539]), .FEAT_BELOW(feature_belows[1539])) ac1539(.scan_win(scan_win1539), .scan_win_std_dev(scan_win_std_dev[1539]), .feature_accum(feature_accums[1539]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1540]), .RECT1_Y(rectangle1_ys[1540]), .RECT1_WIDTH(rectangle1_widths[1540]), .RECT1_HEIGHT(rectangle1_heights[1540]), .RECT1_WEIGHT(rectangle1_weights[1540]), .RECT2_X(rectangle2_xs[1540]), .RECT2_Y(rectangle2_ys[1540]), .RECT2_WIDTH(rectangle2_widths[1540]), .RECT2_HEIGHT(rectangle2_heights[1540]), .RECT2_WEIGHT(rectangle2_weights[1540]), .RECT3_X(rectangle3_xs[1540]), .RECT3_Y(rectangle3_ys[1540]), .RECT3_WIDTH(rectangle3_widths[1540]), .RECT3_HEIGHT(rectangle3_heights[1540]), .RECT3_WEIGHT(rectangle3_weights[1540]), .FEAT_THRES(feature_thresholds[1540]), .FEAT_ABOVE(feature_aboves[1540]), .FEAT_BELOW(feature_belows[1540])) ac1540(.scan_win(scan_win1540), .scan_win_std_dev(scan_win_std_dev[1540]), .feature_accum(feature_accums[1540]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1541]), .RECT1_Y(rectangle1_ys[1541]), .RECT1_WIDTH(rectangle1_widths[1541]), .RECT1_HEIGHT(rectangle1_heights[1541]), .RECT1_WEIGHT(rectangle1_weights[1541]), .RECT2_X(rectangle2_xs[1541]), .RECT2_Y(rectangle2_ys[1541]), .RECT2_WIDTH(rectangle2_widths[1541]), .RECT2_HEIGHT(rectangle2_heights[1541]), .RECT2_WEIGHT(rectangle2_weights[1541]), .RECT3_X(rectangle3_xs[1541]), .RECT3_Y(rectangle3_ys[1541]), .RECT3_WIDTH(rectangle3_widths[1541]), .RECT3_HEIGHT(rectangle3_heights[1541]), .RECT3_WEIGHT(rectangle3_weights[1541]), .FEAT_THRES(feature_thresholds[1541]), .FEAT_ABOVE(feature_aboves[1541]), .FEAT_BELOW(feature_belows[1541])) ac1541(.scan_win(scan_win1541), .scan_win_std_dev(scan_win_std_dev[1541]), .feature_accum(feature_accums[1541]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1542]), .RECT1_Y(rectangle1_ys[1542]), .RECT1_WIDTH(rectangle1_widths[1542]), .RECT1_HEIGHT(rectangle1_heights[1542]), .RECT1_WEIGHT(rectangle1_weights[1542]), .RECT2_X(rectangle2_xs[1542]), .RECT2_Y(rectangle2_ys[1542]), .RECT2_WIDTH(rectangle2_widths[1542]), .RECT2_HEIGHT(rectangle2_heights[1542]), .RECT2_WEIGHT(rectangle2_weights[1542]), .RECT3_X(rectangle3_xs[1542]), .RECT3_Y(rectangle3_ys[1542]), .RECT3_WIDTH(rectangle3_widths[1542]), .RECT3_HEIGHT(rectangle3_heights[1542]), .RECT3_WEIGHT(rectangle3_weights[1542]), .FEAT_THRES(feature_thresholds[1542]), .FEAT_ABOVE(feature_aboves[1542]), .FEAT_BELOW(feature_belows[1542])) ac1542(.scan_win(scan_win1542), .scan_win_std_dev(scan_win_std_dev[1542]), .feature_accum(feature_accums[1542]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1543]), .RECT1_Y(rectangle1_ys[1543]), .RECT1_WIDTH(rectangle1_widths[1543]), .RECT1_HEIGHT(rectangle1_heights[1543]), .RECT1_WEIGHT(rectangle1_weights[1543]), .RECT2_X(rectangle2_xs[1543]), .RECT2_Y(rectangle2_ys[1543]), .RECT2_WIDTH(rectangle2_widths[1543]), .RECT2_HEIGHT(rectangle2_heights[1543]), .RECT2_WEIGHT(rectangle2_weights[1543]), .RECT3_X(rectangle3_xs[1543]), .RECT3_Y(rectangle3_ys[1543]), .RECT3_WIDTH(rectangle3_widths[1543]), .RECT3_HEIGHT(rectangle3_heights[1543]), .RECT3_WEIGHT(rectangle3_weights[1543]), .FEAT_THRES(feature_thresholds[1543]), .FEAT_ABOVE(feature_aboves[1543]), .FEAT_BELOW(feature_belows[1543])) ac1543(.scan_win(scan_win1543), .scan_win_std_dev(scan_win_std_dev[1543]), .feature_accum(feature_accums[1543]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1544]), .RECT1_Y(rectangle1_ys[1544]), .RECT1_WIDTH(rectangle1_widths[1544]), .RECT1_HEIGHT(rectangle1_heights[1544]), .RECT1_WEIGHT(rectangle1_weights[1544]), .RECT2_X(rectangle2_xs[1544]), .RECT2_Y(rectangle2_ys[1544]), .RECT2_WIDTH(rectangle2_widths[1544]), .RECT2_HEIGHT(rectangle2_heights[1544]), .RECT2_WEIGHT(rectangle2_weights[1544]), .RECT3_X(rectangle3_xs[1544]), .RECT3_Y(rectangle3_ys[1544]), .RECT3_WIDTH(rectangle3_widths[1544]), .RECT3_HEIGHT(rectangle3_heights[1544]), .RECT3_WEIGHT(rectangle3_weights[1544]), .FEAT_THRES(feature_thresholds[1544]), .FEAT_ABOVE(feature_aboves[1544]), .FEAT_BELOW(feature_belows[1544])) ac1544(.scan_win(scan_win1544), .scan_win_std_dev(scan_win_std_dev[1544]), .feature_accum(feature_accums[1544]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1545]), .RECT1_Y(rectangle1_ys[1545]), .RECT1_WIDTH(rectangle1_widths[1545]), .RECT1_HEIGHT(rectangle1_heights[1545]), .RECT1_WEIGHT(rectangle1_weights[1545]), .RECT2_X(rectangle2_xs[1545]), .RECT2_Y(rectangle2_ys[1545]), .RECT2_WIDTH(rectangle2_widths[1545]), .RECT2_HEIGHT(rectangle2_heights[1545]), .RECT2_WEIGHT(rectangle2_weights[1545]), .RECT3_X(rectangle3_xs[1545]), .RECT3_Y(rectangle3_ys[1545]), .RECT3_WIDTH(rectangle3_widths[1545]), .RECT3_HEIGHT(rectangle3_heights[1545]), .RECT3_WEIGHT(rectangle3_weights[1545]), .FEAT_THRES(feature_thresholds[1545]), .FEAT_ABOVE(feature_aboves[1545]), .FEAT_BELOW(feature_belows[1545])) ac1545(.scan_win(scan_win1545), .scan_win_std_dev(scan_win_std_dev[1545]), .feature_accum(feature_accums[1545]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1546]), .RECT1_Y(rectangle1_ys[1546]), .RECT1_WIDTH(rectangle1_widths[1546]), .RECT1_HEIGHT(rectangle1_heights[1546]), .RECT1_WEIGHT(rectangle1_weights[1546]), .RECT2_X(rectangle2_xs[1546]), .RECT2_Y(rectangle2_ys[1546]), .RECT2_WIDTH(rectangle2_widths[1546]), .RECT2_HEIGHT(rectangle2_heights[1546]), .RECT2_WEIGHT(rectangle2_weights[1546]), .RECT3_X(rectangle3_xs[1546]), .RECT3_Y(rectangle3_ys[1546]), .RECT3_WIDTH(rectangle3_widths[1546]), .RECT3_HEIGHT(rectangle3_heights[1546]), .RECT3_WEIGHT(rectangle3_weights[1546]), .FEAT_THRES(feature_thresholds[1546]), .FEAT_ABOVE(feature_aboves[1546]), .FEAT_BELOW(feature_belows[1546])) ac1546(.scan_win(scan_win1546), .scan_win_std_dev(scan_win_std_dev[1546]), .feature_accum(feature_accums[1546]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1547]), .RECT1_Y(rectangle1_ys[1547]), .RECT1_WIDTH(rectangle1_widths[1547]), .RECT1_HEIGHT(rectangle1_heights[1547]), .RECT1_WEIGHT(rectangle1_weights[1547]), .RECT2_X(rectangle2_xs[1547]), .RECT2_Y(rectangle2_ys[1547]), .RECT2_WIDTH(rectangle2_widths[1547]), .RECT2_HEIGHT(rectangle2_heights[1547]), .RECT2_WEIGHT(rectangle2_weights[1547]), .RECT3_X(rectangle3_xs[1547]), .RECT3_Y(rectangle3_ys[1547]), .RECT3_WIDTH(rectangle3_widths[1547]), .RECT3_HEIGHT(rectangle3_heights[1547]), .RECT3_WEIGHT(rectangle3_weights[1547]), .FEAT_THRES(feature_thresholds[1547]), .FEAT_ABOVE(feature_aboves[1547]), .FEAT_BELOW(feature_belows[1547])) ac1547(.scan_win(scan_win1547), .scan_win_std_dev(scan_win_std_dev[1547]), .feature_accum(feature_accums[1547]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1548]), .RECT1_Y(rectangle1_ys[1548]), .RECT1_WIDTH(rectangle1_widths[1548]), .RECT1_HEIGHT(rectangle1_heights[1548]), .RECT1_WEIGHT(rectangle1_weights[1548]), .RECT2_X(rectangle2_xs[1548]), .RECT2_Y(rectangle2_ys[1548]), .RECT2_WIDTH(rectangle2_widths[1548]), .RECT2_HEIGHT(rectangle2_heights[1548]), .RECT2_WEIGHT(rectangle2_weights[1548]), .RECT3_X(rectangle3_xs[1548]), .RECT3_Y(rectangle3_ys[1548]), .RECT3_WIDTH(rectangle3_widths[1548]), .RECT3_HEIGHT(rectangle3_heights[1548]), .RECT3_WEIGHT(rectangle3_weights[1548]), .FEAT_THRES(feature_thresholds[1548]), .FEAT_ABOVE(feature_aboves[1548]), .FEAT_BELOW(feature_belows[1548])) ac1548(.scan_win(scan_win1548), .scan_win_std_dev(scan_win_std_dev[1548]), .feature_accum(feature_accums[1548]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1549]), .RECT1_Y(rectangle1_ys[1549]), .RECT1_WIDTH(rectangle1_widths[1549]), .RECT1_HEIGHT(rectangle1_heights[1549]), .RECT1_WEIGHT(rectangle1_weights[1549]), .RECT2_X(rectangle2_xs[1549]), .RECT2_Y(rectangle2_ys[1549]), .RECT2_WIDTH(rectangle2_widths[1549]), .RECT2_HEIGHT(rectangle2_heights[1549]), .RECT2_WEIGHT(rectangle2_weights[1549]), .RECT3_X(rectangle3_xs[1549]), .RECT3_Y(rectangle3_ys[1549]), .RECT3_WIDTH(rectangle3_widths[1549]), .RECT3_HEIGHT(rectangle3_heights[1549]), .RECT3_WEIGHT(rectangle3_weights[1549]), .FEAT_THRES(feature_thresholds[1549]), .FEAT_ABOVE(feature_aboves[1549]), .FEAT_BELOW(feature_belows[1549])) ac1549(.scan_win(scan_win1549), .scan_win_std_dev(scan_win_std_dev[1549]), .feature_accum(feature_accums[1549]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1550]), .RECT1_Y(rectangle1_ys[1550]), .RECT1_WIDTH(rectangle1_widths[1550]), .RECT1_HEIGHT(rectangle1_heights[1550]), .RECT1_WEIGHT(rectangle1_weights[1550]), .RECT2_X(rectangle2_xs[1550]), .RECT2_Y(rectangle2_ys[1550]), .RECT2_WIDTH(rectangle2_widths[1550]), .RECT2_HEIGHT(rectangle2_heights[1550]), .RECT2_WEIGHT(rectangle2_weights[1550]), .RECT3_X(rectangle3_xs[1550]), .RECT3_Y(rectangle3_ys[1550]), .RECT3_WIDTH(rectangle3_widths[1550]), .RECT3_HEIGHT(rectangle3_heights[1550]), .RECT3_WEIGHT(rectangle3_weights[1550]), .FEAT_THRES(feature_thresholds[1550]), .FEAT_ABOVE(feature_aboves[1550]), .FEAT_BELOW(feature_belows[1550])) ac1550(.scan_win(scan_win1550), .scan_win_std_dev(scan_win_std_dev[1550]), .feature_accum(feature_accums[1550]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1551]), .RECT1_Y(rectangle1_ys[1551]), .RECT1_WIDTH(rectangle1_widths[1551]), .RECT1_HEIGHT(rectangle1_heights[1551]), .RECT1_WEIGHT(rectangle1_weights[1551]), .RECT2_X(rectangle2_xs[1551]), .RECT2_Y(rectangle2_ys[1551]), .RECT2_WIDTH(rectangle2_widths[1551]), .RECT2_HEIGHT(rectangle2_heights[1551]), .RECT2_WEIGHT(rectangle2_weights[1551]), .RECT3_X(rectangle3_xs[1551]), .RECT3_Y(rectangle3_ys[1551]), .RECT3_WIDTH(rectangle3_widths[1551]), .RECT3_HEIGHT(rectangle3_heights[1551]), .RECT3_WEIGHT(rectangle3_weights[1551]), .FEAT_THRES(feature_thresholds[1551]), .FEAT_ABOVE(feature_aboves[1551]), .FEAT_BELOW(feature_belows[1551])) ac1551(.scan_win(scan_win1551), .scan_win_std_dev(scan_win_std_dev[1551]), .feature_accum(feature_accums[1551]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1552]), .RECT1_Y(rectangle1_ys[1552]), .RECT1_WIDTH(rectangle1_widths[1552]), .RECT1_HEIGHT(rectangle1_heights[1552]), .RECT1_WEIGHT(rectangle1_weights[1552]), .RECT2_X(rectangle2_xs[1552]), .RECT2_Y(rectangle2_ys[1552]), .RECT2_WIDTH(rectangle2_widths[1552]), .RECT2_HEIGHT(rectangle2_heights[1552]), .RECT2_WEIGHT(rectangle2_weights[1552]), .RECT3_X(rectangle3_xs[1552]), .RECT3_Y(rectangle3_ys[1552]), .RECT3_WIDTH(rectangle3_widths[1552]), .RECT3_HEIGHT(rectangle3_heights[1552]), .RECT3_WEIGHT(rectangle3_weights[1552]), .FEAT_THRES(feature_thresholds[1552]), .FEAT_ABOVE(feature_aboves[1552]), .FEAT_BELOW(feature_belows[1552])) ac1552(.scan_win(scan_win1552), .scan_win_std_dev(scan_win_std_dev[1552]), .feature_accum(feature_accums[1552]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1553]), .RECT1_Y(rectangle1_ys[1553]), .RECT1_WIDTH(rectangle1_widths[1553]), .RECT1_HEIGHT(rectangle1_heights[1553]), .RECT1_WEIGHT(rectangle1_weights[1553]), .RECT2_X(rectangle2_xs[1553]), .RECT2_Y(rectangle2_ys[1553]), .RECT2_WIDTH(rectangle2_widths[1553]), .RECT2_HEIGHT(rectangle2_heights[1553]), .RECT2_WEIGHT(rectangle2_weights[1553]), .RECT3_X(rectangle3_xs[1553]), .RECT3_Y(rectangle3_ys[1553]), .RECT3_WIDTH(rectangle3_widths[1553]), .RECT3_HEIGHT(rectangle3_heights[1553]), .RECT3_WEIGHT(rectangle3_weights[1553]), .FEAT_THRES(feature_thresholds[1553]), .FEAT_ABOVE(feature_aboves[1553]), .FEAT_BELOW(feature_belows[1553])) ac1553(.scan_win(scan_win1553), .scan_win_std_dev(scan_win_std_dev[1553]), .feature_accum(feature_accums[1553]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1554]), .RECT1_Y(rectangle1_ys[1554]), .RECT1_WIDTH(rectangle1_widths[1554]), .RECT1_HEIGHT(rectangle1_heights[1554]), .RECT1_WEIGHT(rectangle1_weights[1554]), .RECT2_X(rectangle2_xs[1554]), .RECT2_Y(rectangle2_ys[1554]), .RECT2_WIDTH(rectangle2_widths[1554]), .RECT2_HEIGHT(rectangle2_heights[1554]), .RECT2_WEIGHT(rectangle2_weights[1554]), .RECT3_X(rectangle3_xs[1554]), .RECT3_Y(rectangle3_ys[1554]), .RECT3_WIDTH(rectangle3_widths[1554]), .RECT3_HEIGHT(rectangle3_heights[1554]), .RECT3_WEIGHT(rectangle3_weights[1554]), .FEAT_THRES(feature_thresholds[1554]), .FEAT_ABOVE(feature_aboves[1554]), .FEAT_BELOW(feature_belows[1554])) ac1554(.scan_win(scan_win1554), .scan_win_std_dev(scan_win_std_dev[1554]), .feature_accum(feature_accums[1554]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1555]), .RECT1_Y(rectangle1_ys[1555]), .RECT1_WIDTH(rectangle1_widths[1555]), .RECT1_HEIGHT(rectangle1_heights[1555]), .RECT1_WEIGHT(rectangle1_weights[1555]), .RECT2_X(rectangle2_xs[1555]), .RECT2_Y(rectangle2_ys[1555]), .RECT2_WIDTH(rectangle2_widths[1555]), .RECT2_HEIGHT(rectangle2_heights[1555]), .RECT2_WEIGHT(rectangle2_weights[1555]), .RECT3_X(rectangle3_xs[1555]), .RECT3_Y(rectangle3_ys[1555]), .RECT3_WIDTH(rectangle3_widths[1555]), .RECT3_HEIGHT(rectangle3_heights[1555]), .RECT3_WEIGHT(rectangle3_weights[1555]), .FEAT_THRES(feature_thresholds[1555]), .FEAT_ABOVE(feature_aboves[1555]), .FEAT_BELOW(feature_belows[1555])) ac1555(.scan_win(scan_win1555), .scan_win_std_dev(scan_win_std_dev[1555]), .feature_accum(feature_accums[1555]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1556]), .RECT1_Y(rectangle1_ys[1556]), .RECT1_WIDTH(rectangle1_widths[1556]), .RECT1_HEIGHT(rectangle1_heights[1556]), .RECT1_WEIGHT(rectangle1_weights[1556]), .RECT2_X(rectangle2_xs[1556]), .RECT2_Y(rectangle2_ys[1556]), .RECT2_WIDTH(rectangle2_widths[1556]), .RECT2_HEIGHT(rectangle2_heights[1556]), .RECT2_WEIGHT(rectangle2_weights[1556]), .RECT3_X(rectangle3_xs[1556]), .RECT3_Y(rectangle3_ys[1556]), .RECT3_WIDTH(rectangle3_widths[1556]), .RECT3_HEIGHT(rectangle3_heights[1556]), .RECT3_WEIGHT(rectangle3_weights[1556]), .FEAT_THRES(feature_thresholds[1556]), .FEAT_ABOVE(feature_aboves[1556]), .FEAT_BELOW(feature_belows[1556])) ac1556(.scan_win(scan_win1556), .scan_win_std_dev(scan_win_std_dev[1556]), .feature_accum(feature_accums[1556]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1557]), .RECT1_Y(rectangle1_ys[1557]), .RECT1_WIDTH(rectangle1_widths[1557]), .RECT1_HEIGHT(rectangle1_heights[1557]), .RECT1_WEIGHT(rectangle1_weights[1557]), .RECT2_X(rectangle2_xs[1557]), .RECT2_Y(rectangle2_ys[1557]), .RECT2_WIDTH(rectangle2_widths[1557]), .RECT2_HEIGHT(rectangle2_heights[1557]), .RECT2_WEIGHT(rectangle2_weights[1557]), .RECT3_X(rectangle3_xs[1557]), .RECT3_Y(rectangle3_ys[1557]), .RECT3_WIDTH(rectangle3_widths[1557]), .RECT3_HEIGHT(rectangle3_heights[1557]), .RECT3_WEIGHT(rectangle3_weights[1557]), .FEAT_THRES(feature_thresholds[1557]), .FEAT_ABOVE(feature_aboves[1557]), .FEAT_BELOW(feature_belows[1557])) ac1557(.scan_win(scan_win1557), .scan_win_std_dev(scan_win_std_dev[1557]), .feature_accum(feature_accums[1557]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1558]), .RECT1_Y(rectangle1_ys[1558]), .RECT1_WIDTH(rectangle1_widths[1558]), .RECT1_HEIGHT(rectangle1_heights[1558]), .RECT1_WEIGHT(rectangle1_weights[1558]), .RECT2_X(rectangle2_xs[1558]), .RECT2_Y(rectangle2_ys[1558]), .RECT2_WIDTH(rectangle2_widths[1558]), .RECT2_HEIGHT(rectangle2_heights[1558]), .RECT2_WEIGHT(rectangle2_weights[1558]), .RECT3_X(rectangle3_xs[1558]), .RECT3_Y(rectangle3_ys[1558]), .RECT3_WIDTH(rectangle3_widths[1558]), .RECT3_HEIGHT(rectangle3_heights[1558]), .RECT3_WEIGHT(rectangle3_weights[1558]), .FEAT_THRES(feature_thresholds[1558]), .FEAT_ABOVE(feature_aboves[1558]), .FEAT_BELOW(feature_belows[1558])) ac1558(.scan_win(scan_win1558), .scan_win_std_dev(scan_win_std_dev[1558]), .feature_accum(feature_accums[1558]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1559]), .RECT1_Y(rectangle1_ys[1559]), .RECT1_WIDTH(rectangle1_widths[1559]), .RECT1_HEIGHT(rectangle1_heights[1559]), .RECT1_WEIGHT(rectangle1_weights[1559]), .RECT2_X(rectangle2_xs[1559]), .RECT2_Y(rectangle2_ys[1559]), .RECT2_WIDTH(rectangle2_widths[1559]), .RECT2_HEIGHT(rectangle2_heights[1559]), .RECT2_WEIGHT(rectangle2_weights[1559]), .RECT3_X(rectangle3_xs[1559]), .RECT3_Y(rectangle3_ys[1559]), .RECT3_WIDTH(rectangle3_widths[1559]), .RECT3_HEIGHT(rectangle3_heights[1559]), .RECT3_WEIGHT(rectangle3_weights[1559]), .FEAT_THRES(feature_thresholds[1559]), .FEAT_ABOVE(feature_aboves[1559]), .FEAT_BELOW(feature_belows[1559])) ac1559(.scan_win(scan_win1559), .scan_win_std_dev(scan_win_std_dev[1559]), .feature_accum(feature_accums[1559]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1560]), .RECT1_Y(rectangle1_ys[1560]), .RECT1_WIDTH(rectangle1_widths[1560]), .RECT1_HEIGHT(rectangle1_heights[1560]), .RECT1_WEIGHT(rectangle1_weights[1560]), .RECT2_X(rectangle2_xs[1560]), .RECT2_Y(rectangle2_ys[1560]), .RECT2_WIDTH(rectangle2_widths[1560]), .RECT2_HEIGHT(rectangle2_heights[1560]), .RECT2_WEIGHT(rectangle2_weights[1560]), .RECT3_X(rectangle3_xs[1560]), .RECT3_Y(rectangle3_ys[1560]), .RECT3_WIDTH(rectangle3_widths[1560]), .RECT3_HEIGHT(rectangle3_heights[1560]), .RECT3_WEIGHT(rectangle3_weights[1560]), .FEAT_THRES(feature_thresholds[1560]), .FEAT_ABOVE(feature_aboves[1560]), .FEAT_BELOW(feature_belows[1560])) ac1560(.scan_win(scan_win1560), .scan_win_std_dev(scan_win_std_dev[1560]), .feature_accum(feature_accums[1560]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1561]), .RECT1_Y(rectangle1_ys[1561]), .RECT1_WIDTH(rectangle1_widths[1561]), .RECT1_HEIGHT(rectangle1_heights[1561]), .RECT1_WEIGHT(rectangle1_weights[1561]), .RECT2_X(rectangle2_xs[1561]), .RECT2_Y(rectangle2_ys[1561]), .RECT2_WIDTH(rectangle2_widths[1561]), .RECT2_HEIGHT(rectangle2_heights[1561]), .RECT2_WEIGHT(rectangle2_weights[1561]), .RECT3_X(rectangle3_xs[1561]), .RECT3_Y(rectangle3_ys[1561]), .RECT3_WIDTH(rectangle3_widths[1561]), .RECT3_HEIGHT(rectangle3_heights[1561]), .RECT3_WEIGHT(rectangle3_weights[1561]), .FEAT_THRES(feature_thresholds[1561]), .FEAT_ABOVE(feature_aboves[1561]), .FEAT_BELOW(feature_belows[1561])) ac1561(.scan_win(scan_win1561), .scan_win_std_dev(scan_win_std_dev[1561]), .feature_accum(feature_accums[1561]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1562]), .RECT1_Y(rectangle1_ys[1562]), .RECT1_WIDTH(rectangle1_widths[1562]), .RECT1_HEIGHT(rectangle1_heights[1562]), .RECT1_WEIGHT(rectangle1_weights[1562]), .RECT2_X(rectangle2_xs[1562]), .RECT2_Y(rectangle2_ys[1562]), .RECT2_WIDTH(rectangle2_widths[1562]), .RECT2_HEIGHT(rectangle2_heights[1562]), .RECT2_WEIGHT(rectangle2_weights[1562]), .RECT3_X(rectangle3_xs[1562]), .RECT3_Y(rectangle3_ys[1562]), .RECT3_WIDTH(rectangle3_widths[1562]), .RECT3_HEIGHT(rectangle3_heights[1562]), .RECT3_WEIGHT(rectangle3_weights[1562]), .FEAT_THRES(feature_thresholds[1562]), .FEAT_ABOVE(feature_aboves[1562]), .FEAT_BELOW(feature_belows[1562])) ac1562(.scan_win(scan_win1562), .scan_win_std_dev(scan_win_std_dev[1562]), .feature_accum(feature_accums[1562]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1563]), .RECT1_Y(rectangle1_ys[1563]), .RECT1_WIDTH(rectangle1_widths[1563]), .RECT1_HEIGHT(rectangle1_heights[1563]), .RECT1_WEIGHT(rectangle1_weights[1563]), .RECT2_X(rectangle2_xs[1563]), .RECT2_Y(rectangle2_ys[1563]), .RECT2_WIDTH(rectangle2_widths[1563]), .RECT2_HEIGHT(rectangle2_heights[1563]), .RECT2_WEIGHT(rectangle2_weights[1563]), .RECT3_X(rectangle3_xs[1563]), .RECT3_Y(rectangle3_ys[1563]), .RECT3_WIDTH(rectangle3_widths[1563]), .RECT3_HEIGHT(rectangle3_heights[1563]), .RECT3_WEIGHT(rectangle3_weights[1563]), .FEAT_THRES(feature_thresholds[1563]), .FEAT_ABOVE(feature_aboves[1563]), .FEAT_BELOW(feature_belows[1563])) ac1563(.scan_win(scan_win1563), .scan_win_std_dev(scan_win_std_dev[1563]), .feature_accum(feature_accums[1563]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1564]), .RECT1_Y(rectangle1_ys[1564]), .RECT1_WIDTH(rectangle1_widths[1564]), .RECT1_HEIGHT(rectangle1_heights[1564]), .RECT1_WEIGHT(rectangle1_weights[1564]), .RECT2_X(rectangle2_xs[1564]), .RECT2_Y(rectangle2_ys[1564]), .RECT2_WIDTH(rectangle2_widths[1564]), .RECT2_HEIGHT(rectangle2_heights[1564]), .RECT2_WEIGHT(rectangle2_weights[1564]), .RECT3_X(rectangle3_xs[1564]), .RECT3_Y(rectangle3_ys[1564]), .RECT3_WIDTH(rectangle3_widths[1564]), .RECT3_HEIGHT(rectangle3_heights[1564]), .RECT3_WEIGHT(rectangle3_weights[1564]), .FEAT_THRES(feature_thresholds[1564]), .FEAT_ABOVE(feature_aboves[1564]), .FEAT_BELOW(feature_belows[1564])) ac1564(.scan_win(scan_win1564), .scan_win_std_dev(scan_win_std_dev[1564]), .feature_accum(feature_accums[1564]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1565]), .RECT1_Y(rectangle1_ys[1565]), .RECT1_WIDTH(rectangle1_widths[1565]), .RECT1_HEIGHT(rectangle1_heights[1565]), .RECT1_WEIGHT(rectangle1_weights[1565]), .RECT2_X(rectangle2_xs[1565]), .RECT2_Y(rectangle2_ys[1565]), .RECT2_WIDTH(rectangle2_widths[1565]), .RECT2_HEIGHT(rectangle2_heights[1565]), .RECT2_WEIGHT(rectangle2_weights[1565]), .RECT3_X(rectangle3_xs[1565]), .RECT3_Y(rectangle3_ys[1565]), .RECT3_WIDTH(rectangle3_widths[1565]), .RECT3_HEIGHT(rectangle3_heights[1565]), .RECT3_WEIGHT(rectangle3_weights[1565]), .FEAT_THRES(feature_thresholds[1565]), .FEAT_ABOVE(feature_aboves[1565]), .FEAT_BELOW(feature_belows[1565])) ac1565(.scan_win(scan_win1565), .scan_win_std_dev(scan_win_std_dev[1565]), .feature_accum(feature_accums[1565]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1566]), .RECT1_Y(rectangle1_ys[1566]), .RECT1_WIDTH(rectangle1_widths[1566]), .RECT1_HEIGHT(rectangle1_heights[1566]), .RECT1_WEIGHT(rectangle1_weights[1566]), .RECT2_X(rectangle2_xs[1566]), .RECT2_Y(rectangle2_ys[1566]), .RECT2_WIDTH(rectangle2_widths[1566]), .RECT2_HEIGHT(rectangle2_heights[1566]), .RECT2_WEIGHT(rectangle2_weights[1566]), .RECT3_X(rectangle3_xs[1566]), .RECT3_Y(rectangle3_ys[1566]), .RECT3_WIDTH(rectangle3_widths[1566]), .RECT3_HEIGHT(rectangle3_heights[1566]), .RECT3_WEIGHT(rectangle3_weights[1566]), .FEAT_THRES(feature_thresholds[1566]), .FEAT_ABOVE(feature_aboves[1566]), .FEAT_BELOW(feature_belows[1566])) ac1566(.scan_win(scan_win1566), .scan_win_std_dev(scan_win_std_dev[1566]), .feature_accum(feature_accums[1566]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1567]), .RECT1_Y(rectangle1_ys[1567]), .RECT1_WIDTH(rectangle1_widths[1567]), .RECT1_HEIGHT(rectangle1_heights[1567]), .RECT1_WEIGHT(rectangle1_weights[1567]), .RECT2_X(rectangle2_xs[1567]), .RECT2_Y(rectangle2_ys[1567]), .RECT2_WIDTH(rectangle2_widths[1567]), .RECT2_HEIGHT(rectangle2_heights[1567]), .RECT2_WEIGHT(rectangle2_weights[1567]), .RECT3_X(rectangle3_xs[1567]), .RECT3_Y(rectangle3_ys[1567]), .RECT3_WIDTH(rectangle3_widths[1567]), .RECT3_HEIGHT(rectangle3_heights[1567]), .RECT3_WEIGHT(rectangle3_weights[1567]), .FEAT_THRES(feature_thresholds[1567]), .FEAT_ABOVE(feature_aboves[1567]), .FEAT_BELOW(feature_belows[1567])) ac1567(.scan_win(scan_win1567), .scan_win_std_dev(scan_win_std_dev[1567]), .feature_accum(feature_accums[1567]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1568]), .RECT1_Y(rectangle1_ys[1568]), .RECT1_WIDTH(rectangle1_widths[1568]), .RECT1_HEIGHT(rectangle1_heights[1568]), .RECT1_WEIGHT(rectangle1_weights[1568]), .RECT2_X(rectangle2_xs[1568]), .RECT2_Y(rectangle2_ys[1568]), .RECT2_WIDTH(rectangle2_widths[1568]), .RECT2_HEIGHT(rectangle2_heights[1568]), .RECT2_WEIGHT(rectangle2_weights[1568]), .RECT3_X(rectangle3_xs[1568]), .RECT3_Y(rectangle3_ys[1568]), .RECT3_WIDTH(rectangle3_widths[1568]), .RECT3_HEIGHT(rectangle3_heights[1568]), .RECT3_WEIGHT(rectangle3_weights[1568]), .FEAT_THRES(feature_thresholds[1568]), .FEAT_ABOVE(feature_aboves[1568]), .FEAT_BELOW(feature_belows[1568])) ac1568(.scan_win(scan_win1568), .scan_win_std_dev(scan_win_std_dev[1568]), .feature_accum(feature_accums[1568]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1569]), .RECT1_Y(rectangle1_ys[1569]), .RECT1_WIDTH(rectangle1_widths[1569]), .RECT1_HEIGHT(rectangle1_heights[1569]), .RECT1_WEIGHT(rectangle1_weights[1569]), .RECT2_X(rectangle2_xs[1569]), .RECT2_Y(rectangle2_ys[1569]), .RECT2_WIDTH(rectangle2_widths[1569]), .RECT2_HEIGHT(rectangle2_heights[1569]), .RECT2_WEIGHT(rectangle2_weights[1569]), .RECT3_X(rectangle3_xs[1569]), .RECT3_Y(rectangle3_ys[1569]), .RECT3_WIDTH(rectangle3_widths[1569]), .RECT3_HEIGHT(rectangle3_heights[1569]), .RECT3_WEIGHT(rectangle3_weights[1569]), .FEAT_THRES(feature_thresholds[1569]), .FEAT_ABOVE(feature_aboves[1569]), .FEAT_BELOW(feature_belows[1569])) ac1569(.scan_win(scan_win1569), .scan_win_std_dev(scan_win_std_dev[1569]), .feature_accum(feature_accums[1569]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1570]), .RECT1_Y(rectangle1_ys[1570]), .RECT1_WIDTH(rectangle1_widths[1570]), .RECT1_HEIGHT(rectangle1_heights[1570]), .RECT1_WEIGHT(rectangle1_weights[1570]), .RECT2_X(rectangle2_xs[1570]), .RECT2_Y(rectangle2_ys[1570]), .RECT2_WIDTH(rectangle2_widths[1570]), .RECT2_HEIGHT(rectangle2_heights[1570]), .RECT2_WEIGHT(rectangle2_weights[1570]), .RECT3_X(rectangle3_xs[1570]), .RECT3_Y(rectangle3_ys[1570]), .RECT3_WIDTH(rectangle3_widths[1570]), .RECT3_HEIGHT(rectangle3_heights[1570]), .RECT3_WEIGHT(rectangle3_weights[1570]), .FEAT_THRES(feature_thresholds[1570]), .FEAT_ABOVE(feature_aboves[1570]), .FEAT_BELOW(feature_belows[1570])) ac1570(.scan_win(scan_win1570), .scan_win_std_dev(scan_win_std_dev[1570]), .feature_accum(feature_accums[1570]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1571]), .RECT1_Y(rectangle1_ys[1571]), .RECT1_WIDTH(rectangle1_widths[1571]), .RECT1_HEIGHT(rectangle1_heights[1571]), .RECT1_WEIGHT(rectangle1_weights[1571]), .RECT2_X(rectangle2_xs[1571]), .RECT2_Y(rectangle2_ys[1571]), .RECT2_WIDTH(rectangle2_widths[1571]), .RECT2_HEIGHT(rectangle2_heights[1571]), .RECT2_WEIGHT(rectangle2_weights[1571]), .RECT3_X(rectangle3_xs[1571]), .RECT3_Y(rectangle3_ys[1571]), .RECT3_WIDTH(rectangle3_widths[1571]), .RECT3_HEIGHT(rectangle3_heights[1571]), .RECT3_WEIGHT(rectangle3_weights[1571]), .FEAT_THRES(feature_thresholds[1571]), .FEAT_ABOVE(feature_aboves[1571]), .FEAT_BELOW(feature_belows[1571])) ac1571(.scan_win(scan_win1571), .scan_win_std_dev(scan_win_std_dev[1571]), .feature_accum(feature_accums[1571]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1572]), .RECT1_Y(rectangle1_ys[1572]), .RECT1_WIDTH(rectangle1_widths[1572]), .RECT1_HEIGHT(rectangle1_heights[1572]), .RECT1_WEIGHT(rectangle1_weights[1572]), .RECT2_X(rectangle2_xs[1572]), .RECT2_Y(rectangle2_ys[1572]), .RECT2_WIDTH(rectangle2_widths[1572]), .RECT2_HEIGHT(rectangle2_heights[1572]), .RECT2_WEIGHT(rectangle2_weights[1572]), .RECT3_X(rectangle3_xs[1572]), .RECT3_Y(rectangle3_ys[1572]), .RECT3_WIDTH(rectangle3_widths[1572]), .RECT3_HEIGHT(rectangle3_heights[1572]), .RECT3_WEIGHT(rectangle3_weights[1572]), .FEAT_THRES(feature_thresholds[1572]), .FEAT_ABOVE(feature_aboves[1572]), .FEAT_BELOW(feature_belows[1572])) ac1572(.scan_win(scan_win1572), .scan_win_std_dev(scan_win_std_dev[1572]), .feature_accum(feature_accums[1572]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1573]), .RECT1_Y(rectangle1_ys[1573]), .RECT1_WIDTH(rectangle1_widths[1573]), .RECT1_HEIGHT(rectangle1_heights[1573]), .RECT1_WEIGHT(rectangle1_weights[1573]), .RECT2_X(rectangle2_xs[1573]), .RECT2_Y(rectangle2_ys[1573]), .RECT2_WIDTH(rectangle2_widths[1573]), .RECT2_HEIGHT(rectangle2_heights[1573]), .RECT2_WEIGHT(rectangle2_weights[1573]), .RECT3_X(rectangle3_xs[1573]), .RECT3_Y(rectangle3_ys[1573]), .RECT3_WIDTH(rectangle3_widths[1573]), .RECT3_HEIGHT(rectangle3_heights[1573]), .RECT3_WEIGHT(rectangle3_weights[1573]), .FEAT_THRES(feature_thresholds[1573]), .FEAT_ABOVE(feature_aboves[1573]), .FEAT_BELOW(feature_belows[1573])) ac1573(.scan_win(scan_win1573), .scan_win_std_dev(scan_win_std_dev[1573]), .feature_accum(feature_accums[1573]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1574]), .RECT1_Y(rectangle1_ys[1574]), .RECT1_WIDTH(rectangle1_widths[1574]), .RECT1_HEIGHT(rectangle1_heights[1574]), .RECT1_WEIGHT(rectangle1_weights[1574]), .RECT2_X(rectangle2_xs[1574]), .RECT2_Y(rectangle2_ys[1574]), .RECT2_WIDTH(rectangle2_widths[1574]), .RECT2_HEIGHT(rectangle2_heights[1574]), .RECT2_WEIGHT(rectangle2_weights[1574]), .RECT3_X(rectangle3_xs[1574]), .RECT3_Y(rectangle3_ys[1574]), .RECT3_WIDTH(rectangle3_widths[1574]), .RECT3_HEIGHT(rectangle3_heights[1574]), .RECT3_WEIGHT(rectangle3_weights[1574]), .FEAT_THRES(feature_thresholds[1574]), .FEAT_ABOVE(feature_aboves[1574]), .FEAT_BELOW(feature_belows[1574])) ac1574(.scan_win(scan_win1574), .scan_win_std_dev(scan_win_std_dev[1574]), .feature_accum(feature_accums[1574]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1575]), .RECT1_Y(rectangle1_ys[1575]), .RECT1_WIDTH(rectangle1_widths[1575]), .RECT1_HEIGHT(rectangle1_heights[1575]), .RECT1_WEIGHT(rectangle1_weights[1575]), .RECT2_X(rectangle2_xs[1575]), .RECT2_Y(rectangle2_ys[1575]), .RECT2_WIDTH(rectangle2_widths[1575]), .RECT2_HEIGHT(rectangle2_heights[1575]), .RECT2_WEIGHT(rectangle2_weights[1575]), .RECT3_X(rectangle3_xs[1575]), .RECT3_Y(rectangle3_ys[1575]), .RECT3_WIDTH(rectangle3_widths[1575]), .RECT3_HEIGHT(rectangle3_heights[1575]), .RECT3_WEIGHT(rectangle3_weights[1575]), .FEAT_THRES(feature_thresholds[1575]), .FEAT_ABOVE(feature_aboves[1575]), .FEAT_BELOW(feature_belows[1575])) ac1575(.scan_win(scan_win1575), .scan_win_std_dev(scan_win_std_dev[1575]), .feature_accum(feature_accums[1575]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1576]), .RECT1_Y(rectangle1_ys[1576]), .RECT1_WIDTH(rectangle1_widths[1576]), .RECT1_HEIGHT(rectangle1_heights[1576]), .RECT1_WEIGHT(rectangle1_weights[1576]), .RECT2_X(rectangle2_xs[1576]), .RECT2_Y(rectangle2_ys[1576]), .RECT2_WIDTH(rectangle2_widths[1576]), .RECT2_HEIGHT(rectangle2_heights[1576]), .RECT2_WEIGHT(rectangle2_weights[1576]), .RECT3_X(rectangle3_xs[1576]), .RECT3_Y(rectangle3_ys[1576]), .RECT3_WIDTH(rectangle3_widths[1576]), .RECT3_HEIGHT(rectangle3_heights[1576]), .RECT3_WEIGHT(rectangle3_weights[1576]), .FEAT_THRES(feature_thresholds[1576]), .FEAT_ABOVE(feature_aboves[1576]), .FEAT_BELOW(feature_belows[1576])) ac1576(.scan_win(scan_win1576), .scan_win_std_dev(scan_win_std_dev[1576]), .feature_accum(feature_accums[1576]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1577]), .RECT1_Y(rectangle1_ys[1577]), .RECT1_WIDTH(rectangle1_widths[1577]), .RECT1_HEIGHT(rectangle1_heights[1577]), .RECT1_WEIGHT(rectangle1_weights[1577]), .RECT2_X(rectangle2_xs[1577]), .RECT2_Y(rectangle2_ys[1577]), .RECT2_WIDTH(rectangle2_widths[1577]), .RECT2_HEIGHT(rectangle2_heights[1577]), .RECT2_WEIGHT(rectangle2_weights[1577]), .RECT3_X(rectangle3_xs[1577]), .RECT3_Y(rectangle3_ys[1577]), .RECT3_WIDTH(rectangle3_widths[1577]), .RECT3_HEIGHT(rectangle3_heights[1577]), .RECT3_WEIGHT(rectangle3_weights[1577]), .FEAT_THRES(feature_thresholds[1577]), .FEAT_ABOVE(feature_aboves[1577]), .FEAT_BELOW(feature_belows[1577])) ac1577(.scan_win(scan_win1577), .scan_win_std_dev(scan_win_std_dev[1577]), .feature_accum(feature_accums[1577]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1578]), .RECT1_Y(rectangle1_ys[1578]), .RECT1_WIDTH(rectangle1_widths[1578]), .RECT1_HEIGHT(rectangle1_heights[1578]), .RECT1_WEIGHT(rectangle1_weights[1578]), .RECT2_X(rectangle2_xs[1578]), .RECT2_Y(rectangle2_ys[1578]), .RECT2_WIDTH(rectangle2_widths[1578]), .RECT2_HEIGHT(rectangle2_heights[1578]), .RECT2_WEIGHT(rectangle2_weights[1578]), .RECT3_X(rectangle3_xs[1578]), .RECT3_Y(rectangle3_ys[1578]), .RECT3_WIDTH(rectangle3_widths[1578]), .RECT3_HEIGHT(rectangle3_heights[1578]), .RECT3_WEIGHT(rectangle3_weights[1578]), .FEAT_THRES(feature_thresholds[1578]), .FEAT_ABOVE(feature_aboves[1578]), .FEAT_BELOW(feature_belows[1578])) ac1578(.scan_win(scan_win1578), .scan_win_std_dev(scan_win_std_dev[1578]), .feature_accum(feature_accums[1578]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1579]), .RECT1_Y(rectangle1_ys[1579]), .RECT1_WIDTH(rectangle1_widths[1579]), .RECT1_HEIGHT(rectangle1_heights[1579]), .RECT1_WEIGHT(rectangle1_weights[1579]), .RECT2_X(rectangle2_xs[1579]), .RECT2_Y(rectangle2_ys[1579]), .RECT2_WIDTH(rectangle2_widths[1579]), .RECT2_HEIGHT(rectangle2_heights[1579]), .RECT2_WEIGHT(rectangle2_weights[1579]), .RECT3_X(rectangle3_xs[1579]), .RECT3_Y(rectangle3_ys[1579]), .RECT3_WIDTH(rectangle3_widths[1579]), .RECT3_HEIGHT(rectangle3_heights[1579]), .RECT3_WEIGHT(rectangle3_weights[1579]), .FEAT_THRES(feature_thresholds[1579]), .FEAT_ABOVE(feature_aboves[1579]), .FEAT_BELOW(feature_belows[1579])) ac1579(.scan_win(scan_win1579), .scan_win_std_dev(scan_win_std_dev[1579]), .feature_accum(feature_accums[1579]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1580]), .RECT1_Y(rectangle1_ys[1580]), .RECT1_WIDTH(rectangle1_widths[1580]), .RECT1_HEIGHT(rectangle1_heights[1580]), .RECT1_WEIGHT(rectangle1_weights[1580]), .RECT2_X(rectangle2_xs[1580]), .RECT2_Y(rectangle2_ys[1580]), .RECT2_WIDTH(rectangle2_widths[1580]), .RECT2_HEIGHT(rectangle2_heights[1580]), .RECT2_WEIGHT(rectangle2_weights[1580]), .RECT3_X(rectangle3_xs[1580]), .RECT3_Y(rectangle3_ys[1580]), .RECT3_WIDTH(rectangle3_widths[1580]), .RECT3_HEIGHT(rectangle3_heights[1580]), .RECT3_WEIGHT(rectangle3_weights[1580]), .FEAT_THRES(feature_thresholds[1580]), .FEAT_ABOVE(feature_aboves[1580]), .FEAT_BELOW(feature_belows[1580])) ac1580(.scan_win(scan_win1580), .scan_win_std_dev(scan_win_std_dev[1580]), .feature_accum(feature_accums[1580]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1581]), .RECT1_Y(rectangle1_ys[1581]), .RECT1_WIDTH(rectangle1_widths[1581]), .RECT1_HEIGHT(rectangle1_heights[1581]), .RECT1_WEIGHT(rectangle1_weights[1581]), .RECT2_X(rectangle2_xs[1581]), .RECT2_Y(rectangle2_ys[1581]), .RECT2_WIDTH(rectangle2_widths[1581]), .RECT2_HEIGHT(rectangle2_heights[1581]), .RECT2_WEIGHT(rectangle2_weights[1581]), .RECT3_X(rectangle3_xs[1581]), .RECT3_Y(rectangle3_ys[1581]), .RECT3_WIDTH(rectangle3_widths[1581]), .RECT3_HEIGHT(rectangle3_heights[1581]), .RECT3_WEIGHT(rectangle3_weights[1581]), .FEAT_THRES(feature_thresholds[1581]), .FEAT_ABOVE(feature_aboves[1581]), .FEAT_BELOW(feature_belows[1581])) ac1581(.scan_win(scan_win1581), .scan_win_std_dev(scan_win_std_dev[1581]), .feature_accum(feature_accums[1581]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1582]), .RECT1_Y(rectangle1_ys[1582]), .RECT1_WIDTH(rectangle1_widths[1582]), .RECT1_HEIGHT(rectangle1_heights[1582]), .RECT1_WEIGHT(rectangle1_weights[1582]), .RECT2_X(rectangle2_xs[1582]), .RECT2_Y(rectangle2_ys[1582]), .RECT2_WIDTH(rectangle2_widths[1582]), .RECT2_HEIGHT(rectangle2_heights[1582]), .RECT2_WEIGHT(rectangle2_weights[1582]), .RECT3_X(rectangle3_xs[1582]), .RECT3_Y(rectangle3_ys[1582]), .RECT3_WIDTH(rectangle3_widths[1582]), .RECT3_HEIGHT(rectangle3_heights[1582]), .RECT3_WEIGHT(rectangle3_weights[1582]), .FEAT_THRES(feature_thresholds[1582]), .FEAT_ABOVE(feature_aboves[1582]), .FEAT_BELOW(feature_belows[1582])) ac1582(.scan_win(scan_win1582), .scan_win_std_dev(scan_win_std_dev[1582]), .feature_accum(feature_accums[1582]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1583]), .RECT1_Y(rectangle1_ys[1583]), .RECT1_WIDTH(rectangle1_widths[1583]), .RECT1_HEIGHT(rectangle1_heights[1583]), .RECT1_WEIGHT(rectangle1_weights[1583]), .RECT2_X(rectangle2_xs[1583]), .RECT2_Y(rectangle2_ys[1583]), .RECT2_WIDTH(rectangle2_widths[1583]), .RECT2_HEIGHT(rectangle2_heights[1583]), .RECT2_WEIGHT(rectangle2_weights[1583]), .RECT3_X(rectangle3_xs[1583]), .RECT3_Y(rectangle3_ys[1583]), .RECT3_WIDTH(rectangle3_widths[1583]), .RECT3_HEIGHT(rectangle3_heights[1583]), .RECT3_WEIGHT(rectangle3_weights[1583]), .FEAT_THRES(feature_thresholds[1583]), .FEAT_ABOVE(feature_aboves[1583]), .FEAT_BELOW(feature_belows[1583])) ac1583(.scan_win(scan_win1583), .scan_win_std_dev(scan_win_std_dev[1583]), .feature_accum(feature_accums[1583]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1584]), .RECT1_Y(rectangle1_ys[1584]), .RECT1_WIDTH(rectangle1_widths[1584]), .RECT1_HEIGHT(rectangle1_heights[1584]), .RECT1_WEIGHT(rectangle1_weights[1584]), .RECT2_X(rectangle2_xs[1584]), .RECT2_Y(rectangle2_ys[1584]), .RECT2_WIDTH(rectangle2_widths[1584]), .RECT2_HEIGHT(rectangle2_heights[1584]), .RECT2_WEIGHT(rectangle2_weights[1584]), .RECT3_X(rectangle3_xs[1584]), .RECT3_Y(rectangle3_ys[1584]), .RECT3_WIDTH(rectangle3_widths[1584]), .RECT3_HEIGHT(rectangle3_heights[1584]), .RECT3_WEIGHT(rectangle3_weights[1584]), .FEAT_THRES(feature_thresholds[1584]), .FEAT_ABOVE(feature_aboves[1584]), .FEAT_BELOW(feature_belows[1584])) ac1584(.scan_win(scan_win1584), .scan_win_std_dev(scan_win_std_dev[1584]), .feature_accum(feature_accums[1584]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1585]), .RECT1_Y(rectangle1_ys[1585]), .RECT1_WIDTH(rectangle1_widths[1585]), .RECT1_HEIGHT(rectangle1_heights[1585]), .RECT1_WEIGHT(rectangle1_weights[1585]), .RECT2_X(rectangle2_xs[1585]), .RECT2_Y(rectangle2_ys[1585]), .RECT2_WIDTH(rectangle2_widths[1585]), .RECT2_HEIGHT(rectangle2_heights[1585]), .RECT2_WEIGHT(rectangle2_weights[1585]), .RECT3_X(rectangle3_xs[1585]), .RECT3_Y(rectangle3_ys[1585]), .RECT3_WIDTH(rectangle3_widths[1585]), .RECT3_HEIGHT(rectangle3_heights[1585]), .RECT3_WEIGHT(rectangle3_weights[1585]), .FEAT_THRES(feature_thresholds[1585]), .FEAT_ABOVE(feature_aboves[1585]), .FEAT_BELOW(feature_belows[1585])) ac1585(.scan_win(scan_win1585), .scan_win_std_dev(scan_win_std_dev[1585]), .feature_accum(feature_accums[1585]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1586]), .RECT1_Y(rectangle1_ys[1586]), .RECT1_WIDTH(rectangle1_widths[1586]), .RECT1_HEIGHT(rectangle1_heights[1586]), .RECT1_WEIGHT(rectangle1_weights[1586]), .RECT2_X(rectangle2_xs[1586]), .RECT2_Y(rectangle2_ys[1586]), .RECT2_WIDTH(rectangle2_widths[1586]), .RECT2_HEIGHT(rectangle2_heights[1586]), .RECT2_WEIGHT(rectangle2_weights[1586]), .RECT3_X(rectangle3_xs[1586]), .RECT3_Y(rectangle3_ys[1586]), .RECT3_WIDTH(rectangle3_widths[1586]), .RECT3_HEIGHT(rectangle3_heights[1586]), .RECT3_WEIGHT(rectangle3_weights[1586]), .FEAT_THRES(feature_thresholds[1586]), .FEAT_ABOVE(feature_aboves[1586]), .FEAT_BELOW(feature_belows[1586])) ac1586(.scan_win(scan_win1586), .scan_win_std_dev(scan_win_std_dev[1586]), .feature_accum(feature_accums[1586]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1587]), .RECT1_Y(rectangle1_ys[1587]), .RECT1_WIDTH(rectangle1_widths[1587]), .RECT1_HEIGHT(rectangle1_heights[1587]), .RECT1_WEIGHT(rectangle1_weights[1587]), .RECT2_X(rectangle2_xs[1587]), .RECT2_Y(rectangle2_ys[1587]), .RECT2_WIDTH(rectangle2_widths[1587]), .RECT2_HEIGHT(rectangle2_heights[1587]), .RECT2_WEIGHT(rectangle2_weights[1587]), .RECT3_X(rectangle3_xs[1587]), .RECT3_Y(rectangle3_ys[1587]), .RECT3_WIDTH(rectangle3_widths[1587]), .RECT3_HEIGHT(rectangle3_heights[1587]), .RECT3_WEIGHT(rectangle3_weights[1587]), .FEAT_THRES(feature_thresholds[1587]), .FEAT_ABOVE(feature_aboves[1587]), .FEAT_BELOW(feature_belows[1587])) ac1587(.scan_win(scan_win1587), .scan_win_std_dev(scan_win_std_dev[1587]), .feature_accum(feature_accums[1587]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1588]), .RECT1_Y(rectangle1_ys[1588]), .RECT1_WIDTH(rectangle1_widths[1588]), .RECT1_HEIGHT(rectangle1_heights[1588]), .RECT1_WEIGHT(rectangle1_weights[1588]), .RECT2_X(rectangle2_xs[1588]), .RECT2_Y(rectangle2_ys[1588]), .RECT2_WIDTH(rectangle2_widths[1588]), .RECT2_HEIGHT(rectangle2_heights[1588]), .RECT2_WEIGHT(rectangle2_weights[1588]), .RECT3_X(rectangle3_xs[1588]), .RECT3_Y(rectangle3_ys[1588]), .RECT3_WIDTH(rectangle3_widths[1588]), .RECT3_HEIGHT(rectangle3_heights[1588]), .RECT3_WEIGHT(rectangle3_weights[1588]), .FEAT_THRES(feature_thresholds[1588]), .FEAT_ABOVE(feature_aboves[1588]), .FEAT_BELOW(feature_belows[1588])) ac1588(.scan_win(scan_win1588), .scan_win_std_dev(scan_win_std_dev[1588]), .feature_accum(feature_accums[1588]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1589]), .RECT1_Y(rectangle1_ys[1589]), .RECT1_WIDTH(rectangle1_widths[1589]), .RECT1_HEIGHT(rectangle1_heights[1589]), .RECT1_WEIGHT(rectangle1_weights[1589]), .RECT2_X(rectangle2_xs[1589]), .RECT2_Y(rectangle2_ys[1589]), .RECT2_WIDTH(rectangle2_widths[1589]), .RECT2_HEIGHT(rectangle2_heights[1589]), .RECT2_WEIGHT(rectangle2_weights[1589]), .RECT3_X(rectangle3_xs[1589]), .RECT3_Y(rectangle3_ys[1589]), .RECT3_WIDTH(rectangle3_widths[1589]), .RECT3_HEIGHT(rectangle3_heights[1589]), .RECT3_WEIGHT(rectangle3_weights[1589]), .FEAT_THRES(feature_thresholds[1589]), .FEAT_ABOVE(feature_aboves[1589]), .FEAT_BELOW(feature_belows[1589])) ac1589(.scan_win(scan_win1589), .scan_win_std_dev(scan_win_std_dev[1589]), .feature_accum(feature_accums[1589]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1590]), .RECT1_Y(rectangle1_ys[1590]), .RECT1_WIDTH(rectangle1_widths[1590]), .RECT1_HEIGHT(rectangle1_heights[1590]), .RECT1_WEIGHT(rectangle1_weights[1590]), .RECT2_X(rectangle2_xs[1590]), .RECT2_Y(rectangle2_ys[1590]), .RECT2_WIDTH(rectangle2_widths[1590]), .RECT2_HEIGHT(rectangle2_heights[1590]), .RECT2_WEIGHT(rectangle2_weights[1590]), .RECT3_X(rectangle3_xs[1590]), .RECT3_Y(rectangle3_ys[1590]), .RECT3_WIDTH(rectangle3_widths[1590]), .RECT3_HEIGHT(rectangle3_heights[1590]), .RECT3_WEIGHT(rectangle3_weights[1590]), .FEAT_THRES(feature_thresholds[1590]), .FEAT_ABOVE(feature_aboves[1590]), .FEAT_BELOW(feature_belows[1590])) ac1590(.scan_win(scan_win1590), .scan_win_std_dev(scan_win_std_dev[1590]), .feature_accum(feature_accums[1590]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1591]), .RECT1_Y(rectangle1_ys[1591]), .RECT1_WIDTH(rectangle1_widths[1591]), .RECT1_HEIGHT(rectangle1_heights[1591]), .RECT1_WEIGHT(rectangle1_weights[1591]), .RECT2_X(rectangle2_xs[1591]), .RECT2_Y(rectangle2_ys[1591]), .RECT2_WIDTH(rectangle2_widths[1591]), .RECT2_HEIGHT(rectangle2_heights[1591]), .RECT2_WEIGHT(rectangle2_weights[1591]), .RECT3_X(rectangle3_xs[1591]), .RECT3_Y(rectangle3_ys[1591]), .RECT3_WIDTH(rectangle3_widths[1591]), .RECT3_HEIGHT(rectangle3_heights[1591]), .RECT3_WEIGHT(rectangle3_weights[1591]), .FEAT_THRES(feature_thresholds[1591]), .FEAT_ABOVE(feature_aboves[1591]), .FEAT_BELOW(feature_belows[1591])) ac1591(.scan_win(scan_win1591), .scan_win_std_dev(scan_win_std_dev[1591]), .feature_accum(feature_accums[1591]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1592]), .RECT1_Y(rectangle1_ys[1592]), .RECT1_WIDTH(rectangle1_widths[1592]), .RECT1_HEIGHT(rectangle1_heights[1592]), .RECT1_WEIGHT(rectangle1_weights[1592]), .RECT2_X(rectangle2_xs[1592]), .RECT2_Y(rectangle2_ys[1592]), .RECT2_WIDTH(rectangle2_widths[1592]), .RECT2_HEIGHT(rectangle2_heights[1592]), .RECT2_WEIGHT(rectangle2_weights[1592]), .RECT3_X(rectangle3_xs[1592]), .RECT3_Y(rectangle3_ys[1592]), .RECT3_WIDTH(rectangle3_widths[1592]), .RECT3_HEIGHT(rectangle3_heights[1592]), .RECT3_WEIGHT(rectangle3_weights[1592]), .FEAT_THRES(feature_thresholds[1592]), .FEAT_ABOVE(feature_aboves[1592]), .FEAT_BELOW(feature_belows[1592])) ac1592(.scan_win(scan_win1592), .scan_win_std_dev(scan_win_std_dev[1592]), .feature_accum(feature_accums[1592]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1593]), .RECT1_Y(rectangle1_ys[1593]), .RECT1_WIDTH(rectangle1_widths[1593]), .RECT1_HEIGHT(rectangle1_heights[1593]), .RECT1_WEIGHT(rectangle1_weights[1593]), .RECT2_X(rectangle2_xs[1593]), .RECT2_Y(rectangle2_ys[1593]), .RECT2_WIDTH(rectangle2_widths[1593]), .RECT2_HEIGHT(rectangle2_heights[1593]), .RECT2_WEIGHT(rectangle2_weights[1593]), .RECT3_X(rectangle3_xs[1593]), .RECT3_Y(rectangle3_ys[1593]), .RECT3_WIDTH(rectangle3_widths[1593]), .RECT3_HEIGHT(rectangle3_heights[1593]), .RECT3_WEIGHT(rectangle3_weights[1593]), .FEAT_THRES(feature_thresholds[1593]), .FEAT_ABOVE(feature_aboves[1593]), .FEAT_BELOW(feature_belows[1593])) ac1593(.scan_win(scan_win1593), .scan_win_std_dev(scan_win_std_dev[1593]), .feature_accum(feature_accums[1593]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1594]), .RECT1_Y(rectangle1_ys[1594]), .RECT1_WIDTH(rectangle1_widths[1594]), .RECT1_HEIGHT(rectangle1_heights[1594]), .RECT1_WEIGHT(rectangle1_weights[1594]), .RECT2_X(rectangle2_xs[1594]), .RECT2_Y(rectangle2_ys[1594]), .RECT2_WIDTH(rectangle2_widths[1594]), .RECT2_HEIGHT(rectangle2_heights[1594]), .RECT2_WEIGHT(rectangle2_weights[1594]), .RECT3_X(rectangle3_xs[1594]), .RECT3_Y(rectangle3_ys[1594]), .RECT3_WIDTH(rectangle3_widths[1594]), .RECT3_HEIGHT(rectangle3_heights[1594]), .RECT3_WEIGHT(rectangle3_weights[1594]), .FEAT_THRES(feature_thresholds[1594]), .FEAT_ABOVE(feature_aboves[1594]), .FEAT_BELOW(feature_belows[1594])) ac1594(.scan_win(scan_win1594), .scan_win_std_dev(scan_win_std_dev[1594]), .feature_accum(feature_accums[1594]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1595]), .RECT1_Y(rectangle1_ys[1595]), .RECT1_WIDTH(rectangle1_widths[1595]), .RECT1_HEIGHT(rectangle1_heights[1595]), .RECT1_WEIGHT(rectangle1_weights[1595]), .RECT2_X(rectangle2_xs[1595]), .RECT2_Y(rectangle2_ys[1595]), .RECT2_WIDTH(rectangle2_widths[1595]), .RECT2_HEIGHT(rectangle2_heights[1595]), .RECT2_WEIGHT(rectangle2_weights[1595]), .RECT3_X(rectangle3_xs[1595]), .RECT3_Y(rectangle3_ys[1595]), .RECT3_WIDTH(rectangle3_widths[1595]), .RECT3_HEIGHT(rectangle3_heights[1595]), .RECT3_WEIGHT(rectangle3_weights[1595]), .FEAT_THRES(feature_thresholds[1595]), .FEAT_ABOVE(feature_aboves[1595]), .FEAT_BELOW(feature_belows[1595])) ac1595(.scan_win(scan_win1595), .scan_win_std_dev(scan_win_std_dev[1595]), .feature_accum(feature_accums[1595]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1596]), .RECT1_Y(rectangle1_ys[1596]), .RECT1_WIDTH(rectangle1_widths[1596]), .RECT1_HEIGHT(rectangle1_heights[1596]), .RECT1_WEIGHT(rectangle1_weights[1596]), .RECT2_X(rectangle2_xs[1596]), .RECT2_Y(rectangle2_ys[1596]), .RECT2_WIDTH(rectangle2_widths[1596]), .RECT2_HEIGHT(rectangle2_heights[1596]), .RECT2_WEIGHT(rectangle2_weights[1596]), .RECT3_X(rectangle3_xs[1596]), .RECT3_Y(rectangle3_ys[1596]), .RECT3_WIDTH(rectangle3_widths[1596]), .RECT3_HEIGHT(rectangle3_heights[1596]), .RECT3_WEIGHT(rectangle3_weights[1596]), .FEAT_THRES(feature_thresholds[1596]), .FEAT_ABOVE(feature_aboves[1596]), .FEAT_BELOW(feature_belows[1596])) ac1596(.scan_win(scan_win1596), .scan_win_std_dev(scan_win_std_dev[1596]), .feature_accum(feature_accums[1596]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1597]), .RECT1_Y(rectangle1_ys[1597]), .RECT1_WIDTH(rectangle1_widths[1597]), .RECT1_HEIGHT(rectangle1_heights[1597]), .RECT1_WEIGHT(rectangle1_weights[1597]), .RECT2_X(rectangle2_xs[1597]), .RECT2_Y(rectangle2_ys[1597]), .RECT2_WIDTH(rectangle2_widths[1597]), .RECT2_HEIGHT(rectangle2_heights[1597]), .RECT2_WEIGHT(rectangle2_weights[1597]), .RECT3_X(rectangle3_xs[1597]), .RECT3_Y(rectangle3_ys[1597]), .RECT3_WIDTH(rectangle3_widths[1597]), .RECT3_HEIGHT(rectangle3_heights[1597]), .RECT3_WEIGHT(rectangle3_weights[1597]), .FEAT_THRES(feature_thresholds[1597]), .FEAT_ABOVE(feature_aboves[1597]), .FEAT_BELOW(feature_belows[1597])) ac1597(.scan_win(scan_win1597), .scan_win_std_dev(scan_win_std_dev[1597]), .feature_accum(feature_accums[1597]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1598]), .RECT1_Y(rectangle1_ys[1598]), .RECT1_WIDTH(rectangle1_widths[1598]), .RECT1_HEIGHT(rectangle1_heights[1598]), .RECT1_WEIGHT(rectangle1_weights[1598]), .RECT2_X(rectangle2_xs[1598]), .RECT2_Y(rectangle2_ys[1598]), .RECT2_WIDTH(rectangle2_widths[1598]), .RECT2_HEIGHT(rectangle2_heights[1598]), .RECT2_WEIGHT(rectangle2_weights[1598]), .RECT3_X(rectangle3_xs[1598]), .RECT3_Y(rectangle3_ys[1598]), .RECT3_WIDTH(rectangle3_widths[1598]), .RECT3_HEIGHT(rectangle3_heights[1598]), .RECT3_WEIGHT(rectangle3_weights[1598]), .FEAT_THRES(feature_thresholds[1598]), .FEAT_ABOVE(feature_aboves[1598]), .FEAT_BELOW(feature_belows[1598])) ac1598(.scan_win(scan_win1598), .scan_win_std_dev(scan_win_std_dev[1598]), .feature_accum(feature_accums[1598]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1599]), .RECT1_Y(rectangle1_ys[1599]), .RECT1_WIDTH(rectangle1_widths[1599]), .RECT1_HEIGHT(rectangle1_heights[1599]), .RECT1_WEIGHT(rectangle1_weights[1599]), .RECT2_X(rectangle2_xs[1599]), .RECT2_Y(rectangle2_ys[1599]), .RECT2_WIDTH(rectangle2_widths[1599]), .RECT2_HEIGHT(rectangle2_heights[1599]), .RECT2_WEIGHT(rectangle2_weights[1599]), .RECT3_X(rectangle3_xs[1599]), .RECT3_Y(rectangle3_ys[1599]), .RECT3_WIDTH(rectangle3_widths[1599]), .RECT3_HEIGHT(rectangle3_heights[1599]), .RECT3_WEIGHT(rectangle3_weights[1599]), .FEAT_THRES(feature_thresholds[1599]), .FEAT_ABOVE(feature_aboves[1599]), .FEAT_BELOW(feature_belows[1599])) ac1599(.scan_win(scan_win1599), .scan_win_std_dev(scan_win_std_dev[1599]), .feature_accum(feature_accums[1599]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1600]), .RECT1_Y(rectangle1_ys[1600]), .RECT1_WIDTH(rectangle1_widths[1600]), .RECT1_HEIGHT(rectangle1_heights[1600]), .RECT1_WEIGHT(rectangle1_weights[1600]), .RECT2_X(rectangle2_xs[1600]), .RECT2_Y(rectangle2_ys[1600]), .RECT2_WIDTH(rectangle2_widths[1600]), .RECT2_HEIGHT(rectangle2_heights[1600]), .RECT2_WEIGHT(rectangle2_weights[1600]), .RECT3_X(rectangle3_xs[1600]), .RECT3_Y(rectangle3_ys[1600]), .RECT3_WIDTH(rectangle3_widths[1600]), .RECT3_HEIGHT(rectangle3_heights[1600]), .RECT3_WEIGHT(rectangle3_weights[1600]), .FEAT_THRES(feature_thresholds[1600]), .FEAT_ABOVE(feature_aboves[1600]), .FEAT_BELOW(feature_belows[1600])) ac1600(.scan_win(scan_win1600), .scan_win_std_dev(scan_win_std_dev[1600]), .feature_accum(feature_accums[1600]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1601]), .RECT1_Y(rectangle1_ys[1601]), .RECT1_WIDTH(rectangle1_widths[1601]), .RECT1_HEIGHT(rectangle1_heights[1601]), .RECT1_WEIGHT(rectangle1_weights[1601]), .RECT2_X(rectangle2_xs[1601]), .RECT2_Y(rectangle2_ys[1601]), .RECT2_WIDTH(rectangle2_widths[1601]), .RECT2_HEIGHT(rectangle2_heights[1601]), .RECT2_WEIGHT(rectangle2_weights[1601]), .RECT3_X(rectangle3_xs[1601]), .RECT3_Y(rectangle3_ys[1601]), .RECT3_WIDTH(rectangle3_widths[1601]), .RECT3_HEIGHT(rectangle3_heights[1601]), .RECT3_WEIGHT(rectangle3_weights[1601]), .FEAT_THRES(feature_thresholds[1601]), .FEAT_ABOVE(feature_aboves[1601]), .FEAT_BELOW(feature_belows[1601])) ac1601(.scan_win(scan_win1601), .scan_win_std_dev(scan_win_std_dev[1601]), .feature_accum(feature_accums[1601]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1602]), .RECT1_Y(rectangle1_ys[1602]), .RECT1_WIDTH(rectangle1_widths[1602]), .RECT1_HEIGHT(rectangle1_heights[1602]), .RECT1_WEIGHT(rectangle1_weights[1602]), .RECT2_X(rectangle2_xs[1602]), .RECT2_Y(rectangle2_ys[1602]), .RECT2_WIDTH(rectangle2_widths[1602]), .RECT2_HEIGHT(rectangle2_heights[1602]), .RECT2_WEIGHT(rectangle2_weights[1602]), .RECT3_X(rectangle3_xs[1602]), .RECT3_Y(rectangle3_ys[1602]), .RECT3_WIDTH(rectangle3_widths[1602]), .RECT3_HEIGHT(rectangle3_heights[1602]), .RECT3_WEIGHT(rectangle3_weights[1602]), .FEAT_THRES(feature_thresholds[1602]), .FEAT_ABOVE(feature_aboves[1602]), .FEAT_BELOW(feature_belows[1602])) ac1602(.scan_win(scan_win1602), .scan_win_std_dev(scan_win_std_dev[1602]), .feature_accum(feature_accums[1602]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1603]), .RECT1_Y(rectangle1_ys[1603]), .RECT1_WIDTH(rectangle1_widths[1603]), .RECT1_HEIGHT(rectangle1_heights[1603]), .RECT1_WEIGHT(rectangle1_weights[1603]), .RECT2_X(rectangle2_xs[1603]), .RECT2_Y(rectangle2_ys[1603]), .RECT2_WIDTH(rectangle2_widths[1603]), .RECT2_HEIGHT(rectangle2_heights[1603]), .RECT2_WEIGHT(rectangle2_weights[1603]), .RECT3_X(rectangle3_xs[1603]), .RECT3_Y(rectangle3_ys[1603]), .RECT3_WIDTH(rectangle3_widths[1603]), .RECT3_HEIGHT(rectangle3_heights[1603]), .RECT3_WEIGHT(rectangle3_weights[1603]), .FEAT_THRES(feature_thresholds[1603]), .FEAT_ABOVE(feature_aboves[1603]), .FEAT_BELOW(feature_belows[1603])) ac1603(.scan_win(scan_win1603), .scan_win_std_dev(scan_win_std_dev[1603]), .feature_accum(feature_accums[1603]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1604]), .RECT1_Y(rectangle1_ys[1604]), .RECT1_WIDTH(rectangle1_widths[1604]), .RECT1_HEIGHT(rectangle1_heights[1604]), .RECT1_WEIGHT(rectangle1_weights[1604]), .RECT2_X(rectangle2_xs[1604]), .RECT2_Y(rectangle2_ys[1604]), .RECT2_WIDTH(rectangle2_widths[1604]), .RECT2_HEIGHT(rectangle2_heights[1604]), .RECT2_WEIGHT(rectangle2_weights[1604]), .RECT3_X(rectangle3_xs[1604]), .RECT3_Y(rectangle3_ys[1604]), .RECT3_WIDTH(rectangle3_widths[1604]), .RECT3_HEIGHT(rectangle3_heights[1604]), .RECT3_WEIGHT(rectangle3_weights[1604]), .FEAT_THRES(feature_thresholds[1604]), .FEAT_ABOVE(feature_aboves[1604]), .FEAT_BELOW(feature_belows[1604])) ac1604(.scan_win(scan_win1604), .scan_win_std_dev(scan_win_std_dev[1604]), .feature_accum(feature_accums[1604]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1605]), .RECT1_Y(rectangle1_ys[1605]), .RECT1_WIDTH(rectangle1_widths[1605]), .RECT1_HEIGHT(rectangle1_heights[1605]), .RECT1_WEIGHT(rectangle1_weights[1605]), .RECT2_X(rectangle2_xs[1605]), .RECT2_Y(rectangle2_ys[1605]), .RECT2_WIDTH(rectangle2_widths[1605]), .RECT2_HEIGHT(rectangle2_heights[1605]), .RECT2_WEIGHT(rectangle2_weights[1605]), .RECT3_X(rectangle3_xs[1605]), .RECT3_Y(rectangle3_ys[1605]), .RECT3_WIDTH(rectangle3_widths[1605]), .RECT3_HEIGHT(rectangle3_heights[1605]), .RECT3_WEIGHT(rectangle3_weights[1605]), .FEAT_THRES(feature_thresholds[1605]), .FEAT_ABOVE(feature_aboves[1605]), .FEAT_BELOW(feature_belows[1605])) ac1605(.scan_win(scan_win1605), .scan_win_std_dev(scan_win_std_dev[1605]), .feature_accum(feature_accums[1605]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1606]), .RECT1_Y(rectangle1_ys[1606]), .RECT1_WIDTH(rectangle1_widths[1606]), .RECT1_HEIGHT(rectangle1_heights[1606]), .RECT1_WEIGHT(rectangle1_weights[1606]), .RECT2_X(rectangle2_xs[1606]), .RECT2_Y(rectangle2_ys[1606]), .RECT2_WIDTH(rectangle2_widths[1606]), .RECT2_HEIGHT(rectangle2_heights[1606]), .RECT2_WEIGHT(rectangle2_weights[1606]), .RECT3_X(rectangle3_xs[1606]), .RECT3_Y(rectangle3_ys[1606]), .RECT3_WIDTH(rectangle3_widths[1606]), .RECT3_HEIGHT(rectangle3_heights[1606]), .RECT3_WEIGHT(rectangle3_weights[1606]), .FEAT_THRES(feature_thresholds[1606]), .FEAT_ABOVE(feature_aboves[1606]), .FEAT_BELOW(feature_belows[1606])) ac1606(.scan_win(scan_win1606), .scan_win_std_dev(scan_win_std_dev[1606]), .feature_accum(feature_accums[1606]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1607]), .RECT1_Y(rectangle1_ys[1607]), .RECT1_WIDTH(rectangle1_widths[1607]), .RECT1_HEIGHT(rectangle1_heights[1607]), .RECT1_WEIGHT(rectangle1_weights[1607]), .RECT2_X(rectangle2_xs[1607]), .RECT2_Y(rectangle2_ys[1607]), .RECT2_WIDTH(rectangle2_widths[1607]), .RECT2_HEIGHT(rectangle2_heights[1607]), .RECT2_WEIGHT(rectangle2_weights[1607]), .RECT3_X(rectangle3_xs[1607]), .RECT3_Y(rectangle3_ys[1607]), .RECT3_WIDTH(rectangle3_widths[1607]), .RECT3_HEIGHT(rectangle3_heights[1607]), .RECT3_WEIGHT(rectangle3_weights[1607]), .FEAT_THRES(feature_thresholds[1607]), .FEAT_ABOVE(feature_aboves[1607]), .FEAT_BELOW(feature_belows[1607])) ac1607(.scan_win(scan_win1607), .scan_win_std_dev(scan_win_std_dev[1607]), .feature_accum(feature_accums[1607]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1608]), .RECT1_Y(rectangle1_ys[1608]), .RECT1_WIDTH(rectangle1_widths[1608]), .RECT1_HEIGHT(rectangle1_heights[1608]), .RECT1_WEIGHT(rectangle1_weights[1608]), .RECT2_X(rectangle2_xs[1608]), .RECT2_Y(rectangle2_ys[1608]), .RECT2_WIDTH(rectangle2_widths[1608]), .RECT2_HEIGHT(rectangle2_heights[1608]), .RECT2_WEIGHT(rectangle2_weights[1608]), .RECT3_X(rectangle3_xs[1608]), .RECT3_Y(rectangle3_ys[1608]), .RECT3_WIDTH(rectangle3_widths[1608]), .RECT3_HEIGHT(rectangle3_heights[1608]), .RECT3_WEIGHT(rectangle3_weights[1608]), .FEAT_THRES(feature_thresholds[1608]), .FEAT_ABOVE(feature_aboves[1608]), .FEAT_BELOW(feature_belows[1608])) ac1608(.scan_win(scan_win1608), .scan_win_std_dev(scan_win_std_dev[1608]), .feature_accum(feature_accums[1608]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1609]), .RECT1_Y(rectangle1_ys[1609]), .RECT1_WIDTH(rectangle1_widths[1609]), .RECT1_HEIGHT(rectangle1_heights[1609]), .RECT1_WEIGHT(rectangle1_weights[1609]), .RECT2_X(rectangle2_xs[1609]), .RECT2_Y(rectangle2_ys[1609]), .RECT2_WIDTH(rectangle2_widths[1609]), .RECT2_HEIGHT(rectangle2_heights[1609]), .RECT2_WEIGHT(rectangle2_weights[1609]), .RECT3_X(rectangle3_xs[1609]), .RECT3_Y(rectangle3_ys[1609]), .RECT3_WIDTH(rectangle3_widths[1609]), .RECT3_HEIGHT(rectangle3_heights[1609]), .RECT3_WEIGHT(rectangle3_weights[1609]), .FEAT_THRES(feature_thresholds[1609]), .FEAT_ABOVE(feature_aboves[1609]), .FEAT_BELOW(feature_belows[1609])) ac1609(.scan_win(scan_win1609), .scan_win_std_dev(scan_win_std_dev[1609]), .feature_accum(feature_accums[1609]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1610]), .RECT1_Y(rectangle1_ys[1610]), .RECT1_WIDTH(rectangle1_widths[1610]), .RECT1_HEIGHT(rectangle1_heights[1610]), .RECT1_WEIGHT(rectangle1_weights[1610]), .RECT2_X(rectangle2_xs[1610]), .RECT2_Y(rectangle2_ys[1610]), .RECT2_WIDTH(rectangle2_widths[1610]), .RECT2_HEIGHT(rectangle2_heights[1610]), .RECT2_WEIGHT(rectangle2_weights[1610]), .RECT3_X(rectangle3_xs[1610]), .RECT3_Y(rectangle3_ys[1610]), .RECT3_WIDTH(rectangle3_widths[1610]), .RECT3_HEIGHT(rectangle3_heights[1610]), .RECT3_WEIGHT(rectangle3_weights[1610]), .FEAT_THRES(feature_thresholds[1610]), .FEAT_ABOVE(feature_aboves[1610]), .FEAT_BELOW(feature_belows[1610])) ac1610(.scan_win(scan_win1610), .scan_win_std_dev(scan_win_std_dev[1610]), .feature_accum(feature_accums[1610]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1611]), .RECT1_Y(rectangle1_ys[1611]), .RECT1_WIDTH(rectangle1_widths[1611]), .RECT1_HEIGHT(rectangle1_heights[1611]), .RECT1_WEIGHT(rectangle1_weights[1611]), .RECT2_X(rectangle2_xs[1611]), .RECT2_Y(rectangle2_ys[1611]), .RECT2_WIDTH(rectangle2_widths[1611]), .RECT2_HEIGHT(rectangle2_heights[1611]), .RECT2_WEIGHT(rectangle2_weights[1611]), .RECT3_X(rectangle3_xs[1611]), .RECT3_Y(rectangle3_ys[1611]), .RECT3_WIDTH(rectangle3_widths[1611]), .RECT3_HEIGHT(rectangle3_heights[1611]), .RECT3_WEIGHT(rectangle3_weights[1611]), .FEAT_THRES(feature_thresholds[1611]), .FEAT_ABOVE(feature_aboves[1611]), .FEAT_BELOW(feature_belows[1611])) ac1611(.scan_win(scan_win1611), .scan_win_std_dev(scan_win_std_dev[1611]), .feature_accum(feature_accums[1611]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1612]), .RECT1_Y(rectangle1_ys[1612]), .RECT1_WIDTH(rectangle1_widths[1612]), .RECT1_HEIGHT(rectangle1_heights[1612]), .RECT1_WEIGHT(rectangle1_weights[1612]), .RECT2_X(rectangle2_xs[1612]), .RECT2_Y(rectangle2_ys[1612]), .RECT2_WIDTH(rectangle2_widths[1612]), .RECT2_HEIGHT(rectangle2_heights[1612]), .RECT2_WEIGHT(rectangle2_weights[1612]), .RECT3_X(rectangle3_xs[1612]), .RECT3_Y(rectangle3_ys[1612]), .RECT3_WIDTH(rectangle3_widths[1612]), .RECT3_HEIGHT(rectangle3_heights[1612]), .RECT3_WEIGHT(rectangle3_weights[1612]), .FEAT_THRES(feature_thresholds[1612]), .FEAT_ABOVE(feature_aboves[1612]), .FEAT_BELOW(feature_belows[1612])) ac1612(.scan_win(scan_win1612), .scan_win_std_dev(scan_win_std_dev[1612]), .feature_accum(feature_accums[1612]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1613]), .RECT1_Y(rectangle1_ys[1613]), .RECT1_WIDTH(rectangle1_widths[1613]), .RECT1_HEIGHT(rectangle1_heights[1613]), .RECT1_WEIGHT(rectangle1_weights[1613]), .RECT2_X(rectangle2_xs[1613]), .RECT2_Y(rectangle2_ys[1613]), .RECT2_WIDTH(rectangle2_widths[1613]), .RECT2_HEIGHT(rectangle2_heights[1613]), .RECT2_WEIGHT(rectangle2_weights[1613]), .RECT3_X(rectangle3_xs[1613]), .RECT3_Y(rectangle3_ys[1613]), .RECT3_WIDTH(rectangle3_widths[1613]), .RECT3_HEIGHT(rectangle3_heights[1613]), .RECT3_WEIGHT(rectangle3_weights[1613]), .FEAT_THRES(feature_thresholds[1613]), .FEAT_ABOVE(feature_aboves[1613]), .FEAT_BELOW(feature_belows[1613])) ac1613(.scan_win(scan_win1613), .scan_win_std_dev(scan_win_std_dev[1613]), .feature_accum(feature_accums[1613]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1614]), .RECT1_Y(rectangle1_ys[1614]), .RECT1_WIDTH(rectangle1_widths[1614]), .RECT1_HEIGHT(rectangle1_heights[1614]), .RECT1_WEIGHT(rectangle1_weights[1614]), .RECT2_X(rectangle2_xs[1614]), .RECT2_Y(rectangle2_ys[1614]), .RECT2_WIDTH(rectangle2_widths[1614]), .RECT2_HEIGHT(rectangle2_heights[1614]), .RECT2_WEIGHT(rectangle2_weights[1614]), .RECT3_X(rectangle3_xs[1614]), .RECT3_Y(rectangle3_ys[1614]), .RECT3_WIDTH(rectangle3_widths[1614]), .RECT3_HEIGHT(rectangle3_heights[1614]), .RECT3_WEIGHT(rectangle3_weights[1614]), .FEAT_THRES(feature_thresholds[1614]), .FEAT_ABOVE(feature_aboves[1614]), .FEAT_BELOW(feature_belows[1614])) ac1614(.scan_win(scan_win1614), .scan_win_std_dev(scan_win_std_dev[1614]), .feature_accum(feature_accums[1614]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1615]), .RECT1_Y(rectangle1_ys[1615]), .RECT1_WIDTH(rectangle1_widths[1615]), .RECT1_HEIGHT(rectangle1_heights[1615]), .RECT1_WEIGHT(rectangle1_weights[1615]), .RECT2_X(rectangle2_xs[1615]), .RECT2_Y(rectangle2_ys[1615]), .RECT2_WIDTH(rectangle2_widths[1615]), .RECT2_HEIGHT(rectangle2_heights[1615]), .RECT2_WEIGHT(rectangle2_weights[1615]), .RECT3_X(rectangle3_xs[1615]), .RECT3_Y(rectangle3_ys[1615]), .RECT3_WIDTH(rectangle3_widths[1615]), .RECT3_HEIGHT(rectangle3_heights[1615]), .RECT3_WEIGHT(rectangle3_weights[1615]), .FEAT_THRES(feature_thresholds[1615]), .FEAT_ABOVE(feature_aboves[1615]), .FEAT_BELOW(feature_belows[1615])) ac1615(.scan_win(scan_win1615), .scan_win_std_dev(scan_win_std_dev[1615]), .feature_accum(feature_accums[1615]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1616]), .RECT1_Y(rectangle1_ys[1616]), .RECT1_WIDTH(rectangle1_widths[1616]), .RECT1_HEIGHT(rectangle1_heights[1616]), .RECT1_WEIGHT(rectangle1_weights[1616]), .RECT2_X(rectangle2_xs[1616]), .RECT2_Y(rectangle2_ys[1616]), .RECT2_WIDTH(rectangle2_widths[1616]), .RECT2_HEIGHT(rectangle2_heights[1616]), .RECT2_WEIGHT(rectangle2_weights[1616]), .RECT3_X(rectangle3_xs[1616]), .RECT3_Y(rectangle3_ys[1616]), .RECT3_WIDTH(rectangle3_widths[1616]), .RECT3_HEIGHT(rectangle3_heights[1616]), .RECT3_WEIGHT(rectangle3_weights[1616]), .FEAT_THRES(feature_thresholds[1616]), .FEAT_ABOVE(feature_aboves[1616]), .FEAT_BELOW(feature_belows[1616])) ac1616(.scan_win(scan_win1616), .scan_win_std_dev(scan_win_std_dev[1616]), .feature_accum(feature_accums[1616]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1617]), .RECT1_Y(rectangle1_ys[1617]), .RECT1_WIDTH(rectangle1_widths[1617]), .RECT1_HEIGHT(rectangle1_heights[1617]), .RECT1_WEIGHT(rectangle1_weights[1617]), .RECT2_X(rectangle2_xs[1617]), .RECT2_Y(rectangle2_ys[1617]), .RECT2_WIDTH(rectangle2_widths[1617]), .RECT2_HEIGHT(rectangle2_heights[1617]), .RECT2_WEIGHT(rectangle2_weights[1617]), .RECT3_X(rectangle3_xs[1617]), .RECT3_Y(rectangle3_ys[1617]), .RECT3_WIDTH(rectangle3_widths[1617]), .RECT3_HEIGHT(rectangle3_heights[1617]), .RECT3_WEIGHT(rectangle3_weights[1617]), .FEAT_THRES(feature_thresholds[1617]), .FEAT_ABOVE(feature_aboves[1617]), .FEAT_BELOW(feature_belows[1617])) ac1617(.scan_win(scan_win1617), .scan_win_std_dev(scan_win_std_dev[1617]), .feature_accum(feature_accums[1617]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1618]), .RECT1_Y(rectangle1_ys[1618]), .RECT1_WIDTH(rectangle1_widths[1618]), .RECT1_HEIGHT(rectangle1_heights[1618]), .RECT1_WEIGHT(rectangle1_weights[1618]), .RECT2_X(rectangle2_xs[1618]), .RECT2_Y(rectangle2_ys[1618]), .RECT2_WIDTH(rectangle2_widths[1618]), .RECT2_HEIGHT(rectangle2_heights[1618]), .RECT2_WEIGHT(rectangle2_weights[1618]), .RECT3_X(rectangle3_xs[1618]), .RECT3_Y(rectangle3_ys[1618]), .RECT3_WIDTH(rectangle3_widths[1618]), .RECT3_HEIGHT(rectangle3_heights[1618]), .RECT3_WEIGHT(rectangle3_weights[1618]), .FEAT_THRES(feature_thresholds[1618]), .FEAT_ABOVE(feature_aboves[1618]), .FEAT_BELOW(feature_belows[1618])) ac1618(.scan_win(scan_win1618), .scan_win_std_dev(scan_win_std_dev[1618]), .feature_accum(feature_accums[1618]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1619]), .RECT1_Y(rectangle1_ys[1619]), .RECT1_WIDTH(rectangle1_widths[1619]), .RECT1_HEIGHT(rectangle1_heights[1619]), .RECT1_WEIGHT(rectangle1_weights[1619]), .RECT2_X(rectangle2_xs[1619]), .RECT2_Y(rectangle2_ys[1619]), .RECT2_WIDTH(rectangle2_widths[1619]), .RECT2_HEIGHT(rectangle2_heights[1619]), .RECT2_WEIGHT(rectangle2_weights[1619]), .RECT3_X(rectangle3_xs[1619]), .RECT3_Y(rectangle3_ys[1619]), .RECT3_WIDTH(rectangle3_widths[1619]), .RECT3_HEIGHT(rectangle3_heights[1619]), .RECT3_WEIGHT(rectangle3_weights[1619]), .FEAT_THRES(feature_thresholds[1619]), .FEAT_ABOVE(feature_aboves[1619]), .FEAT_BELOW(feature_belows[1619])) ac1619(.scan_win(scan_win1619), .scan_win_std_dev(scan_win_std_dev[1619]), .feature_accum(feature_accums[1619]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1620]), .RECT1_Y(rectangle1_ys[1620]), .RECT1_WIDTH(rectangle1_widths[1620]), .RECT1_HEIGHT(rectangle1_heights[1620]), .RECT1_WEIGHT(rectangle1_weights[1620]), .RECT2_X(rectangle2_xs[1620]), .RECT2_Y(rectangle2_ys[1620]), .RECT2_WIDTH(rectangle2_widths[1620]), .RECT2_HEIGHT(rectangle2_heights[1620]), .RECT2_WEIGHT(rectangle2_weights[1620]), .RECT3_X(rectangle3_xs[1620]), .RECT3_Y(rectangle3_ys[1620]), .RECT3_WIDTH(rectangle3_widths[1620]), .RECT3_HEIGHT(rectangle3_heights[1620]), .RECT3_WEIGHT(rectangle3_weights[1620]), .FEAT_THRES(feature_thresholds[1620]), .FEAT_ABOVE(feature_aboves[1620]), .FEAT_BELOW(feature_belows[1620])) ac1620(.scan_win(scan_win1620), .scan_win_std_dev(scan_win_std_dev[1620]), .feature_accum(feature_accums[1620]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1621]), .RECT1_Y(rectangle1_ys[1621]), .RECT1_WIDTH(rectangle1_widths[1621]), .RECT1_HEIGHT(rectangle1_heights[1621]), .RECT1_WEIGHT(rectangle1_weights[1621]), .RECT2_X(rectangle2_xs[1621]), .RECT2_Y(rectangle2_ys[1621]), .RECT2_WIDTH(rectangle2_widths[1621]), .RECT2_HEIGHT(rectangle2_heights[1621]), .RECT2_WEIGHT(rectangle2_weights[1621]), .RECT3_X(rectangle3_xs[1621]), .RECT3_Y(rectangle3_ys[1621]), .RECT3_WIDTH(rectangle3_widths[1621]), .RECT3_HEIGHT(rectangle3_heights[1621]), .RECT3_WEIGHT(rectangle3_weights[1621]), .FEAT_THRES(feature_thresholds[1621]), .FEAT_ABOVE(feature_aboves[1621]), .FEAT_BELOW(feature_belows[1621])) ac1621(.scan_win(scan_win1621), .scan_win_std_dev(scan_win_std_dev[1621]), .feature_accum(feature_accums[1621]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1622]), .RECT1_Y(rectangle1_ys[1622]), .RECT1_WIDTH(rectangle1_widths[1622]), .RECT1_HEIGHT(rectangle1_heights[1622]), .RECT1_WEIGHT(rectangle1_weights[1622]), .RECT2_X(rectangle2_xs[1622]), .RECT2_Y(rectangle2_ys[1622]), .RECT2_WIDTH(rectangle2_widths[1622]), .RECT2_HEIGHT(rectangle2_heights[1622]), .RECT2_WEIGHT(rectangle2_weights[1622]), .RECT3_X(rectangle3_xs[1622]), .RECT3_Y(rectangle3_ys[1622]), .RECT3_WIDTH(rectangle3_widths[1622]), .RECT3_HEIGHT(rectangle3_heights[1622]), .RECT3_WEIGHT(rectangle3_weights[1622]), .FEAT_THRES(feature_thresholds[1622]), .FEAT_ABOVE(feature_aboves[1622]), .FEAT_BELOW(feature_belows[1622])) ac1622(.scan_win(scan_win1622), .scan_win_std_dev(scan_win_std_dev[1622]), .feature_accum(feature_accums[1622]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1623]), .RECT1_Y(rectangle1_ys[1623]), .RECT1_WIDTH(rectangle1_widths[1623]), .RECT1_HEIGHT(rectangle1_heights[1623]), .RECT1_WEIGHT(rectangle1_weights[1623]), .RECT2_X(rectangle2_xs[1623]), .RECT2_Y(rectangle2_ys[1623]), .RECT2_WIDTH(rectangle2_widths[1623]), .RECT2_HEIGHT(rectangle2_heights[1623]), .RECT2_WEIGHT(rectangle2_weights[1623]), .RECT3_X(rectangle3_xs[1623]), .RECT3_Y(rectangle3_ys[1623]), .RECT3_WIDTH(rectangle3_widths[1623]), .RECT3_HEIGHT(rectangle3_heights[1623]), .RECT3_WEIGHT(rectangle3_weights[1623]), .FEAT_THRES(feature_thresholds[1623]), .FEAT_ABOVE(feature_aboves[1623]), .FEAT_BELOW(feature_belows[1623])) ac1623(.scan_win(scan_win1623), .scan_win_std_dev(scan_win_std_dev[1623]), .feature_accum(feature_accums[1623]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1624]), .RECT1_Y(rectangle1_ys[1624]), .RECT1_WIDTH(rectangle1_widths[1624]), .RECT1_HEIGHT(rectangle1_heights[1624]), .RECT1_WEIGHT(rectangle1_weights[1624]), .RECT2_X(rectangle2_xs[1624]), .RECT2_Y(rectangle2_ys[1624]), .RECT2_WIDTH(rectangle2_widths[1624]), .RECT2_HEIGHT(rectangle2_heights[1624]), .RECT2_WEIGHT(rectangle2_weights[1624]), .RECT3_X(rectangle3_xs[1624]), .RECT3_Y(rectangle3_ys[1624]), .RECT3_WIDTH(rectangle3_widths[1624]), .RECT3_HEIGHT(rectangle3_heights[1624]), .RECT3_WEIGHT(rectangle3_weights[1624]), .FEAT_THRES(feature_thresholds[1624]), .FEAT_ABOVE(feature_aboves[1624]), .FEAT_BELOW(feature_belows[1624])) ac1624(.scan_win(scan_win1624), .scan_win_std_dev(scan_win_std_dev[1624]), .feature_accum(feature_accums[1624]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1625]), .RECT1_Y(rectangle1_ys[1625]), .RECT1_WIDTH(rectangle1_widths[1625]), .RECT1_HEIGHT(rectangle1_heights[1625]), .RECT1_WEIGHT(rectangle1_weights[1625]), .RECT2_X(rectangle2_xs[1625]), .RECT2_Y(rectangle2_ys[1625]), .RECT2_WIDTH(rectangle2_widths[1625]), .RECT2_HEIGHT(rectangle2_heights[1625]), .RECT2_WEIGHT(rectangle2_weights[1625]), .RECT3_X(rectangle3_xs[1625]), .RECT3_Y(rectangle3_ys[1625]), .RECT3_WIDTH(rectangle3_widths[1625]), .RECT3_HEIGHT(rectangle3_heights[1625]), .RECT3_WEIGHT(rectangle3_weights[1625]), .FEAT_THRES(feature_thresholds[1625]), .FEAT_ABOVE(feature_aboves[1625]), .FEAT_BELOW(feature_belows[1625])) ac1625(.scan_win(scan_win1625), .scan_win_std_dev(scan_win_std_dev[1625]), .feature_accum(feature_accums[1625]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1626]), .RECT1_Y(rectangle1_ys[1626]), .RECT1_WIDTH(rectangle1_widths[1626]), .RECT1_HEIGHT(rectangle1_heights[1626]), .RECT1_WEIGHT(rectangle1_weights[1626]), .RECT2_X(rectangle2_xs[1626]), .RECT2_Y(rectangle2_ys[1626]), .RECT2_WIDTH(rectangle2_widths[1626]), .RECT2_HEIGHT(rectangle2_heights[1626]), .RECT2_WEIGHT(rectangle2_weights[1626]), .RECT3_X(rectangle3_xs[1626]), .RECT3_Y(rectangle3_ys[1626]), .RECT3_WIDTH(rectangle3_widths[1626]), .RECT3_HEIGHT(rectangle3_heights[1626]), .RECT3_WEIGHT(rectangle3_weights[1626]), .FEAT_THRES(feature_thresholds[1626]), .FEAT_ABOVE(feature_aboves[1626]), .FEAT_BELOW(feature_belows[1626])) ac1626(.scan_win(scan_win1626), .scan_win_std_dev(scan_win_std_dev[1626]), .feature_accum(feature_accums[1626]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1627]), .RECT1_Y(rectangle1_ys[1627]), .RECT1_WIDTH(rectangle1_widths[1627]), .RECT1_HEIGHT(rectangle1_heights[1627]), .RECT1_WEIGHT(rectangle1_weights[1627]), .RECT2_X(rectangle2_xs[1627]), .RECT2_Y(rectangle2_ys[1627]), .RECT2_WIDTH(rectangle2_widths[1627]), .RECT2_HEIGHT(rectangle2_heights[1627]), .RECT2_WEIGHT(rectangle2_weights[1627]), .RECT3_X(rectangle3_xs[1627]), .RECT3_Y(rectangle3_ys[1627]), .RECT3_WIDTH(rectangle3_widths[1627]), .RECT3_HEIGHT(rectangle3_heights[1627]), .RECT3_WEIGHT(rectangle3_weights[1627]), .FEAT_THRES(feature_thresholds[1627]), .FEAT_ABOVE(feature_aboves[1627]), .FEAT_BELOW(feature_belows[1627])) ac1627(.scan_win(scan_win1627), .scan_win_std_dev(scan_win_std_dev[1627]), .feature_accum(feature_accums[1627]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1628]), .RECT1_Y(rectangle1_ys[1628]), .RECT1_WIDTH(rectangle1_widths[1628]), .RECT1_HEIGHT(rectangle1_heights[1628]), .RECT1_WEIGHT(rectangle1_weights[1628]), .RECT2_X(rectangle2_xs[1628]), .RECT2_Y(rectangle2_ys[1628]), .RECT2_WIDTH(rectangle2_widths[1628]), .RECT2_HEIGHT(rectangle2_heights[1628]), .RECT2_WEIGHT(rectangle2_weights[1628]), .RECT3_X(rectangle3_xs[1628]), .RECT3_Y(rectangle3_ys[1628]), .RECT3_WIDTH(rectangle3_widths[1628]), .RECT3_HEIGHT(rectangle3_heights[1628]), .RECT3_WEIGHT(rectangle3_weights[1628]), .FEAT_THRES(feature_thresholds[1628]), .FEAT_ABOVE(feature_aboves[1628]), .FEAT_BELOW(feature_belows[1628])) ac1628(.scan_win(scan_win1628), .scan_win_std_dev(scan_win_std_dev[1628]), .feature_accum(feature_accums[1628]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1629]), .RECT1_Y(rectangle1_ys[1629]), .RECT1_WIDTH(rectangle1_widths[1629]), .RECT1_HEIGHT(rectangle1_heights[1629]), .RECT1_WEIGHT(rectangle1_weights[1629]), .RECT2_X(rectangle2_xs[1629]), .RECT2_Y(rectangle2_ys[1629]), .RECT2_WIDTH(rectangle2_widths[1629]), .RECT2_HEIGHT(rectangle2_heights[1629]), .RECT2_WEIGHT(rectangle2_weights[1629]), .RECT3_X(rectangle3_xs[1629]), .RECT3_Y(rectangle3_ys[1629]), .RECT3_WIDTH(rectangle3_widths[1629]), .RECT3_HEIGHT(rectangle3_heights[1629]), .RECT3_WEIGHT(rectangle3_weights[1629]), .FEAT_THRES(feature_thresholds[1629]), .FEAT_ABOVE(feature_aboves[1629]), .FEAT_BELOW(feature_belows[1629])) ac1629(.scan_win(scan_win1629), .scan_win_std_dev(scan_win_std_dev[1629]), .feature_accum(feature_accums[1629]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1630]), .RECT1_Y(rectangle1_ys[1630]), .RECT1_WIDTH(rectangle1_widths[1630]), .RECT1_HEIGHT(rectangle1_heights[1630]), .RECT1_WEIGHT(rectangle1_weights[1630]), .RECT2_X(rectangle2_xs[1630]), .RECT2_Y(rectangle2_ys[1630]), .RECT2_WIDTH(rectangle2_widths[1630]), .RECT2_HEIGHT(rectangle2_heights[1630]), .RECT2_WEIGHT(rectangle2_weights[1630]), .RECT3_X(rectangle3_xs[1630]), .RECT3_Y(rectangle3_ys[1630]), .RECT3_WIDTH(rectangle3_widths[1630]), .RECT3_HEIGHT(rectangle3_heights[1630]), .RECT3_WEIGHT(rectangle3_weights[1630]), .FEAT_THRES(feature_thresholds[1630]), .FEAT_ABOVE(feature_aboves[1630]), .FEAT_BELOW(feature_belows[1630])) ac1630(.scan_win(scan_win1630), .scan_win_std_dev(scan_win_std_dev[1630]), .feature_accum(feature_accums[1630]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1631]), .RECT1_Y(rectangle1_ys[1631]), .RECT1_WIDTH(rectangle1_widths[1631]), .RECT1_HEIGHT(rectangle1_heights[1631]), .RECT1_WEIGHT(rectangle1_weights[1631]), .RECT2_X(rectangle2_xs[1631]), .RECT2_Y(rectangle2_ys[1631]), .RECT2_WIDTH(rectangle2_widths[1631]), .RECT2_HEIGHT(rectangle2_heights[1631]), .RECT2_WEIGHT(rectangle2_weights[1631]), .RECT3_X(rectangle3_xs[1631]), .RECT3_Y(rectangle3_ys[1631]), .RECT3_WIDTH(rectangle3_widths[1631]), .RECT3_HEIGHT(rectangle3_heights[1631]), .RECT3_WEIGHT(rectangle3_weights[1631]), .FEAT_THRES(feature_thresholds[1631]), .FEAT_ABOVE(feature_aboves[1631]), .FEAT_BELOW(feature_belows[1631])) ac1631(.scan_win(scan_win1631), .scan_win_std_dev(scan_win_std_dev[1631]), .feature_accum(feature_accums[1631]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1632]), .RECT1_Y(rectangle1_ys[1632]), .RECT1_WIDTH(rectangle1_widths[1632]), .RECT1_HEIGHT(rectangle1_heights[1632]), .RECT1_WEIGHT(rectangle1_weights[1632]), .RECT2_X(rectangle2_xs[1632]), .RECT2_Y(rectangle2_ys[1632]), .RECT2_WIDTH(rectangle2_widths[1632]), .RECT2_HEIGHT(rectangle2_heights[1632]), .RECT2_WEIGHT(rectangle2_weights[1632]), .RECT3_X(rectangle3_xs[1632]), .RECT3_Y(rectangle3_ys[1632]), .RECT3_WIDTH(rectangle3_widths[1632]), .RECT3_HEIGHT(rectangle3_heights[1632]), .RECT3_WEIGHT(rectangle3_weights[1632]), .FEAT_THRES(feature_thresholds[1632]), .FEAT_ABOVE(feature_aboves[1632]), .FEAT_BELOW(feature_belows[1632])) ac1632(.scan_win(scan_win1632), .scan_win_std_dev(scan_win_std_dev[1632]), .feature_accum(feature_accums[1632]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1633]), .RECT1_Y(rectangle1_ys[1633]), .RECT1_WIDTH(rectangle1_widths[1633]), .RECT1_HEIGHT(rectangle1_heights[1633]), .RECT1_WEIGHT(rectangle1_weights[1633]), .RECT2_X(rectangle2_xs[1633]), .RECT2_Y(rectangle2_ys[1633]), .RECT2_WIDTH(rectangle2_widths[1633]), .RECT2_HEIGHT(rectangle2_heights[1633]), .RECT2_WEIGHT(rectangle2_weights[1633]), .RECT3_X(rectangle3_xs[1633]), .RECT3_Y(rectangle3_ys[1633]), .RECT3_WIDTH(rectangle3_widths[1633]), .RECT3_HEIGHT(rectangle3_heights[1633]), .RECT3_WEIGHT(rectangle3_weights[1633]), .FEAT_THRES(feature_thresholds[1633]), .FEAT_ABOVE(feature_aboves[1633]), .FEAT_BELOW(feature_belows[1633])) ac1633(.scan_win(scan_win1633), .scan_win_std_dev(scan_win_std_dev[1633]), .feature_accum(feature_accums[1633]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1634]), .RECT1_Y(rectangle1_ys[1634]), .RECT1_WIDTH(rectangle1_widths[1634]), .RECT1_HEIGHT(rectangle1_heights[1634]), .RECT1_WEIGHT(rectangle1_weights[1634]), .RECT2_X(rectangle2_xs[1634]), .RECT2_Y(rectangle2_ys[1634]), .RECT2_WIDTH(rectangle2_widths[1634]), .RECT2_HEIGHT(rectangle2_heights[1634]), .RECT2_WEIGHT(rectangle2_weights[1634]), .RECT3_X(rectangle3_xs[1634]), .RECT3_Y(rectangle3_ys[1634]), .RECT3_WIDTH(rectangle3_widths[1634]), .RECT3_HEIGHT(rectangle3_heights[1634]), .RECT3_WEIGHT(rectangle3_weights[1634]), .FEAT_THRES(feature_thresholds[1634]), .FEAT_ABOVE(feature_aboves[1634]), .FEAT_BELOW(feature_belows[1634])) ac1634(.scan_win(scan_win1634), .scan_win_std_dev(scan_win_std_dev[1634]), .feature_accum(feature_accums[1634]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1635]), .RECT1_Y(rectangle1_ys[1635]), .RECT1_WIDTH(rectangle1_widths[1635]), .RECT1_HEIGHT(rectangle1_heights[1635]), .RECT1_WEIGHT(rectangle1_weights[1635]), .RECT2_X(rectangle2_xs[1635]), .RECT2_Y(rectangle2_ys[1635]), .RECT2_WIDTH(rectangle2_widths[1635]), .RECT2_HEIGHT(rectangle2_heights[1635]), .RECT2_WEIGHT(rectangle2_weights[1635]), .RECT3_X(rectangle3_xs[1635]), .RECT3_Y(rectangle3_ys[1635]), .RECT3_WIDTH(rectangle3_widths[1635]), .RECT3_HEIGHT(rectangle3_heights[1635]), .RECT3_WEIGHT(rectangle3_weights[1635]), .FEAT_THRES(feature_thresholds[1635]), .FEAT_ABOVE(feature_aboves[1635]), .FEAT_BELOW(feature_belows[1635])) ac1635(.scan_win(scan_win1635), .scan_win_std_dev(scan_win_std_dev[1635]), .feature_accum(feature_accums[1635]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1636]), .RECT1_Y(rectangle1_ys[1636]), .RECT1_WIDTH(rectangle1_widths[1636]), .RECT1_HEIGHT(rectangle1_heights[1636]), .RECT1_WEIGHT(rectangle1_weights[1636]), .RECT2_X(rectangle2_xs[1636]), .RECT2_Y(rectangle2_ys[1636]), .RECT2_WIDTH(rectangle2_widths[1636]), .RECT2_HEIGHT(rectangle2_heights[1636]), .RECT2_WEIGHT(rectangle2_weights[1636]), .RECT3_X(rectangle3_xs[1636]), .RECT3_Y(rectangle3_ys[1636]), .RECT3_WIDTH(rectangle3_widths[1636]), .RECT3_HEIGHT(rectangle3_heights[1636]), .RECT3_WEIGHT(rectangle3_weights[1636]), .FEAT_THRES(feature_thresholds[1636]), .FEAT_ABOVE(feature_aboves[1636]), .FEAT_BELOW(feature_belows[1636])) ac1636(.scan_win(scan_win1636), .scan_win_std_dev(scan_win_std_dev[1636]), .feature_accum(feature_accums[1636]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1637]), .RECT1_Y(rectangle1_ys[1637]), .RECT1_WIDTH(rectangle1_widths[1637]), .RECT1_HEIGHT(rectangle1_heights[1637]), .RECT1_WEIGHT(rectangle1_weights[1637]), .RECT2_X(rectangle2_xs[1637]), .RECT2_Y(rectangle2_ys[1637]), .RECT2_WIDTH(rectangle2_widths[1637]), .RECT2_HEIGHT(rectangle2_heights[1637]), .RECT2_WEIGHT(rectangle2_weights[1637]), .RECT3_X(rectangle3_xs[1637]), .RECT3_Y(rectangle3_ys[1637]), .RECT3_WIDTH(rectangle3_widths[1637]), .RECT3_HEIGHT(rectangle3_heights[1637]), .RECT3_WEIGHT(rectangle3_weights[1637]), .FEAT_THRES(feature_thresholds[1637]), .FEAT_ABOVE(feature_aboves[1637]), .FEAT_BELOW(feature_belows[1637])) ac1637(.scan_win(scan_win1637), .scan_win_std_dev(scan_win_std_dev[1637]), .feature_accum(feature_accums[1637]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1638]), .RECT1_Y(rectangle1_ys[1638]), .RECT1_WIDTH(rectangle1_widths[1638]), .RECT1_HEIGHT(rectangle1_heights[1638]), .RECT1_WEIGHT(rectangle1_weights[1638]), .RECT2_X(rectangle2_xs[1638]), .RECT2_Y(rectangle2_ys[1638]), .RECT2_WIDTH(rectangle2_widths[1638]), .RECT2_HEIGHT(rectangle2_heights[1638]), .RECT2_WEIGHT(rectangle2_weights[1638]), .RECT3_X(rectangle3_xs[1638]), .RECT3_Y(rectangle3_ys[1638]), .RECT3_WIDTH(rectangle3_widths[1638]), .RECT3_HEIGHT(rectangle3_heights[1638]), .RECT3_WEIGHT(rectangle3_weights[1638]), .FEAT_THRES(feature_thresholds[1638]), .FEAT_ABOVE(feature_aboves[1638]), .FEAT_BELOW(feature_belows[1638])) ac1638(.scan_win(scan_win1638), .scan_win_std_dev(scan_win_std_dev[1638]), .feature_accum(feature_accums[1638]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1639]), .RECT1_Y(rectangle1_ys[1639]), .RECT1_WIDTH(rectangle1_widths[1639]), .RECT1_HEIGHT(rectangle1_heights[1639]), .RECT1_WEIGHT(rectangle1_weights[1639]), .RECT2_X(rectangle2_xs[1639]), .RECT2_Y(rectangle2_ys[1639]), .RECT2_WIDTH(rectangle2_widths[1639]), .RECT2_HEIGHT(rectangle2_heights[1639]), .RECT2_WEIGHT(rectangle2_weights[1639]), .RECT3_X(rectangle3_xs[1639]), .RECT3_Y(rectangle3_ys[1639]), .RECT3_WIDTH(rectangle3_widths[1639]), .RECT3_HEIGHT(rectangle3_heights[1639]), .RECT3_WEIGHT(rectangle3_weights[1639]), .FEAT_THRES(feature_thresholds[1639]), .FEAT_ABOVE(feature_aboves[1639]), .FEAT_BELOW(feature_belows[1639])) ac1639(.scan_win(scan_win1639), .scan_win_std_dev(scan_win_std_dev[1639]), .feature_accum(feature_accums[1639]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1640]), .RECT1_Y(rectangle1_ys[1640]), .RECT1_WIDTH(rectangle1_widths[1640]), .RECT1_HEIGHT(rectangle1_heights[1640]), .RECT1_WEIGHT(rectangle1_weights[1640]), .RECT2_X(rectangle2_xs[1640]), .RECT2_Y(rectangle2_ys[1640]), .RECT2_WIDTH(rectangle2_widths[1640]), .RECT2_HEIGHT(rectangle2_heights[1640]), .RECT2_WEIGHT(rectangle2_weights[1640]), .RECT3_X(rectangle3_xs[1640]), .RECT3_Y(rectangle3_ys[1640]), .RECT3_WIDTH(rectangle3_widths[1640]), .RECT3_HEIGHT(rectangle3_heights[1640]), .RECT3_WEIGHT(rectangle3_weights[1640]), .FEAT_THRES(feature_thresholds[1640]), .FEAT_ABOVE(feature_aboves[1640]), .FEAT_BELOW(feature_belows[1640])) ac1640(.scan_win(scan_win1640), .scan_win_std_dev(scan_win_std_dev[1640]), .feature_accum(feature_accums[1640]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1641]), .RECT1_Y(rectangle1_ys[1641]), .RECT1_WIDTH(rectangle1_widths[1641]), .RECT1_HEIGHT(rectangle1_heights[1641]), .RECT1_WEIGHT(rectangle1_weights[1641]), .RECT2_X(rectangle2_xs[1641]), .RECT2_Y(rectangle2_ys[1641]), .RECT2_WIDTH(rectangle2_widths[1641]), .RECT2_HEIGHT(rectangle2_heights[1641]), .RECT2_WEIGHT(rectangle2_weights[1641]), .RECT3_X(rectangle3_xs[1641]), .RECT3_Y(rectangle3_ys[1641]), .RECT3_WIDTH(rectangle3_widths[1641]), .RECT3_HEIGHT(rectangle3_heights[1641]), .RECT3_WEIGHT(rectangle3_weights[1641]), .FEAT_THRES(feature_thresholds[1641]), .FEAT_ABOVE(feature_aboves[1641]), .FEAT_BELOW(feature_belows[1641])) ac1641(.scan_win(scan_win1641), .scan_win_std_dev(scan_win_std_dev[1641]), .feature_accum(feature_accums[1641]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1642]), .RECT1_Y(rectangle1_ys[1642]), .RECT1_WIDTH(rectangle1_widths[1642]), .RECT1_HEIGHT(rectangle1_heights[1642]), .RECT1_WEIGHT(rectangle1_weights[1642]), .RECT2_X(rectangle2_xs[1642]), .RECT2_Y(rectangle2_ys[1642]), .RECT2_WIDTH(rectangle2_widths[1642]), .RECT2_HEIGHT(rectangle2_heights[1642]), .RECT2_WEIGHT(rectangle2_weights[1642]), .RECT3_X(rectangle3_xs[1642]), .RECT3_Y(rectangle3_ys[1642]), .RECT3_WIDTH(rectangle3_widths[1642]), .RECT3_HEIGHT(rectangle3_heights[1642]), .RECT3_WEIGHT(rectangle3_weights[1642]), .FEAT_THRES(feature_thresholds[1642]), .FEAT_ABOVE(feature_aboves[1642]), .FEAT_BELOW(feature_belows[1642])) ac1642(.scan_win(scan_win1642), .scan_win_std_dev(scan_win_std_dev[1642]), .feature_accum(feature_accums[1642]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1643]), .RECT1_Y(rectangle1_ys[1643]), .RECT1_WIDTH(rectangle1_widths[1643]), .RECT1_HEIGHT(rectangle1_heights[1643]), .RECT1_WEIGHT(rectangle1_weights[1643]), .RECT2_X(rectangle2_xs[1643]), .RECT2_Y(rectangle2_ys[1643]), .RECT2_WIDTH(rectangle2_widths[1643]), .RECT2_HEIGHT(rectangle2_heights[1643]), .RECT2_WEIGHT(rectangle2_weights[1643]), .RECT3_X(rectangle3_xs[1643]), .RECT3_Y(rectangle3_ys[1643]), .RECT3_WIDTH(rectangle3_widths[1643]), .RECT3_HEIGHT(rectangle3_heights[1643]), .RECT3_WEIGHT(rectangle3_weights[1643]), .FEAT_THRES(feature_thresholds[1643]), .FEAT_ABOVE(feature_aboves[1643]), .FEAT_BELOW(feature_belows[1643])) ac1643(.scan_win(scan_win1643), .scan_win_std_dev(scan_win_std_dev[1643]), .feature_accum(feature_accums[1643]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1644]), .RECT1_Y(rectangle1_ys[1644]), .RECT1_WIDTH(rectangle1_widths[1644]), .RECT1_HEIGHT(rectangle1_heights[1644]), .RECT1_WEIGHT(rectangle1_weights[1644]), .RECT2_X(rectangle2_xs[1644]), .RECT2_Y(rectangle2_ys[1644]), .RECT2_WIDTH(rectangle2_widths[1644]), .RECT2_HEIGHT(rectangle2_heights[1644]), .RECT2_WEIGHT(rectangle2_weights[1644]), .RECT3_X(rectangle3_xs[1644]), .RECT3_Y(rectangle3_ys[1644]), .RECT3_WIDTH(rectangle3_widths[1644]), .RECT3_HEIGHT(rectangle3_heights[1644]), .RECT3_WEIGHT(rectangle3_weights[1644]), .FEAT_THRES(feature_thresholds[1644]), .FEAT_ABOVE(feature_aboves[1644]), .FEAT_BELOW(feature_belows[1644])) ac1644(.scan_win(scan_win1644), .scan_win_std_dev(scan_win_std_dev[1644]), .feature_accum(feature_accums[1644]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1645]), .RECT1_Y(rectangle1_ys[1645]), .RECT1_WIDTH(rectangle1_widths[1645]), .RECT1_HEIGHT(rectangle1_heights[1645]), .RECT1_WEIGHT(rectangle1_weights[1645]), .RECT2_X(rectangle2_xs[1645]), .RECT2_Y(rectangle2_ys[1645]), .RECT2_WIDTH(rectangle2_widths[1645]), .RECT2_HEIGHT(rectangle2_heights[1645]), .RECT2_WEIGHT(rectangle2_weights[1645]), .RECT3_X(rectangle3_xs[1645]), .RECT3_Y(rectangle3_ys[1645]), .RECT3_WIDTH(rectangle3_widths[1645]), .RECT3_HEIGHT(rectangle3_heights[1645]), .RECT3_WEIGHT(rectangle3_weights[1645]), .FEAT_THRES(feature_thresholds[1645]), .FEAT_ABOVE(feature_aboves[1645]), .FEAT_BELOW(feature_belows[1645])) ac1645(.scan_win(scan_win1645), .scan_win_std_dev(scan_win_std_dev[1645]), .feature_accum(feature_accums[1645]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1646]), .RECT1_Y(rectangle1_ys[1646]), .RECT1_WIDTH(rectangle1_widths[1646]), .RECT1_HEIGHT(rectangle1_heights[1646]), .RECT1_WEIGHT(rectangle1_weights[1646]), .RECT2_X(rectangle2_xs[1646]), .RECT2_Y(rectangle2_ys[1646]), .RECT2_WIDTH(rectangle2_widths[1646]), .RECT2_HEIGHT(rectangle2_heights[1646]), .RECT2_WEIGHT(rectangle2_weights[1646]), .RECT3_X(rectangle3_xs[1646]), .RECT3_Y(rectangle3_ys[1646]), .RECT3_WIDTH(rectangle3_widths[1646]), .RECT3_HEIGHT(rectangle3_heights[1646]), .RECT3_WEIGHT(rectangle3_weights[1646]), .FEAT_THRES(feature_thresholds[1646]), .FEAT_ABOVE(feature_aboves[1646]), .FEAT_BELOW(feature_belows[1646])) ac1646(.scan_win(scan_win1646), .scan_win_std_dev(scan_win_std_dev[1646]), .feature_accum(feature_accums[1646]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1647]), .RECT1_Y(rectangle1_ys[1647]), .RECT1_WIDTH(rectangle1_widths[1647]), .RECT1_HEIGHT(rectangle1_heights[1647]), .RECT1_WEIGHT(rectangle1_weights[1647]), .RECT2_X(rectangle2_xs[1647]), .RECT2_Y(rectangle2_ys[1647]), .RECT2_WIDTH(rectangle2_widths[1647]), .RECT2_HEIGHT(rectangle2_heights[1647]), .RECT2_WEIGHT(rectangle2_weights[1647]), .RECT3_X(rectangle3_xs[1647]), .RECT3_Y(rectangle3_ys[1647]), .RECT3_WIDTH(rectangle3_widths[1647]), .RECT3_HEIGHT(rectangle3_heights[1647]), .RECT3_WEIGHT(rectangle3_weights[1647]), .FEAT_THRES(feature_thresholds[1647]), .FEAT_ABOVE(feature_aboves[1647]), .FEAT_BELOW(feature_belows[1647])) ac1647(.scan_win(scan_win1647), .scan_win_std_dev(scan_win_std_dev[1647]), .feature_accum(feature_accums[1647]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1648]), .RECT1_Y(rectangle1_ys[1648]), .RECT1_WIDTH(rectangle1_widths[1648]), .RECT1_HEIGHT(rectangle1_heights[1648]), .RECT1_WEIGHT(rectangle1_weights[1648]), .RECT2_X(rectangle2_xs[1648]), .RECT2_Y(rectangle2_ys[1648]), .RECT2_WIDTH(rectangle2_widths[1648]), .RECT2_HEIGHT(rectangle2_heights[1648]), .RECT2_WEIGHT(rectangle2_weights[1648]), .RECT3_X(rectangle3_xs[1648]), .RECT3_Y(rectangle3_ys[1648]), .RECT3_WIDTH(rectangle3_widths[1648]), .RECT3_HEIGHT(rectangle3_heights[1648]), .RECT3_WEIGHT(rectangle3_weights[1648]), .FEAT_THRES(feature_thresholds[1648]), .FEAT_ABOVE(feature_aboves[1648]), .FEAT_BELOW(feature_belows[1648])) ac1648(.scan_win(scan_win1648), .scan_win_std_dev(scan_win_std_dev[1648]), .feature_accum(feature_accums[1648]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1649]), .RECT1_Y(rectangle1_ys[1649]), .RECT1_WIDTH(rectangle1_widths[1649]), .RECT1_HEIGHT(rectangle1_heights[1649]), .RECT1_WEIGHT(rectangle1_weights[1649]), .RECT2_X(rectangle2_xs[1649]), .RECT2_Y(rectangle2_ys[1649]), .RECT2_WIDTH(rectangle2_widths[1649]), .RECT2_HEIGHT(rectangle2_heights[1649]), .RECT2_WEIGHT(rectangle2_weights[1649]), .RECT3_X(rectangle3_xs[1649]), .RECT3_Y(rectangle3_ys[1649]), .RECT3_WIDTH(rectangle3_widths[1649]), .RECT3_HEIGHT(rectangle3_heights[1649]), .RECT3_WEIGHT(rectangle3_weights[1649]), .FEAT_THRES(feature_thresholds[1649]), .FEAT_ABOVE(feature_aboves[1649]), .FEAT_BELOW(feature_belows[1649])) ac1649(.scan_win(scan_win1649), .scan_win_std_dev(scan_win_std_dev[1649]), .feature_accum(feature_accums[1649]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1650]), .RECT1_Y(rectangle1_ys[1650]), .RECT1_WIDTH(rectangle1_widths[1650]), .RECT1_HEIGHT(rectangle1_heights[1650]), .RECT1_WEIGHT(rectangle1_weights[1650]), .RECT2_X(rectangle2_xs[1650]), .RECT2_Y(rectangle2_ys[1650]), .RECT2_WIDTH(rectangle2_widths[1650]), .RECT2_HEIGHT(rectangle2_heights[1650]), .RECT2_WEIGHT(rectangle2_weights[1650]), .RECT3_X(rectangle3_xs[1650]), .RECT3_Y(rectangle3_ys[1650]), .RECT3_WIDTH(rectangle3_widths[1650]), .RECT3_HEIGHT(rectangle3_heights[1650]), .RECT3_WEIGHT(rectangle3_weights[1650]), .FEAT_THRES(feature_thresholds[1650]), .FEAT_ABOVE(feature_aboves[1650]), .FEAT_BELOW(feature_belows[1650])) ac1650(.scan_win(scan_win1650), .scan_win_std_dev(scan_win_std_dev[1650]), .feature_accum(feature_accums[1650]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1651]), .RECT1_Y(rectangle1_ys[1651]), .RECT1_WIDTH(rectangle1_widths[1651]), .RECT1_HEIGHT(rectangle1_heights[1651]), .RECT1_WEIGHT(rectangle1_weights[1651]), .RECT2_X(rectangle2_xs[1651]), .RECT2_Y(rectangle2_ys[1651]), .RECT2_WIDTH(rectangle2_widths[1651]), .RECT2_HEIGHT(rectangle2_heights[1651]), .RECT2_WEIGHT(rectangle2_weights[1651]), .RECT3_X(rectangle3_xs[1651]), .RECT3_Y(rectangle3_ys[1651]), .RECT3_WIDTH(rectangle3_widths[1651]), .RECT3_HEIGHT(rectangle3_heights[1651]), .RECT3_WEIGHT(rectangle3_weights[1651]), .FEAT_THRES(feature_thresholds[1651]), .FEAT_ABOVE(feature_aboves[1651]), .FEAT_BELOW(feature_belows[1651])) ac1651(.scan_win(scan_win1651), .scan_win_std_dev(scan_win_std_dev[1651]), .feature_accum(feature_accums[1651]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1652]), .RECT1_Y(rectangle1_ys[1652]), .RECT1_WIDTH(rectangle1_widths[1652]), .RECT1_HEIGHT(rectangle1_heights[1652]), .RECT1_WEIGHT(rectangle1_weights[1652]), .RECT2_X(rectangle2_xs[1652]), .RECT2_Y(rectangle2_ys[1652]), .RECT2_WIDTH(rectangle2_widths[1652]), .RECT2_HEIGHT(rectangle2_heights[1652]), .RECT2_WEIGHT(rectangle2_weights[1652]), .RECT3_X(rectangle3_xs[1652]), .RECT3_Y(rectangle3_ys[1652]), .RECT3_WIDTH(rectangle3_widths[1652]), .RECT3_HEIGHT(rectangle3_heights[1652]), .RECT3_WEIGHT(rectangle3_weights[1652]), .FEAT_THRES(feature_thresholds[1652]), .FEAT_ABOVE(feature_aboves[1652]), .FEAT_BELOW(feature_belows[1652])) ac1652(.scan_win(scan_win1652), .scan_win_std_dev(scan_win_std_dev[1652]), .feature_accum(feature_accums[1652]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1653]), .RECT1_Y(rectangle1_ys[1653]), .RECT1_WIDTH(rectangle1_widths[1653]), .RECT1_HEIGHT(rectangle1_heights[1653]), .RECT1_WEIGHT(rectangle1_weights[1653]), .RECT2_X(rectangle2_xs[1653]), .RECT2_Y(rectangle2_ys[1653]), .RECT2_WIDTH(rectangle2_widths[1653]), .RECT2_HEIGHT(rectangle2_heights[1653]), .RECT2_WEIGHT(rectangle2_weights[1653]), .RECT3_X(rectangle3_xs[1653]), .RECT3_Y(rectangle3_ys[1653]), .RECT3_WIDTH(rectangle3_widths[1653]), .RECT3_HEIGHT(rectangle3_heights[1653]), .RECT3_WEIGHT(rectangle3_weights[1653]), .FEAT_THRES(feature_thresholds[1653]), .FEAT_ABOVE(feature_aboves[1653]), .FEAT_BELOW(feature_belows[1653])) ac1653(.scan_win(scan_win1653), .scan_win_std_dev(scan_win_std_dev[1653]), .feature_accum(feature_accums[1653]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1654]), .RECT1_Y(rectangle1_ys[1654]), .RECT1_WIDTH(rectangle1_widths[1654]), .RECT1_HEIGHT(rectangle1_heights[1654]), .RECT1_WEIGHT(rectangle1_weights[1654]), .RECT2_X(rectangle2_xs[1654]), .RECT2_Y(rectangle2_ys[1654]), .RECT2_WIDTH(rectangle2_widths[1654]), .RECT2_HEIGHT(rectangle2_heights[1654]), .RECT2_WEIGHT(rectangle2_weights[1654]), .RECT3_X(rectangle3_xs[1654]), .RECT3_Y(rectangle3_ys[1654]), .RECT3_WIDTH(rectangle3_widths[1654]), .RECT3_HEIGHT(rectangle3_heights[1654]), .RECT3_WEIGHT(rectangle3_weights[1654]), .FEAT_THRES(feature_thresholds[1654]), .FEAT_ABOVE(feature_aboves[1654]), .FEAT_BELOW(feature_belows[1654])) ac1654(.scan_win(scan_win1654), .scan_win_std_dev(scan_win_std_dev[1654]), .feature_accum(feature_accums[1654]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1655]), .RECT1_Y(rectangle1_ys[1655]), .RECT1_WIDTH(rectangle1_widths[1655]), .RECT1_HEIGHT(rectangle1_heights[1655]), .RECT1_WEIGHT(rectangle1_weights[1655]), .RECT2_X(rectangle2_xs[1655]), .RECT2_Y(rectangle2_ys[1655]), .RECT2_WIDTH(rectangle2_widths[1655]), .RECT2_HEIGHT(rectangle2_heights[1655]), .RECT2_WEIGHT(rectangle2_weights[1655]), .RECT3_X(rectangle3_xs[1655]), .RECT3_Y(rectangle3_ys[1655]), .RECT3_WIDTH(rectangle3_widths[1655]), .RECT3_HEIGHT(rectangle3_heights[1655]), .RECT3_WEIGHT(rectangle3_weights[1655]), .FEAT_THRES(feature_thresholds[1655]), .FEAT_ABOVE(feature_aboves[1655]), .FEAT_BELOW(feature_belows[1655])) ac1655(.scan_win(scan_win1655), .scan_win_std_dev(scan_win_std_dev[1655]), .feature_accum(feature_accums[1655]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1656]), .RECT1_Y(rectangle1_ys[1656]), .RECT1_WIDTH(rectangle1_widths[1656]), .RECT1_HEIGHT(rectangle1_heights[1656]), .RECT1_WEIGHT(rectangle1_weights[1656]), .RECT2_X(rectangle2_xs[1656]), .RECT2_Y(rectangle2_ys[1656]), .RECT2_WIDTH(rectangle2_widths[1656]), .RECT2_HEIGHT(rectangle2_heights[1656]), .RECT2_WEIGHT(rectangle2_weights[1656]), .RECT3_X(rectangle3_xs[1656]), .RECT3_Y(rectangle3_ys[1656]), .RECT3_WIDTH(rectangle3_widths[1656]), .RECT3_HEIGHT(rectangle3_heights[1656]), .RECT3_WEIGHT(rectangle3_weights[1656]), .FEAT_THRES(feature_thresholds[1656]), .FEAT_ABOVE(feature_aboves[1656]), .FEAT_BELOW(feature_belows[1656])) ac1656(.scan_win(scan_win1656), .scan_win_std_dev(scan_win_std_dev[1656]), .feature_accum(feature_accums[1656]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1657]), .RECT1_Y(rectangle1_ys[1657]), .RECT1_WIDTH(rectangle1_widths[1657]), .RECT1_HEIGHT(rectangle1_heights[1657]), .RECT1_WEIGHT(rectangle1_weights[1657]), .RECT2_X(rectangle2_xs[1657]), .RECT2_Y(rectangle2_ys[1657]), .RECT2_WIDTH(rectangle2_widths[1657]), .RECT2_HEIGHT(rectangle2_heights[1657]), .RECT2_WEIGHT(rectangle2_weights[1657]), .RECT3_X(rectangle3_xs[1657]), .RECT3_Y(rectangle3_ys[1657]), .RECT3_WIDTH(rectangle3_widths[1657]), .RECT3_HEIGHT(rectangle3_heights[1657]), .RECT3_WEIGHT(rectangle3_weights[1657]), .FEAT_THRES(feature_thresholds[1657]), .FEAT_ABOVE(feature_aboves[1657]), .FEAT_BELOW(feature_belows[1657])) ac1657(.scan_win(scan_win1657), .scan_win_std_dev(scan_win_std_dev[1657]), .feature_accum(feature_accums[1657]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1658]), .RECT1_Y(rectangle1_ys[1658]), .RECT1_WIDTH(rectangle1_widths[1658]), .RECT1_HEIGHT(rectangle1_heights[1658]), .RECT1_WEIGHT(rectangle1_weights[1658]), .RECT2_X(rectangle2_xs[1658]), .RECT2_Y(rectangle2_ys[1658]), .RECT2_WIDTH(rectangle2_widths[1658]), .RECT2_HEIGHT(rectangle2_heights[1658]), .RECT2_WEIGHT(rectangle2_weights[1658]), .RECT3_X(rectangle3_xs[1658]), .RECT3_Y(rectangle3_ys[1658]), .RECT3_WIDTH(rectangle3_widths[1658]), .RECT3_HEIGHT(rectangle3_heights[1658]), .RECT3_WEIGHT(rectangle3_weights[1658]), .FEAT_THRES(feature_thresholds[1658]), .FEAT_ABOVE(feature_aboves[1658]), .FEAT_BELOW(feature_belows[1658])) ac1658(.scan_win(scan_win1658), .scan_win_std_dev(scan_win_std_dev[1658]), .feature_accum(feature_accums[1658]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1659]), .RECT1_Y(rectangle1_ys[1659]), .RECT1_WIDTH(rectangle1_widths[1659]), .RECT1_HEIGHT(rectangle1_heights[1659]), .RECT1_WEIGHT(rectangle1_weights[1659]), .RECT2_X(rectangle2_xs[1659]), .RECT2_Y(rectangle2_ys[1659]), .RECT2_WIDTH(rectangle2_widths[1659]), .RECT2_HEIGHT(rectangle2_heights[1659]), .RECT2_WEIGHT(rectangle2_weights[1659]), .RECT3_X(rectangle3_xs[1659]), .RECT3_Y(rectangle3_ys[1659]), .RECT3_WIDTH(rectangle3_widths[1659]), .RECT3_HEIGHT(rectangle3_heights[1659]), .RECT3_WEIGHT(rectangle3_weights[1659]), .FEAT_THRES(feature_thresholds[1659]), .FEAT_ABOVE(feature_aboves[1659]), .FEAT_BELOW(feature_belows[1659])) ac1659(.scan_win(scan_win1659), .scan_win_std_dev(scan_win_std_dev[1659]), .feature_accum(feature_accums[1659]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1660]), .RECT1_Y(rectangle1_ys[1660]), .RECT1_WIDTH(rectangle1_widths[1660]), .RECT1_HEIGHT(rectangle1_heights[1660]), .RECT1_WEIGHT(rectangle1_weights[1660]), .RECT2_X(rectangle2_xs[1660]), .RECT2_Y(rectangle2_ys[1660]), .RECT2_WIDTH(rectangle2_widths[1660]), .RECT2_HEIGHT(rectangle2_heights[1660]), .RECT2_WEIGHT(rectangle2_weights[1660]), .RECT3_X(rectangle3_xs[1660]), .RECT3_Y(rectangle3_ys[1660]), .RECT3_WIDTH(rectangle3_widths[1660]), .RECT3_HEIGHT(rectangle3_heights[1660]), .RECT3_WEIGHT(rectangle3_weights[1660]), .FEAT_THRES(feature_thresholds[1660]), .FEAT_ABOVE(feature_aboves[1660]), .FEAT_BELOW(feature_belows[1660])) ac1660(.scan_win(scan_win1660), .scan_win_std_dev(scan_win_std_dev[1660]), .feature_accum(feature_accums[1660]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1661]), .RECT1_Y(rectangle1_ys[1661]), .RECT1_WIDTH(rectangle1_widths[1661]), .RECT1_HEIGHT(rectangle1_heights[1661]), .RECT1_WEIGHT(rectangle1_weights[1661]), .RECT2_X(rectangle2_xs[1661]), .RECT2_Y(rectangle2_ys[1661]), .RECT2_WIDTH(rectangle2_widths[1661]), .RECT2_HEIGHT(rectangle2_heights[1661]), .RECT2_WEIGHT(rectangle2_weights[1661]), .RECT3_X(rectangle3_xs[1661]), .RECT3_Y(rectangle3_ys[1661]), .RECT3_WIDTH(rectangle3_widths[1661]), .RECT3_HEIGHT(rectangle3_heights[1661]), .RECT3_WEIGHT(rectangle3_weights[1661]), .FEAT_THRES(feature_thresholds[1661]), .FEAT_ABOVE(feature_aboves[1661]), .FEAT_BELOW(feature_belows[1661])) ac1661(.scan_win(scan_win1661), .scan_win_std_dev(scan_win_std_dev[1661]), .feature_accum(feature_accums[1661]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1662]), .RECT1_Y(rectangle1_ys[1662]), .RECT1_WIDTH(rectangle1_widths[1662]), .RECT1_HEIGHT(rectangle1_heights[1662]), .RECT1_WEIGHT(rectangle1_weights[1662]), .RECT2_X(rectangle2_xs[1662]), .RECT2_Y(rectangle2_ys[1662]), .RECT2_WIDTH(rectangle2_widths[1662]), .RECT2_HEIGHT(rectangle2_heights[1662]), .RECT2_WEIGHT(rectangle2_weights[1662]), .RECT3_X(rectangle3_xs[1662]), .RECT3_Y(rectangle3_ys[1662]), .RECT3_WIDTH(rectangle3_widths[1662]), .RECT3_HEIGHT(rectangle3_heights[1662]), .RECT3_WEIGHT(rectangle3_weights[1662]), .FEAT_THRES(feature_thresholds[1662]), .FEAT_ABOVE(feature_aboves[1662]), .FEAT_BELOW(feature_belows[1662])) ac1662(.scan_win(scan_win1662), .scan_win_std_dev(scan_win_std_dev[1662]), .feature_accum(feature_accums[1662]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1663]), .RECT1_Y(rectangle1_ys[1663]), .RECT1_WIDTH(rectangle1_widths[1663]), .RECT1_HEIGHT(rectangle1_heights[1663]), .RECT1_WEIGHT(rectangle1_weights[1663]), .RECT2_X(rectangle2_xs[1663]), .RECT2_Y(rectangle2_ys[1663]), .RECT2_WIDTH(rectangle2_widths[1663]), .RECT2_HEIGHT(rectangle2_heights[1663]), .RECT2_WEIGHT(rectangle2_weights[1663]), .RECT3_X(rectangle3_xs[1663]), .RECT3_Y(rectangle3_ys[1663]), .RECT3_WIDTH(rectangle3_widths[1663]), .RECT3_HEIGHT(rectangle3_heights[1663]), .RECT3_WEIGHT(rectangle3_weights[1663]), .FEAT_THRES(feature_thresholds[1663]), .FEAT_ABOVE(feature_aboves[1663]), .FEAT_BELOW(feature_belows[1663])) ac1663(.scan_win(scan_win1663), .scan_win_std_dev(scan_win_std_dev[1663]), .feature_accum(feature_accums[1663]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1664]), .RECT1_Y(rectangle1_ys[1664]), .RECT1_WIDTH(rectangle1_widths[1664]), .RECT1_HEIGHT(rectangle1_heights[1664]), .RECT1_WEIGHT(rectangle1_weights[1664]), .RECT2_X(rectangle2_xs[1664]), .RECT2_Y(rectangle2_ys[1664]), .RECT2_WIDTH(rectangle2_widths[1664]), .RECT2_HEIGHT(rectangle2_heights[1664]), .RECT2_WEIGHT(rectangle2_weights[1664]), .RECT3_X(rectangle3_xs[1664]), .RECT3_Y(rectangle3_ys[1664]), .RECT3_WIDTH(rectangle3_widths[1664]), .RECT3_HEIGHT(rectangle3_heights[1664]), .RECT3_WEIGHT(rectangle3_weights[1664]), .FEAT_THRES(feature_thresholds[1664]), .FEAT_ABOVE(feature_aboves[1664]), .FEAT_BELOW(feature_belows[1664])) ac1664(.scan_win(scan_win1664), .scan_win_std_dev(scan_win_std_dev[1664]), .feature_accum(feature_accums[1664]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1665]), .RECT1_Y(rectangle1_ys[1665]), .RECT1_WIDTH(rectangle1_widths[1665]), .RECT1_HEIGHT(rectangle1_heights[1665]), .RECT1_WEIGHT(rectangle1_weights[1665]), .RECT2_X(rectangle2_xs[1665]), .RECT2_Y(rectangle2_ys[1665]), .RECT2_WIDTH(rectangle2_widths[1665]), .RECT2_HEIGHT(rectangle2_heights[1665]), .RECT2_WEIGHT(rectangle2_weights[1665]), .RECT3_X(rectangle3_xs[1665]), .RECT3_Y(rectangle3_ys[1665]), .RECT3_WIDTH(rectangle3_widths[1665]), .RECT3_HEIGHT(rectangle3_heights[1665]), .RECT3_WEIGHT(rectangle3_weights[1665]), .FEAT_THRES(feature_thresholds[1665]), .FEAT_ABOVE(feature_aboves[1665]), .FEAT_BELOW(feature_belows[1665])) ac1665(.scan_win(scan_win1665), .scan_win_std_dev(scan_win_std_dev[1665]), .feature_accum(feature_accums[1665]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1666]), .RECT1_Y(rectangle1_ys[1666]), .RECT1_WIDTH(rectangle1_widths[1666]), .RECT1_HEIGHT(rectangle1_heights[1666]), .RECT1_WEIGHT(rectangle1_weights[1666]), .RECT2_X(rectangle2_xs[1666]), .RECT2_Y(rectangle2_ys[1666]), .RECT2_WIDTH(rectangle2_widths[1666]), .RECT2_HEIGHT(rectangle2_heights[1666]), .RECT2_WEIGHT(rectangle2_weights[1666]), .RECT3_X(rectangle3_xs[1666]), .RECT3_Y(rectangle3_ys[1666]), .RECT3_WIDTH(rectangle3_widths[1666]), .RECT3_HEIGHT(rectangle3_heights[1666]), .RECT3_WEIGHT(rectangle3_weights[1666]), .FEAT_THRES(feature_thresholds[1666]), .FEAT_ABOVE(feature_aboves[1666]), .FEAT_BELOW(feature_belows[1666])) ac1666(.scan_win(scan_win1666), .scan_win_std_dev(scan_win_std_dev[1666]), .feature_accum(feature_accums[1666]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1667]), .RECT1_Y(rectangle1_ys[1667]), .RECT1_WIDTH(rectangle1_widths[1667]), .RECT1_HEIGHT(rectangle1_heights[1667]), .RECT1_WEIGHT(rectangle1_weights[1667]), .RECT2_X(rectangle2_xs[1667]), .RECT2_Y(rectangle2_ys[1667]), .RECT2_WIDTH(rectangle2_widths[1667]), .RECT2_HEIGHT(rectangle2_heights[1667]), .RECT2_WEIGHT(rectangle2_weights[1667]), .RECT3_X(rectangle3_xs[1667]), .RECT3_Y(rectangle3_ys[1667]), .RECT3_WIDTH(rectangle3_widths[1667]), .RECT3_HEIGHT(rectangle3_heights[1667]), .RECT3_WEIGHT(rectangle3_weights[1667]), .FEAT_THRES(feature_thresholds[1667]), .FEAT_ABOVE(feature_aboves[1667]), .FEAT_BELOW(feature_belows[1667])) ac1667(.scan_win(scan_win1667), .scan_win_std_dev(scan_win_std_dev[1667]), .feature_accum(feature_accums[1667]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1668]), .RECT1_Y(rectangle1_ys[1668]), .RECT1_WIDTH(rectangle1_widths[1668]), .RECT1_HEIGHT(rectangle1_heights[1668]), .RECT1_WEIGHT(rectangle1_weights[1668]), .RECT2_X(rectangle2_xs[1668]), .RECT2_Y(rectangle2_ys[1668]), .RECT2_WIDTH(rectangle2_widths[1668]), .RECT2_HEIGHT(rectangle2_heights[1668]), .RECT2_WEIGHT(rectangle2_weights[1668]), .RECT3_X(rectangle3_xs[1668]), .RECT3_Y(rectangle3_ys[1668]), .RECT3_WIDTH(rectangle3_widths[1668]), .RECT3_HEIGHT(rectangle3_heights[1668]), .RECT3_WEIGHT(rectangle3_weights[1668]), .FEAT_THRES(feature_thresholds[1668]), .FEAT_ABOVE(feature_aboves[1668]), .FEAT_BELOW(feature_belows[1668])) ac1668(.scan_win(scan_win1668), .scan_win_std_dev(scan_win_std_dev[1668]), .feature_accum(feature_accums[1668]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1669]), .RECT1_Y(rectangle1_ys[1669]), .RECT1_WIDTH(rectangle1_widths[1669]), .RECT1_HEIGHT(rectangle1_heights[1669]), .RECT1_WEIGHT(rectangle1_weights[1669]), .RECT2_X(rectangle2_xs[1669]), .RECT2_Y(rectangle2_ys[1669]), .RECT2_WIDTH(rectangle2_widths[1669]), .RECT2_HEIGHT(rectangle2_heights[1669]), .RECT2_WEIGHT(rectangle2_weights[1669]), .RECT3_X(rectangle3_xs[1669]), .RECT3_Y(rectangle3_ys[1669]), .RECT3_WIDTH(rectangle3_widths[1669]), .RECT3_HEIGHT(rectangle3_heights[1669]), .RECT3_WEIGHT(rectangle3_weights[1669]), .FEAT_THRES(feature_thresholds[1669]), .FEAT_ABOVE(feature_aboves[1669]), .FEAT_BELOW(feature_belows[1669])) ac1669(.scan_win(scan_win1669), .scan_win_std_dev(scan_win_std_dev[1669]), .feature_accum(feature_accums[1669]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1670]), .RECT1_Y(rectangle1_ys[1670]), .RECT1_WIDTH(rectangle1_widths[1670]), .RECT1_HEIGHT(rectangle1_heights[1670]), .RECT1_WEIGHT(rectangle1_weights[1670]), .RECT2_X(rectangle2_xs[1670]), .RECT2_Y(rectangle2_ys[1670]), .RECT2_WIDTH(rectangle2_widths[1670]), .RECT2_HEIGHT(rectangle2_heights[1670]), .RECT2_WEIGHT(rectangle2_weights[1670]), .RECT3_X(rectangle3_xs[1670]), .RECT3_Y(rectangle3_ys[1670]), .RECT3_WIDTH(rectangle3_widths[1670]), .RECT3_HEIGHT(rectangle3_heights[1670]), .RECT3_WEIGHT(rectangle3_weights[1670]), .FEAT_THRES(feature_thresholds[1670]), .FEAT_ABOVE(feature_aboves[1670]), .FEAT_BELOW(feature_belows[1670])) ac1670(.scan_win(scan_win1670), .scan_win_std_dev(scan_win_std_dev[1670]), .feature_accum(feature_accums[1670]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1671]), .RECT1_Y(rectangle1_ys[1671]), .RECT1_WIDTH(rectangle1_widths[1671]), .RECT1_HEIGHT(rectangle1_heights[1671]), .RECT1_WEIGHT(rectangle1_weights[1671]), .RECT2_X(rectangle2_xs[1671]), .RECT2_Y(rectangle2_ys[1671]), .RECT2_WIDTH(rectangle2_widths[1671]), .RECT2_HEIGHT(rectangle2_heights[1671]), .RECT2_WEIGHT(rectangle2_weights[1671]), .RECT3_X(rectangle3_xs[1671]), .RECT3_Y(rectangle3_ys[1671]), .RECT3_WIDTH(rectangle3_widths[1671]), .RECT3_HEIGHT(rectangle3_heights[1671]), .RECT3_WEIGHT(rectangle3_weights[1671]), .FEAT_THRES(feature_thresholds[1671]), .FEAT_ABOVE(feature_aboves[1671]), .FEAT_BELOW(feature_belows[1671])) ac1671(.scan_win(scan_win1671), .scan_win_std_dev(scan_win_std_dev[1671]), .feature_accum(feature_accums[1671]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1672]), .RECT1_Y(rectangle1_ys[1672]), .RECT1_WIDTH(rectangle1_widths[1672]), .RECT1_HEIGHT(rectangle1_heights[1672]), .RECT1_WEIGHT(rectangle1_weights[1672]), .RECT2_X(rectangle2_xs[1672]), .RECT2_Y(rectangle2_ys[1672]), .RECT2_WIDTH(rectangle2_widths[1672]), .RECT2_HEIGHT(rectangle2_heights[1672]), .RECT2_WEIGHT(rectangle2_weights[1672]), .RECT3_X(rectangle3_xs[1672]), .RECT3_Y(rectangle3_ys[1672]), .RECT3_WIDTH(rectangle3_widths[1672]), .RECT3_HEIGHT(rectangle3_heights[1672]), .RECT3_WEIGHT(rectangle3_weights[1672]), .FEAT_THRES(feature_thresholds[1672]), .FEAT_ABOVE(feature_aboves[1672]), .FEAT_BELOW(feature_belows[1672])) ac1672(.scan_win(scan_win1672), .scan_win_std_dev(scan_win_std_dev[1672]), .feature_accum(feature_accums[1672]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1673]), .RECT1_Y(rectangle1_ys[1673]), .RECT1_WIDTH(rectangle1_widths[1673]), .RECT1_HEIGHT(rectangle1_heights[1673]), .RECT1_WEIGHT(rectangle1_weights[1673]), .RECT2_X(rectangle2_xs[1673]), .RECT2_Y(rectangle2_ys[1673]), .RECT2_WIDTH(rectangle2_widths[1673]), .RECT2_HEIGHT(rectangle2_heights[1673]), .RECT2_WEIGHT(rectangle2_weights[1673]), .RECT3_X(rectangle3_xs[1673]), .RECT3_Y(rectangle3_ys[1673]), .RECT3_WIDTH(rectangle3_widths[1673]), .RECT3_HEIGHT(rectangle3_heights[1673]), .RECT3_WEIGHT(rectangle3_weights[1673]), .FEAT_THRES(feature_thresholds[1673]), .FEAT_ABOVE(feature_aboves[1673]), .FEAT_BELOW(feature_belows[1673])) ac1673(.scan_win(scan_win1673), .scan_win_std_dev(scan_win_std_dev[1673]), .feature_accum(feature_accums[1673]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1674]), .RECT1_Y(rectangle1_ys[1674]), .RECT1_WIDTH(rectangle1_widths[1674]), .RECT1_HEIGHT(rectangle1_heights[1674]), .RECT1_WEIGHT(rectangle1_weights[1674]), .RECT2_X(rectangle2_xs[1674]), .RECT2_Y(rectangle2_ys[1674]), .RECT2_WIDTH(rectangle2_widths[1674]), .RECT2_HEIGHT(rectangle2_heights[1674]), .RECT2_WEIGHT(rectangle2_weights[1674]), .RECT3_X(rectangle3_xs[1674]), .RECT3_Y(rectangle3_ys[1674]), .RECT3_WIDTH(rectangle3_widths[1674]), .RECT3_HEIGHT(rectangle3_heights[1674]), .RECT3_WEIGHT(rectangle3_weights[1674]), .FEAT_THRES(feature_thresholds[1674]), .FEAT_ABOVE(feature_aboves[1674]), .FEAT_BELOW(feature_belows[1674])) ac1674(.scan_win(scan_win1674), .scan_win_std_dev(scan_win_std_dev[1674]), .feature_accum(feature_accums[1674]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1675]), .RECT1_Y(rectangle1_ys[1675]), .RECT1_WIDTH(rectangle1_widths[1675]), .RECT1_HEIGHT(rectangle1_heights[1675]), .RECT1_WEIGHT(rectangle1_weights[1675]), .RECT2_X(rectangle2_xs[1675]), .RECT2_Y(rectangle2_ys[1675]), .RECT2_WIDTH(rectangle2_widths[1675]), .RECT2_HEIGHT(rectangle2_heights[1675]), .RECT2_WEIGHT(rectangle2_weights[1675]), .RECT3_X(rectangle3_xs[1675]), .RECT3_Y(rectangle3_ys[1675]), .RECT3_WIDTH(rectangle3_widths[1675]), .RECT3_HEIGHT(rectangle3_heights[1675]), .RECT3_WEIGHT(rectangle3_weights[1675]), .FEAT_THRES(feature_thresholds[1675]), .FEAT_ABOVE(feature_aboves[1675]), .FEAT_BELOW(feature_belows[1675])) ac1675(.scan_win(scan_win1675), .scan_win_std_dev(scan_win_std_dev[1675]), .feature_accum(feature_accums[1675]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1676]), .RECT1_Y(rectangle1_ys[1676]), .RECT1_WIDTH(rectangle1_widths[1676]), .RECT1_HEIGHT(rectangle1_heights[1676]), .RECT1_WEIGHT(rectangle1_weights[1676]), .RECT2_X(rectangle2_xs[1676]), .RECT2_Y(rectangle2_ys[1676]), .RECT2_WIDTH(rectangle2_widths[1676]), .RECT2_HEIGHT(rectangle2_heights[1676]), .RECT2_WEIGHT(rectangle2_weights[1676]), .RECT3_X(rectangle3_xs[1676]), .RECT3_Y(rectangle3_ys[1676]), .RECT3_WIDTH(rectangle3_widths[1676]), .RECT3_HEIGHT(rectangle3_heights[1676]), .RECT3_WEIGHT(rectangle3_weights[1676]), .FEAT_THRES(feature_thresholds[1676]), .FEAT_ABOVE(feature_aboves[1676]), .FEAT_BELOW(feature_belows[1676])) ac1676(.scan_win(scan_win1676), .scan_win_std_dev(scan_win_std_dev[1676]), .feature_accum(feature_accums[1676]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1677]), .RECT1_Y(rectangle1_ys[1677]), .RECT1_WIDTH(rectangle1_widths[1677]), .RECT1_HEIGHT(rectangle1_heights[1677]), .RECT1_WEIGHT(rectangle1_weights[1677]), .RECT2_X(rectangle2_xs[1677]), .RECT2_Y(rectangle2_ys[1677]), .RECT2_WIDTH(rectangle2_widths[1677]), .RECT2_HEIGHT(rectangle2_heights[1677]), .RECT2_WEIGHT(rectangle2_weights[1677]), .RECT3_X(rectangle3_xs[1677]), .RECT3_Y(rectangle3_ys[1677]), .RECT3_WIDTH(rectangle3_widths[1677]), .RECT3_HEIGHT(rectangle3_heights[1677]), .RECT3_WEIGHT(rectangle3_weights[1677]), .FEAT_THRES(feature_thresholds[1677]), .FEAT_ABOVE(feature_aboves[1677]), .FEAT_BELOW(feature_belows[1677])) ac1677(.scan_win(scan_win1677), .scan_win_std_dev(scan_win_std_dev[1677]), .feature_accum(feature_accums[1677]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1678]), .RECT1_Y(rectangle1_ys[1678]), .RECT1_WIDTH(rectangle1_widths[1678]), .RECT1_HEIGHT(rectangle1_heights[1678]), .RECT1_WEIGHT(rectangle1_weights[1678]), .RECT2_X(rectangle2_xs[1678]), .RECT2_Y(rectangle2_ys[1678]), .RECT2_WIDTH(rectangle2_widths[1678]), .RECT2_HEIGHT(rectangle2_heights[1678]), .RECT2_WEIGHT(rectangle2_weights[1678]), .RECT3_X(rectangle3_xs[1678]), .RECT3_Y(rectangle3_ys[1678]), .RECT3_WIDTH(rectangle3_widths[1678]), .RECT3_HEIGHT(rectangle3_heights[1678]), .RECT3_WEIGHT(rectangle3_weights[1678]), .FEAT_THRES(feature_thresholds[1678]), .FEAT_ABOVE(feature_aboves[1678]), .FEAT_BELOW(feature_belows[1678])) ac1678(.scan_win(scan_win1678), .scan_win_std_dev(scan_win_std_dev[1678]), .feature_accum(feature_accums[1678]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1679]), .RECT1_Y(rectangle1_ys[1679]), .RECT1_WIDTH(rectangle1_widths[1679]), .RECT1_HEIGHT(rectangle1_heights[1679]), .RECT1_WEIGHT(rectangle1_weights[1679]), .RECT2_X(rectangle2_xs[1679]), .RECT2_Y(rectangle2_ys[1679]), .RECT2_WIDTH(rectangle2_widths[1679]), .RECT2_HEIGHT(rectangle2_heights[1679]), .RECT2_WEIGHT(rectangle2_weights[1679]), .RECT3_X(rectangle3_xs[1679]), .RECT3_Y(rectangle3_ys[1679]), .RECT3_WIDTH(rectangle3_widths[1679]), .RECT3_HEIGHT(rectangle3_heights[1679]), .RECT3_WEIGHT(rectangle3_weights[1679]), .FEAT_THRES(feature_thresholds[1679]), .FEAT_ABOVE(feature_aboves[1679]), .FEAT_BELOW(feature_belows[1679])) ac1679(.scan_win(scan_win1679), .scan_win_std_dev(scan_win_std_dev[1679]), .feature_accum(feature_accums[1679]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1680]), .RECT1_Y(rectangle1_ys[1680]), .RECT1_WIDTH(rectangle1_widths[1680]), .RECT1_HEIGHT(rectangle1_heights[1680]), .RECT1_WEIGHT(rectangle1_weights[1680]), .RECT2_X(rectangle2_xs[1680]), .RECT2_Y(rectangle2_ys[1680]), .RECT2_WIDTH(rectangle2_widths[1680]), .RECT2_HEIGHT(rectangle2_heights[1680]), .RECT2_WEIGHT(rectangle2_weights[1680]), .RECT3_X(rectangle3_xs[1680]), .RECT3_Y(rectangle3_ys[1680]), .RECT3_WIDTH(rectangle3_widths[1680]), .RECT3_HEIGHT(rectangle3_heights[1680]), .RECT3_WEIGHT(rectangle3_weights[1680]), .FEAT_THRES(feature_thresholds[1680]), .FEAT_ABOVE(feature_aboves[1680]), .FEAT_BELOW(feature_belows[1680])) ac1680(.scan_win(scan_win1680), .scan_win_std_dev(scan_win_std_dev[1680]), .feature_accum(feature_accums[1680]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1681]), .RECT1_Y(rectangle1_ys[1681]), .RECT1_WIDTH(rectangle1_widths[1681]), .RECT1_HEIGHT(rectangle1_heights[1681]), .RECT1_WEIGHT(rectangle1_weights[1681]), .RECT2_X(rectangle2_xs[1681]), .RECT2_Y(rectangle2_ys[1681]), .RECT2_WIDTH(rectangle2_widths[1681]), .RECT2_HEIGHT(rectangle2_heights[1681]), .RECT2_WEIGHT(rectangle2_weights[1681]), .RECT3_X(rectangle3_xs[1681]), .RECT3_Y(rectangle3_ys[1681]), .RECT3_WIDTH(rectangle3_widths[1681]), .RECT3_HEIGHT(rectangle3_heights[1681]), .RECT3_WEIGHT(rectangle3_weights[1681]), .FEAT_THRES(feature_thresholds[1681]), .FEAT_ABOVE(feature_aboves[1681]), .FEAT_BELOW(feature_belows[1681])) ac1681(.scan_win(scan_win1681), .scan_win_std_dev(scan_win_std_dev[1681]), .feature_accum(feature_accums[1681]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1682]), .RECT1_Y(rectangle1_ys[1682]), .RECT1_WIDTH(rectangle1_widths[1682]), .RECT1_HEIGHT(rectangle1_heights[1682]), .RECT1_WEIGHT(rectangle1_weights[1682]), .RECT2_X(rectangle2_xs[1682]), .RECT2_Y(rectangle2_ys[1682]), .RECT2_WIDTH(rectangle2_widths[1682]), .RECT2_HEIGHT(rectangle2_heights[1682]), .RECT2_WEIGHT(rectangle2_weights[1682]), .RECT3_X(rectangle3_xs[1682]), .RECT3_Y(rectangle3_ys[1682]), .RECT3_WIDTH(rectangle3_widths[1682]), .RECT3_HEIGHT(rectangle3_heights[1682]), .RECT3_WEIGHT(rectangle3_weights[1682]), .FEAT_THRES(feature_thresholds[1682]), .FEAT_ABOVE(feature_aboves[1682]), .FEAT_BELOW(feature_belows[1682])) ac1682(.scan_win(scan_win1682), .scan_win_std_dev(scan_win_std_dev[1682]), .feature_accum(feature_accums[1682]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1683]), .RECT1_Y(rectangle1_ys[1683]), .RECT1_WIDTH(rectangle1_widths[1683]), .RECT1_HEIGHT(rectangle1_heights[1683]), .RECT1_WEIGHT(rectangle1_weights[1683]), .RECT2_X(rectangle2_xs[1683]), .RECT2_Y(rectangle2_ys[1683]), .RECT2_WIDTH(rectangle2_widths[1683]), .RECT2_HEIGHT(rectangle2_heights[1683]), .RECT2_WEIGHT(rectangle2_weights[1683]), .RECT3_X(rectangle3_xs[1683]), .RECT3_Y(rectangle3_ys[1683]), .RECT3_WIDTH(rectangle3_widths[1683]), .RECT3_HEIGHT(rectangle3_heights[1683]), .RECT3_WEIGHT(rectangle3_weights[1683]), .FEAT_THRES(feature_thresholds[1683]), .FEAT_ABOVE(feature_aboves[1683]), .FEAT_BELOW(feature_belows[1683])) ac1683(.scan_win(scan_win1683), .scan_win_std_dev(scan_win_std_dev[1683]), .feature_accum(feature_accums[1683]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1684]), .RECT1_Y(rectangle1_ys[1684]), .RECT1_WIDTH(rectangle1_widths[1684]), .RECT1_HEIGHT(rectangle1_heights[1684]), .RECT1_WEIGHT(rectangle1_weights[1684]), .RECT2_X(rectangle2_xs[1684]), .RECT2_Y(rectangle2_ys[1684]), .RECT2_WIDTH(rectangle2_widths[1684]), .RECT2_HEIGHT(rectangle2_heights[1684]), .RECT2_WEIGHT(rectangle2_weights[1684]), .RECT3_X(rectangle3_xs[1684]), .RECT3_Y(rectangle3_ys[1684]), .RECT3_WIDTH(rectangle3_widths[1684]), .RECT3_HEIGHT(rectangle3_heights[1684]), .RECT3_WEIGHT(rectangle3_weights[1684]), .FEAT_THRES(feature_thresholds[1684]), .FEAT_ABOVE(feature_aboves[1684]), .FEAT_BELOW(feature_belows[1684])) ac1684(.scan_win(scan_win1684), .scan_win_std_dev(scan_win_std_dev[1684]), .feature_accum(feature_accums[1684]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1685]), .RECT1_Y(rectangle1_ys[1685]), .RECT1_WIDTH(rectangle1_widths[1685]), .RECT1_HEIGHT(rectangle1_heights[1685]), .RECT1_WEIGHT(rectangle1_weights[1685]), .RECT2_X(rectangle2_xs[1685]), .RECT2_Y(rectangle2_ys[1685]), .RECT2_WIDTH(rectangle2_widths[1685]), .RECT2_HEIGHT(rectangle2_heights[1685]), .RECT2_WEIGHT(rectangle2_weights[1685]), .RECT3_X(rectangle3_xs[1685]), .RECT3_Y(rectangle3_ys[1685]), .RECT3_WIDTH(rectangle3_widths[1685]), .RECT3_HEIGHT(rectangle3_heights[1685]), .RECT3_WEIGHT(rectangle3_weights[1685]), .FEAT_THRES(feature_thresholds[1685]), .FEAT_ABOVE(feature_aboves[1685]), .FEAT_BELOW(feature_belows[1685])) ac1685(.scan_win(scan_win1685), .scan_win_std_dev(scan_win_std_dev[1685]), .feature_accum(feature_accums[1685]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1686]), .RECT1_Y(rectangle1_ys[1686]), .RECT1_WIDTH(rectangle1_widths[1686]), .RECT1_HEIGHT(rectangle1_heights[1686]), .RECT1_WEIGHT(rectangle1_weights[1686]), .RECT2_X(rectangle2_xs[1686]), .RECT2_Y(rectangle2_ys[1686]), .RECT2_WIDTH(rectangle2_widths[1686]), .RECT2_HEIGHT(rectangle2_heights[1686]), .RECT2_WEIGHT(rectangle2_weights[1686]), .RECT3_X(rectangle3_xs[1686]), .RECT3_Y(rectangle3_ys[1686]), .RECT3_WIDTH(rectangle3_widths[1686]), .RECT3_HEIGHT(rectangle3_heights[1686]), .RECT3_WEIGHT(rectangle3_weights[1686]), .FEAT_THRES(feature_thresholds[1686]), .FEAT_ABOVE(feature_aboves[1686]), .FEAT_BELOW(feature_belows[1686])) ac1686(.scan_win(scan_win1686), .scan_win_std_dev(scan_win_std_dev[1686]), .feature_accum(feature_accums[1686]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1687]), .RECT1_Y(rectangle1_ys[1687]), .RECT1_WIDTH(rectangle1_widths[1687]), .RECT1_HEIGHT(rectangle1_heights[1687]), .RECT1_WEIGHT(rectangle1_weights[1687]), .RECT2_X(rectangle2_xs[1687]), .RECT2_Y(rectangle2_ys[1687]), .RECT2_WIDTH(rectangle2_widths[1687]), .RECT2_HEIGHT(rectangle2_heights[1687]), .RECT2_WEIGHT(rectangle2_weights[1687]), .RECT3_X(rectangle3_xs[1687]), .RECT3_Y(rectangle3_ys[1687]), .RECT3_WIDTH(rectangle3_widths[1687]), .RECT3_HEIGHT(rectangle3_heights[1687]), .RECT3_WEIGHT(rectangle3_weights[1687]), .FEAT_THRES(feature_thresholds[1687]), .FEAT_ABOVE(feature_aboves[1687]), .FEAT_BELOW(feature_belows[1687])) ac1687(.scan_win(scan_win1687), .scan_win_std_dev(scan_win_std_dev[1687]), .feature_accum(feature_accums[1687]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1688]), .RECT1_Y(rectangle1_ys[1688]), .RECT1_WIDTH(rectangle1_widths[1688]), .RECT1_HEIGHT(rectangle1_heights[1688]), .RECT1_WEIGHT(rectangle1_weights[1688]), .RECT2_X(rectangle2_xs[1688]), .RECT2_Y(rectangle2_ys[1688]), .RECT2_WIDTH(rectangle2_widths[1688]), .RECT2_HEIGHT(rectangle2_heights[1688]), .RECT2_WEIGHT(rectangle2_weights[1688]), .RECT3_X(rectangle3_xs[1688]), .RECT3_Y(rectangle3_ys[1688]), .RECT3_WIDTH(rectangle3_widths[1688]), .RECT3_HEIGHT(rectangle3_heights[1688]), .RECT3_WEIGHT(rectangle3_weights[1688]), .FEAT_THRES(feature_thresholds[1688]), .FEAT_ABOVE(feature_aboves[1688]), .FEAT_BELOW(feature_belows[1688])) ac1688(.scan_win(scan_win1688), .scan_win_std_dev(scan_win_std_dev[1688]), .feature_accum(feature_accums[1688]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1689]), .RECT1_Y(rectangle1_ys[1689]), .RECT1_WIDTH(rectangle1_widths[1689]), .RECT1_HEIGHT(rectangle1_heights[1689]), .RECT1_WEIGHT(rectangle1_weights[1689]), .RECT2_X(rectangle2_xs[1689]), .RECT2_Y(rectangle2_ys[1689]), .RECT2_WIDTH(rectangle2_widths[1689]), .RECT2_HEIGHT(rectangle2_heights[1689]), .RECT2_WEIGHT(rectangle2_weights[1689]), .RECT3_X(rectangle3_xs[1689]), .RECT3_Y(rectangle3_ys[1689]), .RECT3_WIDTH(rectangle3_widths[1689]), .RECT3_HEIGHT(rectangle3_heights[1689]), .RECT3_WEIGHT(rectangle3_weights[1689]), .FEAT_THRES(feature_thresholds[1689]), .FEAT_ABOVE(feature_aboves[1689]), .FEAT_BELOW(feature_belows[1689])) ac1689(.scan_win(scan_win1689), .scan_win_std_dev(scan_win_std_dev[1689]), .feature_accum(feature_accums[1689]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1690]), .RECT1_Y(rectangle1_ys[1690]), .RECT1_WIDTH(rectangle1_widths[1690]), .RECT1_HEIGHT(rectangle1_heights[1690]), .RECT1_WEIGHT(rectangle1_weights[1690]), .RECT2_X(rectangle2_xs[1690]), .RECT2_Y(rectangle2_ys[1690]), .RECT2_WIDTH(rectangle2_widths[1690]), .RECT2_HEIGHT(rectangle2_heights[1690]), .RECT2_WEIGHT(rectangle2_weights[1690]), .RECT3_X(rectangle3_xs[1690]), .RECT3_Y(rectangle3_ys[1690]), .RECT3_WIDTH(rectangle3_widths[1690]), .RECT3_HEIGHT(rectangle3_heights[1690]), .RECT3_WEIGHT(rectangle3_weights[1690]), .FEAT_THRES(feature_thresholds[1690]), .FEAT_ABOVE(feature_aboves[1690]), .FEAT_BELOW(feature_belows[1690])) ac1690(.scan_win(scan_win1690), .scan_win_std_dev(scan_win_std_dev[1690]), .feature_accum(feature_accums[1690]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1691]), .RECT1_Y(rectangle1_ys[1691]), .RECT1_WIDTH(rectangle1_widths[1691]), .RECT1_HEIGHT(rectangle1_heights[1691]), .RECT1_WEIGHT(rectangle1_weights[1691]), .RECT2_X(rectangle2_xs[1691]), .RECT2_Y(rectangle2_ys[1691]), .RECT2_WIDTH(rectangle2_widths[1691]), .RECT2_HEIGHT(rectangle2_heights[1691]), .RECT2_WEIGHT(rectangle2_weights[1691]), .RECT3_X(rectangle3_xs[1691]), .RECT3_Y(rectangle3_ys[1691]), .RECT3_WIDTH(rectangle3_widths[1691]), .RECT3_HEIGHT(rectangle3_heights[1691]), .RECT3_WEIGHT(rectangle3_weights[1691]), .FEAT_THRES(feature_thresholds[1691]), .FEAT_ABOVE(feature_aboves[1691]), .FEAT_BELOW(feature_belows[1691])) ac1691(.scan_win(scan_win1691), .scan_win_std_dev(scan_win_std_dev[1691]), .feature_accum(feature_accums[1691]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1692]), .RECT1_Y(rectangle1_ys[1692]), .RECT1_WIDTH(rectangle1_widths[1692]), .RECT1_HEIGHT(rectangle1_heights[1692]), .RECT1_WEIGHT(rectangle1_weights[1692]), .RECT2_X(rectangle2_xs[1692]), .RECT2_Y(rectangle2_ys[1692]), .RECT2_WIDTH(rectangle2_widths[1692]), .RECT2_HEIGHT(rectangle2_heights[1692]), .RECT2_WEIGHT(rectangle2_weights[1692]), .RECT3_X(rectangle3_xs[1692]), .RECT3_Y(rectangle3_ys[1692]), .RECT3_WIDTH(rectangle3_widths[1692]), .RECT3_HEIGHT(rectangle3_heights[1692]), .RECT3_WEIGHT(rectangle3_weights[1692]), .FEAT_THRES(feature_thresholds[1692]), .FEAT_ABOVE(feature_aboves[1692]), .FEAT_BELOW(feature_belows[1692])) ac1692(.scan_win(scan_win1692), .scan_win_std_dev(scan_win_std_dev[1692]), .feature_accum(feature_accums[1692]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1693]), .RECT1_Y(rectangle1_ys[1693]), .RECT1_WIDTH(rectangle1_widths[1693]), .RECT1_HEIGHT(rectangle1_heights[1693]), .RECT1_WEIGHT(rectangle1_weights[1693]), .RECT2_X(rectangle2_xs[1693]), .RECT2_Y(rectangle2_ys[1693]), .RECT2_WIDTH(rectangle2_widths[1693]), .RECT2_HEIGHT(rectangle2_heights[1693]), .RECT2_WEIGHT(rectangle2_weights[1693]), .RECT3_X(rectangle3_xs[1693]), .RECT3_Y(rectangle3_ys[1693]), .RECT3_WIDTH(rectangle3_widths[1693]), .RECT3_HEIGHT(rectangle3_heights[1693]), .RECT3_WEIGHT(rectangle3_weights[1693]), .FEAT_THRES(feature_thresholds[1693]), .FEAT_ABOVE(feature_aboves[1693]), .FEAT_BELOW(feature_belows[1693])) ac1693(.scan_win(scan_win1693), .scan_win_std_dev(scan_win_std_dev[1693]), .feature_accum(feature_accums[1693]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1694]), .RECT1_Y(rectangle1_ys[1694]), .RECT1_WIDTH(rectangle1_widths[1694]), .RECT1_HEIGHT(rectangle1_heights[1694]), .RECT1_WEIGHT(rectangle1_weights[1694]), .RECT2_X(rectangle2_xs[1694]), .RECT2_Y(rectangle2_ys[1694]), .RECT2_WIDTH(rectangle2_widths[1694]), .RECT2_HEIGHT(rectangle2_heights[1694]), .RECT2_WEIGHT(rectangle2_weights[1694]), .RECT3_X(rectangle3_xs[1694]), .RECT3_Y(rectangle3_ys[1694]), .RECT3_WIDTH(rectangle3_widths[1694]), .RECT3_HEIGHT(rectangle3_heights[1694]), .RECT3_WEIGHT(rectangle3_weights[1694]), .FEAT_THRES(feature_thresholds[1694]), .FEAT_ABOVE(feature_aboves[1694]), .FEAT_BELOW(feature_belows[1694])) ac1694(.scan_win(scan_win1694), .scan_win_std_dev(scan_win_std_dev[1694]), .feature_accum(feature_accums[1694]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1695]), .RECT1_Y(rectangle1_ys[1695]), .RECT1_WIDTH(rectangle1_widths[1695]), .RECT1_HEIGHT(rectangle1_heights[1695]), .RECT1_WEIGHT(rectangle1_weights[1695]), .RECT2_X(rectangle2_xs[1695]), .RECT2_Y(rectangle2_ys[1695]), .RECT2_WIDTH(rectangle2_widths[1695]), .RECT2_HEIGHT(rectangle2_heights[1695]), .RECT2_WEIGHT(rectangle2_weights[1695]), .RECT3_X(rectangle3_xs[1695]), .RECT3_Y(rectangle3_ys[1695]), .RECT3_WIDTH(rectangle3_widths[1695]), .RECT3_HEIGHT(rectangle3_heights[1695]), .RECT3_WEIGHT(rectangle3_weights[1695]), .FEAT_THRES(feature_thresholds[1695]), .FEAT_ABOVE(feature_aboves[1695]), .FEAT_BELOW(feature_belows[1695])) ac1695(.scan_win(scan_win1695), .scan_win_std_dev(scan_win_std_dev[1695]), .feature_accum(feature_accums[1695]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1696]), .RECT1_Y(rectangle1_ys[1696]), .RECT1_WIDTH(rectangle1_widths[1696]), .RECT1_HEIGHT(rectangle1_heights[1696]), .RECT1_WEIGHT(rectangle1_weights[1696]), .RECT2_X(rectangle2_xs[1696]), .RECT2_Y(rectangle2_ys[1696]), .RECT2_WIDTH(rectangle2_widths[1696]), .RECT2_HEIGHT(rectangle2_heights[1696]), .RECT2_WEIGHT(rectangle2_weights[1696]), .RECT3_X(rectangle3_xs[1696]), .RECT3_Y(rectangle3_ys[1696]), .RECT3_WIDTH(rectangle3_widths[1696]), .RECT3_HEIGHT(rectangle3_heights[1696]), .RECT3_WEIGHT(rectangle3_weights[1696]), .FEAT_THRES(feature_thresholds[1696]), .FEAT_ABOVE(feature_aboves[1696]), .FEAT_BELOW(feature_belows[1696])) ac1696(.scan_win(scan_win1696), .scan_win_std_dev(scan_win_std_dev[1696]), .feature_accum(feature_accums[1696]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1697]), .RECT1_Y(rectangle1_ys[1697]), .RECT1_WIDTH(rectangle1_widths[1697]), .RECT1_HEIGHT(rectangle1_heights[1697]), .RECT1_WEIGHT(rectangle1_weights[1697]), .RECT2_X(rectangle2_xs[1697]), .RECT2_Y(rectangle2_ys[1697]), .RECT2_WIDTH(rectangle2_widths[1697]), .RECT2_HEIGHT(rectangle2_heights[1697]), .RECT2_WEIGHT(rectangle2_weights[1697]), .RECT3_X(rectangle3_xs[1697]), .RECT3_Y(rectangle3_ys[1697]), .RECT3_WIDTH(rectangle3_widths[1697]), .RECT3_HEIGHT(rectangle3_heights[1697]), .RECT3_WEIGHT(rectangle3_weights[1697]), .FEAT_THRES(feature_thresholds[1697]), .FEAT_ABOVE(feature_aboves[1697]), .FEAT_BELOW(feature_belows[1697])) ac1697(.scan_win(scan_win1697), .scan_win_std_dev(scan_win_std_dev[1697]), .feature_accum(feature_accums[1697]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1698]), .RECT1_Y(rectangle1_ys[1698]), .RECT1_WIDTH(rectangle1_widths[1698]), .RECT1_HEIGHT(rectangle1_heights[1698]), .RECT1_WEIGHT(rectangle1_weights[1698]), .RECT2_X(rectangle2_xs[1698]), .RECT2_Y(rectangle2_ys[1698]), .RECT2_WIDTH(rectangle2_widths[1698]), .RECT2_HEIGHT(rectangle2_heights[1698]), .RECT2_WEIGHT(rectangle2_weights[1698]), .RECT3_X(rectangle3_xs[1698]), .RECT3_Y(rectangle3_ys[1698]), .RECT3_WIDTH(rectangle3_widths[1698]), .RECT3_HEIGHT(rectangle3_heights[1698]), .RECT3_WEIGHT(rectangle3_weights[1698]), .FEAT_THRES(feature_thresholds[1698]), .FEAT_ABOVE(feature_aboves[1698]), .FEAT_BELOW(feature_belows[1698])) ac1698(.scan_win(scan_win1698), .scan_win_std_dev(scan_win_std_dev[1698]), .feature_accum(feature_accums[1698]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1699]), .RECT1_Y(rectangle1_ys[1699]), .RECT1_WIDTH(rectangle1_widths[1699]), .RECT1_HEIGHT(rectangle1_heights[1699]), .RECT1_WEIGHT(rectangle1_weights[1699]), .RECT2_X(rectangle2_xs[1699]), .RECT2_Y(rectangle2_ys[1699]), .RECT2_WIDTH(rectangle2_widths[1699]), .RECT2_HEIGHT(rectangle2_heights[1699]), .RECT2_WEIGHT(rectangle2_weights[1699]), .RECT3_X(rectangle3_xs[1699]), .RECT3_Y(rectangle3_ys[1699]), .RECT3_WIDTH(rectangle3_widths[1699]), .RECT3_HEIGHT(rectangle3_heights[1699]), .RECT3_WEIGHT(rectangle3_weights[1699]), .FEAT_THRES(feature_thresholds[1699]), .FEAT_ABOVE(feature_aboves[1699]), .FEAT_BELOW(feature_belows[1699])) ac1699(.scan_win(scan_win1699), .scan_win_std_dev(scan_win_std_dev[1699]), .feature_accum(feature_accums[1699]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1700]), .RECT1_Y(rectangle1_ys[1700]), .RECT1_WIDTH(rectangle1_widths[1700]), .RECT1_HEIGHT(rectangle1_heights[1700]), .RECT1_WEIGHT(rectangle1_weights[1700]), .RECT2_X(rectangle2_xs[1700]), .RECT2_Y(rectangle2_ys[1700]), .RECT2_WIDTH(rectangle2_widths[1700]), .RECT2_HEIGHT(rectangle2_heights[1700]), .RECT2_WEIGHT(rectangle2_weights[1700]), .RECT3_X(rectangle3_xs[1700]), .RECT3_Y(rectangle3_ys[1700]), .RECT3_WIDTH(rectangle3_widths[1700]), .RECT3_HEIGHT(rectangle3_heights[1700]), .RECT3_WEIGHT(rectangle3_weights[1700]), .FEAT_THRES(feature_thresholds[1700]), .FEAT_ABOVE(feature_aboves[1700]), .FEAT_BELOW(feature_belows[1700])) ac1700(.scan_win(scan_win1700), .scan_win_std_dev(scan_win_std_dev[1700]), .feature_accum(feature_accums[1700]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1701]), .RECT1_Y(rectangle1_ys[1701]), .RECT1_WIDTH(rectangle1_widths[1701]), .RECT1_HEIGHT(rectangle1_heights[1701]), .RECT1_WEIGHT(rectangle1_weights[1701]), .RECT2_X(rectangle2_xs[1701]), .RECT2_Y(rectangle2_ys[1701]), .RECT2_WIDTH(rectangle2_widths[1701]), .RECT2_HEIGHT(rectangle2_heights[1701]), .RECT2_WEIGHT(rectangle2_weights[1701]), .RECT3_X(rectangle3_xs[1701]), .RECT3_Y(rectangle3_ys[1701]), .RECT3_WIDTH(rectangle3_widths[1701]), .RECT3_HEIGHT(rectangle3_heights[1701]), .RECT3_WEIGHT(rectangle3_weights[1701]), .FEAT_THRES(feature_thresholds[1701]), .FEAT_ABOVE(feature_aboves[1701]), .FEAT_BELOW(feature_belows[1701])) ac1701(.scan_win(scan_win1701), .scan_win_std_dev(scan_win_std_dev[1701]), .feature_accum(feature_accums[1701]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1702]), .RECT1_Y(rectangle1_ys[1702]), .RECT1_WIDTH(rectangle1_widths[1702]), .RECT1_HEIGHT(rectangle1_heights[1702]), .RECT1_WEIGHT(rectangle1_weights[1702]), .RECT2_X(rectangle2_xs[1702]), .RECT2_Y(rectangle2_ys[1702]), .RECT2_WIDTH(rectangle2_widths[1702]), .RECT2_HEIGHT(rectangle2_heights[1702]), .RECT2_WEIGHT(rectangle2_weights[1702]), .RECT3_X(rectangle3_xs[1702]), .RECT3_Y(rectangle3_ys[1702]), .RECT3_WIDTH(rectangle3_widths[1702]), .RECT3_HEIGHT(rectangle3_heights[1702]), .RECT3_WEIGHT(rectangle3_weights[1702]), .FEAT_THRES(feature_thresholds[1702]), .FEAT_ABOVE(feature_aboves[1702]), .FEAT_BELOW(feature_belows[1702])) ac1702(.scan_win(scan_win1702), .scan_win_std_dev(scan_win_std_dev[1702]), .feature_accum(feature_accums[1702]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1703]), .RECT1_Y(rectangle1_ys[1703]), .RECT1_WIDTH(rectangle1_widths[1703]), .RECT1_HEIGHT(rectangle1_heights[1703]), .RECT1_WEIGHT(rectangle1_weights[1703]), .RECT2_X(rectangle2_xs[1703]), .RECT2_Y(rectangle2_ys[1703]), .RECT2_WIDTH(rectangle2_widths[1703]), .RECT2_HEIGHT(rectangle2_heights[1703]), .RECT2_WEIGHT(rectangle2_weights[1703]), .RECT3_X(rectangle3_xs[1703]), .RECT3_Y(rectangle3_ys[1703]), .RECT3_WIDTH(rectangle3_widths[1703]), .RECT3_HEIGHT(rectangle3_heights[1703]), .RECT3_WEIGHT(rectangle3_weights[1703]), .FEAT_THRES(feature_thresholds[1703]), .FEAT_ABOVE(feature_aboves[1703]), .FEAT_BELOW(feature_belows[1703])) ac1703(.scan_win(scan_win1703), .scan_win_std_dev(scan_win_std_dev[1703]), .feature_accum(feature_accums[1703]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1704]), .RECT1_Y(rectangle1_ys[1704]), .RECT1_WIDTH(rectangle1_widths[1704]), .RECT1_HEIGHT(rectangle1_heights[1704]), .RECT1_WEIGHT(rectangle1_weights[1704]), .RECT2_X(rectangle2_xs[1704]), .RECT2_Y(rectangle2_ys[1704]), .RECT2_WIDTH(rectangle2_widths[1704]), .RECT2_HEIGHT(rectangle2_heights[1704]), .RECT2_WEIGHT(rectangle2_weights[1704]), .RECT3_X(rectangle3_xs[1704]), .RECT3_Y(rectangle3_ys[1704]), .RECT3_WIDTH(rectangle3_widths[1704]), .RECT3_HEIGHT(rectangle3_heights[1704]), .RECT3_WEIGHT(rectangle3_weights[1704]), .FEAT_THRES(feature_thresholds[1704]), .FEAT_ABOVE(feature_aboves[1704]), .FEAT_BELOW(feature_belows[1704])) ac1704(.scan_win(scan_win1704), .scan_win_std_dev(scan_win_std_dev[1704]), .feature_accum(feature_accums[1704]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1705]), .RECT1_Y(rectangle1_ys[1705]), .RECT1_WIDTH(rectangle1_widths[1705]), .RECT1_HEIGHT(rectangle1_heights[1705]), .RECT1_WEIGHT(rectangle1_weights[1705]), .RECT2_X(rectangle2_xs[1705]), .RECT2_Y(rectangle2_ys[1705]), .RECT2_WIDTH(rectangle2_widths[1705]), .RECT2_HEIGHT(rectangle2_heights[1705]), .RECT2_WEIGHT(rectangle2_weights[1705]), .RECT3_X(rectangle3_xs[1705]), .RECT3_Y(rectangle3_ys[1705]), .RECT3_WIDTH(rectangle3_widths[1705]), .RECT3_HEIGHT(rectangle3_heights[1705]), .RECT3_WEIGHT(rectangle3_weights[1705]), .FEAT_THRES(feature_thresholds[1705]), .FEAT_ABOVE(feature_aboves[1705]), .FEAT_BELOW(feature_belows[1705])) ac1705(.scan_win(scan_win1705), .scan_win_std_dev(scan_win_std_dev[1705]), .feature_accum(feature_accums[1705]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1706]), .RECT1_Y(rectangle1_ys[1706]), .RECT1_WIDTH(rectangle1_widths[1706]), .RECT1_HEIGHT(rectangle1_heights[1706]), .RECT1_WEIGHT(rectangle1_weights[1706]), .RECT2_X(rectangle2_xs[1706]), .RECT2_Y(rectangle2_ys[1706]), .RECT2_WIDTH(rectangle2_widths[1706]), .RECT2_HEIGHT(rectangle2_heights[1706]), .RECT2_WEIGHT(rectangle2_weights[1706]), .RECT3_X(rectangle3_xs[1706]), .RECT3_Y(rectangle3_ys[1706]), .RECT3_WIDTH(rectangle3_widths[1706]), .RECT3_HEIGHT(rectangle3_heights[1706]), .RECT3_WEIGHT(rectangle3_weights[1706]), .FEAT_THRES(feature_thresholds[1706]), .FEAT_ABOVE(feature_aboves[1706]), .FEAT_BELOW(feature_belows[1706])) ac1706(.scan_win(scan_win1706), .scan_win_std_dev(scan_win_std_dev[1706]), .feature_accum(feature_accums[1706]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1707]), .RECT1_Y(rectangle1_ys[1707]), .RECT1_WIDTH(rectangle1_widths[1707]), .RECT1_HEIGHT(rectangle1_heights[1707]), .RECT1_WEIGHT(rectangle1_weights[1707]), .RECT2_X(rectangle2_xs[1707]), .RECT2_Y(rectangle2_ys[1707]), .RECT2_WIDTH(rectangle2_widths[1707]), .RECT2_HEIGHT(rectangle2_heights[1707]), .RECT2_WEIGHT(rectangle2_weights[1707]), .RECT3_X(rectangle3_xs[1707]), .RECT3_Y(rectangle3_ys[1707]), .RECT3_WIDTH(rectangle3_widths[1707]), .RECT3_HEIGHT(rectangle3_heights[1707]), .RECT3_WEIGHT(rectangle3_weights[1707]), .FEAT_THRES(feature_thresholds[1707]), .FEAT_ABOVE(feature_aboves[1707]), .FEAT_BELOW(feature_belows[1707])) ac1707(.scan_win(scan_win1707), .scan_win_std_dev(scan_win_std_dev[1707]), .feature_accum(feature_accums[1707]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1708]), .RECT1_Y(rectangle1_ys[1708]), .RECT1_WIDTH(rectangle1_widths[1708]), .RECT1_HEIGHT(rectangle1_heights[1708]), .RECT1_WEIGHT(rectangle1_weights[1708]), .RECT2_X(rectangle2_xs[1708]), .RECT2_Y(rectangle2_ys[1708]), .RECT2_WIDTH(rectangle2_widths[1708]), .RECT2_HEIGHT(rectangle2_heights[1708]), .RECT2_WEIGHT(rectangle2_weights[1708]), .RECT3_X(rectangle3_xs[1708]), .RECT3_Y(rectangle3_ys[1708]), .RECT3_WIDTH(rectangle3_widths[1708]), .RECT3_HEIGHT(rectangle3_heights[1708]), .RECT3_WEIGHT(rectangle3_weights[1708]), .FEAT_THRES(feature_thresholds[1708]), .FEAT_ABOVE(feature_aboves[1708]), .FEAT_BELOW(feature_belows[1708])) ac1708(.scan_win(scan_win1708), .scan_win_std_dev(scan_win_std_dev[1708]), .feature_accum(feature_accums[1708]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1709]), .RECT1_Y(rectangle1_ys[1709]), .RECT1_WIDTH(rectangle1_widths[1709]), .RECT1_HEIGHT(rectangle1_heights[1709]), .RECT1_WEIGHT(rectangle1_weights[1709]), .RECT2_X(rectangle2_xs[1709]), .RECT2_Y(rectangle2_ys[1709]), .RECT2_WIDTH(rectangle2_widths[1709]), .RECT2_HEIGHT(rectangle2_heights[1709]), .RECT2_WEIGHT(rectangle2_weights[1709]), .RECT3_X(rectangle3_xs[1709]), .RECT3_Y(rectangle3_ys[1709]), .RECT3_WIDTH(rectangle3_widths[1709]), .RECT3_HEIGHT(rectangle3_heights[1709]), .RECT3_WEIGHT(rectangle3_weights[1709]), .FEAT_THRES(feature_thresholds[1709]), .FEAT_ABOVE(feature_aboves[1709]), .FEAT_BELOW(feature_belows[1709])) ac1709(.scan_win(scan_win1709), .scan_win_std_dev(scan_win_std_dev[1709]), .feature_accum(feature_accums[1709]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1710]), .RECT1_Y(rectangle1_ys[1710]), .RECT1_WIDTH(rectangle1_widths[1710]), .RECT1_HEIGHT(rectangle1_heights[1710]), .RECT1_WEIGHT(rectangle1_weights[1710]), .RECT2_X(rectangle2_xs[1710]), .RECT2_Y(rectangle2_ys[1710]), .RECT2_WIDTH(rectangle2_widths[1710]), .RECT2_HEIGHT(rectangle2_heights[1710]), .RECT2_WEIGHT(rectangle2_weights[1710]), .RECT3_X(rectangle3_xs[1710]), .RECT3_Y(rectangle3_ys[1710]), .RECT3_WIDTH(rectangle3_widths[1710]), .RECT3_HEIGHT(rectangle3_heights[1710]), .RECT3_WEIGHT(rectangle3_weights[1710]), .FEAT_THRES(feature_thresholds[1710]), .FEAT_ABOVE(feature_aboves[1710]), .FEAT_BELOW(feature_belows[1710])) ac1710(.scan_win(scan_win1710), .scan_win_std_dev(scan_win_std_dev[1710]), .feature_accum(feature_accums[1710]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1711]), .RECT1_Y(rectangle1_ys[1711]), .RECT1_WIDTH(rectangle1_widths[1711]), .RECT1_HEIGHT(rectangle1_heights[1711]), .RECT1_WEIGHT(rectangle1_weights[1711]), .RECT2_X(rectangle2_xs[1711]), .RECT2_Y(rectangle2_ys[1711]), .RECT2_WIDTH(rectangle2_widths[1711]), .RECT2_HEIGHT(rectangle2_heights[1711]), .RECT2_WEIGHT(rectangle2_weights[1711]), .RECT3_X(rectangle3_xs[1711]), .RECT3_Y(rectangle3_ys[1711]), .RECT3_WIDTH(rectangle3_widths[1711]), .RECT3_HEIGHT(rectangle3_heights[1711]), .RECT3_WEIGHT(rectangle3_weights[1711]), .FEAT_THRES(feature_thresholds[1711]), .FEAT_ABOVE(feature_aboves[1711]), .FEAT_BELOW(feature_belows[1711])) ac1711(.scan_win(scan_win1711), .scan_win_std_dev(scan_win_std_dev[1711]), .feature_accum(feature_accums[1711]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1712]), .RECT1_Y(rectangle1_ys[1712]), .RECT1_WIDTH(rectangle1_widths[1712]), .RECT1_HEIGHT(rectangle1_heights[1712]), .RECT1_WEIGHT(rectangle1_weights[1712]), .RECT2_X(rectangle2_xs[1712]), .RECT2_Y(rectangle2_ys[1712]), .RECT2_WIDTH(rectangle2_widths[1712]), .RECT2_HEIGHT(rectangle2_heights[1712]), .RECT2_WEIGHT(rectangle2_weights[1712]), .RECT3_X(rectangle3_xs[1712]), .RECT3_Y(rectangle3_ys[1712]), .RECT3_WIDTH(rectangle3_widths[1712]), .RECT3_HEIGHT(rectangle3_heights[1712]), .RECT3_WEIGHT(rectangle3_weights[1712]), .FEAT_THRES(feature_thresholds[1712]), .FEAT_ABOVE(feature_aboves[1712]), .FEAT_BELOW(feature_belows[1712])) ac1712(.scan_win(scan_win1712), .scan_win_std_dev(scan_win_std_dev[1712]), .feature_accum(feature_accums[1712]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1713]), .RECT1_Y(rectangle1_ys[1713]), .RECT1_WIDTH(rectangle1_widths[1713]), .RECT1_HEIGHT(rectangle1_heights[1713]), .RECT1_WEIGHT(rectangle1_weights[1713]), .RECT2_X(rectangle2_xs[1713]), .RECT2_Y(rectangle2_ys[1713]), .RECT2_WIDTH(rectangle2_widths[1713]), .RECT2_HEIGHT(rectangle2_heights[1713]), .RECT2_WEIGHT(rectangle2_weights[1713]), .RECT3_X(rectangle3_xs[1713]), .RECT3_Y(rectangle3_ys[1713]), .RECT3_WIDTH(rectangle3_widths[1713]), .RECT3_HEIGHT(rectangle3_heights[1713]), .RECT3_WEIGHT(rectangle3_weights[1713]), .FEAT_THRES(feature_thresholds[1713]), .FEAT_ABOVE(feature_aboves[1713]), .FEAT_BELOW(feature_belows[1713])) ac1713(.scan_win(scan_win1713), .scan_win_std_dev(scan_win_std_dev[1713]), .feature_accum(feature_accums[1713]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1714]), .RECT1_Y(rectangle1_ys[1714]), .RECT1_WIDTH(rectangle1_widths[1714]), .RECT1_HEIGHT(rectangle1_heights[1714]), .RECT1_WEIGHT(rectangle1_weights[1714]), .RECT2_X(rectangle2_xs[1714]), .RECT2_Y(rectangle2_ys[1714]), .RECT2_WIDTH(rectangle2_widths[1714]), .RECT2_HEIGHT(rectangle2_heights[1714]), .RECT2_WEIGHT(rectangle2_weights[1714]), .RECT3_X(rectangle3_xs[1714]), .RECT3_Y(rectangle3_ys[1714]), .RECT3_WIDTH(rectangle3_widths[1714]), .RECT3_HEIGHT(rectangle3_heights[1714]), .RECT3_WEIGHT(rectangle3_weights[1714]), .FEAT_THRES(feature_thresholds[1714]), .FEAT_ABOVE(feature_aboves[1714]), .FEAT_BELOW(feature_belows[1714])) ac1714(.scan_win(scan_win1714), .scan_win_std_dev(scan_win_std_dev[1714]), .feature_accum(feature_accums[1714]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1715]), .RECT1_Y(rectangle1_ys[1715]), .RECT1_WIDTH(rectangle1_widths[1715]), .RECT1_HEIGHT(rectangle1_heights[1715]), .RECT1_WEIGHT(rectangle1_weights[1715]), .RECT2_X(rectangle2_xs[1715]), .RECT2_Y(rectangle2_ys[1715]), .RECT2_WIDTH(rectangle2_widths[1715]), .RECT2_HEIGHT(rectangle2_heights[1715]), .RECT2_WEIGHT(rectangle2_weights[1715]), .RECT3_X(rectangle3_xs[1715]), .RECT3_Y(rectangle3_ys[1715]), .RECT3_WIDTH(rectangle3_widths[1715]), .RECT3_HEIGHT(rectangle3_heights[1715]), .RECT3_WEIGHT(rectangle3_weights[1715]), .FEAT_THRES(feature_thresholds[1715]), .FEAT_ABOVE(feature_aboves[1715]), .FEAT_BELOW(feature_belows[1715])) ac1715(.scan_win(scan_win1715), .scan_win_std_dev(scan_win_std_dev[1715]), .feature_accum(feature_accums[1715]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1716]), .RECT1_Y(rectangle1_ys[1716]), .RECT1_WIDTH(rectangle1_widths[1716]), .RECT1_HEIGHT(rectangle1_heights[1716]), .RECT1_WEIGHT(rectangle1_weights[1716]), .RECT2_X(rectangle2_xs[1716]), .RECT2_Y(rectangle2_ys[1716]), .RECT2_WIDTH(rectangle2_widths[1716]), .RECT2_HEIGHT(rectangle2_heights[1716]), .RECT2_WEIGHT(rectangle2_weights[1716]), .RECT3_X(rectangle3_xs[1716]), .RECT3_Y(rectangle3_ys[1716]), .RECT3_WIDTH(rectangle3_widths[1716]), .RECT3_HEIGHT(rectangle3_heights[1716]), .RECT3_WEIGHT(rectangle3_weights[1716]), .FEAT_THRES(feature_thresholds[1716]), .FEAT_ABOVE(feature_aboves[1716]), .FEAT_BELOW(feature_belows[1716])) ac1716(.scan_win(scan_win1716), .scan_win_std_dev(scan_win_std_dev[1716]), .feature_accum(feature_accums[1716]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1717]), .RECT1_Y(rectangle1_ys[1717]), .RECT1_WIDTH(rectangle1_widths[1717]), .RECT1_HEIGHT(rectangle1_heights[1717]), .RECT1_WEIGHT(rectangle1_weights[1717]), .RECT2_X(rectangle2_xs[1717]), .RECT2_Y(rectangle2_ys[1717]), .RECT2_WIDTH(rectangle2_widths[1717]), .RECT2_HEIGHT(rectangle2_heights[1717]), .RECT2_WEIGHT(rectangle2_weights[1717]), .RECT3_X(rectangle3_xs[1717]), .RECT3_Y(rectangle3_ys[1717]), .RECT3_WIDTH(rectangle3_widths[1717]), .RECT3_HEIGHT(rectangle3_heights[1717]), .RECT3_WEIGHT(rectangle3_weights[1717]), .FEAT_THRES(feature_thresholds[1717]), .FEAT_ABOVE(feature_aboves[1717]), .FEAT_BELOW(feature_belows[1717])) ac1717(.scan_win(scan_win1717), .scan_win_std_dev(scan_win_std_dev[1717]), .feature_accum(feature_accums[1717]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1718]), .RECT1_Y(rectangle1_ys[1718]), .RECT1_WIDTH(rectangle1_widths[1718]), .RECT1_HEIGHT(rectangle1_heights[1718]), .RECT1_WEIGHT(rectangle1_weights[1718]), .RECT2_X(rectangle2_xs[1718]), .RECT2_Y(rectangle2_ys[1718]), .RECT2_WIDTH(rectangle2_widths[1718]), .RECT2_HEIGHT(rectangle2_heights[1718]), .RECT2_WEIGHT(rectangle2_weights[1718]), .RECT3_X(rectangle3_xs[1718]), .RECT3_Y(rectangle3_ys[1718]), .RECT3_WIDTH(rectangle3_widths[1718]), .RECT3_HEIGHT(rectangle3_heights[1718]), .RECT3_WEIGHT(rectangle3_weights[1718]), .FEAT_THRES(feature_thresholds[1718]), .FEAT_ABOVE(feature_aboves[1718]), .FEAT_BELOW(feature_belows[1718])) ac1718(.scan_win(scan_win1718), .scan_win_std_dev(scan_win_std_dev[1718]), .feature_accum(feature_accums[1718]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1719]), .RECT1_Y(rectangle1_ys[1719]), .RECT1_WIDTH(rectangle1_widths[1719]), .RECT1_HEIGHT(rectangle1_heights[1719]), .RECT1_WEIGHT(rectangle1_weights[1719]), .RECT2_X(rectangle2_xs[1719]), .RECT2_Y(rectangle2_ys[1719]), .RECT2_WIDTH(rectangle2_widths[1719]), .RECT2_HEIGHT(rectangle2_heights[1719]), .RECT2_WEIGHT(rectangle2_weights[1719]), .RECT3_X(rectangle3_xs[1719]), .RECT3_Y(rectangle3_ys[1719]), .RECT3_WIDTH(rectangle3_widths[1719]), .RECT3_HEIGHT(rectangle3_heights[1719]), .RECT3_WEIGHT(rectangle3_weights[1719]), .FEAT_THRES(feature_thresholds[1719]), .FEAT_ABOVE(feature_aboves[1719]), .FEAT_BELOW(feature_belows[1719])) ac1719(.scan_win(scan_win1719), .scan_win_std_dev(scan_win_std_dev[1719]), .feature_accum(feature_accums[1719]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1720]), .RECT1_Y(rectangle1_ys[1720]), .RECT1_WIDTH(rectangle1_widths[1720]), .RECT1_HEIGHT(rectangle1_heights[1720]), .RECT1_WEIGHT(rectangle1_weights[1720]), .RECT2_X(rectangle2_xs[1720]), .RECT2_Y(rectangle2_ys[1720]), .RECT2_WIDTH(rectangle2_widths[1720]), .RECT2_HEIGHT(rectangle2_heights[1720]), .RECT2_WEIGHT(rectangle2_weights[1720]), .RECT3_X(rectangle3_xs[1720]), .RECT3_Y(rectangle3_ys[1720]), .RECT3_WIDTH(rectangle3_widths[1720]), .RECT3_HEIGHT(rectangle3_heights[1720]), .RECT3_WEIGHT(rectangle3_weights[1720]), .FEAT_THRES(feature_thresholds[1720]), .FEAT_ABOVE(feature_aboves[1720]), .FEAT_BELOW(feature_belows[1720])) ac1720(.scan_win(scan_win1720), .scan_win_std_dev(scan_win_std_dev[1720]), .feature_accum(feature_accums[1720]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1721]), .RECT1_Y(rectangle1_ys[1721]), .RECT1_WIDTH(rectangle1_widths[1721]), .RECT1_HEIGHT(rectangle1_heights[1721]), .RECT1_WEIGHT(rectangle1_weights[1721]), .RECT2_X(rectangle2_xs[1721]), .RECT2_Y(rectangle2_ys[1721]), .RECT2_WIDTH(rectangle2_widths[1721]), .RECT2_HEIGHT(rectangle2_heights[1721]), .RECT2_WEIGHT(rectangle2_weights[1721]), .RECT3_X(rectangle3_xs[1721]), .RECT3_Y(rectangle3_ys[1721]), .RECT3_WIDTH(rectangle3_widths[1721]), .RECT3_HEIGHT(rectangle3_heights[1721]), .RECT3_WEIGHT(rectangle3_weights[1721]), .FEAT_THRES(feature_thresholds[1721]), .FEAT_ABOVE(feature_aboves[1721]), .FEAT_BELOW(feature_belows[1721])) ac1721(.scan_win(scan_win1721), .scan_win_std_dev(scan_win_std_dev[1721]), .feature_accum(feature_accums[1721]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1722]), .RECT1_Y(rectangle1_ys[1722]), .RECT1_WIDTH(rectangle1_widths[1722]), .RECT1_HEIGHT(rectangle1_heights[1722]), .RECT1_WEIGHT(rectangle1_weights[1722]), .RECT2_X(rectangle2_xs[1722]), .RECT2_Y(rectangle2_ys[1722]), .RECT2_WIDTH(rectangle2_widths[1722]), .RECT2_HEIGHT(rectangle2_heights[1722]), .RECT2_WEIGHT(rectangle2_weights[1722]), .RECT3_X(rectangle3_xs[1722]), .RECT3_Y(rectangle3_ys[1722]), .RECT3_WIDTH(rectangle3_widths[1722]), .RECT3_HEIGHT(rectangle3_heights[1722]), .RECT3_WEIGHT(rectangle3_weights[1722]), .FEAT_THRES(feature_thresholds[1722]), .FEAT_ABOVE(feature_aboves[1722]), .FEAT_BELOW(feature_belows[1722])) ac1722(.scan_win(scan_win1722), .scan_win_std_dev(scan_win_std_dev[1722]), .feature_accum(feature_accums[1722]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1723]), .RECT1_Y(rectangle1_ys[1723]), .RECT1_WIDTH(rectangle1_widths[1723]), .RECT1_HEIGHT(rectangle1_heights[1723]), .RECT1_WEIGHT(rectangle1_weights[1723]), .RECT2_X(rectangle2_xs[1723]), .RECT2_Y(rectangle2_ys[1723]), .RECT2_WIDTH(rectangle2_widths[1723]), .RECT2_HEIGHT(rectangle2_heights[1723]), .RECT2_WEIGHT(rectangle2_weights[1723]), .RECT3_X(rectangle3_xs[1723]), .RECT3_Y(rectangle3_ys[1723]), .RECT3_WIDTH(rectangle3_widths[1723]), .RECT3_HEIGHT(rectangle3_heights[1723]), .RECT3_WEIGHT(rectangle3_weights[1723]), .FEAT_THRES(feature_thresholds[1723]), .FEAT_ABOVE(feature_aboves[1723]), .FEAT_BELOW(feature_belows[1723])) ac1723(.scan_win(scan_win1723), .scan_win_std_dev(scan_win_std_dev[1723]), .feature_accum(feature_accums[1723]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1724]), .RECT1_Y(rectangle1_ys[1724]), .RECT1_WIDTH(rectangle1_widths[1724]), .RECT1_HEIGHT(rectangle1_heights[1724]), .RECT1_WEIGHT(rectangle1_weights[1724]), .RECT2_X(rectangle2_xs[1724]), .RECT2_Y(rectangle2_ys[1724]), .RECT2_WIDTH(rectangle2_widths[1724]), .RECT2_HEIGHT(rectangle2_heights[1724]), .RECT2_WEIGHT(rectangle2_weights[1724]), .RECT3_X(rectangle3_xs[1724]), .RECT3_Y(rectangle3_ys[1724]), .RECT3_WIDTH(rectangle3_widths[1724]), .RECT3_HEIGHT(rectangle3_heights[1724]), .RECT3_WEIGHT(rectangle3_weights[1724]), .FEAT_THRES(feature_thresholds[1724]), .FEAT_ABOVE(feature_aboves[1724]), .FEAT_BELOW(feature_belows[1724])) ac1724(.scan_win(scan_win1724), .scan_win_std_dev(scan_win_std_dev[1724]), .feature_accum(feature_accums[1724]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1725]), .RECT1_Y(rectangle1_ys[1725]), .RECT1_WIDTH(rectangle1_widths[1725]), .RECT1_HEIGHT(rectangle1_heights[1725]), .RECT1_WEIGHT(rectangle1_weights[1725]), .RECT2_X(rectangle2_xs[1725]), .RECT2_Y(rectangle2_ys[1725]), .RECT2_WIDTH(rectangle2_widths[1725]), .RECT2_HEIGHT(rectangle2_heights[1725]), .RECT2_WEIGHT(rectangle2_weights[1725]), .RECT3_X(rectangle3_xs[1725]), .RECT3_Y(rectangle3_ys[1725]), .RECT3_WIDTH(rectangle3_widths[1725]), .RECT3_HEIGHT(rectangle3_heights[1725]), .RECT3_WEIGHT(rectangle3_weights[1725]), .FEAT_THRES(feature_thresholds[1725]), .FEAT_ABOVE(feature_aboves[1725]), .FEAT_BELOW(feature_belows[1725])) ac1725(.scan_win(scan_win1725), .scan_win_std_dev(scan_win_std_dev[1725]), .feature_accum(feature_accums[1725]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1726]), .RECT1_Y(rectangle1_ys[1726]), .RECT1_WIDTH(rectangle1_widths[1726]), .RECT1_HEIGHT(rectangle1_heights[1726]), .RECT1_WEIGHT(rectangle1_weights[1726]), .RECT2_X(rectangle2_xs[1726]), .RECT2_Y(rectangle2_ys[1726]), .RECT2_WIDTH(rectangle2_widths[1726]), .RECT2_HEIGHT(rectangle2_heights[1726]), .RECT2_WEIGHT(rectangle2_weights[1726]), .RECT3_X(rectangle3_xs[1726]), .RECT3_Y(rectangle3_ys[1726]), .RECT3_WIDTH(rectangle3_widths[1726]), .RECT3_HEIGHT(rectangle3_heights[1726]), .RECT3_WEIGHT(rectangle3_weights[1726]), .FEAT_THRES(feature_thresholds[1726]), .FEAT_ABOVE(feature_aboves[1726]), .FEAT_BELOW(feature_belows[1726])) ac1726(.scan_win(scan_win1726), .scan_win_std_dev(scan_win_std_dev[1726]), .feature_accum(feature_accums[1726]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1727]), .RECT1_Y(rectangle1_ys[1727]), .RECT1_WIDTH(rectangle1_widths[1727]), .RECT1_HEIGHT(rectangle1_heights[1727]), .RECT1_WEIGHT(rectangle1_weights[1727]), .RECT2_X(rectangle2_xs[1727]), .RECT2_Y(rectangle2_ys[1727]), .RECT2_WIDTH(rectangle2_widths[1727]), .RECT2_HEIGHT(rectangle2_heights[1727]), .RECT2_WEIGHT(rectangle2_weights[1727]), .RECT3_X(rectangle3_xs[1727]), .RECT3_Y(rectangle3_ys[1727]), .RECT3_WIDTH(rectangle3_widths[1727]), .RECT3_HEIGHT(rectangle3_heights[1727]), .RECT3_WEIGHT(rectangle3_weights[1727]), .FEAT_THRES(feature_thresholds[1727]), .FEAT_ABOVE(feature_aboves[1727]), .FEAT_BELOW(feature_belows[1727])) ac1727(.scan_win(scan_win1727), .scan_win_std_dev(scan_win_std_dev[1727]), .feature_accum(feature_accums[1727]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1728]), .RECT1_Y(rectangle1_ys[1728]), .RECT1_WIDTH(rectangle1_widths[1728]), .RECT1_HEIGHT(rectangle1_heights[1728]), .RECT1_WEIGHT(rectangle1_weights[1728]), .RECT2_X(rectangle2_xs[1728]), .RECT2_Y(rectangle2_ys[1728]), .RECT2_WIDTH(rectangle2_widths[1728]), .RECT2_HEIGHT(rectangle2_heights[1728]), .RECT2_WEIGHT(rectangle2_weights[1728]), .RECT3_X(rectangle3_xs[1728]), .RECT3_Y(rectangle3_ys[1728]), .RECT3_WIDTH(rectangle3_widths[1728]), .RECT3_HEIGHT(rectangle3_heights[1728]), .RECT3_WEIGHT(rectangle3_weights[1728]), .FEAT_THRES(feature_thresholds[1728]), .FEAT_ABOVE(feature_aboves[1728]), .FEAT_BELOW(feature_belows[1728])) ac1728(.scan_win(scan_win1728), .scan_win_std_dev(scan_win_std_dev[1728]), .feature_accum(feature_accums[1728]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1729]), .RECT1_Y(rectangle1_ys[1729]), .RECT1_WIDTH(rectangle1_widths[1729]), .RECT1_HEIGHT(rectangle1_heights[1729]), .RECT1_WEIGHT(rectangle1_weights[1729]), .RECT2_X(rectangle2_xs[1729]), .RECT2_Y(rectangle2_ys[1729]), .RECT2_WIDTH(rectangle2_widths[1729]), .RECT2_HEIGHT(rectangle2_heights[1729]), .RECT2_WEIGHT(rectangle2_weights[1729]), .RECT3_X(rectangle3_xs[1729]), .RECT3_Y(rectangle3_ys[1729]), .RECT3_WIDTH(rectangle3_widths[1729]), .RECT3_HEIGHT(rectangle3_heights[1729]), .RECT3_WEIGHT(rectangle3_weights[1729]), .FEAT_THRES(feature_thresholds[1729]), .FEAT_ABOVE(feature_aboves[1729]), .FEAT_BELOW(feature_belows[1729])) ac1729(.scan_win(scan_win1729), .scan_win_std_dev(scan_win_std_dev[1729]), .feature_accum(feature_accums[1729]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1730]), .RECT1_Y(rectangle1_ys[1730]), .RECT1_WIDTH(rectangle1_widths[1730]), .RECT1_HEIGHT(rectangle1_heights[1730]), .RECT1_WEIGHT(rectangle1_weights[1730]), .RECT2_X(rectangle2_xs[1730]), .RECT2_Y(rectangle2_ys[1730]), .RECT2_WIDTH(rectangle2_widths[1730]), .RECT2_HEIGHT(rectangle2_heights[1730]), .RECT2_WEIGHT(rectangle2_weights[1730]), .RECT3_X(rectangle3_xs[1730]), .RECT3_Y(rectangle3_ys[1730]), .RECT3_WIDTH(rectangle3_widths[1730]), .RECT3_HEIGHT(rectangle3_heights[1730]), .RECT3_WEIGHT(rectangle3_weights[1730]), .FEAT_THRES(feature_thresholds[1730]), .FEAT_ABOVE(feature_aboves[1730]), .FEAT_BELOW(feature_belows[1730])) ac1730(.scan_win(scan_win1730), .scan_win_std_dev(scan_win_std_dev[1730]), .feature_accum(feature_accums[1730]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1731]), .RECT1_Y(rectangle1_ys[1731]), .RECT1_WIDTH(rectangle1_widths[1731]), .RECT1_HEIGHT(rectangle1_heights[1731]), .RECT1_WEIGHT(rectangle1_weights[1731]), .RECT2_X(rectangle2_xs[1731]), .RECT2_Y(rectangle2_ys[1731]), .RECT2_WIDTH(rectangle2_widths[1731]), .RECT2_HEIGHT(rectangle2_heights[1731]), .RECT2_WEIGHT(rectangle2_weights[1731]), .RECT3_X(rectangle3_xs[1731]), .RECT3_Y(rectangle3_ys[1731]), .RECT3_WIDTH(rectangle3_widths[1731]), .RECT3_HEIGHT(rectangle3_heights[1731]), .RECT3_WEIGHT(rectangle3_weights[1731]), .FEAT_THRES(feature_thresholds[1731]), .FEAT_ABOVE(feature_aboves[1731]), .FEAT_BELOW(feature_belows[1731])) ac1731(.scan_win(scan_win1731), .scan_win_std_dev(scan_win_std_dev[1731]), .feature_accum(feature_accums[1731]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1732]), .RECT1_Y(rectangle1_ys[1732]), .RECT1_WIDTH(rectangle1_widths[1732]), .RECT1_HEIGHT(rectangle1_heights[1732]), .RECT1_WEIGHT(rectangle1_weights[1732]), .RECT2_X(rectangle2_xs[1732]), .RECT2_Y(rectangle2_ys[1732]), .RECT2_WIDTH(rectangle2_widths[1732]), .RECT2_HEIGHT(rectangle2_heights[1732]), .RECT2_WEIGHT(rectangle2_weights[1732]), .RECT3_X(rectangle3_xs[1732]), .RECT3_Y(rectangle3_ys[1732]), .RECT3_WIDTH(rectangle3_widths[1732]), .RECT3_HEIGHT(rectangle3_heights[1732]), .RECT3_WEIGHT(rectangle3_weights[1732]), .FEAT_THRES(feature_thresholds[1732]), .FEAT_ABOVE(feature_aboves[1732]), .FEAT_BELOW(feature_belows[1732])) ac1732(.scan_win(scan_win1732), .scan_win_std_dev(scan_win_std_dev[1732]), .feature_accum(feature_accums[1732]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1733]), .RECT1_Y(rectangle1_ys[1733]), .RECT1_WIDTH(rectangle1_widths[1733]), .RECT1_HEIGHT(rectangle1_heights[1733]), .RECT1_WEIGHT(rectangle1_weights[1733]), .RECT2_X(rectangle2_xs[1733]), .RECT2_Y(rectangle2_ys[1733]), .RECT2_WIDTH(rectangle2_widths[1733]), .RECT2_HEIGHT(rectangle2_heights[1733]), .RECT2_WEIGHT(rectangle2_weights[1733]), .RECT3_X(rectangle3_xs[1733]), .RECT3_Y(rectangle3_ys[1733]), .RECT3_WIDTH(rectangle3_widths[1733]), .RECT3_HEIGHT(rectangle3_heights[1733]), .RECT3_WEIGHT(rectangle3_weights[1733]), .FEAT_THRES(feature_thresholds[1733]), .FEAT_ABOVE(feature_aboves[1733]), .FEAT_BELOW(feature_belows[1733])) ac1733(.scan_win(scan_win1733), .scan_win_std_dev(scan_win_std_dev[1733]), .feature_accum(feature_accums[1733]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1734]), .RECT1_Y(rectangle1_ys[1734]), .RECT1_WIDTH(rectangle1_widths[1734]), .RECT1_HEIGHT(rectangle1_heights[1734]), .RECT1_WEIGHT(rectangle1_weights[1734]), .RECT2_X(rectangle2_xs[1734]), .RECT2_Y(rectangle2_ys[1734]), .RECT2_WIDTH(rectangle2_widths[1734]), .RECT2_HEIGHT(rectangle2_heights[1734]), .RECT2_WEIGHT(rectangle2_weights[1734]), .RECT3_X(rectangle3_xs[1734]), .RECT3_Y(rectangle3_ys[1734]), .RECT3_WIDTH(rectangle3_widths[1734]), .RECT3_HEIGHT(rectangle3_heights[1734]), .RECT3_WEIGHT(rectangle3_weights[1734]), .FEAT_THRES(feature_thresholds[1734]), .FEAT_ABOVE(feature_aboves[1734]), .FEAT_BELOW(feature_belows[1734])) ac1734(.scan_win(scan_win1734), .scan_win_std_dev(scan_win_std_dev[1734]), .feature_accum(feature_accums[1734]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1735]), .RECT1_Y(rectangle1_ys[1735]), .RECT1_WIDTH(rectangle1_widths[1735]), .RECT1_HEIGHT(rectangle1_heights[1735]), .RECT1_WEIGHT(rectangle1_weights[1735]), .RECT2_X(rectangle2_xs[1735]), .RECT2_Y(rectangle2_ys[1735]), .RECT2_WIDTH(rectangle2_widths[1735]), .RECT2_HEIGHT(rectangle2_heights[1735]), .RECT2_WEIGHT(rectangle2_weights[1735]), .RECT3_X(rectangle3_xs[1735]), .RECT3_Y(rectangle3_ys[1735]), .RECT3_WIDTH(rectangle3_widths[1735]), .RECT3_HEIGHT(rectangle3_heights[1735]), .RECT3_WEIGHT(rectangle3_weights[1735]), .FEAT_THRES(feature_thresholds[1735]), .FEAT_ABOVE(feature_aboves[1735]), .FEAT_BELOW(feature_belows[1735])) ac1735(.scan_win(scan_win1735), .scan_win_std_dev(scan_win_std_dev[1735]), .feature_accum(feature_accums[1735]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1736]), .RECT1_Y(rectangle1_ys[1736]), .RECT1_WIDTH(rectangle1_widths[1736]), .RECT1_HEIGHT(rectangle1_heights[1736]), .RECT1_WEIGHT(rectangle1_weights[1736]), .RECT2_X(rectangle2_xs[1736]), .RECT2_Y(rectangle2_ys[1736]), .RECT2_WIDTH(rectangle2_widths[1736]), .RECT2_HEIGHT(rectangle2_heights[1736]), .RECT2_WEIGHT(rectangle2_weights[1736]), .RECT3_X(rectangle3_xs[1736]), .RECT3_Y(rectangle3_ys[1736]), .RECT3_WIDTH(rectangle3_widths[1736]), .RECT3_HEIGHT(rectangle3_heights[1736]), .RECT3_WEIGHT(rectangle3_weights[1736]), .FEAT_THRES(feature_thresholds[1736]), .FEAT_ABOVE(feature_aboves[1736]), .FEAT_BELOW(feature_belows[1736])) ac1736(.scan_win(scan_win1736), .scan_win_std_dev(scan_win_std_dev[1736]), .feature_accum(feature_accums[1736]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1737]), .RECT1_Y(rectangle1_ys[1737]), .RECT1_WIDTH(rectangle1_widths[1737]), .RECT1_HEIGHT(rectangle1_heights[1737]), .RECT1_WEIGHT(rectangle1_weights[1737]), .RECT2_X(rectangle2_xs[1737]), .RECT2_Y(rectangle2_ys[1737]), .RECT2_WIDTH(rectangle2_widths[1737]), .RECT2_HEIGHT(rectangle2_heights[1737]), .RECT2_WEIGHT(rectangle2_weights[1737]), .RECT3_X(rectangle3_xs[1737]), .RECT3_Y(rectangle3_ys[1737]), .RECT3_WIDTH(rectangle3_widths[1737]), .RECT3_HEIGHT(rectangle3_heights[1737]), .RECT3_WEIGHT(rectangle3_weights[1737]), .FEAT_THRES(feature_thresholds[1737]), .FEAT_ABOVE(feature_aboves[1737]), .FEAT_BELOW(feature_belows[1737])) ac1737(.scan_win(scan_win1737), .scan_win_std_dev(scan_win_std_dev[1737]), .feature_accum(feature_accums[1737]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1738]), .RECT1_Y(rectangle1_ys[1738]), .RECT1_WIDTH(rectangle1_widths[1738]), .RECT1_HEIGHT(rectangle1_heights[1738]), .RECT1_WEIGHT(rectangle1_weights[1738]), .RECT2_X(rectangle2_xs[1738]), .RECT2_Y(rectangle2_ys[1738]), .RECT2_WIDTH(rectangle2_widths[1738]), .RECT2_HEIGHT(rectangle2_heights[1738]), .RECT2_WEIGHT(rectangle2_weights[1738]), .RECT3_X(rectangle3_xs[1738]), .RECT3_Y(rectangle3_ys[1738]), .RECT3_WIDTH(rectangle3_widths[1738]), .RECT3_HEIGHT(rectangle3_heights[1738]), .RECT3_WEIGHT(rectangle3_weights[1738]), .FEAT_THRES(feature_thresholds[1738]), .FEAT_ABOVE(feature_aboves[1738]), .FEAT_BELOW(feature_belows[1738])) ac1738(.scan_win(scan_win1738), .scan_win_std_dev(scan_win_std_dev[1738]), .feature_accum(feature_accums[1738]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1739]), .RECT1_Y(rectangle1_ys[1739]), .RECT1_WIDTH(rectangle1_widths[1739]), .RECT1_HEIGHT(rectangle1_heights[1739]), .RECT1_WEIGHT(rectangle1_weights[1739]), .RECT2_X(rectangle2_xs[1739]), .RECT2_Y(rectangle2_ys[1739]), .RECT2_WIDTH(rectangle2_widths[1739]), .RECT2_HEIGHT(rectangle2_heights[1739]), .RECT2_WEIGHT(rectangle2_weights[1739]), .RECT3_X(rectangle3_xs[1739]), .RECT3_Y(rectangle3_ys[1739]), .RECT3_WIDTH(rectangle3_widths[1739]), .RECT3_HEIGHT(rectangle3_heights[1739]), .RECT3_WEIGHT(rectangle3_weights[1739]), .FEAT_THRES(feature_thresholds[1739]), .FEAT_ABOVE(feature_aboves[1739]), .FEAT_BELOW(feature_belows[1739])) ac1739(.scan_win(scan_win1739), .scan_win_std_dev(scan_win_std_dev[1739]), .feature_accum(feature_accums[1739]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1740]), .RECT1_Y(rectangle1_ys[1740]), .RECT1_WIDTH(rectangle1_widths[1740]), .RECT1_HEIGHT(rectangle1_heights[1740]), .RECT1_WEIGHT(rectangle1_weights[1740]), .RECT2_X(rectangle2_xs[1740]), .RECT2_Y(rectangle2_ys[1740]), .RECT2_WIDTH(rectangle2_widths[1740]), .RECT2_HEIGHT(rectangle2_heights[1740]), .RECT2_WEIGHT(rectangle2_weights[1740]), .RECT3_X(rectangle3_xs[1740]), .RECT3_Y(rectangle3_ys[1740]), .RECT3_WIDTH(rectangle3_widths[1740]), .RECT3_HEIGHT(rectangle3_heights[1740]), .RECT3_WEIGHT(rectangle3_weights[1740]), .FEAT_THRES(feature_thresholds[1740]), .FEAT_ABOVE(feature_aboves[1740]), .FEAT_BELOW(feature_belows[1740])) ac1740(.scan_win(scan_win1740), .scan_win_std_dev(scan_win_std_dev[1740]), .feature_accum(feature_accums[1740]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1741]), .RECT1_Y(rectangle1_ys[1741]), .RECT1_WIDTH(rectangle1_widths[1741]), .RECT1_HEIGHT(rectangle1_heights[1741]), .RECT1_WEIGHT(rectangle1_weights[1741]), .RECT2_X(rectangle2_xs[1741]), .RECT2_Y(rectangle2_ys[1741]), .RECT2_WIDTH(rectangle2_widths[1741]), .RECT2_HEIGHT(rectangle2_heights[1741]), .RECT2_WEIGHT(rectangle2_weights[1741]), .RECT3_X(rectangle3_xs[1741]), .RECT3_Y(rectangle3_ys[1741]), .RECT3_WIDTH(rectangle3_widths[1741]), .RECT3_HEIGHT(rectangle3_heights[1741]), .RECT3_WEIGHT(rectangle3_weights[1741]), .FEAT_THRES(feature_thresholds[1741]), .FEAT_ABOVE(feature_aboves[1741]), .FEAT_BELOW(feature_belows[1741])) ac1741(.scan_win(scan_win1741), .scan_win_std_dev(scan_win_std_dev[1741]), .feature_accum(feature_accums[1741]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1742]), .RECT1_Y(rectangle1_ys[1742]), .RECT1_WIDTH(rectangle1_widths[1742]), .RECT1_HEIGHT(rectangle1_heights[1742]), .RECT1_WEIGHT(rectangle1_weights[1742]), .RECT2_X(rectangle2_xs[1742]), .RECT2_Y(rectangle2_ys[1742]), .RECT2_WIDTH(rectangle2_widths[1742]), .RECT2_HEIGHT(rectangle2_heights[1742]), .RECT2_WEIGHT(rectangle2_weights[1742]), .RECT3_X(rectangle3_xs[1742]), .RECT3_Y(rectangle3_ys[1742]), .RECT3_WIDTH(rectangle3_widths[1742]), .RECT3_HEIGHT(rectangle3_heights[1742]), .RECT3_WEIGHT(rectangle3_weights[1742]), .FEAT_THRES(feature_thresholds[1742]), .FEAT_ABOVE(feature_aboves[1742]), .FEAT_BELOW(feature_belows[1742])) ac1742(.scan_win(scan_win1742), .scan_win_std_dev(scan_win_std_dev[1742]), .feature_accum(feature_accums[1742]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1743]), .RECT1_Y(rectangle1_ys[1743]), .RECT1_WIDTH(rectangle1_widths[1743]), .RECT1_HEIGHT(rectangle1_heights[1743]), .RECT1_WEIGHT(rectangle1_weights[1743]), .RECT2_X(rectangle2_xs[1743]), .RECT2_Y(rectangle2_ys[1743]), .RECT2_WIDTH(rectangle2_widths[1743]), .RECT2_HEIGHT(rectangle2_heights[1743]), .RECT2_WEIGHT(rectangle2_weights[1743]), .RECT3_X(rectangle3_xs[1743]), .RECT3_Y(rectangle3_ys[1743]), .RECT3_WIDTH(rectangle3_widths[1743]), .RECT3_HEIGHT(rectangle3_heights[1743]), .RECT3_WEIGHT(rectangle3_weights[1743]), .FEAT_THRES(feature_thresholds[1743]), .FEAT_ABOVE(feature_aboves[1743]), .FEAT_BELOW(feature_belows[1743])) ac1743(.scan_win(scan_win1743), .scan_win_std_dev(scan_win_std_dev[1743]), .feature_accum(feature_accums[1743]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1744]), .RECT1_Y(rectangle1_ys[1744]), .RECT1_WIDTH(rectangle1_widths[1744]), .RECT1_HEIGHT(rectangle1_heights[1744]), .RECT1_WEIGHT(rectangle1_weights[1744]), .RECT2_X(rectangle2_xs[1744]), .RECT2_Y(rectangle2_ys[1744]), .RECT2_WIDTH(rectangle2_widths[1744]), .RECT2_HEIGHT(rectangle2_heights[1744]), .RECT2_WEIGHT(rectangle2_weights[1744]), .RECT3_X(rectangle3_xs[1744]), .RECT3_Y(rectangle3_ys[1744]), .RECT3_WIDTH(rectangle3_widths[1744]), .RECT3_HEIGHT(rectangle3_heights[1744]), .RECT3_WEIGHT(rectangle3_weights[1744]), .FEAT_THRES(feature_thresholds[1744]), .FEAT_ABOVE(feature_aboves[1744]), .FEAT_BELOW(feature_belows[1744])) ac1744(.scan_win(scan_win1744), .scan_win_std_dev(scan_win_std_dev[1744]), .feature_accum(feature_accums[1744]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1745]), .RECT1_Y(rectangle1_ys[1745]), .RECT1_WIDTH(rectangle1_widths[1745]), .RECT1_HEIGHT(rectangle1_heights[1745]), .RECT1_WEIGHT(rectangle1_weights[1745]), .RECT2_X(rectangle2_xs[1745]), .RECT2_Y(rectangle2_ys[1745]), .RECT2_WIDTH(rectangle2_widths[1745]), .RECT2_HEIGHT(rectangle2_heights[1745]), .RECT2_WEIGHT(rectangle2_weights[1745]), .RECT3_X(rectangle3_xs[1745]), .RECT3_Y(rectangle3_ys[1745]), .RECT3_WIDTH(rectangle3_widths[1745]), .RECT3_HEIGHT(rectangle3_heights[1745]), .RECT3_WEIGHT(rectangle3_weights[1745]), .FEAT_THRES(feature_thresholds[1745]), .FEAT_ABOVE(feature_aboves[1745]), .FEAT_BELOW(feature_belows[1745])) ac1745(.scan_win(scan_win1745), .scan_win_std_dev(scan_win_std_dev[1745]), .feature_accum(feature_accums[1745]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1746]), .RECT1_Y(rectangle1_ys[1746]), .RECT1_WIDTH(rectangle1_widths[1746]), .RECT1_HEIGHT(rectangle1_heights[1746]), .RECT1_WEIGHT(rectangle1_weights[1746]), .RECT2_X(rectangle2_xs[1746]), .RECT2_Y(rectangle2_ys[1746]), .RECT2_WIDTH(rectangle2_widths[1746]), .RECT2_HEIGHT(rectangle2_heights[1746]), .RECT2_WEIGHT(rectangle2_weights[1746]), .RECT3_X(rectangle3_xs[1746]), .RECT3_Y(rectangle3_ys[1746]), .RECT3_WIDTH(rectangle3_widths[1746]), .RECT3_HEIGHT(rectangle3_heights[1746]), .RECT3_WEIGHT(rectangle3_weights[1746]), .FEAT_THRES(feature_thresholds[1746]), .FEAT_ABOVE(feature_aboves[1746]), .FEAT_BELOW(feature_belows[1746])) ac1746(.scan_win(scan_win1746), .scan_win_std_dev(scan_win_std_dev[1746]), .feature_accum(feature_accums[1746]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1747]), .RECT1_Y(rectangle1_ys[1747]), .RECT1_WIDTH(rectangle1_widths[1747]), .RECT1_HEIGHT(rectangle1_heights[1747]), .RECT1_WEIGHT(rectangle1_weights[1747]), .RECT2_X(rectangle2_xs[1747]), .RECT2_Y(rectangle2_ys[1747]), .RECT2_WIDTH(rectangle2_widths[1747]), .RECT2_HEIGHT(rectangle2_heights[1747]), .RECT2_WEIGHT(rectangle2_weights[1747]), .RECT3_X(rectangle3_xs[1747]), .RECT3_Y(rectangle3_ys[1747]), .RECT3_WIDTH(rectangle3_widths[1747]), .RECT3_HEIGHT(rectangle3_heights[1747]), .RECT3_WEIGHT(rectangle3_weights[1747]), .FEAT_THRES(feature_thresholds[1747]), .FEAT_ABOVE(feature_aboves[1747]), .FEAT_BELOW(feature_belows[1747])) ac1747(.scan_win(scan_win1747), .scan_win_std_dev(scan_win_std_dev[1747]), .feature_accum(feature_accums[1747]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1748]), .RECT1_Y(rectangle1_ys[1748]), .RECT1_WIDTH(rectangle1_widths[1748]), .RECT1_HEIGHT(rectangle1_heights[1748]), .RECT1_WEIGHT(rectangle1_weights[1748]), .RECT2_X(rectangle2_xs[1748]), .RECT2_Y(rectangle2_ys[1748]), .RECT2_WIDTH(rectangle2_widths[1748]), .RECT2_HEIGHT(rectangle2_heights[1748]), .RECT2_WEIGHT(rectangle2_weights[1748]), .RECT3_X(rectangle3_xs[1748]), .RECT3_Y(rectangle3_ys[1748]), .RECT3_WIDTH(rectangle3_widths[1748]), .RECT3_HEIGHT(rectangle3_heights[1748]), .RECT3_WEIGHT(rectangle3_weights[1748]), .FEAT_THRES(feature_thresholds[1748]), .FEAT_ABOVE(feature_aboves[1748]), .FEAT_BELOW(feature_belows[1748])) ac1748(.scan_win(scan_win1748), .scan_win_std_dev(scan_win_std_dev[1748]), .feature_accum(feature_accums[1748]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1749]), .RECT1_Y(rectangle1_ys[1749]), .RECT1_WIDTH(rectangle1_widths[1749]), .RECT1_HEIGHT(rectangle1_heights[1749]), .RECT1_WEIGHT(rectangle1_weights[1749]), .RECT2_X(rectangle2_xs[1749]), .RECT2_Y(rectangle2_ys[1749]), .RECT2_WIDTH(rectangle2_widths[1749]), .RECT2_HEIGHT(rectangle2_heights[1749]), .RECT2_WEIGHT(rectangle2_weights[1749]), .RECT3_X(rectangle3_xs[1749]), .RECT3_Y(rectangle3_ys[1749]), .RECT3_WIDTH(rectangle3_widths[1749]), .RECT3_HEIGHT(rectangle3_heights[1749]), .RECT3_WEIGHT(rectangle3_weights[1749]), .FEAT_THRES(feature_thresholds[1749]), .FEAT_ABOVE(feature_aboves[1749]), .FEAT_BELOW(feature_belows[1749])) ac1749(.scan_win(scan_win1749), .scan_win_std_dev(scan_win_std_dev[1749]), .feature_accum(feature_accums[1749]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1750]), .RECT1_Y(rectangle1_ys[1750]), .RECT1_WIDTH(rectangle1_widths[1750]), .RECT1_HEIGHT(rectangle1_heights[1750]), .RECT1_WEIGHT(rectangle1_weights[1750]), .RECT2_X(rectangle2_xs[1750]), .RECT2_Y(rectangle2_ys[1750]), .RECT2_WIDTH(rectangle2_widths[1750]), .RECT2_HEIGHT(rectangle2_heights[1750]), .RECT2_WEIGHT(rectangle2_weights[1750]), .RECT3_X(rectangle3_xs[1750]), .RECT3_Y(rectangle3_ys[1750]), .RECT3_WIDTH(rectangle3_widths[1750]), .RECT3_HEIGHT(rectangle3_heights[1750]), .RECT3_WEIGHT(rectangle3_weights[1750]), .FEAT_THRES(feature_thresholds[1750]), .FEAT_ABOVE(feature_aboves[1750]), .FEAT_BELOW(feature_belows[1750])) ac1750(.scan_win(scan_win1750), .scan_win_std_dev(scan_win_std_dev[1750]), .feature_accum(feature_accums[1750]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1751]), .RECT1_Y(rectangle1_ys[1751]), .RECT1_WIDTH(rectangle1_widths[1751]), .RECT1_HEIGHT(rectangle1_heights[1751]), .RECT1_WEIGHT(rectangle1_weights[1751]), .RECT2_X(rectangle2_xs[1751]), .RECT2_Y(rectangle2_ys[1751]), .RECT2_WIDTH(rectangle2_widths[1751]), .RECT2_HEIGHT(rectangle2_heights[1751]), .RECT2_WEIGHT(rectangle2_weights[1751]), .RECT3_X(rectangle3_xs[1751]), .RECT3_Y(rectangle3_ys[1751]), .RECT3_WIDTH(rectangle3_widths[1751]), .RECT3_HEIGHT(rectangle3_heights[1751]), .RECT3_WEIGHT(rectangle3_weights[1751]), .FEAT_THRES(feature_thresholds[1751]), .FEAT_ABOVE(feature_aboves[1751]), .FEAT_BELOW(feature_belows[1751])) ac1751(.scan_win(scan_win1751), .scan_win_std_dev(scan_win_std_dev[1751]), .feature_accum(feature_accums[1751]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1752]), .RECT1_Y(rectangle1_ys[1752]), .RECT1_WIDTH(rectangle1_widths[1752]), .RECT1_HEIGHT(rectangle1_heights[1752]), .RECT1_WEIGHT(rectangle1_weights[1752]), .RECT2_X(rectangle2_xs[1752]), .RECT2_Y(rectangle2_ys[1752]), .RECT2_WIDTH(rectangle2_widths[1752]), .RECT2_HEIGHT(rectangle2_heights[1752]), .RECT2_WEIGHT(rectangle2_weights[1752]), .RECT3_X(rectangle3_xs[1752]), .RECT3_Y(rectangle3_ys[1752]), .RECT3_WIDTH(rectangle3_widths[1752]), .RECT3_HEIGHT(rectangle3_heights[1752]), .RECT3_WEIGHT(rectangle3_weights[1752]), .FEAT_THRES(feature_thresholds[1752]), .FEAT_ABOVE(feature_aboves[1752]), .FEAT_BELOW(feature_belows[1752])) ac1752(.scan_win(scan_win1752), .scan_win_std_dev(scan_win_std_dev[1752]), .feature_accum(feature_accums[1752]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1753]), .RECT1_Y(rectangle1_ys[1753]), .RECT1_WIDTH(rectangle1_widths[1753]), .RECT1_HEIGHT(rectangle1_heights[1753]), .RECT1_WEIGHT(rectangle1_weights[1753]), .RECT2_X(rectangle2_xs[1753]), .RECT2_Y(rectangle2_ys[1753]), .RECT2_WIDTH(rectangle2_widths[1753]), .RECT2_HEIGHT(rectangle2_heights[1753]), .RECT2_WEIGHT(rectangle2_weights[1753]), .RECT3_X(rectangle3_xs[1753]), .RECT3_Y(rectangle3_ys[1753]), .RECT3_WIDTH(rectangle3_widths[1753]), .RECT3_HEIGHT(rectangle3_heights[1753]), .RECT3_WEIGHT(rectangle3_weights[1753]), .FEAT_THRES(feature_thresholds[1753]), .FEAT_ABOVE(feature_aboves[1753]), .FEAT_BELOW(feature_belows[1753])) ac1753(.scan_win(scan_win1753), .scan_win_std_dev(scan_win_std_dev[1753]), .feature_accum(feature_accums[1753]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1754]), .RECT1_Y(rectangle1_ys[1754]), .RECT1_WIDTH(rectangle1_widths[1754]), .RECT1_HEIGHT(rectangle1_heights[1754]), .RECT1_WEIGHT(rectangle1_weights[1754]), .RECT2_X(rectangle2_xs[1754]), .RECT2_Y(rectangle2_ys[1754]), .RECT2_WIDTH(rectangle2_widths[1754]), .RECT2_HEIGHT(rectangle2_heights[1754]), .RECT2_WEIGHT(rectangle2_weights[1754]), .RECT3_X(rectangle3_xs[1754]), .RECT3_Y(rectangle3_ys[1754]), .RECT3_WIDTH(rectangle3_widths[1754]), .RECT3_HEIGHT(rectangle3_heights[1754]), .RECT3_WEIGHT(rectangle3_weights[1754]), .FEAT_THRES(feature_thresholds[1754]), .FEAT_ABOVE(feature_aboves[1754]), .FEAT_BELOW(feature_belows[1754])) ac1754(.scan_win(scan_win1754), .scan_win_std_dev(scan_win_std_dev[1754]), .feature_accum(feature_accums[1754]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1755]), .RECT1_Y(rectangle1_ys[1755]), .RECT1_WIDTH(rectangle1_widths[1755]), .RECT1_HEIGHT(rectangle1_heights[1755]), .RECT1_WEIGHT(rectangle1_weights[1755]), .RECT2_X(rectangle2_xs[1755]), .RECT2_Y(rectangle2_ys[1755]), .RECT2_WIDTH(rectangle2_widths[1755]), .RECT2_HEIGHT(rectangle2_heights[1755]), .RECT2_WEIGHT(rectangle2_weights[1755]), .RECT3_X(rectangle3_xs[1755]), .RECT3_Y(rectangle3_ys[1755]), .RECT3_WIDTH(rectangle3_widths[1755]), .RECT3_HEIGHT(rectangle3_heights[1755]), .RECT3_WEIGHT(rectangle3_weights[1755]), .FEAT_THRES(feature_thresholds[1755]), .FEAT_ABOVE(feature_aboves[1755]), .FEAT_BELOW(feature_belows[1755])) ac1755(.scan_win(scan_win1755), .scan_win_std_dev(scan_win_std_dev[1755]), .feature_accum(feature_accums[1755]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1756]), .RECT1_Y(rectangle1_ys[1756]), .RECT1_WIDTH(rectangle1_widths[1756]), .RECT1_HEIGHT(rectangle1_heights[1756]), .RECT1_WEIGHT(rectangle1_weights[1756]), .RECT2_X(rectangle2_xs[1756]), .RECT2_Y(rectangle2_ys[1756]), .RECT2_WIDTH(rectangle2_widths[1756]), .RECT2_HEIGHT(rectangle2_heights[1756]), .RECT2_WEIGHT(rectangle2_weights[1756]), .RECT3_X(rectangle3_xs[1756]), .RECT3_Y(rectangle3_ys[1756]), .RECT3_WIDTH(rectangle3_widths[1756]), .RECT3_HEIGHT(rectangle3_heights[1756]), .RECT3_WEIGHT(rectangle3_weights[1756]), .FEAT_THRES(feature_thresholds[1756]), .FEAT_ABOVE(feature_aboves[1756]), .FEAT_BELOW(feature_belows[1756])) ac1756(.scan_win(scan_win1756), .scan_win_std_dev(scan_win_std_dev[1756]), .feature_accum(feature_accums[1756]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1757]), .RECT1_Y(rectangle1_ys[1757]), .RECT1_WIDTH(rectangle1_widths[1757]), .RECT1_HEIGHT(rectangle1_heights[1757]), .RECT1_WEIGHT(rectangle1_weights[1757]), .RECT2_X(rectangle2_xs[1757]), .RECT2_Y(rectangle2_ys[1757]), .RECT2_WIDTH(rectangle2_widths[1757]), .RECT2_HEIGHT(rectangle2_heights[1757]), .RECT2_WEIGHT(rectangle2_weights[1757]), .RECT3_X(rectangle3_xs[1757]), .RECT3_Y(rectangle3_ys[1757]), .RECT3_WIDTH(rectangle3_widths[1757]), .RECT3_HEIGHT(rectangle3_heights[1757]), .RECT3_WEIGHT(rectangle3_weights[1757]), .FEAT_THRES(feature_thresholds[1757]), .FEAT_ABOVE(feature_aboves[1757]), .FEAT_BELOW(feature_belows[1757])) ac1757(.scan_win(scan_win1757), .scan_win_std_dev(scan_win_std_dev[1757]), .feature_accum(feature_accums[1757]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1758]), .RECT1_Y(rectangle1_ys[1758]), .RECT1_WIDTH(rectangle1_widths[1758]), .RECT1_HEIGHT(rectangle1_heights[1758]), .RECT1_WEIGHT(rectangle1_weights[1758]), .RECT2_X(rectangle2_xs[1758]), .RECT2_Y(rectangle2_ys[1758]), .RECT2_WIDTH(rectangle2_widths[1758]), .RECT2_HEIGHT(rectangle2_heights[1758]), .RECT2_WEIGHT(rectangle2_weights[1758]), .RECT3_X(rectangle3_xs[1758]), .RECT3_Y(rectangle3_ys[1758]), .RECT3_WIDTH(rectangle3_widths[1758]), .RECT3_HEIGHT(rectangle3_heights[1758]), .RECT3_WEIGHT(rectangle3_weights[1758]), .FEAT_THRES(feature_thresholds[1758]), .FEAT_ABOVE(feature_aboves[1758]), .FEAT_BELOW(feature_belows[1758])) ac1758(.scan_win(scan_win1758), .scan_win_std_dev(scan_win_std_dev[1758]), .feature_accum(feature_accums[1758]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1759]), .RECT1_Y(rectangle1_ys[1759]), .RECT1_WIDTH(rectangle1_widths[1759]), .RECT1_HEIGHT(rectangle1_heights[1759]), .RECT1_WEIGHT(rectangle1_weights[1759]), .RECT2_X(rectangle2_xs[1759]), .RECT2_Y(rectangle2_ys[1759]), .RECT2_WIDTH(rectangle2_widths[1759]), .RECT2_HEIGHT(rectangle2_heights[1759]), .RECT2_WEIGHT(rectangle2_weights[1759]), .RECT3_X(rectangle3_xs[1759]), .RECT3_Y(rectangle3_ys[1759]), .RECT3_WIDTH(rectangle3_widths[1759]), .RECT3_HEIGHT(rectangle3_heights[1759]), .RECT3_WEIGHT(rectangle3_weights[1759]), .FEAT_THRES(feature_thresholds[1759]), .FEAT_ABOVE(feature_aboves[1759]), .FEAT_BELOW(feature_belows[1759])) ac1759(.scan_win(scan_win1759), .scan_win_std_dev(scan_win_std_dev[1759]), .feature_accum(feature_accums[1759]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1760]), .RECT1_Y(rectangle1_ys[1760]), .RECT1_WIDTH(rectangle1_widths[1760]), .RECT1_HEIGHT(rectangle1_heights[1760]), .RECT1_WEIGHT(rectangle1_weights[1760]), .RECT2_X(rectangle2_xs[1760]), .RECT2_Y(rectangle2_ys[1760]), .RECT2_WIDTH(rectangle2_widths[1760]), .RECT2_HEIGHT(rectangle2_heights[1760]), .RECT2_WEIGHT(rectangle2_weights[1760]), .RECT3_X(rectangle3_xs[1760]), .RECT3_Y(rectangle3_ys[1760]), .RECT3_WIDTH(rectangle3_widths[1760]), .RECT3_HEIGHT(rectangle3_heights[1760]), .RECT3_WEIGHT(rectangle3_weights[1760]), .FEAT_THRES(feature_thresholds[1760]), .FEAT_ABOVE(feature_aboves[1760]), .FEAT_BELOW(feature_belows[1760])) ac1760(.scan_win(scan_win1760), .scan_win_std_dev(scan_win_std_dev[1760]), .feature_accum(feature_accums[1760]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1761]), .RECT1_Y(rectangle1_ys[1761]), .RECT1_WIDTH(rectangle1_widths[1761]), .RECT1_HEIGHT(rectangle1_heights[1761]), .RECT1_WEIGHT(rectangle1_weights[1761]), .RECT2_X(rectangle2_xs[1761]), .RECT2_Y(rectangle2_ys[1761]), .RECT2_WIDTH(rectangle2_widths[1761]), .RECT2_HEIGHT(rectangle2_heights[1761]), .RECT2_WEIGHT(rectangle2_weights[1761]), .RECT3_X(rectangle3_xs[1761]), .RECT3_Y(rectangle3_ys[1761]), .RECT3_WIDTH(rectangle3_widths[1761]), .RECT3_HEIGHT(rectangle3_heights[1761]), .RECT3_WEIGHT(rectangle3_weights[1761]), .FEAT_THRES(feature_thresholds[1761]), .FEAT_ABOVE(feature_aboves[1761]), .FEAT_BELOW(feature_belows[1761])) ac1761(.scan_win(scan_win1761), .scan_win_std_dev(scan_win_std_dev[1761]), .feature_accum(feature_accums[1761]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1762]), .RECT1_Y(rectangle1_ys[1762]), .RECT1_WIDTH(rectangle1_widths[1762]), .RECT1_HEIGHT(rectangle1_heights[1762]), .RECT1_WEIGHT(rectangle1_weights[1762]), .RECT2_X(rectangle2_xs[1762]), .RECT2_Y(rectangle2_ys[1762]), .RECT2_WIDTH(rectangle2_widths[1762]), .RECT2_HEIGHT(rectangle2_heights[1762]), .RECT2_WEIGHT(rectangle2_weights[1762]), .RECT3_X(rectangle3_xs[1762]), .RECT3_Y(rectangle3_ys[1762]), .RECT3_WIDTH(rectangle3_widths[1762]), .RECT3_HEIGHT(rectangle3_heights[1762]), .RECT3_WEIGHT(rectangle3_weights[1762]), .FEAT_THRES(feature_thresholds[1762]), .FEAT_ABOVE(feature_aboves[1762]), .FEAT_BELOW(feature_belows[1762])) ac1762(.scan_win(scan_win1762), .scan_win_std_dev(scan_win_std_dev[1762]), .feature_accum(feature_accums[1762]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1763]), .RECT1_Y(rectangle1_ys[1763]), .RECT1_WIDTH(rectangle1_widths[1763]), .RECT1_HEIGHT(rectangle1_heights[1763]), .RECT1_WEIGHT(rectangle1_weights[1763]), .RECT2_X(rectangle2_xs[1763]), .RECT2_Y(rectangle2_ys[1763]), .RECT2_WIDTH(rectangle2_widths[1763]), .RECT2_HEIGHT(rectangle2_heights[1763]), .RECT2_WEIGHT(rectangle2_weights[1763]), .RECT3_X(rectangle3_xs[1763]), .RECT3_Y(rectangle3_ys[1763]), .RECT3_WIDTH(rectangle3_widths[1763]), .RECT3_HEIGHT(rectangle3_heights[1763]), .RECT3_WEIGHT(rectangle3_weights[1763]), .FEAT_THRES(feature_thresholds[1763]), .FEAT_ABOVE(feature_aboves[1763]), .FEAT_BELOW(feature_belows[1763])) ac1763(.scan_win(scan_win1763), .scan_win_std_dev(scan_win_std_dev[1763]), .feature_accum(feature_accums[1763]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1764]), .RECT1_Y(rectangle1_ys[1764]), .RECT1_WIDTH(rectangle1_widths[1764]), .RECT1_HEIGHT(rectangle1_heights[1764]), .RECT1_WEIGHT(rectangle1_weights[1764]), .RECT2_X(rectangle2_xs[1764]), .RECT2_Y(rectangle2_ys[1764]), .RECT2_WIDTH(rectangle2_widths[1764]), .RECT2_HEIGHT(rectangle2_heights[1764]), .RECT2_WEIGHT(rectangle2_weights[1764]), .RECT3_X(rectangle3_xs[1764]), .RECT3_Y(rectangle3_ys[1764]), .RECT3_WIDTH(rectangle3_widths[1764]), .RECT3_HEIGHT(rectangle3_heights[1764]), .RECT3_WEIGHT(rectangle3_weights[1764]), .FEAT_THRES(feature_thresholds[1764]), .FEAT_ABOVE(feature_aboves[1764]), .FEAT_BELOW(feature_belows[1764])) ac1764(.scan_win(scan_win1764), .scan_win_std_dev(scan_win_std_dev[1764]), .feature_accum(feature_accums[1764]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1765]), .RECT1_Y(rectangle1_ys[1765]), .RECT1_WIDTH(rectangle1_widths[1765]), .RECT1_HEIGHT(rectangle1_heights[1765]), .RECT1_WEIGHT(rectangle1_weights[1765]), .RECT2_X(rectangle2_xs[1765]), .RECT2_Y(rectangle2_ys[1765]), .RECT2_WIDTH(rectangle2_widths[1765]), .RECT2_HEIGHT(rectangle2_heights[1765]), .RECT2_WEIGHT(rectangle2_weights[1765]), .RECT3_X(rectangle3_xs[1765]), .RECT3_Y(rectangle3_ys[1765]), .RECT3_WIDTH(rectangle3_widths[1765]), .RECT3_HEIGHT(rectangle3_heights[1765]), .RECT3_WEIGHT(rectangle3_weights[1765]), .FEAT_THRES(feature_thresholds[1765]), .FEAT_ABOVE(feature_aboves[1765]), .FEAT_BELOW(feature_belows[1765])) ac1765(.scan_win(scan_win1765), .scan_win_std_dev(scan_win_std_dev[1765]), .feature_accum(feature_accums[1765]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1766]), .RECT1_Y(rectangle1_ys[1766]), .RECT1_WIDTH(rectangle1_widths[1766]), .RECT1_HEIGHT(rectangle1_heights[1766]), .RECT1_WEIGHT(rectangle1_weights[1766]), .RECT2_X(rectangle2_xs[1766]), .RECT2_Y(rectangle2_ys[1766]), .RECT2_WIDTH(rectangle2_widths[1766]), .RECT2_HEIGHT(rectangle2_heights[1766]), .RECT2_WEIGHT(rectangle2_weights[1766]), .RECT3_X(rectangle3_xs[1766]), .RECT3_Y(rectangle3_ys[1766]), .RECT3_WIDTH(rectangle3_widths[1766]), .RECT3_HEIGHT(rectangle3_heights[1766]), .RECT3_WEIGHT(rectangle3_weights[1766]), .FEAT_THRES(feature_thresholds[1766]), .FEAT_ABOVE(feature_aboves[1766]), .FEAT_BELOW(feature_belows[1766])) ac1766(.scan_win(scan_win1766), .scan_win_std_dev(scan_win_std_dev[1766]), .feature_accum(feature_accums[1766]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1767]), .RECT1_Y(rectangle1_ys[1767]), .RECT1_WIDTH(rectangle1_widths[1767]), .RECT1_HEIGHT(rectangle1_heights[1767]), .RECT1_WEIGHT(rectangle1_weights[1767]), .RECT2_X(rectangle2_xs[1767]), .RECT2_Y(rectangle2_ys[1767]), .RECT2_WIDTH(rectangle2_widths[1767]), .RECT2_HEIGHT(rectangle2_heights[1767]), .RECT2_WEIGHT(rectangle2_weights[1767]), .RECT3_X(rectangle3_xs[1767]), .RECT3_Y(rectangle3_ys[1767]), .RECT3_WIDTH(rectangle3_widths[1767]), .RECT3_HEIGHT(rectangle3_heights[1767]), .RECT3_WEIGHT(rectangle3_weights[1767]), .FEAT_THRES(feature_thresholds[1767]), .FEAT_ABOVE(feature_aboves[1767]), .FEAT_BELOW(feature_belows[1767])) ac1767(.scan_win(scan_win1767), .scan_win_std_dev(scan_win_std_dev[1767]), .feature_accum(feature_accums[1767]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1768]), .RECT1_Y(rectangle1_ys[1768]), .RECT1_WIDTH(rectangle1_widths[1768]), .RECT1_HEIGHT(rectangle1_heights[1768]), .RECT1_WEIGHT(rectangle1_weights[1768]), .RECT2_X(rectangle2_xs[1768]), .RECT2_Y(rectangle2_ys[1768]), .RECT2_WIDTH(rectangle2_widths[1768]), .RECT2_HEIGHT(rectangle2_heights[1768]), .RECT2_WEIGHT(rectangle2_weights[1768]), .RECT3_X(rectangle3_xs[1768]), .RECT3_Y(rectangle3_ys[1768]), .RECT3_WIDTH(rectangle3_widths[1768]), .RECT3_HEIGHT(rectangle3_heights[1768]), .RECT3_WEIGHT(rectangle3_weights[1768]), .FEAT_THRES(feature_thresholds[1768]), .FEAT_ABOVE(feature_aboves[1768]), .FEAT_BELOW(feature_belows[1768])) ac1768(.scan_win(scan_win1768), .scan_win_std_dev(scan_win_std_dev[1768]), .feature_accum(feature_accums[1768]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1769]), .RECT1_Y(rectangle1_ys[1769]), .RECT1_WIDTH(rectangle1_widths[1769]), .RECT1_HEIGHT(rectangle1_heights[1769]), .RECT1_WEIGHT(rectangle1_weights[1769]), .RECT2_X(rectangle2_xs[1769]), .RECT2_Y(rectangle2_ys[1769]), .RECT2_WIDTH(rectangle2_widths[1769]), .RECT2_HEIGHT(rectangle2_heights[1769]), .RECT2_WEIGHT(rectangle2_weights[1769]), .RECT3_X(rectangle3_xs[1769]), .RECT3_Y(rectangle3_ys[1769]), .RECT3_WIDTH(rectangle3_widths[1769]), .RECT3_HEIGHT(rectangle3_heights[1769]), .RECT3_WEIGHT(rectangle3_weights[1769]), .FEAT_THRES(feature_thresholds[1769]), .FEAT_ABOVE(feature_aboves[1769]), .FEAT_BELOW(feature_belows[1769])) ac1769(.scan_win(scan_win1769), .scan_win_std_dev(scan_win_std_dev[1769]), .feature_accum(feature_accums[1769]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1770]), .RECT1_Y(rectangle1_ys[1770]), .RECT1_WIDTH(rectangle1_widths[1770]), .RECT1_HEIGHT(rectangle1_heights[1770]), .RECT1_WEIGHT(rectangle1_weights[1770]), .RECT2_X(rectangle2_xs[1770]), .RECT2_Y(rectangle2_ys[1770]), .RECT2_WIDTH(rectangle2_widths[1770]), .RECT2_HEIGHT(rectangle2_heights[1770]), .RECT2_WEIGHT(rectangle2_weights[1770]), .RECT3_X(rectangle3_xs[1770]), .RECT3_Y(rectangle3_ys[1770]), .RECT3_WIDTH(rectangle3_widths[1770]), .RECT3_HEIGHT(rectangle3_heights[1770]), .RECT3_WEIGHT(rectangle3_weights[1770]), .FEAT_THRES(feature_thresholds[1770]), .FEAT_ABOVE(feature_aboves[1770]), .FEAT_BELOW(feature_belows[1770])) ac1770(.scan_win(scan_win1770), .scan_win_std_dev(scan_win_std_dev[1770]), .feature_accum(feature_accums[1770]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1771]), .RECT1_Y(rectangle1_ys[1771]), .RECT1_WIDTH(rectangle1_widths[1771]), .RECT1_HEIGHT(rectangle1_heights[1771]), .RECT1_WEIGHT(rectangle1_weights[1771]), .RECT2_X(rectangle2_xs[1771]), .RECT2_Y(rectangle2_ys[1771]), .RECT2_WIDTH(rectangle2_widths[1771]), .RECT2_HEIGHT(rectangle2_heights[1771]), .RECT2_WEIGHT(rectangle2_weights[1771]), .RECT3_X(rectangle3_xs[1771]), .RECT3_Y(rectangle3_ys[1771]), .RECT3_WIDTH(rectangle3_widths[1771]), .RECT3_HEIGHT(rectangle3_heights[1771]), .RECT3_WEIGHT(rectangle3_weights[1771]), .FEAT_THRES(feature_thresholds[1771]), .FEAT_ABOVE(feature_aboves[1771]), .FEAT_BELOW(feature_belows[1771])) ac1771(.scan_win(scan_win1771), .scan_win_std_dev(scan_win_std_dev[1771]), .feature_accum(feature_accums[1771]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1772]), .RECT1_Y(rectangle1_ys[1772]), .RECT1_WIDTH(rectangle1_widths[1772]), .RECT1_HEIGHT(rectangle1_heights[1772]), .RECT1_WEIGHT(rectangle1_weights[1772]), .RECT2_X(rectangle2_xs[1772]), .RECT2_Y(rectangle2_ys[1772]), .RECT2_WIDTH(rectangle2_widths[1772]), .RECT2_HEIGHT(rectangle2_heights[1772]), .RECT2_WEIGHT(rectangle2_weights[1772]), .RECT3_X(rectangle3_xs[1772]), .RECT3_Y(rectangle3_ys[1772]), .RECT3_WIDTH(rectangle3_widths[1772]), .RECT3_HEIGHT(rectangle3_heights[1772]), .RECT3_WEIGHT(rectangle3_weights[1772]), .FEAT_THRES(feature_thresholds[1772]), .FEAT_ABOVE(feature_aboves[1772]), .FEAT_BELOW(feature_belows[1772])) ac1772(.scan_win(scan_win1772), .scan_win_std_dev(scan_win_std_dev[1772]), .feature_accum(feature_accums[1772]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1773]), .RECT1_Y(rectangle1_ys[1773]), .RECT1_WIDTH(rectangle1_widths[1773]), .RECT1_HEIGHT(rectangle1_heights[1773]), .RECT1_WEIGHT(rectangle1_weights[1773]), .RECT2_X(rectangle2_xs[1773]), .RECT2_Y(rectangle2_ys[1773]), .RECT2_WIDTH(rectangle2_widths[1773]), .RECT2_HEIGHT(rectangle2_heights[1773]), .RECT2_WEIGHT(rectangle2_weights[1773]), .RECT3_X(rectangle3_xs[1773]), .RECT3_Y(rectangle3_ys[1773]), .RECT3_WIDTH(rectangle3_widths[1773]), .RECT3_HEIGHT(rectangle3_heights[1773]), .RECT3_WEIGHT(rectangle3_weights[1773]), .FEAT_THRES(feature_thresholds[1773]), .FEAT_ABOVE(feature_aboves[1773]), .FEAT_BELOW(feature_belows[1773])) ac1773(.scan_win(scan_win1773), .scan_win_std_dev(scan_win_std_dev[1773]), .feature_accum(feature_accums[1773]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1774]), .RECT1_Y(rectangle1_ys[1774]), .RECT1_WIDTH(rectangle1_widths[1774]), .RECT1_HEIGHT(rectangle1_heights[1774]), .RECT1_WEIGHT(rectangle1_weights[1774]), .RECT2_X(rectangle2_xs[1774]), .RECT2_Y(rectangle2_ys[1774]), .RECT2_WIDTH(rectangle2_widths[1774]), .RECT2_HEIGHT(rectangle2_heights[1774]), .RECT2_WEIGHT(rectangle2_weights[1774]), .RECT3_X(rectangle3_xs[1774]), .RECT3_Y(rectangle3_ys[1774]), .RECT3_WIDTH(rectangle3_widths[1774]), .RECT3_HEIGHT(rectangle3_heights[1774]), .RECT3_WEIGHT(rectangle3_weights[1774]), .FEAT_THRES(feature_thresholds[1774]), .FEAT_ABOVE(feature_aboves[1774]), .FEAT_BELOW(feature_belows[1774])) ac1774(.scan_win(scan_win1774), .scan_win_std_dev(scan_win_std_dev[1774]), .feature_accum(feature_accums[1774]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1775]), .RECT1_Y(rectangle1_ys[1775]), .RECT1_WIDTH(rectangle1_widths[1775]), .RECT1_HEIGHT(rectangle1_heights[1775]), .RECT1_WEIGHT(rectangle1_weights[1775]), .RECT2_X(rectangle2_xs[1775]), .RECT2_Y(rectangle2_ys[1775]), .RECT2_WIDTH(rectangle2_widths[1775]), .RECT2_HEIGHT(rectangle2_heights[1775]), .RECT2_WEIGHT(rectangle2_weights[1775]), .RECT3_X(rectangle3_xs[1775]), .RECT3_Y(rectangle3_ys[1775]), .RECT3_WIDTH(rectangle3_widths[1775]), .RECT3_HEIGHT(rectangle3_heights[1775]), .RECT3_WEIGHT(rectangle3_weights[1775]), .FEAT_THRES(feature_thresholds[1775]), .FEAT_ABOVE(feature_aboves[1775]), .FEAT_BELOW(feature_belows[1775])) ac1775(.scan_win(scan_win1775), .scan_win_std_dev(scan_win_std_dev[1775]), .feature_accum(feature_accums[1775]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1776]), .RECT1_Y(rectangle1_ys[1776]), .RECT1_WIDTH(rectangle1_widths[1776]), .RECT1_HEIGHT(rectangle1_heights[1776]), .RECT1_WEIGHT(rectangle1_weights[1776]), .RECT2_X(rectangle2_xs[1776]), .RECT2_Y(rectangle2_ys[1776]), .RECT2_WIDTH(rectangle2_widths[1776]), .RECT2_HEIGHT(rectangle2_heights[1776]), .RECT2_WEIGHT(rectangle2_weights[1776]), .RECT3_X(rectangle3_xs[1776]), .RECT3_Y(rectangle3_ys[1776]), .RECT3_WIDTH(rectangle3_widths[1776]), .RECT3_HEIGHT(rectangle3_heights[1776]), .RECT3_WEIGHT(rectangle3_weights[1776]), .FEAT_THRES(feature_thresholds[1776]), .FEAT_ABOVE(feature_aboves[1776]), .FEAT_BELOW(feature_belows[1776])) ac1776(.scan_win(scan_win1776), .scan_win_std_dev(scan_win_std_dev[1776]), .feature_accum(feature_accums[1776]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1777]), .RECT1_Y(rectangle1_ys[1777]), .RECT1_WIDTH(rectangle1_widths[1777]), .RECT1_HEIGHT(rectangle1_heights[1777]), .RECT1_WEIGHT(rectangle1_weights[1777]), .RECT2_X(rectangle2_xs[1777]), .RECT2_Y(rectangle2_ys[1777]), .RECT2_WIDTH(rectangle2_widths[1777]), .RECT2_HEIGHT(rectangle2_heights[1777]), .RECT2_WEIGHT(rectangle2_weights[1777]), .RECT3_X(rectangle3_xs[1777]), .RECT3_Y(rectangle3_ys[1777]), .RECT3_WIDTH(rectangle3_widths[1777]), .RECT3_HEIGHT(rectangle3_heights[1777]), .RECT3_WEIGHT(rectangle3_weights[1777]), .FEAT_THRES(feature_thresholds[1777]), .FEAT_ABOVE(feature_aboves[1777]), .FEAT_BELOW(feature_belows[1777])) ac1777(.scan_win(scan_win1777), .scan_win_std_dev(scan_win_std_dev[1777]), .feature_accum(feature_accums[1777]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1778]), .RECT1_Y(rectangle1_ys[1778]), .RECT1_WIDTH(rectangle1_widths[1778]), .RECT1_HEIGHT(rectangle1_heights[1778]), .RECT1_WEIGHT(rectangle1_weights[1778]), .RECT2_X(rectangle2_xs[1778]), .RECT2_Y(rectangle2_ys[1778]), .RECT2_WIDTH(rectangle2_widths[1778]), .RECT2_HEIGHT(rectangle2_heights[1778]), .RECT2_WEIGHT(rectangle2_weights[1778]), .RECT3_X(rectangle3_xs[1778]), .RECT3_Y(rectangle3_ys[1778]), .RECT3_WIDTH(rectangle3_widths[1778]), .RECT3_HEIGHT(rectangle3_heights[1778]), .RECT3_WEIGHT(rectangle3_weights[1778]), .FEAT_THRES(feature_thresholds[1778]), .FEAT_ABOVE(feature_aboves[1778]), .FEAT_BELOW(feature_belows[1778])) ac1778(.scan_win(scan_win1778), .scan_win_std_dev(scan_win_std_dev[1778]), .feature_accum(feature_accums[1778]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1779]), .RECT1_Y(rectangle1_ys[1779]), .RECT1_WIDTH(rectangle1_widths[1779]), .RECT1_HEIGHT(rectangle1_heights[1779]), .RECT1_WEIGHT(rectangle1_weights[1779]), .RECT2_X(rectangle2_xs[1779]), .RECT2_Y(rectangle2_ys[1779]), .RECT2_WIDTH(rectangle2_widths[1779]), .RECT2_HEIGHT(rectangle2_heights[1779]), .RECT2_WEIGHT(rectangle2_weights[1779]), .RECT3_X(rectangle3_xs[1779]), .RECT3_Y(rectangle3_ys[1779]), .RECT3_WIDTH(rectangle3_widths[1779]), .RECT3_HEIGHT(rectangle3_heights[1779]), .RECT3_WEIGHT(rectangle3_weights[1779]), .FEAT_THRES(feature_thresholds[1779]), .FEAT_ABOVE(feature_aboves[1779]), .FEAT_BELOW(feature_belows[1779])) ac1779(.scan_win(scan_win1779), .scan_win_std_dev(scan_win_std_dev[1779]), .feature_accum(feature_accums[1779]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1780]), .RECT1_Y(rectangle1_ys[1780]), .RECT1_WIDTH(rectangle1_widths[1780]), .RECT1_HEIGHT(rectangle1_heights[1780]), .RECT1_WEIGHT(rectangle1_weights[1780]), .RECT2_X(rectangle2_xs[1780]), .RECT2_Y(rectangle2_ys[1780]), .RECT2_WIDTH(rectangle2_widths[1780]), .RECT2_HEIGHT(rectangle2_heights[1780]), .RECT2_WEIGHT(rectangle2_weights[1780]), .RECT3_X(rectangle3_xs[1780]), .RECT3_Y(rectangle3_ys[1780]), .RECT3_WIDTH(rectangle3_widths[1780]), .RECT3_HEIGHT(rectangle3_heights[1780]), .RECT3_WEIGHT(rectangle3_weights[1780]), .FEAT_THRES(feature_thresholds[1780]), .FEAT_ABOVE(feature_aboves[1780]), .FEAT_BELOW(feature_belows[1780])) ac1780(.scan_win(scan_win1780), .scan_win_std_dev(scan_win_std_dev[1780]), .feature_accum(feature_accums[1780]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1781]), .RECT1_Y(rectangle1_ys[1781]), .RECT1_WIDTH(rectangle1_widths[1781]), .RECT1_HEIGHT(rectangle1_heights[1781]), .RECT1_WEIGHT(rectangle1_weights[1781]), .RECT2_X(rectangle2_xs[1781]), .RECT2_Y(rectangle2_ys[1781]), .RECT2_WIDTH(rectangle2_widths[1781]), .RECT2_HEIGHT(rectangle2_heights[1781]), .RECT2_WEIGHT(rectangle2_weights[1781]), .RECT3_X(rectangle3_xs[1781]), .RECT3_Y(rectangle3_ys[1781]), .RECT3_WIDTH(rectangle3_widths[1781]), .RECT3_HEIGHT(rectangle3_heights[1781]), .RECT3_WEIGHT(rectangle3_weights[1781]), .FEAT_THRES(feature_thresholds[1781]), .FEAT_ABOVE(feature_aboves[1781]), .FEAT_BELOW(feature_belows[1781])) ac1781(.scan_win(scan_win1781), .scan_win_std_dev(scan_win_std_dev[1781]), .feature_accum(feature_accums[1781]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1782]), .RECT1_Y(rectangle1_ys[1782]), .RECT1_WIDTH(rectangle1_widths[1782]), .RECT1_HEIGHT(rectangle1_heights[1782]), .RECT1_WEIGHT(rectangle1_weights[1782]), .RECT2_X(rectangle2_xs[1782]), .RECT2_Y(rectangle2_ys[1782]), .RECT2_WIDTH(rectangle2_widths[1782]), .RECT2_HEIGHT(rectangle2_heights[1782]), .RECT2_WEIGHT(rectangle2_weights[1782]), .RECT3_X(rectangle3_xs[1782]), .RECT3_Y(rectangle3_ys[1782]), .RECT3_WIDTH(rectangle3_widths[1782]), .RECT3_HEIGHT(rectangle3_heights[1782]), .RECT3_WEIGHT(rectangle3_weights[1782]), .FEAT_THRES(feature_thresholds[1782]), .FEAT_ABOVE(feature_aboves[1782]), .FEAT_BELOW(feature_belows[1782])) ac1782(.scan_win(scan_win1782), .scan_win_std_dev(scan_win_std_dev[1782]), .feature_accum(feature_accums[1782]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1783]), .RECT1_Y(rectangle1_ys[1783]), .RECT1_WIDTH(rectangle1_widths[1783]), .RECT1_HEIGHT(rectangle1_heights[1783]), .RECT1_WEIGHT(rectangle1_weights[1783]), .RECT2_X(rectangle2_xs[1783]), .RECT2_Y(rectangle2_ys[1783]), .RECT2_WIDTH(rectangle2_widths[1783]), .RECT2_HEIGHT(rectangle2_heights[1783]), .RECT2_WEIGHT(rectangle2_weights[1783]), .RECT3_X(rectangle3_xs[1783]), .RECT3_Y(rectangle3_ys[1783]), .RECT3_WIDTH(rectangle3_widths[1783]), .RECT3_HEIGHT(rectangle3_heights[1783]), .RECT3_WEIGHT(rectangle3_weights[1783]), .FEAT_THRES(feature_thresholds[1783]), .FEAT_ABOVE(feature_aboves[1783]), .FEAT_BELOW(feature_belows[1783])) ac1783(.scan_win(scan_win1783), .scan_win_std_dev(scan_win_std_dev[1783]), .feature_accum(feature_accums[1783]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1784]), .RECT1_Y(rectangle1_ys[1784]), .RECT1_WIDTH(rectangle1_widths[1784]), .RECT1_HEIGHT(rectangle1_heights[1784]), .RECT1_WEIGHT(rectangle1_weights[1784]), .RECT2_X(rectangle2_xs[1784]), .RECT2_Y(rectangle2_ys[1784]), .RECT2_WIDTH(rectangle2_widths[1784]), .RECT2_HEIGHT(rectangle2_heights[1784]), .RECT2_WEIGHT(rectangle2_weights[1784]), .RECT3_X(rectangle3_xs[1784]), .RECT3_Y(rectangle3_ys[1784]), .RECT3_WIDTH(rectangle3_widths[1784]), .RECT3_HEIGHT(rectangle3_heights[1784]), .RECT3_WEIGHT(rectangle3_weights[1784]), .FEAT_THRES(feature_thresholds[1784]), .FEAT_ABOVE(feature_aboves[1784]), .FEAT_BELOW(feature_belows[1784])) ac1784(.scan_win(scan_win1784), .scan_win_std_dev(scan_win_std_dev[1784]), .feature_accum(feature_accums[1784]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1785]), .RECT1_Y(rectangle1_ys[1785]), .RECT1_WIDTH(rectangle1_widths[1785]), .RECT1_HEIGHT(rectangle1_heights[1785]), .RECT1_WEIGHT(rectangle1_weights[1785]), .RECT2_X(rectangle2_xs[1785]), .RECT2_Y(rectangle2_ys[1785]), .RECT2_WIDTH(rectangle2_widths[1785]), .RECT2_HEIGHT(rectangle2_heights[1785]), .RECT2_WEIGHT(rectangle2_weights[1785]), .RECT3_X(rectangle3_xs[1785]), .RECT3_Y(rectangle3_ys[1785]), .RECT3_WIDTH(rectangle3_widths[1785]), .RECT3_HEIGHT(rectangle3_heights[1785]), .RECT3_WEIGHT(rectangle3_weights[1785]), .FEAT_THRES(feature_thresholds[1785]), .FEAT_ABOVE(feature_aboves[1785]), .FEAT_BELOW(feature_belows[1785])) ac1785(.scan_win(scan_win1785), .scan_win_std_dev(scan_win_std_dev[1785]), .feature_accum(feature_accums[1785]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1786]), .RECT1_Y(rectangle1_ys[1786]), .RECT1_WIDTH(rectangle1_widths[1786]), .RECT1_HEIGHT(rectangle1_heights[1786]), .RECT1_WEIGHT(rectangle1_weights[1786]), .RECT2_X(rectangle2_xs[1786]), .RECT2_Y(rectangle2_ys[1786]), .RECT2_WIDTH(rectangle2_widths[1786]), .RECT2_HEIGHT(rectangle2_heights[1786]), .RECT2_WEIGHT(rectangle2_weights[1786]), .RECT3_X(rectangle3_xs[1786]), .RECT3_Y(rectangle3_ys[1786]), .RECT3_WIDTH(rectangle3_widths[1786]), .RECT3_HEIGHT(rectangle3_heights[1786]), .RECT3_WEIGHT(rectangle3_weights[1786]), .FEAT_THRES(feature_thresholds[1786]), .FEAT_ABOVE(feature_aboves[1786]), .FEAT_BELOW(feature_belows[1786])) ac1786(.scan_win(scan_win1786), .scan_win_std_dev(scan_win_std_dev[1786]), .feature_accum(feature_accums[1786]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1787]), .RECT1_Y(rectangle1_ys[1787]), .RECT1_WIDTH(rectangle1_widths[1787]), .RECT1_HEIGHT(rectangle1_heights[1787]), .RECT1_WEIGHT(rectangle1_weights[1787]), .RECT2_X(rectangle2_xs[1787]), .RECT2_Y(rectangle2_ys[1787]), .RECT2_WIDTH(rectangle2_widths[1787]), .RECT2_HEIGHT(rectangle2_heights[1787]), .RECT2_WEIGHT(rectangle2_weights[1787]), .RECT3_X(rectangle3_xs[1787]), .RECT3_Y(rectangle3_ys[1787]), .RECT3_WIDTH(rectangle3_widths[1787]), .RECT3_HEIGHT(rectangle3_heights[1787]), .RECT3_WEIGHT(rectangle3_weights[1787]), .FEAT_THRES(feature_thresholds[1787]), .FEAT_ABOVE(feature_aboves[1787]), .FEAT_BELOW(feature_belows[1787])) ac1787(.scan_win(scan_win1787), .scan_win_std_dev(scan_win_std_dev[1787]), .feature_accum(feature_accums[1787]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1788]), .RECT1_Y(rectangle1_ys[1788]), .RECT1_WIDTH(rectangle1_widths[1788]), .RECT1_HEIGHT(rectangle1_heights[1788]), .RECT1_WEIGHT(rectangle1_weights[1788]), .RECT2_X(rectangle2_xs[1788]), .RECT2_Y(rectangle2_ys[1788]), .RECT2_WIDTH(rectangle2_widths[1788]), .RECT2_HEIGHT(rectangle2_heights[1788]), .RECT2_WEIGHT(rectangle2_weights[1788]), .RECT3_X(rectangle3_xs[1788]), .RECT3_Y(rectangle3_ys[1788]), .RECT3_WIDTH(rectangle3_widths[1788]), .RECT3_HEIGHT(rectangle3_heights[1788]), .RECT3_WEIGHT(rectangle3_weights[1788]), .FEAT_THRES(feature_thresholds[1788]), .FEAT_ABOVE(feature_aboves[1788]), .FEAT_BELOW(feature_belows[1788])) ac1788(.scan_win(scan_win1788), .scan_win_std_dev(scan_win_std_dev[1788]), .feature_accum(feature_accums[1788]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1789]), .RECT1_Y(rectangle1_ys[1789]), .RECT1_WIDTH(rectangle1_widths[1789]), .RECT1_HEIGHT(rectangle1_heights[1789]), .RECT1_WEIGHT(rectangle1_weights[1789]), .RECT2_X(rectangle2_xs[1789]), .RECT2_Y(rectangle2_ys[1789]), .RECT2_WIDTH(rectangle2_widths[1789]), .RECT2_HEIGHT(rectangle2_heights[1789]), .RECT2_WEIGHT(rectangle2_weights[1789]), .RECT3_X(rectangle3_xs[1789]), .RECT3_Y(rectangle3_ys[1789]), .RECT3_WIDTH(rectangle3_widths[1789]), .RECT3_HEIGHT(rectangle3_heights[1789]), .RECT3_WEIGHT(rectangle3_weights[1789]), .FEAT_THRES(feature_thresholds[1789]), .FEAT_ABOVE(feature_aboves[1789]), .FEAT_BELOW(feature_belows[1789])) ac1789(.scan_win(scan_win1789), .scan_win_std_dev(scan_win_std_dev[1789]), .feature_accum(feature_accums[1789]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1790]), .RECT1_Y(rectangle1_ys[1790]), .RECT1_WIDTH(rectangle1_widths[1790]), .RECT1_HEIGHT(rectangle1_heights[1790]), .RECT1_WEIGHT(rectangle1_weights[1790]), .RECT2_X(rectangle2_xs[1790]), .RECT2_Y(rectangle2_ys[1790]), .RECT2_WIDTH(rectangle2_widths[1790]), .RECT2_HEIGHT(rectangle2_heights[1790]), .RECT2_WEIGHT(rectangle2_weights[1790]), .RECT3_X(rectangle3_xs[1790]), .RECT3_Y(rectangle3_ys[1790]), .RECT3_WIDTH(rectangle3_widths[1790]), .RECT3_HEIGHT(rectangle3_heights[1790]), .RECT3_WEIGHT(rectangle3_weights[1790]), .FEAT_THRES(feature_thresholds[1790]), .FEAT_ABOVE(feature_aboves[1790]), .FEAT_BELOW(feature_belows[1790])) ac1790(.scan_win(scan_win1790), .scan_win_std_dev(scan_win_std_dev[1790]), .feature_accum(feature_accums[1790]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1791]), .RECT1_Y(rectangle1_ys[1791]), .RECT1_WIDTH(rectangle1_widths[1791]), .RECT1_HEIGHT(rectangle1_heights[1791]), .RECT1_WEIGHT(rectangle1_weights[1791]), .RECT2_X(rectangle2_xs[1791]), .RECT2_Y(rectangle2_ys[1791]), .RECT2_WIDTH(rectangle2_widths[1791]), .RECT2_HEIGHT(rectangle2_heights[1791]), .RECT2_WEIGHT(rectangle2_weights[1791]), .RECT3_X(rectangle3_xs[1791]), .RECT3_Y(rectangle3_ys[1791]), .RECT3_WIDTH(rectangle3_widths[1791]), .RECT3_HEIGHT(rectangle3_heights[1791]), .RECT3_WEIGHT(rectangle3_weights[1791]), .FEAT_THRES(feature_thresholds[1791]), .FEAT_ABOVE(feature_aboves[1791]), .FEAT_BELOW(feature_belows[1791])) ac1791(.scan_win(scan_win1791), .scan_win_std_dev(scan_win_std_dev[1791]), .feature_accum(feature_accums[1791]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1792]), .RECT1_Y(rectangle1_ys[1792]), .RECT1_WIDTH(rectangle1_widths[1792]), .RECT1_HEIGHT(rectangle1_heights[1792]), .RECT1_WEIGHT(rectangle1_weights[1792]), .RECT2_X(rectangle2_xs[1792]), .RECT2_Y(rectangle2_ys[1792]), .RECT2_WIDTH(rectangle2_widths[1792]), .RECT2_HEIGHT(rectangle2_heights[1792]), .RECT2_WEIGHT(rectangle2_weights[1792]), .RECT3_X(rectangle3_xs[1792]), .RECT3_Y(rectangle3_ys[1792]), .RECT3_WIDTH(rectangle3_widths[1792]), .RECT3_HEIGHT(rectangle3_heights[1792]), .RECT3_WEIGHT(rectangle3_weights[1792]), .FEAT_THRES(feature_thresholds[1792]), .FEAT_ABOVE(feature_aboves[1792]), .FEAT_BELOW(feature_belows[1792])) ac1792(.scan_win(scan_win1792), .scan_win_std_dev(scan_win_std_dev[1792]), .feature_accum(feature_accums[1792]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1793]), .RECT1_Y(rectangle1_ys[1793]), .RECT1_WIDTH(rectangle1_widths[1793]), .RECT1_HEIGHT(rectangle1_heights[1793]), .RECT1_WEIGHT(rectangle1_weights[1793]), .RECT2_X(rectangle2_xs[1793]), .RECT2_Y(rectangle2_ys[1793]), .RECT2_WIDTH(rectangle2_widths[1793]), .RECT2_HEIGHT(rectangle2_heights[1793]), .RECT2_WEIGHT(rectangle2_weights[1793]), .RECT3_X(rectangle3_xs[1793]), .RECT3_Y(rectangle3_ys[1793]), .RECT3_WIDTH(rectangle3_widths[1793]), .RECT3_HEIGHT(rectangle3_heights[1793]), .RECT3_WEIGHT(rectangle3_weights[1793]), .FEAT_THRES(feature_thresholds[1793]), .FEAT_ABOVE(feature_aboves[1793]), .FEAT_BELOW(feature_belows[1793])) ac1793(.scan_win(scan_win1793), .scan_win_std_dev(scan_win_std_dev[1793]), .feature_accum(feature_accums[1793]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1794]), .RECT1_Y(rectangle1_ys[1794]), .RECT1_WIDTH(rectangle1_widths[1794]), .RECT1_HEIGHT(rectangle1_heights[1794]), .RECT1_WEIGHT(rectangle1_weights[1794]), .RECT2_X(rectangle2_xs[1794]), .RECT2_Y(rectangle2_ys[1794]), .RECT2_WIDTH(rectangle2_widths[1794]), .RECT2_HEIGHT(rectangle2_heights[1794]), .RECT2_WEIGHT(rectangle2_weights[1794]), .RECT3_X(rectangle3_xs[1794]), .RECT3_Y(rectangle3_ys[1794]), .RECT3_WIDTH(rectangle3_widths[1794]), .RECT3_HEIGHT(rectangle3_heights[1794]), .RECT3_WEIGHT(rectangle3_weights[1794]), .FEAT_THRES(feature_thresholds[1794]), .FEAT_ABOVE(feature_aboves[1794]), .FEAT_BELOW(feature_belows[1794])) ac1794(.scan_win(scan_win1794), .scan_win_std_dev(scan_win_std_dev[1794]), .feature_accum(feature_accums[1794]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1795]), .RECT1_Y(rectangle1_ys[1795]), .RECT1_WIDTH(rectangle1_widths[1795]), .RECT1_HEIGHT(rectangle1_heights[1795]), .RECT1_WEIGHT(rectangle1_weights[1795]), .RECT2_X(rectangle2_xs[1795]), .RECT2_Y(rectangle2_ys[1795]), .RECT2_WIDTH(rectangle2_widths[1795]), .RECT2_HEIGHT(rectangle2_heights[1795]), .RECT2_WEIGHT(rectangle2_weights[1795]), .RECT3_X(rectangle3_xs[1795]), .RECT3_Y(rectangle3_ys[1795]), .RECT3_WIDTH(rectangle3_widths[1795]), .RECT3_HEIGHT(rectangle3_heights[1795]), .RECT3_WEIGHT(rectangle3_weights[1795]), .FEAT_THRES(feature_thresholds[1795]), .FEAT_ABOVE(feature_aboves[1795]), .FEAT_BELOW(feature_belows[1795])) ac1795(.scan_win(scan_win1795), .scan_win_std_dev(scan_win_std_dev[1795]), .feature_accum(feature_accums[1795]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1796]), .RECT1_Y(rectangle1_ys[1796]), .RECT1_WIDTH(rectangle1_widths[1796]), .RECT1_HEIGHT(rectangle1_heights[1796]), .RECT1_WEIGHT(rectangle1_weights[1796]), .RECT2_X(rectangle2_xs[1796]), .RECT2_Y(rectangle2_ys[1796]), .RECT2_WIDTH(rectangle2_widths[1796]), .RECT2_HEIGHT(rectangle2_heights[1796]), .RECT2_WEIGHT(rectangle2_weights[1796]), .RECT3_X(rectangle3_xs[1796]), .RECT3_Y(rectangle3_ys[1796]), .RECT3_WIDTH(rectangle3_widths[1796]), .RECT3_HEIGHT(rectangle3_heights[1796]), .RECT3_WEIGHT(rectangle3_weights[1796]), .FEAT_THRES(feature_thresholds[1796]), .FEAT_ABOVE(feature_aboves[1796]), .FEAT_BELOW(feature_belows[1796])) ac1796(.scan_win(scan_win1796), .scan_win_std_dev(scan_win_std_dev[1796]), .feature_accum(feature_accums[1796]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1797]), .RECT1_Y(rectangle1_ys[1797]), .RECT1_WIDTH(rectangle1_widths[1797]), .RECT1_HEIGHT(rectangle1_heights[1797]), .RECT1_WEIGHT(rectangle1_weights[1797]), .RECT2_X(rectangle2_xs[1797]), .RECT2_Y(rectangle2_ys[1797]), .RECT2_WIDTH(rectangle2_widths[1797]), .RECT2_HEIGHT(rectangle2_heights[1797]), .RECT2_WEIGHT(rectangle2_weights[1797]), .RECT3_X(rectangle3_xs[1797]), .RECT3_Y(rectangle3_ys[1797]), .RECT3_WIDTH(rectangle3_widths[1797]), .RECT3_HEIGHT(rectangle3_heights[1797]), .RECT3_WEIGHT(rectangle3_weights[1797]), .FEAT_THRES(feature_thresholds[1797]), .FEAT_ABOVE(feature_aboves[1797]), .FEAT_BELOW(feature_belows[1797])) ac1797(.scan_win(scan_win1797), .scan_win_std_dev(scan_win_std_dev[1797]), .feature_accum(feature_accums[1797]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1798]), .RECT1_Y(rectangle1_ys[1798]), .RECT1_WIDTH(rectangle1_widths[1798]), .RECT1_HEIGHT(rectangle1_heights[1798]), .RECT1_WEIGHT(rectangle1_weights[1798]), .RECT2_X(rectangle2_xs[1798]), .RECT2_Y(rectangle2_ys[1798]), .RECT2_WIDTH(rectangle2_widths[1798]), .RECT2_HEIGHT(rectangle2_heights[1798]), .RECT2_WEIGHT(rectangle2_weights[1798]), .RECT3_X(rectangle3_xs[1798]), .RECT3_Y(rectangle3_ys[1798]), .RECT3_WIDTH(rectangle3_widths[1798]), .RECT3_HEIGHT(rectangle3_heights[1798]), .RECT3_WEIGHT(rectangle3_weights[1798]), .FEAT_THRES(feature_thresholds[1798]), .FEAT_ABOVE(feature_aboves[1798]), .FEAT_BELOW(feature_belows[1798])) ac1798(.scan_win(scan_win1798), .scan_win_std_dev(scan_win_std_dev[1798]), .feature_accum(feature_accums[1798]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1799]), .RECT1_Y(rectangle1_ys[1799]), .RECT1_WIDTH(rectangle1_widths[1799]), .RECT1_HEIGHT(rectangle1_heights[1799]), .RECT1_WEIGHT(rectangle1_weights[1799]), .RECT2_X(rectangle2_xs[1799]), .RECT2_Y(rectangle2_ys[1799]), .RECT2_WIDTH(rectangle2_widths[1799]), .RECT2_HEIGHT(rectangle2_heights[1799]), .RECT2_WEIGHT(rectangle2_weights[1799]), .RECT3_X(rectangle3_xs[1799]), .RECT3_Y(rectangle3_ys[1799]), .RECT3_WIDTH(rectangle3_widths[1799]), .RECT3_HEIGHT(rectangle3_heights[1799]), .RECT3_WEIGHT(rectangle3_weights[1799]), .FEAT_THRES(feature_thresholds[1799]), .FEAT_ABOVE(feature_aboves[1799]), .FEAT_BELOW(feature_belows[1799])) ac1799(.scan_win(scan_win1799), .scan_win_std_dev(scan_win_std_dev[1799]), .feature_accum(feature_accums[1799]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1800]), .RECT1_Y(rectangle1_ys[1800]), .RECT1_WIDTH(rectangle1_widths[1800]), .RECT1_HEIGHT(rectangle1_heights[1800]), .RECT1_WEIGHT(rectangle1_weights[1800]), .RECT2_X(rectangle2_xs[1800]), .RECT2_Y(rectangle2_ys[1800]), .RECT2_WIDTH(rectangle2_widths[1800]), .RECT2_HEIGHT(rectangle2_heights[1800]), .RECT2_WEIGHT(rectangle2_weights[1800]), .RECT3_X(rectangle3_xs[1800]), .RECT3_Y(rectangle3_ys[1800]), .RECT3_WIDTH(rectangle3_widths[1800]), .RECT3_HEIGHT(rectangle3_heights[1800]), .RECT3_WEIGHT(rectangle3_weights[1800]), .FEAT_THRES(feature_thresholds[1800]), .FEAT_ABOVE(feature_aboves[1800]), .FEAT_BELOW(feature_belows[1800])) ac1800(.scan_win(scan_win1800), .scan_win_std_dev(scan_win_std_dev[1800]), .feature_accum(feature_accums[1800]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1801]), .RECT1_Y(rectangle1_ys[1801]), .RECT1_WIDTH(rectangle1_widths[1801]), .RECT1_HEIGHT(rectangle1_heights[1801]), .RECT1_WEIGHT(rectangle1_weights[1801]), .RECT2_X(rectangle2_xs[1801]), .RECT2_Y(rectangle2_ys[1801]), .RECT2_WIDTH(rectangle2_widths[1801]), .RECT2_HEIGHT(rectangle2_heights[1801]), .RECT2_WEIGHT(rectangle2_weights[1801]), .RECT3_X(rectangle3_xs[1801]), .RECT3_Y(rectangle3_ys[1801]), .RECT3_WIDTH(rectangle3_widths[1801]), .RECT3_HEIGHT(rectangle3_heights[1801]), .RECT3_WEIGHT(rectangle3_weights[1801]), .FEAT_THRES(feature_thresholds[1801]), .FEAT_ABOVE(feature_aboves[1801]), .FEAT_BELOW(feature_belows[1801])) ac1801(.scan_win(scan_win1801), .scan_win_std_dev(scan_win_std_dev[1801]), .feature_accum(feature_accums[1801]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1802]), .RECT1_Y(rectangle1_ys[1802]), .RECT1_WIDTH(rectangle1_widths[1802]), .RECT1_HEIGHT(rectangle1_heights[1802]), .RECT1_WEIGHT(rectangle1_weights[1802]), .RECT2_X(rectangle2_xs[1802]), .RECT2_Y(rectangle2_ys[1802]), .RECT2_WIDTH(rectangle2_widths[1802]), .RECT2_HEIGHT(rectangle2_heights[1802]), .RECT2_WEIGHT(rectangle2_weights[1802]), .RECT3_X(rectangle3_xs[1802]), .RECT3_Y(rectangle3_ys[1802]), .RECT3_WIDTH(rectangle3_widths[1802]), .RECT3_HEIGHT(rectangle3_heights[1802]), .RECT3_WEIGHT(rectangle3_weights[1802]), .FEAT_THRES(feature_thresholds[1802]), .FEAT_ABOVE(feature_aboves[1802]), .FEAT_BELOW(feature_belows[1802])) ac1802(.scan_win(scan_win1802), .scan_win_std_dev(scan_win_std_dev[1802]), .feature_accum(feature_accums[1802]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1803]), .RECT1_Y(rectangle1_ys[1803]), .RECT1_WIDTH(rectangle1_widths[1803]), .RECT1_HEIGHT(rectangle1_heights[1803]), .RECT1_WEIGHT(rectangle1_weights[1803]), .RECT2_X(rectangle2_xs[1803]), .RECT2_Y(rectangle2_ys[1803]), .RECT2_WIDTH(rectangle2_widths[1803]), .RECT2_HEIGHT(rectangle2_heights[1803]), .RECT2_WEIGHT(rectangle2_weights[1803]), .RECT3_X(rectangle3_xs[1803]), .RECT3_Y(rectangle3_ys[1803]), .RECT3_WIDTH(rectangle3_widths[1803]), .RECT3_HEIGHT(rectangle3_heights[1803]), .RECT3_WEIGHT(rectangle3_weights[1803]), .FEAT_THRES(feature_thresholds[1803]), .FEAT_ABOVE(feature_aboves[1803]), .FEAT_BELOW(feature_belows[1803])) ac1803(.scan_win(scan_win1803), .scan_win_std_dev(scan_win_std_dev[1803]), .feature_accum(feature_accums[1803]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1804]), .RECT1_Y(rectangle1_ys[1804]), .RECT1_WIDTH(rectangle1_widths[1804]), .RECT1_HEIGHT(rectangle1_heights[1804]), .RECT1_WEIGHT(rectangle1_weights[1804]), .RECT2_X(rectangle2_xs[1804]), .RECT2_Y(rectangle2_ys[1804]), .RECT2_WIDTH(rectangle2_widths[1804]), .RECT2_HEIGHT(rectangle2_heights[1804]), .RECT2_WEIGHT(rectangle2_weights[1804]), .RECT3_X(rectangle3_xs[1804]), .RECT3_Y(rectangle3_ys[1804]), .RECT3_WIDTH(rectangle3_widths[1804]), .RECT3_HEIGHT(rectangle3_heights[1804]), .RECT3_WEIGHT(rectangle3_weights[1804]), .FEAT_THRES(feature_thresholds[1804]), .FEAT_ABOVE(feature_aboves[1804]), .FEAT_BELOW(feature_belows[1804])) ac1804(.scan_win(scan_win1804), .scan_win_std_dev(scan_win_std_dev[1804]), .feature_accum(feature_accums[1804]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1805]), .RECT1_Y(rectangle1_ys[1805]), .RECT1_WIDTH(rectangle1_widths[1805]), .RECT1_HEIGHT(rectangle1_heights[1805]), .RECT1_WEIGHT(rectangle1_weights[1805]), .RECT2_X(rectangle2_xs[1805]), .RECT2_Y(rectangle2_ys[1805]), .RECT2_WIDTH(rectangle2_widths[1805]), .RECT2_HEIGHT(rectangle2_heights[1805]), .RECT2_WEIGHT(rectangle2_weights[1805]), .RECT3_X(rectangle3_xs[1805]), .RECT3_Y(rectangle3_ys[1805]), .RECT3_WIDTH(rectangle3_widths[1805]), .RECT3_HEIGHT(rectangle3_heights[1805]), .RECT3_WEIGHT(rectangle3_weights[1805]), .FEAT_THRES(feature_thresholds[1805]), .FEAT_ABOVE(feature_aboves[1805]), .FEAT_BELOW(feature_belows[1805])) ac1805(.scan_win(scan_win1805), .scan_win_std_dev(scan_win_std_dev[1805]), .feature_accum(feature_accums[1805]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1806]), .RECT1_Y(rectangle1_ys[1806]), .RECT1_WIDTH(rectangle1_widths[1806]), .RECT1_HEIGHT(rectangle1_heights[1806]), .RECT1_WEIGHT(rectangle1_weights[1806]), .RECT2_X(rectangle2_xs[1806]), .RECT2_Y(rectangle2_ys[1806]), .RECT2_WIDTH(rectangle2_widths[1806]), .RECT2_HEIGHT(rectangle2_heights[1806]), .RECT2_WEIGHT(rectangle2_weights[1806]), .RECT3_X(rectangle3_xs[1806]), .RECT3_Y(rectangle3_ys[1806]), .RECT3_WIDTH(rectangle3_widths[1806]), .RECT3_HEIGHT(rectangle3_heights[1806]), .RECT3_WEIGHT(rectangle3_weights[1806]), .FEAT_THRES(feature_thresholds[1806]), .FEAT_ABOVE(feature_aboves[1806]), .FEAT_BELOW(feature_belows[1806])) ac1806(.scan_win(scan_win1806), .scan_win_std_dev(scan_win_std_dev[1806]), .feature_accum(feature_accums[1806]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1807]), .RECT1_Y(rectangle1_ys[1807]), .RECT1_WIDTH(rectangle1_widths[1807]), .RECT1_HEIGHT(rectangle1_heights[1807]), .RECT1_WEIGHT(rectangle1_weights[1807]), .RECT2_X(rectangle2_xs[1807]), .RECT2_Y(rectangle2_ys[1807]), .RECT2_WIDTH(rectangle2_widths[1807]), .RECT2_HEIGHT(rectangle2_heights[1807]), .RECT2_WEIGHT(rectangle2_weights[1807]), .RECT3_X(rectangle3_xs[1807]), .RECT3_Y(rectangle3_ys[1807]), .RECT3_WIDTH(rectangle3_widths[1807]), .RECT3_HEIGHT(rectangle3_heights[1807]), .RECT3_WEIGHT(rectangle3_weights[1807]), .FEAT_THRES(feature_thresholds[1807]), .FEAT_ABOVE(feature_aboves[1807]), .FEAT_BELOW(feature_belows[1807])) ac1807(.scan_win(scan_win1807), .scan_win_std_dev(scan_win_std_dev[1807]), .feature_accum(feature_accums[1807]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1808]), .RECT1_Y(rectangle1_ys[1808]), .RECT1_WIDTH(rectangle1_widths[1808]), .RECT1_HEIGHT(rectangle1_heights[1808]), .RECT1_WEIGHT(rectangle1_weights[1808]), .RECT2_X(rectangle2_xs[1808]), .RECT2_Y(rectangle2_ys[1808]), .RECT2_WIDTH(rectangle2_widths[1808]), .RECT2_HEIGHT(rectangle2_heights[1808]), .RECT2_WEIGHT(rectangle2_weights[1808]), .RECT3_X(rectangle3_xs[1808]), .RECT3_Y(rectangle3_ys[1808]), .RECT3_WIDTH(rectangle3_widths[1808]), .RECT3_HEIGHT(rectangle3_heights[1808]), .RECT3_WEIGHT(rectangle3_weights[1808]), .FEAT_THRES(feature_thresholds[1808]), .FEAT_ABOVE(feature_aboves[1808]), .FEAT_BELOW(feature_belows[1808])) ac1808(.scan_win(scan_win1808), .scan_win_std_dev(scan_win_std_dev[1808]), .feature_accum(feature_accums[1808]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1809]), .RECT1_Y(rectangle1_ys[1809]), .RECT1_WIDTH(rectangle1_widths[1809]), .RECT1_HEIGHT(rectangle1_heights[1809]), .RECT1_WEIGHT(rectangle1_weights[1809]), .RECT2_X(rectangle2_xs[1809]), .RECT2_Y(rectangle2_ys[1809]), .RECT2_WIDTH(rectangle2_widths[1809]), .RECT2_HEIGHT(rectangle2_heights[1809]), .RECT2_WEIGHT(rectangle2_weights[1809]), .RECT3_X(rectangle3_xs[1809]), .RECT3_Y(rectangle3_ys[1809]), .RECT3_WIDTH(rectangle3_widths[1809]), .RECT3_HEIGHT(rectangle3_heights[1809]), .RECT3_WEIGHT(rectangle3_weights[1809]), .FEAT_THRES(feature_thresholds[1809]), .FEAT_ABOVE(feature_aboves[1809]), .FEAT_BELOW(feature_belows[1809])) ac1809(.scan_win(scan_win1809), .scan_win_std_dev(scan_win_std_dev[1809]), .feature_accum(feature_accums[1809]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1810]), .RECT1_Y(rectangle1_ys[1810]), .RECT1_WIDTH(rectangle1_widths[1810]), .RECT1_HEIGHT(rectangle1_heights[1810]), .RECT1_WEIGHT(rectangle1_weights[1810]), .RECT2_X(rectangle2_xs[1810]), .RECT2_Y(rectangle2_ys[1810]), .RECT2_WIDTH(rectangle2_widths[1810]), .RECT2_HEIGHT(rectangle2_heights[1810]), .RECT2_WEIGHT(rectangle2_weights[1810]), .RECT3_X(rectangle3_xs[1810]), .RECT3_Y(rectangle3_ys[1810]), .RECT3_WIDTH(rectangle3_widths[1810]), .RECT3_HEIGHT(rectangle3_heights[1810]), .RECT3_WEIGHT(rectangle3_weights[1810]), .FEAT_THRES(feature_thresholds[1810]), .FEAT_ABOVE(feature_aboves[1810]), .FEAT_BELOW(feature_belows[1810])) ac1810(.scan_win(scan_win1810), .scan_win_std_dev(scan_win_std_dev[1810]), .feature_accum(feature_accums[1810]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1811]), .RECT1_Y(rectangle1_ys[1811]), .RECT1_WIDTH(rectangle1_widths[1811]), .RECT1_HEIGHT(rectangle1_heights[1811]), .RECT1_WEIGHT(rectangle1_weights[1811]), .RECT2_X(rectangle2_xs[1811]), .RECT2_Y(rectangle2_ys[1811]), .RECT2_WIDTH(rectangle2_widths[1811]), .RECT2_HEIGHT(rectangle2_heights[1811]), .RECT2_WEIGHT(rectangle2_weights[1811]), .RECT3_X(rectangle3_xs[1811]), .RECT3_Y(rectangle3_ys[1811]), .RECT3_WIDTH(rectangle3_widths[1811]), .RECT3_HEIGHT(rectangle3_heights[1811]), .RECT3_WEIGHT(rectangle3_weights[1811]), .FEAT_THRES(feature_thresholds[1811]), .FEAT_ABOVE(feature_aboves[1811]), .FEAT_BELOW(feature_belows[1811])) ac1811(.scan_win(scan_win1811), .scan_win_std_dev(scan_win_std_dev[1811]), .feature_accum(feature_accums[1811]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1812]), .RECT1_Y(rectangle1_ys[1812]), .RECT1_WIDTH(rectangle1_widths[1812]), .RECT1_HEIGHT(rectangle1_heights[1812]), .RECT1_WEIGHT(rectangle1_weights[1812]), .RECT2_X(rectangle2_xs[1812]), .RECT2_Y(rectangle2_ys[1812]), .RECT2_WIDTH(rectangle2_widths[1812]), .RECT2_HEIGHT(rectangle2_heights[1812]), .RECT2_WEIGHT(rectangle2_weights[1812]), .RECT3_X(rectangle3_xs[1812]), .RECT3_Y(rectangle3_ys[1812]), .RECT3_WIDTH(rectangle3_widths[1812]), .RECT3_HEIGHT(rectangle3_heights[1812]), .RECT3_WEIGHT(rectangle3_weights[1812]), .FEAT_THRES(feature_thresholds[1812]), .FEAT_ABOVE(feature_aboves[1812]), .FEAT_BELOW(feature_belows[1812])) ac1812(.scan_win(scan_win1812), .scan_win_std_dev(scan_win_std_dev[1812]), .feature_accum(feature_accums[1812]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1813]), .RECT1_Y(rectangle1_ys[1813]), .RECT1_WIDTH(rectangle1_widths[1813]), .RECT1_HEIGHT(rectangle1_heights[1813]), .RECT1_WEIGHT(rectangle1_weights[1813]), .RECT2_X(rectangle2_xs[1813]), .RECT2_Y(rectangle2_ys[1813]), .RECT2_WIDTH(rectangle2_widths[1813]), .RECT2_HEIGHT(rectangle2_heights[1813]), .RECT2_WEIGHT(rectangle2_weights[1813]), .RECT3_X(rectangle3_xs[1813]), .RECT3_Y(rectangle3_ys[1813]), .RECT3_WIDTH(rectangle3_widths[1813]), .RECT3_HEIGHT(rectangle3_heights[1813]), .RECT3_WEIGHT(rectangle3_weights[1813]), .FEAT_THRES(feature_thresholds[1813]), .FEAT_ABOVE(feature_aboves[1813]), .FEAT_BELOW(feature_belows[1813])) ac1813(.scan_win(scan_win1813), .scan_win_std_dev(scan_win_std_dev[1813]), .feature_accum(feature_accums[1813]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1814]), .RECT1_Y(rectangle1_ys[1814]), .RECT1_WIDTH(rectangle1_widths[1814]), .RECT1_HEIGHT(rectangle1_heights[1814]), .RECT1_WEIGHT(rectangle1_weights[1814]), .RECT2_X(rectangle2_xs[1814]), .RECT2_Y(rectangle2_ys[1814]), .RECT2_WIDTH(rectangle2_widths[1814]), .RECT2_HEIGHT(rectangle2_heights[1814]), .RECT2_WEIGHT(rectangle2_weights[1814]), .RECT3_X(rectangle3_xs[1814]), .RECT3_Y(rectangle3_ys[1814]), .RECT3_WIDTH(rectangle3_widths[1814]), .RECT3_HEIGHT(rectangle3_heights[1814]), .RECT3_WEIGHT(rectangle3_weights[1814]), .FEAT_THRES(feature_thresholds[1814]), .FEAT_ABOVE(feature_aboves[1814]), .FEAT_BELOW(feature_belows[1814])) ac1814(.scan_win(scan_win1814), .scan_win_std_dev(scan_win_std_dev[1814]), .feature_accum(feature_accums[1814]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1815]), .RECT1_Y(rectangle1_ys[1815]), .RECT1_WIDTH(rectangle1_widths[1815]), .RECT1_HEIGHT(rectangle1_heights[1815]), .RECT1_WEIGHT(rectangle1_weights[1815]), .RECT2_X(rectangle2_xs[1815]), .RECT2_Y(rectangle2_ys[1815]), .RECT2_WIDTH(rectangle2_widths[1815]), .RECT2_HEIGHT(rectangle2_heights[1815]), .RECT2_WEIGHT(rectangle2_weights[1815]), .RECT3_X(rectangle3_xs[1815]), .RECT3_Y(rectangle3_ys[1815]), .RECT3_WIDTH(rectangle3_widths[1815]), .RECT3_HEIGHT(rectangle3_heights[1815]), .RECT3_WEIGHT(rectangle3_weights[1815]), .FEAT_THRES(feature_thresholds[1815]), .FEAT_ABOVE(feature_aboves[1815]), .FEAT_BELOW(feature_belows[1815])) ac1815(.scan_win(scan_win1815), .scan_win_std_dev(scan_win_std_dev[1815]), .feature_accum(feature_accums[1815]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1816]), .RECT1_Y(rectangle1_ys[1816]), .RECT1_WIDTH(rectangle1_widths[1816]), .RECT1_HEIGHT(rectangle1_heights[1816]), .RECT1_WEIGHT(rectangle1_weights[1816]), .RECT2_X(rectangle2_xs[1816]), .RECT2_Y(rectangle2_ys[1816]), .RECT2_WIDTH(rectangle2_widths[1816]), .RECT2_HEIGHT(rectangle2_heights[1816]), .RECT2_WEIGHT(rectangle2_weights[1816]), .RECT3_X(rectangle3_xs[1816]), .RECT3_Y(rectangle3_ys[1816]), .RECT3_WIDTH(rectangle3_widths[1816]), .RECT3_HEIGHT(rectangle3_heights[1816]), .RECT3_WEIGHT(rectangle3_weights[1816]), .FEAT_THRES(feature_thresholds[1816]), .FEAT_ABOVE(feature_aboves[1816]), .FEAT_BELOW(feature_belows[1816])) ac1816(.scan_win(scan_win1816), .scan_win_std_dev(scan_win_std_dev[1816]), .feature_accum(feature_accums[1816]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1817]), .RECT1_Y(rectangle1_ys[1817]), .RECT1_WIDTH(rectangle1_widths[1817]), .RECT1_HEIGHT(rectangle1_heights[1817]), .RECT1_WEIGHT(rectangle1_weights[1817]), .RECT2_X(rectangle2_xs[1817]), .RECT2_Y(rectangle2_ys[1817]), .RECT2_WIDTH(rectangle2_widths[1817]), .RECT2_HEIGHT(rectangle2_heights[1817]), .RECT2_WEIGHT(rectangle2_weights[1817]), .RECT3_X(rectangle3_xs[1817]), .RECT3_Y(rectangle3_ys[1817]), .RECT3_WIDTH(rectangle3_widths[1817]), .RECT3_HEIGHT(rectangle3_heights[1817]), .RECT3_WEIGHT(rectangle3_weights[1817]), .FEAT_THRES(feature_thresholds[1817]), .FEAT_ABOVE(feature_aboves[1817]), .FEAT_BELOW(feature_belows[1817])) ac1817(.scan_win(scan_win1817), .scan_win_std_dev(scan_win_std_dev[1817]), .feature_accum(feature_accums[1817]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1818]), .RECT1_Y(rectangle1_ys[1818]), .RECT1_WIDTH(rectangle1_widths[1818]), .RECT1_HEIGHT(rectangle1_heights[1818]), .RECT1_WEIGHT(rectangle1_weights[1818]), .RECT2_X(rectangle2_xs[1818]), .RECT2_Y(rectangle2_ys[1818]), .RECT2_WIDTH(rectangle2_widths[1818]), .RECT2_HEIGHT(rectangle2_heights[1818]), .RECT2_WEIGHT(rectangle2_weights[1818]), .RECT3_X(rectangle3_xs[1818]), .RECT3_Y(rectangle3_ys[1818]), .RECT3_WIDTH(rectangle3_widths[1818]), .RECT3_HEIGHT(rectangle3_heights[1818]), .RECT3_WEIGHT(rectangle3_weights[1818]), .FEAT_THRES(feature_thresholds[1818]), .FEAT_ABOVE(feature_aboves[1818]), .FEAT_BELOW(feature_belows[1818])) ac1818(.scan_win(scan_win1818), .scan_win_std_dev(scan_win_std_dev[1818]), .feature_accum(feature_accums[1818]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1819]), .RECT1_Y(rectangle1_ys[1819]), .RECT1_WIDTH(rectangle1_widths[1819]), .RECT1_HEIGHT(rectangle1_heights[1819]), .RECT1_WEIGHT(rectangle1_weights[1819]), .RECT2_X(rectangle2_xs[1819]), .RECT2_Y(rectangle2_ys[1819]), .RECT2_WIDTH(rectangle2_widths[1819]), .RECT2_HEIGHT(rectangle2_heights[1819]), .RECT2_WEIGHT(rectangle2_weights[1819]), .RECT3_X(rectangle3_xs[1819]), .RECT3_Y(rectangle3_ys[1819]), .RECT3_WIDTH(rectangle3_widths[1819]), .RECT3_HEIGHT(rectangle3_heights[1819]), .RECT3_WEIGHT(rectangle3_weights[1819]), .FEAT_THRES(feature_thresholds[1819]), .FEAT_ABOVE(feature_aboves[1819]), .FEAT_BELOW(feature_belows[1819])) ac1819(.scan_win(scan_win1819), .scan_win_std_dev(scan_win_std_dev[1819]), .feature_accum(feature_accums[1819]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1820]), .RECT1_Y(rectangle1_ys[1820]), .RECT1_WIDTH(rectangle1_widths[1820]), .RECT1_HEIGHT(rectangle1_heights[1820]), .RECT1_WEIGHT(rectangle1_weights[1820]), .RECT2_X(rectangle2_xs[1820]), .RECT2_Y(rectangle2_ys[1820]), .RECT2_WIDTH(rectangle2_widths[1820]), .RECT2_HEIGHT(rectangle2_heights[1820]), .RECT2_WEIGHT(rectangle2_weights[1820]), .RECT3_X(rectangle3_xs[1820]), .RECT3_Y(rectangle3_ys[1820]), .RECT3_WIDTH(rectangle3_widths[1820]), .RECT3_HEIGHT(rectangle3_heights[1820]), .RECT3_WEIGHT(rectangle3_weights[1820]), .FEAT_THRES(feature_thresholds[1820]), .FEAT_ABOVE(feature_aboves[1820]), .FEAT_BELOW(feature_belows[1820])) ac1820(.scan_win(scan_win1820), .scan_win_std_dev(scan_win_std_dev[1820]), .feature_accum(feature_accums[1820]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1821]), .RECT1_Y(rectangle1_ys[1821]), .RECT1_WIDTH(rectangle1_widths[1821]), .RECT1_HEIGHT(rectangle1_heights[1821]), .RECT1_WEIGHT(rectangle1_weights[1821]), .RECT2_X(rectangle2_xs[1821]), .RECT2_Y(rectangle2_ys[1821]), .RECT2_WIDTH(rectangle2_widths[1821]), .RECT2_HEIGHT(rectangle2_heights[1821]), .RECT2_WEIGHT(rectangle2_weights[1821]), .RECT3_X(rectangle3_xs[1821]), .RECT3_Y(rectangle3_ys[1821]), .RECT3_WIDTH(rectangle3_widths[1821]), .RECT3_HEIGHT(rectangle3_heights[1821]), .RECT3_WEIGHT(rectangle3_weights[1821]), .FEAT_THRES(feature_thresholds[1821]), .FEAT_ABOVE(feature_aboves[1821]), .FEAT_BELOW(feature_belows[1821])) ac1821(.scan_win(scan_win1821), .scan_win_std_dev(scan_win_std_dev[1821]), .feature_accum(feature_accums[1821]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1822]), .RECT1_Y(rectangle1_ys[1822]), .RECT1_WIDTH(rectangle1_widths[1822]), .RECT1_HEIGHT(rectangle1_heights[1822]), .RECT1_WEIGHT(rectangle1_weights[1822]), .RECT2_X(rectangle2_xs[1822]), .RECT2_Y(rectangle2_ys[1822]), .RECT2_WIDTH(rectangle2_widths[1822]), .RECT2_HEIGHT(rectangle2_heights[1822]), .RECT2_WEIGHT(rectangle2_weights[1822]), .RECT3_X(rectangle3_xs[1822]), .RECT3_Y(rectangle3_ys[1822]), .RECT3_WIDTH(rectangle3_widths[1822]), .RECT3_HEIGHT(rectangle3_heights[1822]), .RECT3_WEIGHT(rectangle3_weights[1822]), .FEAT_THRES(feature_thresholds[1822]), .FEAT_ABOVE(feature_aboves[1822]), .FEAT_BELOW(feature_belows[1822])) ac1822(.scan_win(scan_win1822), .scan_win_std_dev(scan_win_std_dev[1822]), .feature_accum(feature_accums[1822]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1823]), .RECT1_Y(rectangle1_ys[1823]), .RECT1_WIDTH(rectangle1_widths[1823]), .RECT1_HEIGHT(rectangle1_heights[1823]), .RECT1_WEIGHT(rectangle1_weights[1823]), .RECT2_X(rectangle2_xs[1823]), .RECT2_Y(rectangle2_ys[1823]), .RECT2_WIDTH(rectangle2_widths[1823]), .RECT2_HEIGHT(rectangle2_heights[1823]), .RECT2_WEIGHT(rectangle2_weights[1823]), .RECT3_X(rectangle3_xs[1823]), .RECT3_Y(rectangle3_ys[1823]), .RECT3_WIDTH(rectangle3_widths[1823]), .RECT3_HEIGHT(rectangle3_heights[1823]), .RECT3_WEIGHT(rectangle3_weights[1823]), .FEAT_THRES(feature_thresholds[1823]), .FEAT_ABOVE(feature_aboves[1823]), .FEAT_BELOW(feature_belows[1823])) ac1823(.scan_win(scan_win1823), .scan_win_std_dev(scan_win_std_dev[1823]), .feature_accum(feature_accums[1823]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1824]), .RECT1_Y(rectangle1_ys[1824]), .RECT1_WIDTH(rectangle1_widths[1824]), .RECT1_HEIGHT(rectangle1_heights[1824]), .RECT1_WEIGHT(rectangle1_weights[1824]), .RECT2_X(rectangle2_xs[1824]), .RECT2_Y(rectangle2_ys[1824]), .RECT2_WIDTH(rectangle2_widths[1824]), .RECT2_HEIGHT(rectangle2_heights[1824]), .RECT2_WEIGHT(rectangle2_weights[1824]), .RECT3_X(rectangle3_xs[1824]), .RECT3_Y(rectangle3_ys[1824]), .RECT3_WIDTH(rectangle3_widths[1824]), .RECT3_HEIGHT(rectangle3_heights[1824]), .RECT3_WEIGHT(rectangle3_weights[1824]), .FEAT_THRES(feature_thresholds[1824]), .FEAT_ABOVE(feature_aboves[1824]), .FEAT_BELOW(feature_belows[1824])) ac1824(.scan_win(scan_win1824), .scan_win_std_dev(scan_win_std_dev[1824]), .feature_accum(feature_accums[1824]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1825]), .RECT1_Y(rectangle1_ys[1825]), .RECT1_WIDTH(rectangle1_widths[1825]), .RECT1_HEIGHT(rectangle1_heights[1825]), .RECT1_WEIGHT(rectangle1_weights[1825]), .RECT2_X(rectangle2_xs[1825]), .RECT2_Y(rectangle2_ys[1825]), .RECT2_WIDTH(rectangle2_widths[1825]), .RECT2_HEIGHT(rectangle2_heights[1825]), .RECT2_WEIGHT(rectangle2_weights[1825]), .RECT3_X(rectangle3_xs[1825]), .RECT3_Y(rectangle3_ys[1825]), .RECT3_WIDTH(rectangle3_widths[1825]), .RECT3_HEIGHT(rectangle3_heights[1825]), .RECT3_WEIGHT(rectangle3_weights[1825]), .FEAT_THRES(feature_thresholds[1825]), .FEAT_ABOVE(feature_aboves[1825]), .FEAT_BELOW(feature_belows[1825])) ac1825(.scan_win(scan_win1825), .scan_win_std_dev(scan_win_std_dev[1825]), .feature_accum(feature_accums[1825]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1826]), .RECT1_Y(rectangle1_ys[1826]), .RECT1_WIDTH(rectangle1_widths[1826]), .RECT1_HEIGHT(rectangle1_heights[1826]), .RECT1_WEIGHT(rectangle1_weights[1826]), .RECT2_X(rectangle2_xs[1826]), .RECT2_Y(rectangle2_ys[1826]), .RECT2_WIDTH(rectangle2_widths[1826]), .RECT2_HEIGHT(rectangle2_heights[1826]), .RECT2_WEIGHT(rectangle2_weights[1826]), .RECT3_X(rectangle3_xs[1826]), .RECT3_Y(rectangle3_ys[1826]), .RECT3_WIDTH(rectangle3_widths[1826]), .RECT3_HEIGHT(rectangle3_heights[1826]), .RECT3_WEIGHT(rectangle3_weights[1826]), .FEAT_THRES(feature_thresholds[1826]), .FEAT_ABOVE(feature_aboves[1826]), .FEAT_BELOW(feature_belows[1826])) ac1826(.scan_win(scan_win1826), .scan_win_std_dev(scan_win_std_dev[1826]), .feature_accum(feature_accums[1826]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1827]), .RECT1_Y(rectangle1_ys[1827]), .RECT1_WIDTH(rectangle1_widths[1827]), .RECT1_HEIGHT(rectangle1_heights[1827]), .RECT1_WEIGHT(rectangle1_weights[1827]), .RECT2_X(rectangle2_xs[1827]), .RECT2_Y(rectangle2_ys[1827]), .RECT2_WIDTH(rectangle2_widths[1827]), .RECT2_HEIGHT(rectangle2_heights[1827]), .RECT2_WEIGHT(rectangle2_weights[1827]), .RECT3_X(rectangle3_xs[1827]), .RECT3_Y(rectangle3_ys[1827]), .RECT3_WIDTH(rectangle3_widths[1827]), .RECT3_HEIGHT(rectangle3_heights[1827]), .RECT3_WEIGHT(rectangle3_weights[1827]), .FEAT_THRES(feature_thresholds[1827]), .FEAT_ABOVE(feature_aboves[1827]), .FEAT_BELOW(feature_belows[1827])) ac1827(.scan_win(scan_win1827), .scan_win_std_dev(scan_win_std_dev[1827]), .feature_accum(feature_accums[1827]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1828]), .RECT1_Y(rectangle1_ys[1828]), .RECT1_WIDTH(rectangle1_widths[1828]), .RECT1_HEIGHT(rectangle1_heights[1828]), .RECT1_WEIGHT(rectangle1_weights[1828]), .RECT2_X(rectangle2_xs[1828]), .RECT2_Y(rectangle2_ys[1828]), .RECT2_WIDTH(rectangle2_widths[1828]), .RECT2_HEIGHT(rectangle2_heights[1828]), .RECT2_WEIGHT(rectangle2_weights[1828]), .RECT3_X(rectangle3_xs[1828]), .RECT3_Y(rectangle3_ys[1828]), .RECT3_WIDTH(rectangle3_widths[1828]), .RECT3_HEIGHT(rectangle3_heights[1828]), .RECT3_WEIGHT(rectangle3_weights[1828]), .FEAT_THRES(feature_thresholds[1828]), .FEAT_ABOVE(feature_aboves[1828]), .FEAT_BELOW(feature_belows[1828])) ac1828(.scan_win(scan_win1828), .scan_win_std_dev(scan_win_std_dev[1828]), .feature_accum(feature_accums[1828]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1829]), .RECT1_Y(rectangle1_ys[1829]), .RECT1_WIDTH(rectangle1_widths[1829]), .RECT1_HEIGHT(rectangle1_heights[1829]), .RECT1_WEIGHT(rectangle1_weights[1829]), .RECT2_X(rectangle2_xs[1829]), .RECT2_Y(rectangle2_ys[1829]), .RECT2_WIDTH(rectangle2_widths[1829]), .RECT2_HEIGHT(rectangle2_heights[1829]), .RECT2_WEIGHT(rectangle2_weights[1829]), .RECT3_X(rectangle3_xs[1829]), .RECT3_Y(rectangle3_ys[1829]), .RECT3_WIDTH(rectangle3_widths[1829]), .RECT3_HEIGHT(rectangle3_heights[1829]), .RECT3_WEIGHT(rectangle3_weights[1829]), .FEAT_THRES(feature_thresholds[1829]), .FEAT_ABOVE(feature_aboves[1829]), .FEAT_BELOW(feature_belows[1829])) ac1829(.scan_win(scan_win1829), .scan_win_std_dev(scan_win_std_dev[1829]), .feature_accum(feature_accums[1829]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1830]), .RECT1_Y(rectangle1_ys[1830]), .RECT1_WIDTH(rectangle1_widths[1830]), .RECT1_HEIGHT(rectangle1_heights[1830]), .RECT1_WEIGHT(rectangle1_weights[1830]), .RECT2_X(rectangle2_xs[1830]), .RECT2_Y(rectangle2_ys[1830]), .RECT2_WIDTH(rectangle2_widths[1830]), .RECT2_HEIGHT(rectangle2_heights[1830]), .RECT2_WEIGHT(rectangle2_weights[1830]), .RECT3_X(rectangle3_xs[1830]), .RECT3_Y(rectangle3_ys[1830]), .RECT3_WIDTH(rectangle3_widths[1830]), .RECT3_HEIGHT(rectangle3_heights[1830]), .RECT3_WEIGHT(rectangle3_weights[1830]), .FEAT_THRES(feature_thresholds[1830]), .FEAT_ABOVE(feature_aboves[1830]), .FEAT_BELOW(feature_belows[1830])) ac1830(.scan_win(scan_win1830), .scan_win_std_dev(scan_win_std_dev[1830]), .feature_accum(feature_accums[1830]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1831]), .RECT1_Y(rectangle1_ys[1831]), .RECT1_WIDTH(rectangle1_widths[1831]), .RECT1_HEIGHT(rectangle1_heights[1831]), .RECT1_WEIGHT(rectangle1_weights[1831]), .RECT2_X(rectangle2_xs[1831]), .RECT2_Y(rectangle2_ys[1831]), .RECT2_WIDTH(rectangle2_widths[1831]), .RECT2_HEIGHT(rectangle2_heights[1831]), .RECT2_WEIGHT(rectangle2_weights[1831]), .RECT3_X(rectangle3_xs[1831]), .RECT3_Y(rectangle3_ys[1831]), .RECT3_WIDTH(rectangle3_widths[1831]), .RECT3_HEIGHT(rectangle3_heights[1831]), .RECT3_WEIGHT(rectangle3_weights[1831]), .FEAT_THRES(feature_thresholds[1831]), .FEAT_ABOVE(feature_aboves[1831]), .FEAT_BELOW(feature_belows[1831])) ac1831(.scan_win(scan_win1831), .scan_win_std_dev(scan_win_std_dev[1831]), .feature_accum(feature_accums[1831]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1832]), .RECT1_Y(rectangle1_ys[1832]), .RECT1_WIDTH(rectangle1_widths[1832]), .RECT1_HEIGHT(rectangle1_heights[1832]), .RECT1_WEIGHT(rectangle1_weights[1832]), .RECT2_X(rectangle2_xs[1832]), .RECT2_Y(rectangle2_ys[1832]), .RECT2_WIDTH(rectangle2_widths[1832]), .RECT2_HEIGHT(rectangle2_heights[1832]), .RECT2_WEIGHT(rectangle2_weights[1832]), .RECT3_X(rectangle3_xs[1832]), .RECT3_Y(rectangle3_ys[1832]), .RECT3_WIDTH(rectangle3_widths[1832]), .RECT3_HEIGHT(rectangle3_heights[1832]), .RECT3_WEIGHT(rectangle3_weights[1832]), .FEAT_THRES(feature_thresholds[1832]), .FEAT_ABOVE(feature_aboves[1832]), .FEAT_BELOW(feature_belows[1832])) ac1832(.scan_win(scan_win1832), .scan_win_std_dev(scan_win_std_dev[1832]), .feature_accum(feature_accums[1832]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1833]), .RECT1_Y(rectangle1_ys[1833]), .RECT1_WIDTH(rectangle1_widths[1833]), .RECT1_HEIGHT(rectangle1_heights[1833]), .RECT1_WEIGHT(rectangle1_weights[1833]), .RECT2_X(rectangle2_xs[1833]), .RECT2_Y(rectangle2_ys[1833]), .RECT2_WIDTH(rectangle2_widths[1833]), .RECT2_HEIGHT(rectangle2_heights[1833]), .RECT2_WEIGHT(rectangle2_weights[1833]), .RECT3_X(rectangle3_xs[1833]), .RECT3_Y(rectangle3_ys[1833]), .RECT3_WIDTH(rectangle3_widths[1833]), .RECT3_HEIGHT(rectangle3_heights[1833]), .RECT3_WEIGHT(rectangle3_weights[1833]), .FEAT_THRES(feature_thresholds[1833]), .FEAT_ABOVE(feature_aboves[1833]), .FEAT_BELOW(feature_belows[1833])) ac1833(.scan_win(scan_win1833), .scan_win_std_dev(scan_win_std_dev[1833]), .feature_accum(feature_accums[1833]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1834]), .RECT1_Y(rectangle1_ys[1834]), .RECT1_WIDTH(rectangle1_widths[1834]), .RECT1_HEIGHT(rectangle1_heights[1834]), .RECT1_WEIGHT(rectangle1_weights[1834]), .RECT2_X(rectangle2_xs[1834]), .RECT2_Y(rectangle2_ys[1834]), .RECT2_WIDTH(rectangle2_widths[1834]), .RECT2_HEIGHT(rectangle2_heights[1834]), .RECT2_WEIGHT(rectangle2_weights[1834]), .RECT3_X(rectangle3_xs[1834]), .RECT3_Y(rectangle3_ys[1834]), .RECT3_WIDTH(rectangle3_widths[1834]), .RECT3_HEIGHT(rectangle3_heights[1834]), .RECT3_WEIGHT(rectangle3_weights[1834]), .FEAT_THRES(feature_thresholds[1834]), .FEAT_ABOVE(feature_aboves[1834]), .FEAT_BELOW(feature_belows[1834])) ac1834(.scan_win(scan_win1834), .scan_win_std_dev(scan_win_std_dev[1834]), .feature_accum(feature_accums[1834]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1835]), .RECT1_Y(rectangle1_ys[1835]), .RECT1_WIDTH(rectangle1_widths[1835]), .RECT1_HEIGHT(rectangle1_heights[1835]), .RECT1_WEIGHT(rectangle1_weights[1835]), .RECT2_X(rectangle2_xs[1835]), .RECT2_Y(rectangle2_ys[1835]), .RECT2_WIDTH(rectangle2_widths[1835]), .RECT2_HEIGHT(rectangle2_heights[1835]), .RECT2_WEIGHT(rectangle2_weights[1835]), .RECT3_X(rectangle3_xs[1835]), .RECT3_Y(rectangle3_ys[1835]), .RECT3_WIDTH(rectangle3_widths[1835]), .RECT3_HEIGHT(rectangle3_heights[1835]), .RECT3_WEIGHT(rectangle3_weights[1835]), .FEAT_THRES(feature_thresholds[1835]), .FEAT_ABOVE(feature_aboves[1835]), .FEAT_BELOW(feature_belows[1835])) ac1835(.scan_win(scan_win1835), .scan_win_std_dev(scan_win_std_dev[1835]), .feature_accum(feature_accums[1835]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1836]), .RECT1_Y(rectangle1_ys[1836]), .RECT1_WIDTH(rectangle1_widths[1836]), .RECT1_HEIGHT(rectangle1_heights[1836]), .RECT1_WEIGHT(rectangle1_weights[1836]), .RECT2_X(rectangle2_xs[1836]), .RECT2_Y(rectangle2_ys[1836]), .RECT2_WIDTH(rectangle2_widths[1836]), .RECT2_HEIGHT(rectangle2_heights[1836]), .RECT2_WEIGHT(rectangle2_weights[1836]), .RECT3_X(rectangle3_xs[1836]), .RECT3_Y(rectangle3_ys[1836]), .RECT3_WIDTH(rectangle3_widths[1836]), .RECT3_HEIGHT(rectangle3_heights[1836]), .RECT3_WEIGHT(rectangle3_weights[1836]), .FEAT_THRES(feature_thresholds[1836]), .FEAT_ABOVE(feature_aboves[1836]), .FEAT_BELOW(feature_belows[1836])) ac1836(.scan_win(scan_win1836), .scan_win_std_dev(scan_win_std_dev[1836]), .feature_accum(feature_accums[1836]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1837]), .RECT1_Y(rectangle1_ys[1837]), .RECT1_WIDTH(rectangle1_widths[1837]), .RECT1_HEIGHT(rectangle1_heights[1837]), .RECT1_WEIGHT(rectangle1_weights[1837]), .RECT2_X(rectangle2_xs[1837]), .RECT2_Y(rectangle2_ys[1837]), .RECT2_WIDTH(rectangle2_widths[1837]), .RECT2_HEIGHT(rectangle2_heights[1837]), .RECT2_WEIGHT(rectangle2_weights[1837]), .RECT3_X(rectangle3_xs[1837]), .RECT3_Y(rectangle3_ys[1837]), .RECT3_WIDTH(rectangle3_widths[1837]), .RECT3_HEIGHT(rectangle3_heights[1837]), .RECT3_WEIGHT(rectangle3_weights[1837]), .FEAT_THRES(feature_thresholds[1837]), .FEAT_ABOVE(feature_aboves[1837]), .FEAT_BELOW(feature_belows[1837])) ac1837(.scan_win(scan_win1837), .scan_win_std_dev(scan_win_std_dev[1837]), .feature_accum(feature_accums[1837]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1838]), .RECT1_Y(rectangle1_ys[1838]), .RECT1_WIDTH(rectangle1_widths[1838]), .RECT1_HEIGHT(rectangle1_heights[1838]), .RECT1_WEIGHT(rectangle1_weights[1838]), .RECT2_X(rectangle2_xs[1838]), .RECT2_Y(rectangle2_ys[1838]), .RECT2_WIDTH(rectangle2_widths[1838]), .RECT2_HEIGHT(rectangle2_heights[1838]), .RECT2_WEIGHT(rectangle2_weights[1838]), .RECT3_X(rectangle3_xs[1838]), .RECT3_Y(rectangle3_ys[1838]), .RECT3_WIDTH(rectangle3_widths[1838]), .RECT3_HEIGHT(rectangle3_heights[1838]), .RECT3_WEIGHT(rectangle3_weights[1838]), .FEAT_THRES(feature_thresholds[1838]), .FEAT_ABOVE(feature_aboves[1838]), .FEAT_BELOW(feature_belows[1838])) ac1838(.scan_win(scan_win1838), .scan_win_std_dev(scan_win_std_dev[1838]), .feature_accum(feature_accums[1838]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1839]), .RECT1_Y(rectangle1_ys[1839]), .RECT1_WIDTH(rectangle1_widths[1839]), .RECT1_HEIGHT(rectangle1_heights[1839]), .RECT1_WEIGHT(rectangle1_weights[1839]), .RECT2_X(rectangle2_xs[1839]), .RECT2_Y(rectangle2_ys[1839]), .RECT2_WIDTH(rectangle2_widths[1839]), .RECT2_HEIGHT(rectangle2_heights[1839]), .RECT2_WEIGHT(rectangle2_weights[1839]), .RECT3_X(rectangle3_xs[1839]), .RECT3_Y(rectangle3_ys[1839]), .RECT3_WIDTH(rectangle3_widths[1839]), .RECT3_HEIGHT(rectangle3_heights[1839]), .RECT3_WEIGHT(rectangle3_weights[1839]), .FEAT_THRES(feature_thresholds[1839]), .FEAT_ABOVE(feature_aboves[1839]), .FEAT_BELOW(feature_belows[1839])) ac1839(.scan_win(scan_win1839), .scan_win_std_dev(scan_win_std_dev[1839]), .feature_accum(feature_accums[1839]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1840]), .RECT1_Y(rectangle1_ys[1840]), .RECT1_WIDTH(rectangle1_widths[1840]), .RECT1_HEIGHT(rectangle1_heights[1840]), .RECT1_WEIGHT(rectangle1_weights[1840]), .RECT2_X(rectangle2_xs[1840]), .RECT2_Y(rectangle2_ys[1840]), .RECT2_WIDTH(rectangle2_widths[1840]), .RECT2_HEIGHT(rectangle2_heights[1840]), .RECT2_WEIGHT(rectangle2_weights[1840]), .RECT3_X(rectangle3_xs[1840]), .RECT3_Y(rectangle3_ys[1840]), .RECT3_WIDTH(rectangle3_widths[1840]), .RECT3_HEIGHT(rectangle3_heights[1840]), .RECT3_WEIGHT(rectangle3_weights[1840]), .FEAT_THRES(feature_thresholds[1840]), .FEAT_ABOVE(feature_aboves[1840]), .FEAT_BELOW(feature_belows[1840])) ac1840(.scan_win(scan_win1840), .scan_win_std_dev(scan_win_std_dev[1840]), .feature_accum(feature_accums[1840]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1841]), .RECT1_Y(rectangle1_ys[1841]), .RECT1_WIDTH(rectangle1_widths[1841]), .RECT1_HEIGHT(rectangle1_heights[1841]), .RECT1_WEIGHT(rectangle1_weights[1841]), .RECT2_X(rectangle2_xs[1841]), .RECT2_Y(rectangle2_ys[1841]), .RECT2_WIDTH(rectangle2_widths[1841]), .RECT2_HEIGHT(rectangle2_heights[1841]), .RECT2_WEIGHT(rectangle2_weights[1841]), .RECT3_X(rectangle3_xs[1841]), .RECT3_Y(rectangle3_ys[1841]), .RECT3_WIDTH(rectangle3_widths[1841]), .RECT3_HEIGHT(rectangle3_heights[1841]), .RECT3_WEIGHT(rectangle3_weights[1841]), .FEAT_THRES(feature_thresholds[1841]), .FEAT_ABOVE(feature_aboves[1841]), .FEAT_BELOW(feature_belows[1841])) ac1841(.scan_win(scan_win1841), .scan_win_std_dev(scan_win_std_dev[1841]), .feature_accum(feature_accums[1841]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1842]), .RECT1_Y(rectangle1_ys[1842]), .RECT1_WIDTH(rectangle1_widths[1842]), .RECT1_HEIGHT(rectangle1_heights[1842]), .RECT1_WEIGHT(rectangle1_weights[1842]), .RECT2_X(rectangle2_xs[1842]), .RECT2_Y(rectangle2_ys[1842]), .RECT2_WIDTH(rectangle2_widths[1842]), .RECT2_HEIGHT(rectangle2_heights[1842]), .RECT2_WEIGHT(rectangle2_weights[1842]), .RECT3_X(rectangle3_xs[1842]), .RECT3_Y(rectangle3_ys[1842]), .RECT3_WIDTH(rectangle3_widths[1842]), .RECT3_HEIGHT(rectangle3_heights[1842]), .RECT3_WEIGHT(rectangle3_weights[1842]), .FEAT_THRES(feature_thresholds[1842]), .FEAT_ABOVE(feature_aboves[1842]), .FEAT_BELOW(feature_belows[1842])) ac1842(.scan_win(scan_win1842), .scan_win_std_dev(scan_win_std_dev[1842]), .feature_accum(feature_accums[1842]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1843]), .RECT1_Y(rectangle1_ys[1843]), .RECT1_WIDTH(rectangle1_widths[1843]), .RECT1_HEIGHT(rectangle1_heights[1843]), .RECT1_WEIGHT(rectangle1_weights[1843]), .RECT2_X(rectangle2_xs[1843]), .RECT2_Y(rectangle2_ys[1843]), .RECT2_WIDTH(rectangle2_widths[1843]), .RECT2_HEIGHT(rectangle2_heights[1843]), .RECT2_WEIGHT(rectangle2_weights[1843]), .RECT3_X(rectangle3_xs[1843]), .RECT3_Y(rectangle3_ys[1843]), .RECT3_WIDTH(rectangle3_widths[1843]), .RECT3_HEIGHT(rectangle3_heights[1843]), .RECT3_WEIGHT(rectangle3_weights[1843]), .FEAT_THRES(feature_thresholds[1843]), .FEAT_ABOVE(feature_aboves[1843]), .FEAT_BELOW(feature_belows[1843])) ac1843(.scan_win(scan_win1843), .scan_win_std_dev(scan_win_std_dev[1843]), .feature_accum(feature_accums[1843]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1844]), .RECT1_Y(rectangle1_ys[1844]), .RECT1_WIDTH(rectangle1_widths[1844]), .RECT1_HEIGHT(rectangle1_heights[1844]), .RECT1_WEIGHT(rectangle1_weights[1844]), .RECT2_X(rectangle2_xs[1844]), .RECT2_Y(rectangle2_ys[1844]), .RECT2_WIDTH(rectangle2_widths[1844]), .RECT2_HEIGHT(rectangle2_heights[1844]), .RECT2_WEIGHT(rectangle2_weights[1844]), .RECT3_X(rectangle3_xs[1844]), .RECT3_Y(rectangle3_ys[1844]), .RECT3_WIDTH(rectangle3_widths[1844]), .RECT3_HEIGHT(rectangle3_heights[1844]), .RECT3_WEIGHT(rectangle3_weights[1844]), .FEAT_THRES(feature_thresholds[1844]), .FEAT_ABOVE(feature_aboves[1844]), .FEAT_BELOW(feature_belows[1844])) ac1844(.scan_win(scan_win1844), .scan_win_std_dev(scan_win_std_dev[1844]), .feature_accum(feature_accums[1844]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1845]), .RECT1_Y(rectangle1_ys[1845]), .RECT1_WIDTH(rectangle1_widths[1845]), .RECT1_HEIGHT(rectangle1_heights[1845]), .RECT1_WEIGHT(rectangle1_weights[1845]), .RECT2_X(rectangle2_xs[1845]), .RECT2_Y(rectangle2_ys[1845]), .RECT2_WIDTH(rectangle2_widths[1845]), .RECT2_HEIGHT(rectangle2_heights[1845]), .RECT2_WEIGHT(rectangle2_weights[1845]), .RECT3_X(rectangle3_xs[1845]), .RECT3_Y(rectangle3_ys[1845]), .RECT3_WIDTH(rectangle3_widths[1845]), .RECT3_HEIGHT(rectangle3_heights[1845]), .RECT3_WEIGHT(rectangle3_weights[1845]), .FEAT_THRES(feature_thresholds[1845]), .FEAT_ABOVE(feature_aboves[1845]), .FEAT_BELOW(feature_belows[1845])) ac1845(.scan_win(scan_win1845), .scan_win_std_dev(scan_win_std_dev[1845]), .feature_accum(feature_accums[1845]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1846]), .RECT1_Y(rectangle1_ys[1846]), .RECT1_WIDTH(rectangle1_widths[1846]), .RECT1_HEIGHT(rectangle1_heights[1846]), .RECT1_WEIGHT(rectangle1_weights[1846]), .RECT2_X(rectangle2_xs[1846]), .RECT2_Y(rectangle2_ys[1846]), .RECT2_WIDTH(rectangle2_widths[1846]), .RECT2_HEIGHT(rectangle2_heights[1846]), .RECT2_WEIGHT(rectangle2_weights[1846]), .RECT3_X(rectangle3_xs[1846]), .RECT3_Y(rectangle3_ys[1846]), .RECT3_WIDTH(rectangle3_widths[1846]), .RECT3_HEIGHT(rectangle3_heights[1846]), .RECT3_WEIGHT(rectangle3_weights[1846]), .FEAT_THRES(feature_thresholds[1846]), .FEAT_ABOVE(feature_aboves[1846]), .FEAT_BELOW(feature_belows[1846])) ac1846(.scan_win(scan_win1846), .scan_win_std_dev(scan_win_std_dev[1846]), .feature_accum(feature_accums[1846]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1847]), .RECT1_Y(rectangle1_ys[1847]), .RECT1_WIDTH(rectangle1_widths[1847]), .RECT1_HEIGHT(rectangle1_heights[1847]), .RECT1_WEIGHT(rectangle1_weights[1847]), .RECT2_X(rectangle2_xs[1847]), .RECT2_Y(rectangle2_ys[1847]), .RECT2_WIDTH(rectangle2_widths[1847]), .RECT2_HEIGHT(rectangle2_heights[1847]), .RECT2_WEIGHT(rectangle2_weights[1847]), .RECT3_X(rectangle3_xs[1847]), .RECT3_Y(rectangle3_ys[1847]), .RECT3_WIDTH(rectangle3_widths[1847]), .RECT3_HEIGHT(rectangle3_heights[1847]), .RECT3_WEIGHT(rectangle3_weights[1847]), .FEAT_THRES(feature_thresholds[1847]), .FEAT_ABOVE(feature_aboves[1847]), .FEAT_BELOW(feature_belows[1847])) ac1847(.scan_win(scan_win1847), .scan_win_std_dev(scan_win_std_dev[1847]), .feature_accum(feature_accums[1847]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1848]), .RECT1_Y(rectangle1_ys[1848]), .RECT1_WIDTH(rectangle1_widths[1848]), .RECT1_HEIGHT(rectangle1_heights[1848]), .RECT1_WEIGHT(rectangle1_weights[1848]), .RECT2_X(rectangle2_xs[1848]), .RECT2_Y(rectangle2_ys[1848]), .RECT2_WIDTH(rectangle2_widths[1848]), .RECT2_HEIGHT(rectangle2_heights[1848]), .RECT2_WEIGHT(rectangle2_weights[1848]), .RECT3_X(rectangle3_xs[1848]), .RECT3_Y(rectangle3_ys[1848]), .RECT3_WIDTH(rectangle3_widths[1848]), .RECT3_HEIGHT(rectangle3_heights[1848]), .RECT3_WEIGHT(rectangle3_weights[1848]), .FEAT_THRES(feature_thresholds[1848]), .FEAT_ABOVE(feature_aboves[1848]), .FEAT_BELOW(feature_belows[1848])) ac1848(.scan_win(scan_win1848), .scan_win_std_dev(scan_win_std_dev[1848]), .feature_accum(feature_accums[1848]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1849]), .RECT1_Y(rectangle1_ys[1849]), .RECT1_WIDTH(rectangle1_widths[1849]), .RECT1_HEIGHT(rectangle1_heights[1849]), .RECT1_WEIGHT(rectangle1_weights[1849]), .RECT2_X(rectangle2_xs[1849]), .RECT2_Y(rectangle2_ys[1849]), .RECT2_WIDTH(rectangle2_widths[1849]), .RECT2_HEIGHT(rectangle2_heights[1849]), .RECT2_WEIGHT(rectangle2_weights[1849]), .RECT3_X(rectangle3_xs[1849]), .RECT3_Y(rectangle3_ys[1849]), .RECT3_WIDTH(rectangle3_widths[1849]), .RECT3_HEIGHT(rectangle3_heights[1849]), .RECT3_WEIGHT(rectangle3_weights[1849]), .FEAT_THRES(feature_thresholds[1849]), .FEAT_ABOVE(feature_aboves[1849]), .FEAT_BELOW(feature_belows[1849])) ac1849(.scan_win(scan_win1849), .scan_win_std_dev(scan_win_std_dev[1849]), .feature_accum(feature_accums[1849]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1850]), .RECT1_Y(rectangle1_ys[1850]), .RECT1_WIDTH(rectangle1_widths[1850]), .RECT1_HEIGHT(rectangle1_heights[1850]), .RECT1_WEIGHT(rectangle1_weights[1850]), .RECT2_X(rectangle2_xs[1850]), .RECT2_Y(rectangle2_ys[1850]), .RECT2_WIDTH(rectangle2_widths[1850]), .RECT2_HEIGHT(rectangle2_heights[1850]), .RECT2_WEIGHT(rectangle2_weights[1850]), .RECT3_X(rectangle3_xs[1850]), .RECT3_Y(rectangle3_ys[1850]), .RECT3_WIDTH(rectangle3_widths[1850]), .RECT3_HEIGHT(rectangle3_heights[1850]), .RECT3_WEIGHT(rectangle3_weights[1850]), .FEAT_THRES(feature_thresholds[1850]), .FEAT_ABOVE(feature_aboves[1850]), .FEAT_BELOW(feature_belows[1850])) ac1850(.scan_win(scan_win1850), .scan_win_std_dev(scan_win_std_dev[1850]), .feature_accum(feature_accums[1850]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1851]), .RECT1_Y(rectangle1_ys[1851]), .RECT1_WIDTH(rectangle1_widths[1851]), .RECT1_HEIGHT(rectangle1_heights[1851]), .RECT1_WEIGHT(rectangle1_weights[1851]), .RECT2_X(rectangle2_xs[1851]), .RECT2_Y(rectangle2_ys[1851]), .RECT2_WIDTH(rectangle2_widths[1851]), .RECT2_HEIGHT(rectangle2_heights[1851]), .RECT2_WEIGHT(rectangle2_weights[1851]), .RECT3_X(rectangle3_xs[1851]), .RECT3_Y(rectangle3_ys[1851]), .RECT3_WIDTH(rectangle3_widths[1851]), .RECT3_HEIGHT(rectangle3_heights[1851]), .RECT3_WEIGHT(rectangle3_weights[1851]), .FEAT_THRES(feature_thresholds[1851]), .FEAT_ABOVE(feature_aboves[1851]), .FEAT_BELOW(feature_belows[1851])) ac1851(.scan_win(scan_win1851), .scan_win_std_dev(scan_win_std_dev[1851]), .feature_accum(feature_accums[1851]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1852]), .RECT1_Y(rectangle1_ys[1852]), .RECT1_WIDTH(rectangle1_widths[1852]), .RECT1_HEIGHT(rectangle1_heights[1852]), .RECT1_WEIGHT(rectangle1_weights[1852]), .RECT2_X(rectangle2_xs[1852]), .RECT2_Y(rectangle2_ys[1852]), .RECT2_WIDTH(rectangle2_widths[1852]), .RECT2_HEIGHT(rectangle2_heights[1852]), .RECT2_WEIGHT(rectangle2_weights[1852]), .RECT3_X(rectangle3_xs[1852]), .RECT3_Y(rectangle3_ys[1852]), .RECT3_WIDTH(rectangle3_widths[1852]), .RECT3_HEIGHT(rectangle3_heights[1852]), .RECT3_WEIGHT(rectangle3_weights[1852]), .FEAT_THRES(feature_thresholds[1852]), .FEAT_ABOVE(feature_aboves[1852]), .FEAT_BELOW(feature_belows[1852])) ac1852(.scan_win(scan_win1852), .scan_win_std_dev(scan_win_std_dev[1852]), .feature_accum(feature_accums[1852]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1853]), .RECT1_Y(rectangle1_ys[1853]), .RECT1_WIDTH(rectangle1_widths[1853]), .RECT1_HEIGHT(rectangle1_heights[1853]), .RECT1_WEIGHT(rectangle1_weights[1853]), .RECT2_X(rectangle2_xs[1853]), .RECT2_Y(rectangle2_ys[1853]), .RECT2_WIDTH(rectangle2_widths[1853]), .RECT2_HEIGHT(rectangle2_heights[1853]), .RECT2_WEIGHT(rectangle2_weights[1853]), .RECT3_X(rectangle3_xs[1853]), .RECT3_Y(rectangle3_ys[1853]), .RECT3_WIDTH(rectangle3_widths[1853]), .RECT3_HEIGHT(rectangle3_heights[1853]), .RECT3_WEIGHT(rectangle3_weights[1853]), .FEAT_THRES(feature_thresholds[1853]), .FEAT_ABOVE(feature_aboves[1853]), .FEAT_BELOW(feature_belows[1853])) ac1853(.scan_win(scan_win1853), .scan_win_std_dev(scan_win_std_dev[1853]), .feature_accum(feature_accums[1853]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1854]), .RECT1_Y(rectangle1_ys[1854]), .RECT1_WIDTH(rectangle1_widths[1854]), .RECT1_HEIGHT(rectangle1_heights[1854]), .RECT1_WEIGHT(rectangle1_weights[1854]), .RECT2_X(rectangle2_xs[1854]), .RECT2_Y(rectangle2_ys[1854]), .RECT2_WIDTH(rectangle2_widths[1854]), .RECT2_HEIGHT(rectangle2_heights[1854]), .RECT2_WEIGHT(rectangle2_weights[1854]), .RECT3_X(rectangle3_xs[1854]), .RECT3_Y(rectangle3_ys[1854]), .RECT3_WIDTH(rectangle3_widths[1854]), .RECT3_HEIGHT(rectangle3_heights[1854]), .RECT3_WEIGHT(rectangle3_weights[1854]), .FEAT_THRES(feature_thresholds[1854]), .FEAT_ABOVE(feature_aboves[1854]), .FEAT_BELOW(feature_belows[1854])) ac1854(.scan_win(scan_win1854), .scan_win_std_dev(scan_win_std_dev[1854]), .feature_accum(feature_accums[1854]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1855]), .RECT1_Y(rectangle1_ys[1855]), .RECT1_WIDTH(rectangle1_widths[1855]), .RECT1_HEIGHT(rectangle1_heights[1855]), .RECT1_WEIGHT(rectangle1_weights[1855]), .RECT2_X(rectangle2_xs[1855]), .RECT2_Y(rectangle2_ys[1855]), .RECT2_WIDTH(rectangle2_widths[1855]), .RECT2_HEIGHT(rectangle2_heights[1855]), .RECT2_WEIGHT(rectangle2_weights[1855]), .RECT3_X(rectangle3_xs[1855]), .RECT3_Y(rectangle3_ys[1855]), .RECT3_WIDTH(rectangle3_widths[1855]), .RECT3_HEIGHT(rectangle3_heights[1855]), .RECT3_WEIGHT(rectangle3_weights[1855]), .FEAT_THRES(feature_thresholds[1855]), .FEAT_ABOVE(feature_aboves[1855]), .FEAT_BELOW(feature_belows[1855])) ac1855(.scan_win(scan_win1855), .scan_win_std_dev(scan_win_std_dev[1855]), .feature_accum(feature_accums[1855]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1856]), .RECT1_Y(rectangle1_ys[1856]), .RECT1_WIDTH(rectangle1_widths[1856]), .RECT1_HEIGHT(rectangle1_heights[1856]), .RECT1_WEIGHT(rectangle1_weights[1856]), .RECT2_X(rectangle2_xs[1856]), .RECT2_Y(rectangle2_ys[1856]), .RECT2_WIDTH(rectangle2_widths[1856]), .RECT2_HEIGHT(rectangle2_heights[1856]), .RECT2_WEIGHT(rectangle2_weights[1856]), .RECT3_X(rectangle3_xs[1856]), .RECT3_Y(rectangle3_ys[1856]), .RECT3_WIDTH(rectangle3_widths[1856]), .RECT3_HEIGHT(rectangle3_heights[1856]), .RECT3_WEIGHT(rectangle3_weights[1856]), .FEAT_THRES(feature_thresholds[1856]), .FEAT_ABOVE(feature_aboves[1856]), .FEAT_BELOW(feature_belows[1856])) ac1856(.scan_win(scan_win1856), .scan_win_std_dev(scan_win_std_dev[1856]), .feature_accum(feature_accums[1856]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1857]), .RECT1_Y(rectangle1_ys[1857]), .RECT1_WIDTH(rectangle1_widths[1857]), .RECT1_HEIGHT(rectangle1_heights[1857]), .RECT1_WEIGHT(rectangle1_weights[1857]), .RECT2_X(rectangle2_xs[1857]), .RECT2_Y(rectangle2_ys[1857]), .RECT2_WIDTH(rectangle2_widths[1857]), .RECT2_HEIGHT(rectangle2_heights[1857]), .RECT2_WEIGHT(rectangle2_weights[1857]), .RECT3_X(rectangle3_xs[1857]), .RECT3_Y(rectangle3_ys[1857]), .RECT3_WIDTH(rectangle3_widths[1857]), .RECT3_HEIGHT(rectangle3_heights[1857]), .RECT3_WEIGHT(rectangle3_weights[1857]), .FEAT_THRES(feature_thresholds[1857]), .FEAT_ABOVE(feature_aboves[1857]), .FEAT_BELOW(feature_belows[1857])) ac1857(.scan_win(scan_win1857), .scan_win_std_dev(scan_win_std_dev[1857]), .feature_accum(feature_accums[1857]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1858]), .RECT1_Y(rectangle1_ys[1858]), .RECT1_WIDTH(rectangle1_widths[1858]), .RECT1_HEIGHT(rectangle1_heights[1858]), .RECT1_WEIGHT(rectangle1_weights[1858]), .RECT2_X(rectangle2_xs[1858]), .RECT2_Y(rectangle2_ys[1858]), .RECT2_WIDTH(rectangle2_widths[1858]), .RECT2_HEIGHT(rectangle2_heights[1858]), .RECT2_WEIGHT(rectangle2_weights[1858]), .RECT3_X(rectangle3_xs[1858]), .RECT3_Y(rectangle3_ys[1858]), .RECT3_WIDTH(rectangle3_widths[1858]), .RECT3_HEIGHT(rectangle3_heights[1858]), .RECT3_WEIGHT(rectangle3_weights[1858]), .FEAT_THRES(feature_thresholds[1858]), .FEAT_ABOVE(feature_aboves[1858]), .FEAT_BELOW(feature_belows[1858])) ac1858(.scan_win(scan_win1858), .scan_win_std_dev(scan_win_std_dev[1858]), .feature_accum(feature_accums[1858]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1859]), .RECT1_Y(rectangle1_ys[1859]), .RECT1_WIDTH(rectangle1_widths[1859]), .RECT1_HEIGHT(rectangle1_heights[1859]), .RECT1_WEIGHT(rectangle1_weights[1859]), .RECT2_X(rectangle2_xs[1859]), .RECT2_Y(rectangle2_ys[1859]), .RECT2_WIDTH(rectangle2_widths[1859]), .RECT2_HEIGHT(rectangle2_heights[1859]), .RECT2_WEIGHT(rectangle2_weights[1859]), .RECT3_X(rectangle3_xs[1859]), .RECT3_Y(rectangle3_ys[1859]), .RECT3_WIDTH(rectangle3_widths[1859]), .RECT3_HEIGHT(rectangle3_heights[1859]), .RECT3_WEIGHT(rectangle3_weights[1859]), .FEAT_THRES(feature_thresholds[1859]), .FEAT_ABOVE(feature_aboves[1859]), .FEAT_BELOW(feature_belows[1859])) ac1859(.scan_win(scan_win1859), .scan_win_std_dev(scan_win_std_dev[1859]), .feature_accum(feature_accums[1859]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1860]), .RECT1_Y(rectangle1_ys[1860]), .RECT1_WIDTH(rectangle1_widths[1860]), .RECT1_HEIGHT(rectangle1_heights[1860]), .RECT1_WEIGHT(rectangle1_weights[1860]), .RECT2_X(rectangle2_xs[1860]), .RECT2_Y(rectangle2_ys[1860]), .RECT2_WIDTH(rectangle2_widths[1860]), .RECT2_HEIGHT(rectangle2_heights[1860]), .RECT2_WEIGHT(rectangle2_weights[1860]), .RECT3_X(rectangle3_xs[1860]), .RECT3_Y(rectangle3_ys[1860]), .RECT3_WIDTH(rectangle3_widths[1860]), .RECT3_HEIGHT(rectangle3_heights[1860]), .RECT3_WEIGHT(rectangle3_weights[1860]), .FEAT_THRES(feature_thresholds[1860]), .FEAT_ABOVE(feature_aboves[1860]), .FEAT_BELOW(feature_belows[1860])) ac1860(.scan_win(scan_win1860), .scan_win_std_dev(scan_win_std_dev[1860]), .feature_accum(feature_accums[1860]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1861]), .RECT1_Y(rectangle1_ys[1861]), .RECT1_WIDTH(rectangle1_widths[1861]), .RECT1_HEIGHT(rectangle1_heights[1861]), .RECT1_WEIGHT(rectangle1_weights[1861]), .RECT2_X(rectangle2_xs[1861]), .RECT2_Y(rectangle2_ys[1861]), .RECT2_WIDTH(rectangle2_widths[1861]), .RECT2_HEIGHT(rectangle2_heights[1861]), .RECT2_WEIGHT(rectangle2_weights[1861]), .RECT3_X(rectangle3_xs[1861]), .RECT3_Y(rectangle3_ys[1861]), .RECT3_WIDTH(rectangle3_widths[1861]), .RECT3_HEIGHT(rectangle3_heights[1861]), .RECT3_WEIGHT(rectangle3_weights[1861]), .FEAT_THRES(feature_thresholds[1861]), .FEAT_ABOVE(feature_aboves[1861]), .FEAT_BELOW(feature_belows[1861])) ac1861(.scan_win(scan_win1861), .scan_win_std_dev(scan_win_std_dev[1861]), .feature_accum(feature_accums[1861]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1862]), .RECT1_Y(rectangle1_ys[1862]), .RECT1_WIDTH(rectangle1_widths[1862]), .RECT1_HEIGHT(rectangle1_heights[1862]), .RECT1_WEIGHT(rectangle1_weights[1862]), .RECT2_X(rectangle2_xs[1862]), .RECT2_Y(rectangle2_ys[1862]), .RECT2_WIDTH(rectangle2_widths[1862]), .RECT2_HEIGHT(rectangle2_heights[1862]), .RECT2_WEIGHT(rectangle2_weights[1862]), .RECT3_X(rectangle3_xs[1862]), .RECT3_Y(rectangle3_ys[1862]), .RECT3_WIDTH(rectangle3_widths[1862]), .RECT3_HEIGHT(rectangle3_heights[1862]), .RECT3_WEIGHT(rectangle3_weights[1862]), .FEAT_THRES(feature_thresholds[1862]), .FEAT_ABOVE(feature_aboves[1862]), .FEAT_BELOW(feature_belows[1862])) ac1862(.scan_win(scan_win1862), .scan_win_std_dev(scan_win_std_dev[1862]), .feature_accum(feature_accums[1862]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1863]), .RECT1_Y(rectangle1_ys[1863]), .RECT1_WIDTH(rectangle1_widths[1863]), .RECT1_HEIGHT(rectangle1_heights[1863]), .RECT1_WEIGHT(rectangle1_weights[1863]), .RECT2_X(rectangle2_xs[1863]), .RECT2_Y(rectangle2_ys[1863]), .RECT2_WIDTH(rectangle2_widths[1863]), .RECT2_HEIGHT(rectangle2_heights[1863]), .RECT2_WEIGHT(rectangle2_weights[1863]), .RECT3_X(rectangle3_xs[1863]), .RECT3_Y(rectangle3_ys[1863]), .RECT3_WIDTH(rectangle3_widths[1863]), .RECT3_HEIGHT(rectangle3_heights[1863]), .RECT3_WEIGHT(rectangle3_weights[1863]), .FEAT_THRES(feature_thresholds[1863]), .FEAT_ABOVE(feature_aboves[1863]), .FEAT_BELOW(feature_belows[1863])) ac1863(.scan_win(scan_win1863), .scan_win_std_dev(scan_win_std_dev[1863]), .feature_accum(feature_accums[1863]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1864]), .RECT1_Y(rectangle1_ys[1864]), .RECT1_WIDTH(rectangle1_widths[1864]), .RECT1_HEIGHT(rectangle1_heights[1864]), .RECT1_WEIGHT(rectangle1_weights[1864]), .RECT2_X(rectangle2_xs[1864]), .RECT2_Y(rectangle2_ys[1864]), .RECT2_WIDTH(rectangle2_widths[1864]), .RECT2_HEIGHT(rectangle2_heights[1864]), .RECT2_WEIGHT(rectangle2_weights[1864]), .RECT3_X(rectangle3_xs[1864]), .RECT3_Y(rectangle3_ys[1864]), .RECT3_WIDTH(rectangle3_widths[1864]), .RECT3_HEIGHT(rectangle3_heights[1864]), .RECT3_WEIGHT(rectangle3_weights[1864]), .FEAT_THRES(feature_thresholds[1864]), .FEAT_ABOVE(feature_aboves[1864]), .FEAT_BELOW(feature_belows[1864])) ac1864(.scan_win(scan_win1864), .scan_win_std_dev(scan_win_std_dev[1864]), .feature_accum(feature_accums[1864]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1865]), .RECT1_Y(rectangle1_ys[1865]), .RECT1_WIDTH(rectangle1_widths[1865]), .RECT1_HEIGHT(rectangle1_heights[1865]), .RECT1_WEIGHT(rectangle1_weights[1865]), .RECT2_X(rectangle2_xs[1865]), .RECT2_Y(rectangle2_ys[1865]), .RECT2_WIDTH(rectangle2_widths[1865]), .RECT2_HEIGHT(rectangle2_heights[1865]), .RECT2_WEIGHT(rectangle2_weights[1865]), .RECT3_X(rectangle3_xs[1865]), .RECT3_Y(rectangle3_ys[1865]), .RECT3_WIDTH(rectangle3_widths[1865]), .RECT3_HEIGHT(rectangle3_heights[1865]), .RECT3_WEIGHT(rectangle3_weights[1865]), .FEAT_THRES(feature_thresholds[1865]), .FEAT_ABOVE(feature_aboves[1865]), .FEAT_BELOW(feature_belows[1865])) ac1865(.scan_win(scan_win1865), .scan_win_std_dev(scan_win_std_dev[1865]), .feature_accum(feature_accums[1865]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1866]), .RECT1_Y(rectangle1_ys[1866]), .RECT1_WIDTH(rectangle1_widths[1866]), .RECT1_HEIGHT(rectangle1_heights[1866]), .RECT1_WEIGHT(rectangle1_weights[1866]), .RECT2_X(rectangle2_xs[1866]), .RECT2_Y(rectangle2_ys[1866]), .RECT2_WIDTH(rectangle2_widths[1866]), .RECT2_HEIGHT(rectangle2_heights[1866]), .RECT2_WEIGHT(rectangle2_weights[1866]), .RECT3_X(rectangle3_xs[1866]), .RECT3_Y(rectangle3_ys[1866]), .RECT3_WIDTH(rectangle3_widths[1866]), .RECT3_HEIGHT(rectangle3_heights[1866]), .RECT3_WEIGHT(rectangle3_weights[1866]), .FEAT_THRES(feature_thresholds[1866]), .FEAT_ABOVE(feature_aboves[1866]), .FEAT_BELOW(feature_belows[1866])) ac1866(.scan_win(scan_win1866), .scan_win_std_dev(scan_win_std_dev[1866]), .feature_accum(feature_accums[1866]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1867]), .RECT1_Y(rectangle1_ys[1867]), .RECT1_WIDTH(rectangle1_widths[1867]), .RECT1_HEIGHT(rectangle1_heights[1867]), .RECT1_WEIGHT(rectangle1_weights[1867]), .RECT2_X(rectangle2_xs[1867]), .RECT2_Y(rectangle2_ys[1867]), .RECT2_WIDTH(rectangle2_widths[1867]), .RECT2_HEIGHT(rectangle2_heights[1867]), .RECT2_WEIGHT(rectangle2_weights[1867]), .RECT3_X(rectangle3_xs[1867]), .RECT3_Y(rectangle3_ys[1867]), .RECT3_WIDTH(rectangle3_widths[1867]), .RECT3_HEIGHT(rectangle3_heights[1867]), .RECT3_WEIGHT(rectangle3_weights[1867]), .FEAT_THRES(feature_thresholds[1867]), .FEAT_ABOVE(feature_aboves[1867]), .FEAT_BELOW(feature_belows[1867])) ac1867(.scan_win(scan_win1867), .scan_win_std_dev(scan_win_std_dev[1867]), .feature_accum(feature_accums[1867]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1868]), .RECT1_Y(rectangle1_ys[1868]), .RECT1_WIDTH(rectangle1_widths[1868]), .RECT1_HEIGHT(rectangle1_heights[1868]), .RECT1_WEIGHT(rectangle1_weights[1868]), .RECT2_X(rectangle2_xs[1868]), .RECT2_Y(rectangle2_ys[1868]), .RECT2_WIDTH(rectangle2_widths[1868]), .RECT2_HEIGHT(rectangle2_heights[1868]), .RECT2_WEIGHT(rectangle2_weights[1868]), .RECT3_X(rectangle3_xs[1868]), .RECT3_Y(rectangle3_ys[1868]), .RECT3_WIDTH(rectangle3_widths[1868]), .RECT3_HEIGHT(rectangle3_heights[1868]), .RECT3_WEIGHT(rectangle3_weights[1868]), .FEAT_THRES(feature_thresholds[1868]), .FEAT_ABOVE(feature_aboves[1868]), .FEAT_BELOW(feature_belows[1868])) ac1868(.scan_win(scan_win1868), .scan_win_std_dev(scan_win_std_dev[1868]), .feature_accum(feature_accums[1868]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1869]), .RECT1_Y(rectangle1_ys[1869]), .RECT1_WIDTH(rectangle1_widths[1869]), .RECT1_HEIGHT(rectangle1_heights[1869]), .RECT1_WEIGHT(rectangle1_weights[1869]), .RECT2_X(rectangle2_xs[1869]), .RECT2_Y(rectangle2_ys[1869]), .RECT2_WIDTH(rectangle2_widths[1869]), .RECT2_HEIGHT(rectangle2_heights[1869]), .RECT2_WEIGHT(rectangle2_weights[1869]), .RECT3_X(rectangle3_xs[1869]), .RECT3_Y(rectangle3_ys[1869]), .RECT3_WIDTH(rectangle3_widths[1869]), .RECT3_HEIGHT(rectangle3_heights[1869]), .RECT3_WEIGHT(rectangle3_weights[1869]), .FEAT_THRES(feature_thresholds[1869]), .FEAT_ABOVE(feature_aboves[1869]), .FEAT_BELOW(feature_belows[1869])) ac1869(.scan_win(scan_win1869), .scan_win_std_dev(scan_win_std_dev[1869]), .feature_accum(feature_accums[1869]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1870]), .RECT1_Y(rectangle1_ys[1870]), .RECT1_WIDTH(rectangle1_widths[1870]), .RECT1_HEIGHT(rectangle1_heights[1870]), .RECT1_WEIGHT(rectangle1_weights[1870]), .RECT2_X(rectangle2_xs[1870]), .RECT2_Y(rectangle2_ys[1870]), .RECT2_WIDTH(rectangle2_widths[1870]), .RECT2_HEIGHT(rectangle2_heights[1870]), .RECT2_WEIGHT(rectangle2_weights[1870]), .RECT3_X(rectangle3_xs[1870]), .RECT3_Y(rectangle3_ys[1870]), .RECT3_WIDTH(rectangle3_widths[1870]), .RECT3_HEIGHT(rectangle3_heights[1870]), .RECT3_WEIGHT(rectangle3_weights[1870]), .FEAT_THRES(feature_thresholds[1870]), .FEAT_ABOVE(feature_aboves[1870]), .FEAT_BELOW(feature_belows[1870])) ac1870(.scan_win(scan_win1870), .scan_win_std_dev(scan_win_std_dev[1870]), .feature_accum(feature_accums[1870]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1871]), .RECT1_Y(rectangle1_ys[1871]), .RECT1_WIDTH(rectangle1_widths[1871]), .RECT1_HEIGHT(rectangle1_heights[1871]), .RECT1_WEIGHT(rectangle1_weights[1871]), .RECT2_X(rectangle2_xs[1871]), .RECT2_Y(rectangle2_ys[1871]), .RECT2_WIDTH(rectangle2_widths[1871]), .RECT2_HEIGHT(rectangle2_heights[1871]), .RECT2_WEIGHT(rectangle2_weights[1871]), .RECT3_X(rectangle3_xs[1871]), .RECT3_Y(rectangle3_ys[1871]), .RECT3_WIDTH(rectangle3_widths[1871]), .RECT3_HEIGHT(rectangle3_heights[1871]), .RECT3_WEIGHT(rectangle3_weights[1871]), .FEAT_THRES(feature_thresholds[1871]), .FEAT_ABOVE(feature_aboves[1871]), .FEAT_BELOW(feature_belows[1871])) ac1871(.scan_win(scan_win1871), .scan_win_std_dev(scan_win_std_dev[1871]), .feature_accum(feature_accums[1871]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1872]), .RECT1_Y(rectangle1_ys[1872]), .RECT1_WIDTH(rectangle1_widths[1872]), .RECT1_HEIGHT(rectangle1_heights[1872]), .RECT1_WEIGHT(rectangle1_weights[1872]), .RECT2_X(rectangle2_xs[1872]), .RECT2_Y(rectangle2_ys[1872]), .RECT2_WIDTH(rectangle2_widths[1872]), .RECT2_HEIGHT(rectangle2_heights[1872]), .RECT2_WEIGHT(rectangle2_weights[1872]), .RECT3_X(rectangle3_xs[1872]), .RECT3_Y(rectangle3_ys[1872]), .RECT3_WIDTH(rectangle3_widths[1872]), .RECT3_HEIGHT(rectangle3_heights[1872]), .RECT3_WEIGHT(rectangle3_weights[1872]), .FEAT_THRES(feature_thresholds[1872]), .FEAT_ABOVE(feature_aboves[1872]), .FEAT_BELOW(feature_belows[1872])) ac1872(.scan_win(scan_win1872), .scan_win_std_dev(scan_win_std_dev[1872]), .feature_accum(feature_accums[1872]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1873]), .RECT1_Y(rectangle1_ys[1873]), .RECT1_WIDTH(rectangle1_widths[1873]), .RECT1_HEIGHT(rectangle1_heights[1873]), .RECT1_WEIGHT(rectangle1_weights[1873]), .RECT2_X(rectangle2_xs[1873]), .RECT2_Y(rectangle2_ys[1873]), .RECT2_WIDTH(rectangle2_widths[1873]), .RECT2_HEIGHT(rectangle2_heights[1873]), .RECT2_WEIGHT(rectangle2_weights[1873]), .RECT3_X(rectangle3_xs[1873]), .RECT3_Y(rectangle3_ys[1873]), .RECT3_WIDTH(rectangle3_widths[1873]), .RECT3_HEIGHT(rectangle3_heights[1873]), .RECT3_WEIGHT(rectangle3_weights[1873]), .FEAT_THRES(feature_thresholds[1873]), .FEAT_ABOVE(feature_aboves[1873]), .FEAT_BELOW(feature_belows[1873])) ac1873(.scan_win(scan_win1873), .scan_win_std_dev(scan_win_std_dev[1873]), .feature_accum(feature_accums[1873]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1874]), .RECT1_Y(rectangle1_ys[1874]), .RECT1_WIDTH(rectangle1_widths[1874]), .RECT1_HEIGHT(rectangle1_heights[1874]), .RECT1_WEIGHT(rectangle1_weights[1874]), .RECT2_X(rectangle2_xs[1874]), .RECT2_Y(rectangle2_ys[1874]), .RECT2_WIDTH(rectangle2_widths[1874]), .RECT2_HEIGHT(rectangle2_heights[1874]), .RECT2_WEIGHT(rectangle2_weights[1874]), .RECT3_X(rectangle3_xs[1874]), .RECT3_Y(rectangle3_ys[1874]), .RECT3_WIDTH(rectangle3_widths[1874]), .RECT3_HEIGHT(rectangle3_heights[1874]), .RECT3_WEIGHT(rectangle3_weights[1874]), .FEAT_THRES(feature_thresholds[1874]), .FEAT_ABOVE(feature_aboves[1874]), .FEAT_BELOW(feature_belows[1874])) ac1874(.scan_win(scan_win1874), .scan_win_std_dev(scan_win_std_dev[1874]), .feature_accum(feature_accums[1874]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1875]), .RECT1_Y(rectangle1_ys[1875]), .RECT1_WIDTH(rectangle1_widths[1875]), .RECT1_HEIGHT(rectangle1_heights[1875]), .RECT1_WEIGHT(rectangle1_weights[1875]), .RECT2_X(rectangle2_xs[1875]), .RECT2_Y(rectangle2_ys[1875]), .RECT2_WIDTH(rectangle2_widths[1875]), .RECT2_HEIGHT(rectangle2_heights[1875]), .RECT2_WEIGHT(rectangle2_weights[1875]), .RECT3_X(rectangle3_xs[1875]), .RECT3_Y(rectangle3_ys[1875]), .RECT3_WIDTH(rectangle3_widths[1875]), .RECT3_HEIGHT(rectangle3_heights[1875]), .RECT3_WEIGHT(rectangle3_weights[1875]), .FEAT_THRES(feature_thresholds[1875]), .FEAT_ABOVE(feature_aboves[1875]), .FEAT_BELOW(feature_belows[1875])) ac1875(.scan_win(scan_win1875), .scan_win_std_dev(scan_win_std_dev[1875]), .feature_accum(feature_accums[1875]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1876]), .RECT1_Y(rectangle1_ys[1876]), .RECT1_WIDTH(rectangle1_widths[1876]), .RECT1_HEIGHT(rectangle1_heights[1876]), .RECT1_WEIGHT(rectangle1_weights[1876]), .RECT2_X(rectangle2_xs[1876]), .RECT2_Y(rectangle2_ys[1876]), .RECT2_WIDTH(rectangle2_widths[1876]), .RECT2_HEIGHT(rectangle2_heights[1876]), .RECT2_WEIGHT(rectangle2_weights[1876]), .RECT3_X(rectangle3_xs[1876]), .RECT3_Y(rectangle3_ys[1876]), .RECT3_WIDTH(rectangle3_widths[1876]), .RECT3_HEIGHT(rectangle3_heights[1876]), .RECT3_WEIGHT(rectangle3_weights[1876]), .FEAT_THRES(feature_thresholds[1876]), .FEAT_ABOVE(feature_aboves[1876]), .FEAT_BELOW(feature_belows[1876])) ac1876(.scan_win(scan_win1876), .scan_win_std_dev(scan_win_std_dev[1876]), .feature_accum(feature_accums[1876]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1877]), .RECT1_Y(rectangle1_ys[1877]), .RECT1_WIDTH(rectangle1_widths[1877]), .RECT1_HEIGHT(rectangle1_heights[1877]), .RECT1_WEIGHT(rectangle1_weights[1877]), .RECT2_X(rectangle2_xs[1877]), .RECT2_Y(rectangle2_ys[1877]), .RECT2_WIDTH(rectangle2_widths[1877]), .RECT2_HEIGHT(rectangle2_heights[1877]), .RECT2_WEIGHT(rectangle2_weights[1877]), .RECT3_X(rectangle3_xs[1877]), .RECT3_Y(rectangle3_ys[1877]), .RECT3_WIDTH(rectangle3_widths[1877]), .RECT3_HEIGHT(rectangle3_heights[1877]), .RECT3_WEIGHT(rectangle3_weights[1877]), .FEAT_THRES(feature_thresholds[1877]), .FEAT_ABOVE(feature_aboves[1877]), .FEAT_BELOW(feature_belows[1877])) ac1877(.scan_win(scan_win1877), .scan_win_std_dev(scan_win_std_dev[1877]), .feature_accum(feature_accums[1877]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1878]), .RECT1_Y(rectangle1_ys[1878]), .RECT1_WIDTH(rectangle1_widths[1878]), .RECT1_HEIGHT(rectangle1_heights[1878]), .RECT1_WEIGHT(rectangle1_weights[1878]), .RECT2_X(rectangle2_xs[1878]), .RECT2_Y(rectangle2_ys[1878]), .RECT2_WIDTH(rectangle2_widths[1878]), .RECT2_HEIGHT(rectangle2_heights[1878]), .RECT2_WEIGHT(rectangle2_weights[1878]), .RECT3_X(rectangle3_xs[1878]), .RECT3_Y(rectangle3_ys[1878]), .RECT3_WIDTH(rectangle3_widths[1878]), .RECT3_HEIGHT(rectangle3_heights[1878]), .RECT3_WEIGHT(rectangle3_weights[1878]), .FEAT_THRES(feature_thresholds[1878]), .FEAT_ABOVE(feature_aboves[1878]), .FEAT_BELOW(feature_belows[1878])) ac1878(.scan_win(scan_win1878), .scan_win_std_dev(scan_win_std_dev[1878]), .feature_accum(feature_accums[1878]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1879]), .RECT1_Y(rectangle1_ys[1879]), .RECT1_WIDTH(rectangle1_widths[1879]), .RECT1_HEIGHT(rectangle1_heights[1879]), .RECT1_WEIGHT(rectangle1_weights[1879]), .RECT2_X(rectangle2_xs[1879]), .RECT2_Y(rectangle2_ys[1879]), .RECT2_WIDTH(rectangle2_widths[1879]), .RECT2_HEIGHT(rectangle2_heights[1879]), .RECT2_WEIGHT(rectangle2_weights[1879]), .RECT3_X(rectangle3_xs[1879]), .RECT3_Y(rectangle3_ys[1879]), .RECT3_WIDTH(rectangle3_widths[1879]), .RECT3_HEIGHT(rectangle3_heights[1879]), .RECT3_WEIGHT(rectangle3_weights[1879]), .FEAT_THRES(feature_thresholds[1879]), .FEAT_ABOVE(feature_aboves[1879]), .FEAT_BELOW(feature_belows[1879])) ac1879(.scan_win(scan_win1879), .scan_win_std_dev(scan_win_std_dev[1879]), .feature_accum(feature_accums[1879]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1880]), .RECT1_Y(rectangle1_ys[1880]), .RECT1_WIDTH(rectangle1_widths[1880]), .RECT1_HEIGHT(rectangle1_heights[1880]), .RECT1_WEIGHT(rectangle1_weights[1880]), .RECT2_X(rectangle2_xs[1880]), .RECT2_Y(rectangle2_ys[1880]), .RECT2_WIDTH(rectangle2_widths[1880]), .RECT2_HEIGHT(rectangle2_heights[1880]), .RECT2_WEIGHT(rectangle2_weights[1880]), .RECT3_X(rectangle3_xs[1880]), .RECT3_Y(rectangle3_ys[1880]), .RECT3_WIDTH(rectangle3_widths[1880]), .RECT3_HEIGHT(rectangle3_heights[1880]), .RECT3_WEIGHT(rectangle3_weights[1880]), .FEAT_THRES(feature_thresholds[1880]), .FEAT_ABOVE(feature_aboves[1880]), .FEAT_BELOW(feature_belows[1880])) ac1880(.scan_win(scan_win1880), .scan_win_std_dev(scan_win_std_dev[1880]), .feature_accum(feature_accums[1880]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1881]), .RECT1_Y(rectangle1_ys[1881]), .RECT1_WIDTH(rectangle1_widths[1881]), .RECT1_HEIGHT(rectangle1_heights[1881]), .RECT1_WEIGHT(rectangle1_weights[1881]), .RECT2_X(rectangle2_xs[1881]), .RECT2_Y(rectangle2_ys[1881]), .RECT2_WIDTH(rectangle2_widths[1881]), .RECT2_HEIGHT(rectangle2_heights[1881]), .RECT2_WEIGHT(rectangle2_weights[1881]), .RECT3_X(rectangle3_xs[1881]), .RECT3_Y(rectangle3_ys[1881]), .RECT3_WIDTH(rectangle3_widths[1881]), .RECT3_HEIGHT(rectangle3_heights[1881]), .RECT3_WEIGHT(rectangle3_weights[1881]), .FEAT_THRES(feature_thresholds[1881]), .FEAT_ABOVE(feature_aboves[1881]), .FEAT_BELOW(feature_belows[1881])) ac1881(.scan_win(scan_win1881), .scan_win_std_dev(scan_win_std_dev[1881]), .feature_accum(feature_accums[1881]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1882]), .RECT1_Y(rectangle1_ys[1882]), .RECT1_WIDTH(rectangle1_widths[1882]), .RECT1_HEIGHT(rectangle1_heights[1882]), .RECT1_WEIGHT(rectangle1_weights[1882]), .RECT2_X(rectangle2_xs[1882]), .RECT2_Y(rectangle2_ys[1882]), .RECT2_WIDTH(rectangle2_widths[1882]), .RECT2_HEIGHT(rectangle2_heights[1882]), .RECT2_WEIGHT(rectangle2_weights[1882]), .RECT3_X(rectangle3_xs[1882]), .RECT3_Y(rectangle3_ys[1882]), .RECT3_WIDTH(rectangle3_widths[1882]), .RECT3_HEIGHT(rectangle3_heights[1882]), .RECT3_WEIGHT(rectangle3_weights[1882]), .FEAT_THRES(feature_thresholds[1882]), .FEAT_ABOVE(feature_aboves[1882]), .FEAT_BELOW(feature_belows[1882])) ac1882(.scan_win(scan_win1882), .scan_win_std_dev(scan_win_std_dev[1882]), .feature_accum(feature_accums[1882]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1883]), .RECT1_Y(rectangle1_ys[1883]), .RECT1_WIDTH(rectangle1_widths[1883]), .RECT1_HEIGHT(rectangle1_heights[1883]), .RECT1_WEIGHT(rectangle1_weights[1883]), .RECT2_X(rectangle2_xs[1883]), .RECT2_Y(rectangle2_ys[1883]), .RECT2_WIDTH(rectangle2_widths[1883]), .RECT2_HEIGHT(rectangle2_heights[1883]), .RECT2_WEIGHT(rectangle2_weights[1883]), .RECT3_X(rectangle3_xs[1883]), .RECT3_Y(rectangle3_ys[1883]), .RECT3_WIDTH(rectangle3_widths[1883]), .RECT3_HEIGHT(rectangle3_heights[1883]), .RECT3_WEIGHT(rectangle3_weights[1883]), .FEAT_THRES(feature_thresholds[1883]), .FEAT_ABOVE(feature_aboves[1883]), .FEAT_BELOW(feature_belows[1883])) ac1883(.scan_win(scan_win1883), .scan_win_std_dev(scan_win_std_dev[1883]), .feature_accum(feature_accums[1883]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1884]), .RECT1_Y(rectangle1_ys[1884]), .RECT1_WIDTH(rectangle1_widths[1884]), .RECT1_HEIGHT(rectangle1_heights[1884]), .RECT1_WEIGHT(rectangle1_weights[1884]), .RECT2_X(rectangle2_xs[1884]), .RECT2_Y(rectangle2_ys[1884]), .RECT2_WIDTH(rectangle2_widths[1884]), .RECT2_HEIGHT(rectangle2_heights[1884]), .RECT2_WEIGHT(rectangle2_weights[1884]), .RECT3_X(rectangle3_xs[1884]), .RECT3_Y(rectangle3_ys[1884]), .RECT3_WIDTH(rectangle3_widths[1884]), .RECT3_HEIGHT(rectangle3_heights[1884]), .RECT3_WEIGHT(rectangle3_weights[1884]), .FEAT_THRES(feature_thresholds[1884]), .FEAT_ABOVE(feature_aboves[1884]), .FEAT_BELOW(feature_belows[1884])) ac1884(.scan_win(scan_win1884), .scan_win_std_dev(scan_win_std_dev[1884]), .feature_accum(feature_accums[1884]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1885]), .RECT1_Y(rectangle1_ys[1885]), .RECT1_WIDTH(rectangle1_widths[1885]), .RECT1_HEIGHT(rectangle1_heights[1885]), .RECT1_WEIGHT(rectangle1_weights[1885]), .RECT2_X(rectangle2_xs[1885]), .RECT2_Y(rectangle2_ys[1885]), .RECT2_WIDTH(rectangle2_widths[1885]), .RECT2_HEIGHT(rectangle2_heights[1885]), .RECT2_WEIGHT(rectangle2_weights[1885]), .RECT3_X(rectangle3_xs[1885]), .RECT3_Y(rectangle3_ys[1885]), .RECT3_WIDTH(rectangle3_widths[1885]), .RECT3_HEIGHT(rectangle3_heights[1885]), .RECT3_WEIGHT(rectangle3_weights[1885]), .FEAT_THRES(feature_thresholds[1885]), .FEAT_ABOVE(feature_aboves[1885]), .FEAT_BELOW(feature_belows[1885])) ac1885(.scan_win(scan_win1885), .scan_win_std_dev(scan_win_std_dev[1885]), .feature_accum(feature_accums[1885]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1886]), .RECT1_Y(rectangle1_ys[1886]), .RECT1_WIDTH(rectangle1_widths[1886]), .RECT1_HEIGHT(rectangle1_heights[1886]), .RECT1_WEIGHT(rectangle1_weights[1886]), .RECT2_X(rectangle2_xs[1886]), .RECT2_Y(rectangle2_ys[1886]), .RECT2_WIDTH(rectangle2_widths[1886]), .RECT2_HEIGHT(rectangle2_heights[1886]), .RECT2_WEIGHT(rectangle2_weights[1886]), .RECT3_X(rectangle3_xs[1886]), .RECT3_Y(rectangle3_ys[1886]), .RECT3_WIDTH(rectangle3_widths[1886]), .RECT3_HEIGHT(rectangle3_heights[1886]), .RECT3_WEIGHT(rectangle3_weights[1886]), .FEAT_THRES(feature_thresholds[1886]), .FEAT_ABOVE(feature_aboves[1886]), .FEAT_BELOW(feature_belows[1886])) ac1886(.scan_win(scan_win1886), .scan_win_std_dev(scan_win_std_dev[1886]), .feature_accum(feature_accums[1886]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1887]), .RECT1_Y(rectangle1_ys[1887]), .RECT1_WIDTH(rectangle1_widths[1887]), .RECT1_HEIGHT(rectangle1_heights[1887]), .RECT1_WEIGHT(rectangle1_weights[1887]), .RECT2_X(rectangle2_xs[1887]), .RECT2_Y(rectangle2_ys[1887]), .RECT2_WIDTH(rectangle2_widths[1887]), .RECT2_HEIGHT(rectangle2_heights[1887]), .RECT2_WEIGHT(rectangle2_weights[1887]), .RECT3_X(rectangle3_xs[1887]), .RECT3_Y(rectangle3_ys[1887]), .RECT3_WIDTH(rectangle3_widths[1887]), .RECT3_HEIGHT(rectangle3_heights[1887]), .RECT3_WEIGHT(rectangle3_weights[1887]), .FEAT_THRES(feature_thresholds[1887]), .FEAT_ABOVE(feature_aboves[1887]), .FEAT_BELOW(feature_belows[1887])) ac1887(.scan_win(scan_win1887), .scan_win_std_dev(scan_win_std_dev[1887]), .feature_accum(feature_accums[1887]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1888]), .RECT1_Y(rectangle1_ys[1888]), .RECT1_WIDTH(rectangle1_widths[1888]), .RECT1_HEIGHT(rectangle1_heights[1888]), .RECT1_WEIGHT(rectangle1_weights[1888]), .RECT2_X(rectangle2_xs[1888]), .RECT2_Y(rectangle2_ys[1888]), .RECT2_WIDTH(rectangle2_widths[1888]), .RECT2_HEIGHT(rectangle2_heights[1888]), .RECT2_WEIGHT(rectangle2_weights[1888]), .RECT3_X(rectangle3_xs[1888]), .RECT3_Y(rectangle3_ys[1888]), .RECT3_WIDTH(rectangle3_widths[1888]), .RECT3_HEIGHT(rectangle3_heights[1888]), .RECT3_WEIGHT(rectangle3_weights[1888]), .FEAT_THRES(feature_thresholds[1888]), .FEAT_ABOVE(feature_aboves[1888]), .FEAT_BELOW(feature_belows[1888])) ac1888(.scan_win(scan_win1888), .scan_win_std_dev(scan_win_std_dev[1888]), .feature_accum(feature_accums[1888]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1889]), .RECT1_Y(rectangle1_ys[1889]), .RECT1_WIDTH(rectangle1_widths[1889]), .RECT1_HEIGHT(rectangle1_heights[1889]), .RECT1_WEIGHT(rectangle1_weights[1889]), .RECT2_X(rectangle2_xs[1889]), .RECT2_Y(rectangle2_ys[1889]), .RECT2_WIDTH(rectangle2_widths[1889]), .RECT2_HEIGHT(rectangle2_heights[1889]), .RECT2_WEIGHT(rectangle2_weights[1889]), .RECT3_X(rectangle3_xs[1889]), .RECT3_Y(rectangle3_ys[1889]), .RECT3_WIDTH(rectangle3_widths[1889]), .RECT3_HEIGHT(rectangle3_heights[1889]), .RECT3_WEIGHT(rectangle3_weights[1889]), .FEAT_THRES(feature_thresholds[1889]), .FEAT_ABOVE(feature_aboves[1889]), .FEAT_BELOW(feature_belows[1889])) ac1889(.scan_win(scan_win1889), .scan_win_std_dev(scan_win_std_dev[1889]), .feature_accum(feature_accums[1889]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1890]), .RECT1_Y(rectangle1_ys[1890]), .RECT1_WIDTH(rectangle1_widths[1890]), .RECT1_HEIGHT(rectangle1_heights[1890]), .RECT1_WEIGHT(rectangle1_weights[1890]), .RECT2_X(rectangle2_xs[1890]), .RECT2_Y(rectangle2_ys[1890]), .RECT2_WIDTH(rectangle2_widths[1890]), .RECT2_HEIGHT(rectangle2_heights[1890]), .RECT2_WEIGHT(rectangle2_weights[1890]), .RECT3_X(rectangle3_xs[1890]), .RECT3_Y(rectangle3_ys[1890]), .RECT3_WIDTH(rectangle3_widths[1890]), .RECT3_HEIGHT(rectangle3_heights[1890]), .RECT3_WEIGHT(rectangle3_weights[1890]), .FEAT_THRES(feature_thresholds[1890]), .FEAT_ABOVE(feature_aboves[1890]), .FEAT_BELOW(feature_belows[1890])) ac1890(.scan_win(scan_win1890), .scan_win_std_dev(scan_win_std_dev[1890]), .feature_accum(feature_accums[1890]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1891]), .RECT1_Y(rectangle1_ys[1891]), .RECT1_WIDTH(rectangle1_widths[1891]), .RECT1_HEIGHT(rectangle1_heights[1891]), .RECT1_WEIGHT(rectangle1_weights[1891]), .RECT2_X(rectangle2_xs[1891]), .RECT2_Y(rectangle2_ys[1891]), .RECT2_WIDTH(rectangle2_widths[1891]), .RECT2_HEIGHT(rectangle2_heights[1891]), .RECT2_WEIGHT(rectangle2_weights[1891]), .RECT3_X(rectangle3_xs[1891]), .RECT3_Y(rectangle3_ys[1891]), .RECT3_WIDTH(rectangle3_widths[1891]), .RECT3_HEIGHT(rectangle3_heights[1891]), .RECT3_WEIGHT(rectangle3_weights[1891]), .FEAT_THRES(feature_thresholds[1891]), .FEAT_ABOVE(feature_aboves[1891]), .FEAT_BELOW(feature_belows[1891])) ac1891(.scan_win(scan_win1891), .scan_win_std_dev(scan_win_std_dev[1891]), .feature_accum(feature_accums[1891]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1892]), .RECT1_Y(rectangle1_ys[1892]), .RECT1_WIDTH(rectangle1_widths[1892]), .RECT1_HEIGHT(rectangle1_heights[1892]), .RECT1_WEIGHT(rectangle1_weights[1892]), .RECT2_X(rectangle2_xs[1892]), .RECT2_Y(rectangle2_ys[1892]), .RECT2_WIDTH(rectangle2_widths[1892]), .RECT2_HEIGHT(rectangle2_heights[1892]), .RECT2_WEIGHT(rectangle2_weights[1892]), .RECT3_X(rectangle3_xs[1892]), .RECT3_Y(rectangle3_ys[1892]), .RECT3_WIDTH(rectangle3_widths[1892]), .RECT3_HEIGHT(rectangle3_heights[1892]), .RECT3_WEIGHT(rectangle3_weights[1892]), .FEAT_THRES(feature_thresholds[1892]), .FEAT_ABOVE(feature_aboves[1892]), .FEAT_BELOW(feature_belows[1892])) ac1892(.scan_win(scan_win1892), .scan_win_std_dev(scan_win_std_dev[1892]), .feature_accum(feature_accums[1892]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1893]), .RECT1_Y(rectangle1_ys[1893]), .RECT1_WIDTH(rectangle1_widths[1893]), .RECT1_HEIGHT(rectangle1_heights[1893]), .RECT1_WEIGHT(rectangle1_weights[1893]), .RECT2_X(rectangle2_xs[1893]), .RECT2_Y(rectangle2_ys[1893]), .RECT2_WIDTH(rectangle2_widths[1893]), .RECT2_HEIGHT(rectangle2_heights[1893]), .RECT2_WEIGHT(rectangle2_weights[1893]), .RECT3_X(rectangle3_xs[1893]), .RECT3_Y(rectangle3_ys[1893]), .RECT3_WIDTH(rectangle3_widths[1893]), .RECT3_HEIGHT(rectangle3_heights[1893]), .RECT3_WEIGHT(rectangle3_weights[1893]), .FEAT_THRES(feature_thresholds[1893]), .FEAT_ABOVE(feature_aboves[1893]), .FEAT_BELOW(feature_belows[1893])) ac1893(.scan_win(scan_win1893), .scan_win_std_dev(scan_win_std_dev[1893]), .feature_accum(feature_accums[1893]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1894]), .RECT1_Y(rectangle1_ys[1894]), .RECT1_WIDTH(rectangle1_widths[1894]), .RECT1_HEIGHT(rectangle1_heights[1894]), .RECT1_WEIGHT(rectangle1_weights[1894]), .RECT2_X(rectangle2_xs[1894]), .RECT2_Y(rectangle2_ys[1894]), .RECT2_WIDTH(rectangle2_widths[1894]), .RECT2_HEIGHT(rectangle2_heights[1894]), .RECT2_WEIGHT(rectangle2_weights[1894]), .RECT3_X(rectangle3_xs[1894]), .RECT3_Y(rectangle3_ys[1894]), .RECT3_WIDTH(rectangle3_widths[1894]), .RECT3_HEIGHT(rectangle3_heights[1894]), .RECT3_WEIGHT(rectangle3_weights[1894]), .FEAT_THRES(feature_thresholds[1894]), .FEAT_ABOVE(feature_aboves[1894]), .FEAT_BELOW(feature_belows[1894])) ac1894(.scan_win(scan_win1894), .scan_win_std_dev(scan_win_std_dev[1894]), .feature_accum(feature_accums[1894]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1895]), .RECT1_Y(rectangle1_ys[1895]), .RECT1_WIDTH(rectangle1_widths[1895]), .RECT1_HEIGHT(rectangle1_heights[1895]), .RECT1_WEIGHT(rectangle1_weights[1895]), .RECT2_X(rectangle2_xs[1895]), .RECT2_Y(rectangle2_ys[1895]), .RECT2_WIDTH(rectangle2_widths[1895]), .RECT2_HEIGHT(rectangle2_heights[1895]), .RECT2_WEIGHT(rectangle2_weights[1895]), .RECT3_X(rectangle3_xs[1895]), .RECT3_Y(rectangle3_ys[1895]), .RECT3_WIDTH(rectangle3_widths[1895]), .RECT3_HEIGHT(rectangle3_heights[1895]), .RECT3_WEIGHT(rectangle3_weights[1895]), .FEAT_THRES(feature_thresholds[1895]), .FEAT_ABOVE(feature_aboves[1895]), .FEAT_BELOW(feature_belows[1895])) ac1895(.scan_win(scan_win1895), .scan_win_std_dev(scan_win_std_dev[1895]), .feature_accum(feature_accums[1895]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1896]), .RECT1_Y(rectangle1_ys[1896]), .RECT1_WIDTH(rectangle1_widths[1896]), .RECT1_HEIGHT(rectangle1_heights[1896]), .RECT1_WEIGHT(rectangle1_weights[1896]), .RECT2_X(rectangle2_xs[1896]), .RECT2_Y(rectangle2_ys[1896]), .RECT2_WIDTH(rectangle2_widths[1896]), .RECT2_HEIGHT(rectangle2_heights[1896]), .RECT2_WEIGHT(rectangle2_weights[1896]), .RECT3_X(rectangle3_xs[1896]), .RECT3_Y(rectangle3_ys[1896]), .RECT3_WIDTH(rectangle3_widths[1896]), .RECT3_HEIGHT(rectangle3_heights[1896]), .RECT3_WEIGHT(rectangle3_weights[1896]), .FEAT_THRES(feature_thresholds[1896]), .FEAT_ABOVE(feature_aboves[1896]), .FEAT_BELOW(feature_belows[1896])) ac1896(.scan_win(scan_win1896), .scan_win_std_dev(scan_win_std_dev[1896]), .feature_accum(feature_accums[1896]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1897]), .RECT1_Y(rectangle1_ys[1897]), .RECT1_WIDTH(rectangle1_widths[1897]), .RECT1_HEIGHT(rectangle1_heights[1897]), .RECT1_WEIGHT(rectangle1_weights[1897]), .RECT2_X(rectangle2_xs[1897]), .RECT2_Y(rectangle2_ys[1897]), .RECT2_WIDTH(rectangle2_widths[1897]), .RECT2_HEIGHT(rectangle2_heights[1897]), .RECT2_WEIGHT(rectangle2_weights[1897]), .RECT3_X(rectangle3_xs[1897]), .RECT3_Y(rectangle3_ys[1897]), .RECT3_WIDTH(rectangle3_widths[1897]), .RECT3_HEIGHT(rectangle3_heights[1897]), .RECT3_WEIGHT(rectangle3_weights[1897]), .FEAT_THRES(feature_thresholds[1897]), .FEAT_ABOVE(feature_aboves[1897]), .FEAT_BELOW(feature_belows[1897])) ac1897(.scan_win(scan_win1897), .scan_win_std_dev(scan_win_std_dev[1897]), .feature_accum(feature_accums[1897]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1898]), .RECT1_Y(rectangle1_ys[1898]), .RECT1_WIDTH(rectangle1_widths[1898]), .RECT1_HEIGHT(rectangle1_heights[1898]), .RECT1_WEIGHT(rectangle1_weights[1898]), .RECT2_X(rectangle2_xs[1898]), .RECT2_Y(rectangle2_ys[1898]), .RECT2_WIDTH(rectangle2_widths[1898]), .RECT2_HEIGHT(rectangle2_heights[1898]), .RECT2_WEIGHT(rectangle2_weights[1898]), .RECT3_X(rectangle3_xs[1898]), .RECT3_Y(rectangle3_ys[1898]), .RECT3_WIDTH(rectangle3_widths[1898]), .RECT3_HEIGHT(rectangle3_heights[1898]), .RECT3_WEIGHT(rectangle3_weights[1898]), .FEAT_THRES(feature_thresholds[1898]), .FEAT_ABOVE(feature_aboves[1898]), .FEAT_BELOW(feature_belows[1898])) ac1898(.scan_win(scan_win1898), .scan_win_std_dev(scan_win_std_dev[1898]), .feature_accum(feature_accums[1898]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1899]), .RECT1_Y(rectangle1_ys[1899]), .RECT1_WIDTH(rectangle1_widths[1899]), .RECT1_HEIGHT(rectangle1_heights[1899]), .RECT1_WEIGHT(rectangle1_weights[1899]), .RECT2_X(rectangle2_xs[1899]), .RECT2_Y(rectangle2_ys[1899]), .RECT2_WIDTH(rectangle2_widths[1899]), .RECT2_HEIGHT(rectangle2_heights[1899]), .RECT2_WEIGHT(rectangle2_weights[1899]), .RECT3_X(rectangle3_xs[1899]), .RECT3_Y(rectangle3_ys[1899]), .RECT3_WIDTH(rectangle3_widths[1899]), .RECT3_HEIGHT(rectangle3_heights[1899]), .RECT3_WEIGHT(rectangle3_weights[1899]), .FEAT_THRES(feature_thresholds[1899]), .FEAT_ABOVE(feature_aboves[1899]), .FEAT_BELOW(feature_belows[1899])) ac1899(.scan_win(scan_win1899), .scan_win_std_dev(scan_win_std_dev[1899]), .feature_accum(feature_accums[1899]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1900]), .RECT1_Y(rectangle1_ys[1900]), .RECT1_WIDTH(rectangle1_widths[1900]), .RECT1_HEIGHT(rectangle1_heights[1900]), .RECT1_WEIGHT(rectangle1_weights[1900]), .RECT2_X(rectangle2_xs[1900]), .RECT2_Y(rectangle2_ys[1900]), .RECT2_WIDTH(rectangle2_widths[1900]), .RECT2_HEIGHT(rectangle2_heights[1900]), .RECT2_WEIGHT(rectangle2_weights[1900]), .RECT3_X(rectangle3_xs[1900]), .RECT3_Y(rectangle3_ys[1900]), .RECT3_WIDTH(rectangle3_widths[1900]), .RECT3_HEIGHT(rectangle3_heights[1900]), .RECT3_WEIGHT(rectangle3_weights[1900]), .FEAT_THRES(feature_thresholds[1900]), .FEAT_ABOVE(feature_aboves[1900]), .FEAT_BELOW(feature_belows[1900])) ac1900(.scan_win(scan_win1900), .scan_win_std_dev(scan_win_std_dev[1900]), .feature_accum(feature_accums[1900]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1901]), .RECT1_Y(rectangle1_ys[1901]), .RECT1_WIDTH(rectangle1_widths[1901]), .RECT1_HEIGHT(rectangle1_heights[1901]), .RECT1_WEIGHT(rectangle1_weights[1901]), .RECT2_X(rectangle2_xs[1901]), .RECT2_Y(rectangle2_ys[1901]), .RECT2_WIDTH(rectangle2_widths[1901]), .RECT2_HEIGHT(rectangle2_heights[1901]), .RECT2_WEIGHT(rectangle2_weights[1901]), .RECT3_X(rectangle3_xs[1901]), .RECT3_Y(rectangle3_ys[1901]), .RECT3_WIDTH(rectangle3_widths[1901]), .RECT3_HEIGHT(rectangle3_heights[1901]), .RECT3_WEIGHT(rectangle3_weights[1901]), .FEAT_THRES(feature_thresholds[1901]), .FEAT_ABOVE(feature_aboves[1901]), .FEAT_BELOW(feature_belows[1901])) ac1901(.scan_win(scan_win1901), .scan_win_std_dev(scan_win_std_dev[1901]), .feature_accum(feature_accums[1901]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1902]), .RECT1_Y(rectangle1_ys[1902]), .RECT1_WIDTH(rectangle1_widths[1902]), .RECT1_HEIGHT(rectangle1_heights[1902]), .RECT1_WEIGHT(rectangle1_weights[1902]), .RECT2_X(rectangle2_xs[1902]), .RECT2_Y(rectangle2_ys[1902]), .RECT2_WIDTH(rectangle2_widths[1902]), .RECT2_HEIGHT(rectangle2_heights[1902]), .RECT2_WEIGHT(rectangle2_weights[1902]), .RECT3_X(rectangle3_xs[1902]), .RECT3_Y(rectangle3_ys[1902]), .RECT3_WIDTH(rectangle3_widths[1902]), .RECT3_HEIGHT(rectangle3_heights[1902]), .RECT3_WEIGHT(rectangle3_weights[1902]), .FEAT_THRES(feature_thresholds[1902]), .FEAT_ABOVE(feature_aboves[1902]), .FEAT_BELOW(feature_belows[1902])) ac1902(.scan_win(scan_win1902), .scan_win_std_dev(scan_win_std_dev[1902]), .feature_accum(feature_accums[1902]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1903]), .RECT1_Y(rectangle1_ys[1903]), .RECT1_WIDTH(rectangle1_widths[1903]), .RECT1_HEIGHT(rectangle1_heights[1903]), .RECT1_WEIGHT(rectangle1_weights[1903]), .RECT2_X(rectangle2_xs[1903]), .RECT2_Y(rectangle2_ys[1903]), .RECT2_WIDTH(rectangle2_widths[1903]), .RECT2_HEIGHT(rectangle2_heights[1903]), .RECT2_WEIGHT(rectangle2_weights[1903]), .RECT3_X(rectangle3_xs[1903]), .RECT3_Y(rectangle3_ys[1903]), .RECT3_WIDTH(rectangle3_widths[1903]), .RECT3_HEIGHT(rectangle3_heights[1903]), .RECT3_WEIGHT(rectangle3_weights[1903]), .FEAT_THRES(feature_thresholds[1903]), .FEAT_ABOVE(feature_aboves[1903]), .FEAT_BELOW(feature_belows[1903])) ac1903(.scan_win(scan_win1903), .scan_win_std_dev(scan_win_std_dev[1903]), .feature_accum(feature_accums[1903]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1904]), .RECT1_Y(rectangle1_ys[1904]), .RECT1_WIDTH(rectangle1_widths[1904]), .RECT1_HEIGHT(rectangle1_heights[1904]), .RECT1_WEIGHT(rectangle1_weights[1904]), .RECT2_X(rectangle2_xs[1904]), .RECT2_Y(rectangle2_ys[1904]), .RECT2_WIDTH(rectangle2_widths[1904]), .RECT2_HEIGHT(rectangle2_heights[1904]), .RECT2_WEIGHT(rectangle2_weights[1904]), .RECT3_X(rectangle3_xs[1904]), .RECT3_Y(rectangle3_ys[1904]), .RECT3_WIDTH(rectangle3_widths[1904]), .RECT3_HEIGHT(rectangle3_heights[1904]), .RECT3_WEIGHT(rectangle3_weights[1904]), .FEAT_THRES(feature_thresholds[1904]), .FEAT_ABOVE(feature_aboves[1904]), .FEAT_BELOW(feature_belows[1904])) ac1904(.scan_win(scan_win1904), .scan_win_std_dev(scan_win_std_dev[1904]), .feature_accum(feature_accums[1904]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1905]), .RECT1_Y(rectangle1_ys[1905]), .RECT1_WIDTH(rectangle1_widths[1905]), .RECT1_HEIGHT(rectangle1_heights[1905]), .RECT1_WEIGHT(rectangle1_weights[1905]), .RECT2_X(rectangle2_xs[1905]), .RECT2_Y(rectangle2_ys[1905]), .RECT2_WIDTH(rectangle2_widths[1905]), .RECT2_HEIGHT(rectangle2_heights[1905]), .RECT2_WEIGHT(rectangle2_weights[1905]), .RECT3_X(rectangle3_xs[1905]), .RECT3_Y(rectangle3_ys[1905]), .RECT3_WIDTH(rectangle3_widths[1905]), .RECT3_HEIGHT(rectangle3_heights[1905]), .RECT3_WEIGHT(rectangle3_weights[1905]), .FEAT_THRES(feature_thresholds[1905]), .FEAT_ABOVE(feature_aboves[1905]), .FEAT_BELOW(feature_belows[1905])) ac1905(.scan_win(scan_win1905), .scan_win_std_dev(scan_win_std_dev[1905]), .feature_accum(feature_accums[1905]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1906]), .RECT1_Y(rectangle1_ys[1906]), .RECT1_WIDTH(rectangle1_widths[1906]), .RECT1_HEIGHT(rectangle1_heights[1906]), .RECT1_WEIGHT(rectangle1_weights[1906]), .RECT2_X(rectangle2_xs[1906]), .RECT2_Y(rectangle2_ys[1906]), .RECT2_WIDTH(rectangle2_widths[1906]), .RECT2_HEIGHT(rectangle2_heights[1906]), .RECT2_WEIGHT(rectangle2_weights[1906]), .RECT3_X(rectangle3_xs[1906]), .RECT3_Y(rectangle3_ys[1906]), .RECT3_WIDTH(rectangle3_widths[1906]), .RECT3_HEIGHT(rectangle3_heights[1906]), .RECT3_WEIGHT(rectangle3_weights[1906]), .FEAT_THRES(feature_thresholds[1906]), .FEAT_ABOVE(feature_aboves[1906]), .FEAT_BELOW(feature_belows[1906])) ac1906(.scan_win(scan_win1906), .scan_win_std_dev(scan_win_std_dev[1906]), .feature_accum(feature_accums[1906]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1907]), .RECT1_Y(rectangle1_ys[1907]), .RECT1_WIDTH(rectangle1_widths[1907]), .RECT1_HEIGHT(rectangle1_heights[1907]), .RECT1_WEIGHT(rectangle1_weights[1907]), .RECT2_X(rectangle2_xs[1907]), .RECT2_Y(rectangle2_ys[1907]), .RECT2_WIDTH(rectangle2_widths[1907]), .RECT2_HEIGHT(rectangle2_heights[1907]), .RECT2_WEIGHT(rectangle2_weights[1907]), .RECT3_X(rectangle3_xs[1907]), .RECT3_Y(rectangle3_ys[1907]), .RECT3_WIDTH(rectangle3_widths[1907]), .RECT3_HEIGHT(rectangle3_heights[1907]), .RECT3_WEIGHT(rectangle3_weights[1907]), .FEAT_THRES(feature_thresholds[1907]), .FEAT_ABOVE(feature_aboves[1907]), .FEAT_BELOW(feature_belows[1907])) ac1907(.scan_win(scan_win1907), .scan_win_std_dev(scan_win_std_dev[1907]), .feature_accum(feature_accums[1907]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1908]), .RECT1_Y(rectangle1_ys[1908]), .RECT1_WIDTH(rectangle1_widths[1908]), .RECT1_HEIGHT(rectangle1_heights[1908]), .RECT1_WEIGHT(rectangle1_weights[1908]), .RECT2_X(rectangle2_xs[1908]), .RECT2_Y(rectangle2_ys[1908]), .RECT2_WIDTH(rectangle2_widths[1908]), .RECT2_HEIGHT(rectangle2_heights[1908]), .RECT2_WEIGHT(rectangle2_weights[1908]), .RECT3_X(rectangle3_xs[1908]), .RECT3_Y(rectangle3_ys[1908]), .RECT3_WIDTH(rectangle3_widths[1908]), .RECT3_HEIGHT(rectangle3_heights[1908]), .RECT3_WEIGHT(rectangle3_weights[1908]), .FEAT_THRES(feature_thresholds[1908]), .FEAT_ABOVE(feature_aboves[1908]), .FEAT_BELOW(feature_belows[1908])) ac1908(.scan_win(scan_win1908), .scan_win_std_dev(scan_win_std_dev[1908]), .feature_accum(feature_accums[1908]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1909]), .RECT1_Y(rectangle1_ys[1909]), .RECT1_WIDTH(rectangle1_widths[1909]), .RECT1_HEIGHT(rectangle1_heights[1909]), .RECT1_WEIGHT(rectangle1_weights[1909]), .RECT2_X(rectangle2_xs[1909]), .RECT2_Y(rectangle2_ys[1909]), .RECT2_WIDTH(rectangle2_widths[1909]), .RECT2_HEIGHT(rectangle2_heights[1909]), .RECT2_WEIGHT(rectangle2_weights[1909]), .RECT3_X(rectangle3_xs[1909]), .RECT3_Y(rectangle3_ys[1909]), .RECT3_WIDTH(rectangle3_widths[1909]), .RECT3_HEIGHT(rectangle3_heights[1909]), .RECT3_WEIGHT(rectangle3_weights[1909]), .FEAT_THRES(feature_thresholds[1909]), .FEAT_ABOVE(feature_aboves[1909]), .FEAT_BELOW(feature_belows[1909])) ac1909(.scan_win(scan_win1909), .scan_win_std_dev(scan_win_std_dev[1909]), .feature_accum(feature_accums[1909]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1910]), .RECT1_Y(rectangle1_ys[1910]), .RECT1_WIDTH(rectangle1_widths[1910]), .RECT1_HEIGHT(rectangle1_heights[1910]), .RECT1_WEIGHT(rectangle1_weights[1910]), .RECT2_X(rectangle2_xs[1910]), .RECT2_Y(rectangle2_ys[1910]), .RECT2_WIDTH(rectangle2_widths[1910]), .RECT2_HEIGHT(rectangle2_heights[1910]), .RECT2_WEIGHT(rectangle2_weights[1910]), .RECT3_X(rectangle3_xs[1910]), .RECT3_Y(rectangle3_ys[1910]), .RECT3_WIDTH(rectangle3_widths[1910]), .RECT3_HEIGHT(rectangle3_heights[1910]), .RECT3_WEIGHT(rectangle3_weights[1910]), .FEAT_THRES(feature_thresholds[1910]), .FEAT_ABOVE(feature_aboves[1910]), .FEAT_BELOW(feature_belows[1910])) ac1910(.scan_win(scan_win1910), .scan_win_std_dev(scan_win_std_dev[1910]), .feature_accum(feature_accums[1910]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1911]), .RECT1_Y(rectangle1_ys[1911]), .RECT1_WIDTH(rectangle1_widths[1911]), .RECT1_HEIGHT(rectangle1_heights[1911]), .RECT1_WEIGHT(rectangle1_weights[1911]), .RECT2_X(rectangle2_xs[1911]), .RECT2_Y(rectangle2_ys[1911]), .RECT2_WIDTH(rectangle2_widths[1911]), .RECT2_HEIGHT(rectangle2_heights[1911]), .RECT2_WEIGHT(rectangle2_weights[1911]), .RECT3_X(rectangle3_xs[1911]), .RECT3_Y(rectangle3_ys[1911]), .RECT3_WIDTH(rectangle3_widths[1911]), .RECT3_HEIGHT(rectangle3_heights[1911]), .RECT3_WEIGHT(rectangle3_weights[1911]), .FEAT_THRES(feature_thresholds[1911]), .FEAT_ABOVE(feature_aboves[1911]), .FEAT_BELOW(feature_belows[1911])) ac1911(.scan_win(scan_win1911), .scan_win_std_dev(scan_win_std_dev[1911]), .feature_accum(feature_accums[1911]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1912]), .RECT1_Y(rectangle1_ys[1912]), .RECT1_WIDTH(rectangle1_widths[1912]), .RECT1_HEIGHT(rectangle1_heights[1912]), .RECT1_WEIGHT(rectangle1_weights[1912]), .RECT2_X(rectangle2_xs[1912]), .RECT2_Y(rectangle2_ys[1912]), .RECT2_WIDTH(rectangle2_widths[1912]), .RECT2_HEIGHT(rectangle2_heights[1912]), .RECT2_WEIGHT(rectangle2_weights[1912]), .RECT3_X(rectangle3_xs[1912]), .RECT3_Y(rectangle3_ys[1912]), .RECT3_WIDTH(rectangle3_widths[1912]), .RECT3_HEIGHT(rectangle3_heights[1912]), .RECT3_WEIGHT(rectangle3_weights[1912]), .FEAT_THRES(feature_thresholds[1912]), .FEAT_ABOVE(feature_aboves[1912]), .FEAT_BELOW(feature_belows[1912])) ac1912(.scan_win(scan_win1912), .scan_win_std_dev(scan_win_std_dev[1912]), .feature_accum(feature_accums[1912]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1913]), .RECT1_Y(rectangle1_ys[1913]), .RECT1_WIDTH(rectangle1_widths[1913]), .RECT1_HEIGHT(rectangle1_heights[1913]), .RECT1_WEIGHT(rectangle1_weights[1913]), .RECT2_X(rectangle2_xs[1913]), .RECT2_Y(rectangle2_ys[1913]), .RECT2_WIDTH(rectangle2_widths[1913]), .RECT2_HEIGHT(rectangle2_heights[1913]), .RECT2_WEIGHT(rectangle2_weights[1913]), .RECT3_X(rectangle3_xs[1913]), .RECT3_Y(rectangle3_ys[1913]), .RECT3_WIDTH(rectangle3_widths[1913]), .RECT3_HEIGHT(rectangle3_heights[1913]), .RECT3_WEIGHT(rectangle3_weights[1913]), .FEAT_THRES(feature_thresholds[1913]), .FEAT_ABOVE(feature_aboves[1913]), .FEAT_BELOW(feature_belows[1913])) ac1913(.scan_win(scan_win1913), .scan_win_std_dev(scan_win_std_dev[1913]), .feature_accum(feature_accums[1913]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1914]), .RECT1_Y(rectangle1_ys[1914]), .RECT1_WIDTH(rectangle1_widths[1914]), .RECT1_HEIGHT(rectangle1_heights[1914]), .RECT1_WEIGHT(rectangle1_weights[1914]), .RECT2_X(rectangle2_xs[1914]), .RECT2_Y(rectangle2_ys[1914]), .RECT2_WIDTH(rectangle2_widths[1914]), .RECT2_HEIGHT(rectangle2_heights[1914]), .RECT2_WEIGHT(rectangle2_weights[1914]), .RECT3_X(rectangle3_xs[1914]), .RECT3_Y(rectangle3_ys[1914]), .RECT3_WIDTH(rectangle3_widths[1914]), .RECT3_HEIGHT(rectangle3_heights[1914]), .RECT3_WEIGHT(rectangle3_weights[1914]), .FEAT_THRES(feature_thresholds[1914]), .FEAT_ABOVE(feature_aboves[1914]), .FEAT_BELOW(feature_belows[1914])) ac1914(.scan_win(scan_win1914), .scan_win_std_dev(scan_win_std_dev[1914]), .feature_accum(feature_accums[1914]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1915]), .RECT1_Y(rectangle1_ys[1915]), .RECT1_WIDTH(rectangle1_widths[1915]), .RECT1_HEIGHT(rectangle1_heights[1915]), .RECT1_WEIGHT(rectangle1_weights[1915]), .RECT2_X(rectangle2_xs[1915]), .RECT2_Y(rectangle2_ys[1915]), .RECT2_WIDTH(rectangle2_widths[1915]), .RECT2_HEIGHT(rectangle2_heights[1915]), .RECT2_WEIGHT(rectangle2_weights[1915]), .RECT3_X(rectangle3_xs[1915]), .RECT3_Y(rectangle3_ys[1915]), .RECT3_WIDTH(rectangle3_widths[1915]), .RECT3_HEIGHT(rectangle3_heights[1915]), .RECT3_WEIGHT(rectangle3_weights[1915]), .FEAT_THRES(feature_thresholds[1915]), .FEAT_ABOVE(feature_aboves[1915]), .FEAT_BELOW(feature_belows[1915])) ac1915(.scan_win(scan_win1915), .scan_win_std_dev(scan_win_std_dev[1915]), .feature_accum(feature_accums[1915]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1916]), .RECT1_Y(rectangle1_ys[1916]), .RECT1_WIDTH(rectangle1_widths[1916]), .RECT1_HEIGHT(rectangle1_heights[1916]), .RECT1_WEIGHT(rectangle1_weights[1916]), .RECT2_X(rectangle2_xs[1916]), .RECT2_Y(rectangle2_ys[1916]), .RECT2_WIDTH(rectangle2_widths[1916]), .RECT2_HEIGHT(rectangle2_heights[1916]), .RECT2_WEIGHT(rectangle2_weights[1916]), .RECT3_X(rectangle3_xs[1916]), .RECT3_Y(rectangle3_ys[1916]), .RECT3_WIDTH(rectangle3_widths[1916]), .RECT3_HEIGHT(rectangle3_heights[1916]), .RECT3_WEIGHT(rectangle3_weights[1916]), .FEAT_THRES(feature_thresholds[1916]), .FEAT_ABOVE(feature_aboves[1916]), .FEAT_BELOW(feature_belows[1916])) ac1916(.scan_win(scan_win1916), .scan_win_std_dev(scan_win_std_dev[1916]), .feature_accum(feature_accums[1916]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1917]), .RECT1_Y(rectangle1_ys[1917]), .RECT1_WIDTH(rectangle1_widths[1917]), .RECT1_HEIGHT(rectangle1_heights[1917]), .RECT1_WEIGHT(rectangle1_weights[1917]), .RECT2_X(rectangle2_xs[1917]), .RECT2_Y(rectangle2_ys[1917]), .RECT2_WIDTH(rectangle2_widths[1917]), .RECT2_HEIGHT(rectangle2_heights[1917]), .RECT2_WEIGHT(rectangle2_weights[1917]), .RECT3_X(rectangle3_xs[1917]), .RECT3_Y(rectangle3_ys[1917]), .RECT3_WIDTH(rectangle3_widths[1917]), .RECT3_HEIGHT(rectangle3_heights[1917]), .RECT3_WEIGHT(rectangle3_weights[1917]), .FEAT_THRES(feature_thresholds[1917]), .FEAT_ABOVE(feature_aboves[1917]), .FEAT_BELOW(feature_belows[1917])) ac1917(.scan_win(scan_win1917), .scan_win_std_dev(scan_win_std_dev[1917]), .feature_accum(feature_accums[1917]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1918]), .RECT1_Y(rectangle1_ys[1918]), .RECT1_WIDTH(rectangle1_widths[1918]), .RECT1_HEIGHT(rectangle1_heights[1918]), .RECT1_WEIGHT(rectangle1_weights[1918]), .RECT2_X(rectangle2_xs[1918]), .RECT2_Y(rectangle2_ys[1918]), .RECT2_WIDTH(rectangle2_widths[1918]), .RECT2_HEIGHT(rectangle2_heights[1918]), .RECT2_WEIGHT(rectangle2_weights[1918]), .RECT3_X(rectangle3_xs[1918]), .RECT3_Y(rectangle3_ys[1918]), .RECT3_WIDTH(rectangle3_widths[1918]), .RECT3_HEIGHT(rectangle3_heights[1918]), .RECT3_WEIGHT(rectangle3_weights[1918]), .FEAT_THRES(feature_thresholds[1918]), .FEAT_ABOVE(feature_aboves[1918]), .FEAT_BELOW(feature_belows[1918])) ac1918(.scan_win(scan_win1918), .scan_win_std_dev(scan_win_std_dev[1918]), .feature_accum(feature_accums[1918]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1919]), .RECT1_Y(rectangle1_ys[1919]), .RECT1_WIDTH(rectangle1_widths[1919]), .RECT1_HEIGHT(rectangle1_heights[1919]), .RECT1_WEIGHT(rectangle1_weights[1919]), .RECT2_X(rectangle2_xs[1919]), .RECT2_Y(rectangle2_ys[1919]), .RECT2_WIDTH(rectangle2_widths[1919]), .RECT2_HEIGHT(rectangle2_heights[1919]), .RECT2_WEIGHT(rectangle2_weights[1919]), .RECT3_X(rectangle3_xs[1919]), .RECT3_Y(rectangle3_ys[1919]), .RECT3_WIDTH(rectangle3_widths[1919]), .RECT3_HEIGHT(rectangle3_heights[1919]), .RECT3_WEIGHT(rectangle3_weights[1919]), .FEAT_THRES(feature_thresholds[1919]), .FEAT_ABOVE(feature_aboves[1919]), .FEAT_BELOW(feature_belows[1919])) ac1919(.scan_win(scan_win1919), .scan_win_std_dev(scan_win_std_dev[1919]), .feature_accum(feature_accums[1919]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1920]), .RECT1_Y(rectangle1_ys[1920]), .RECT1_WIDTH(rectangle1_widths[1920]), .RECT1_HEIGHT(rectangle1_heights[1920]), .RECT1_WEIGHT(rectangle1_weights[1920]), .RECT2_X(rectangle2_xs[1920]), .RECT2_Y(rectangle2_ys[1920]), .RECT2_WIDTH(rectangle2_widths[1920]), .RECT2_HEIGHT(rectangle2_heights[1920]), .RECT2_WEIGHT(rectangle2_weights[1920]), .RECT3_X(rectangle3_xs[1920]), .RECT3_Y(rectangle3_ys[1920]), .RECT3_WIDTH(rectangle3_widths[1920]), .RECT3_HEIGHT(rectangle3_heights[1920]), .RECT3_WEIGHT(rectangle3_weights[1920]), .FEAT_THRES(feature_thresholds[1920]), .FEAT_ABOVE(feature_aboves[1920]), .FEAT_BELOW(feature_belows[1920])) ac1920(.scan_win(scan_win1920), .scan_win_std_dev(scan_win_std_dev[1920]), .feature_accum(feature_accums[1920]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1921]), .RECT1_Y(rectangle1_ys[1921]), .RECT1_WIDTH(rectangle1_widths[1921]), .RECT1_HEIGHT(rectangle1_heights[1921]), .RECT1_WEIGHT(rectangle1_weights[1921]), .RECT2_X(rectangle2_xs[1921]), .RECT2_Y(rectangle2_ys[1921]), .RECT2_WIDTH(rectangle2_widths[1921]), .RECT2_HEIGHT(rectangle2_heights[1921]), .RECT2_WEIGHT(rectangle2_weights[1921]), .RECT3_X(rectangle3_xs[1921]), .RECT3_Y(rectangle3_ys[1921]), .RECT3_WIDTH(rectangle3_widths[1921]), .RECT3_HEIGHT(rectangle3_heights[1921]), .RECT3_WEIGHT(rectangle3_weights[1921]), .FEAT_THRES(feature_thresholds[1921]), .FEAT_ABOVE(feature_aboves[1921]), .FEAT_BELOW(feature_belows[1921])) ac1921(.scan_win(scan_win1921), .scan_win_std_dev(scan_win_std_dev[1921]), .feature_accum(feature_accums[1921]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1922]), .RECT1_Y(rectangle1_ys[1922]), .RECT1_WIDTH(rectangle1_widths[1922]), .RECT1_HEIGHT(rectangle1_heights[1922]), .RECT1_WEIGHT(rectangle1_weights[1922]), .RECT2_X(rectangle2_xs[1922]), .RECT2_Y(rectangle2_ys[1922]), .RECT2_WIDTH(rectangle2_widths[1922]), .RECT2_HEIGHT(rectangle2_heights[1922]), .RECT2_WEIGHT(rectangle2_weights[1922]), .RECT3_X(rectangle3_xs[1922]), .RECT3_Y(rectangle3_ys[1922]), .RECT3_WIDTH(rectangle3_widths[1922]), .RECT3_HEIGHT(rectangle3_heights[1922]), .RECT3_WEIGHT(rectangle3_weights[1922]), .FEAT_THRES(feature_thresholds[1922]), .FEAT_ABOVE(feature_aboves[1922]), .FEAT_BELOW(feature_belows[1922])) ac1922(.scan_win(scan_win1922), .scan_win_std_dev(scan_win_std_dev[1922]), .feature_accum(feature_accums[1922]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1923]), .RECT1_Y(rectangle1_ys[1923]), .RECT1_WIDTH(rectangle1_widths[1923]), .RECT1_HEIGHT(rectangle1_heights[1923]), .RECT1_WEIGHT(rectangle1_weights[1923]), .RECT2_X(rectangle2_xs[1923]), .RECT2_Y(rectangle2_ys[1923]), .RECT2_WIDTH(rectangle2_widths[1923]), .RECT2_HEIGHT(rectangle2_heights[1923]), .RECT2_WEIGHT(rectangle2_weights[1923]), .RECT3_X(rectangle3_xs[1923]), .RECT3_Y(rectangle3_ys[1923]), .RECT3_WIDTH(rectangle3_widths[1923]), .RECT3_HEIGHT(rectangle3_heights[1923]), .RECT3_WEIGHT(rectangle3_weights[1923]), .FEAT_THRES(feature_thresholds[1923]), .FEAT_ABOVE(feature_aboves[1923]), .FEAT_BELOW(feature_belows[1923])) ac1923(.scan_win(scan_win1923), .scan_win_std_dev(scan_win_std_dev[1923]), .feature_accum(feature_accums[1923]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1924]), .RECT1_Y(rectangle1_ys[1924]), .RECT1_WIDTH(rectangle1_widths[1924]), .RECT1_HEIGHT(rectangle1_heights[1924]), .RECT1_WEIGHT(rectangle1_weights[1924]), .RECT2_X(rectangle2_xs[1924]), .RECT2_Y(rectangle2_ys[1924]), .RECT2_WIDTH(rectangle2_widths[1924]), .RECT2_HEIGHT(rectangle2_heights[1924]), .RECT2_WEIGHT(rectangle2_weights[1924]), .RECT3_X(rectangle3_xs[1924]), .RECT3_Y(rectangle3_ys[1924]), .RECT3_WIDTH(rectangle3_widths[1924]), .RECT3_HEIGHT(rectangle3_heights[1924]), .RECT3_WEIGHT(rectangle3_weights[1924]), .FEAT_THRES(feature_thresholds[1924]), .FEAT_ABOVE(feature_aboves[1924]), .FEAT_BELOW(feature_belows[1924])) ac1924(.scan_win(scan_win1924), .scan_win_std_dev(scan_win_std_dev[1924]), .feature_accum(feature_accums[1924]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1925]), .RECT1_Y(rectangle1_ys[1925]), .RECT1_WIDTH(rectangle1_widths[1925]), .RECT1_HEIGHT(rectangle1_heights[1925]), .RECT1_WEIGHT(rectangle1_weights[1925]), .RECT2_X(rectangle2_xs[1925]), .RECT2_Y(rectangle2_ys[1925]), .RECT2_WIDTH(rectangle2_widths[1925]), .RECT2_HEIGHT(rectangle2_heights[1925]), .RECT2_WEIGHT(rectangle2_weights[1925]), .RECT3_X(rectangle3_xs[1925]), .RECT3_Y(rectangle3_ys[1925]), .RECT3_WIDTH(rectangle3_widths[1925]), .RECT3_HEIGHT(rectangle3_heights[1925]), .RECT3_WEIGHT(rectangle3_weights[1925]), .FEAT_THRES(feature_thresholds[1925]), .FEAT_ABOVE(feature_aboves[1925]), .FEAT_BELOW(feature_belows[1925])) ac1925(.scan_win(scan_win1925), .scan_win_std_dev(scan_win_std_dev[1925]), .feature_accum(feature_accums[1925]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1926]), .RECT1_Y(rectangle1_ys[1926]), .RECT1_WIDTH(rectangle1_widths[1926]), .RECT1_HEIGHT(rectangle1_heights[1926]), .RECT1_WEIGHT(rectangle1_weights[1926]), .RECT2_X(rectangle2_xs[1926]), .RECT2_Y(rectangle2_ys[1926]), .RECT2_WIDTH(rectangle2_widths[1926]), .RECT2_HEIGHT(rectangle2_heights[1926]), .RECT2_WEIGHT(rectangle2_weights[1926]), .RECT3_X(rectangle3_xs[1926]), .RECT3_Y(rectangle3_ys[1926]), .RECT3_WIDTH(rectangle3_widths[1926]), .RECT3_HEIGHT(rectangle3_heights[1926]), .RECT3_WEIGHT(rectangle3_weights[1926]), .FEAT_THRES(feature_thresholds[1926]), .FEAT_ABOVE(feature_aboves[1926]), .FEAT_BELOW(feature_belows[1926])) ac1926(.scan_win(scan_win1926), .scan_win_std_dev(scan_win_std_dev[1926]), .feature_accum(feature_accums[1926]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1927]), .RECT1_Y(rectangle1_ys[1927]), .RECT1_WIDTH(rectangle1_widths[1927]), .RECT1_HEIGHT(rectangle1_heights[1927]), .RECT1_WEIGHT(rectangle1_weights[1927]), .RECT2_X(rectangle2_xs[1927]), .RECT2_Y(rectangle2_ys[1927]), .RECT2_WIDTH(rectangle2_widths[1927]), .RECT2_HEIGHT(rectangle2_heights[1927]), .RECT2_WEIGHT(rectangle2_weights[1927]), .RECT3_X(rectangle3_xs[1927]), .RECT3_Y(rectangle3_ys[1927]), .RECT3_WIDTH(rectangle3_widths[1927]), .RECT3_HEIGHT(rectangle3_heights[1927]), .RECT3_WEIGHT(rectangle3_weights[1927]), .FEAT_THRES(feature_thresholds[1927]), .FEAT_ABOVE(feature_aboves[1927]), .FEAT_BELOW(feature_belows[1927])) ac1927(.scan_win(scan_win1927), .scan_win_std_dev(scan_win_std_dev[1927]), .feature_accum(feature_accums[1927]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1928]), .RECT1_Y(rectangle1_ys[1928]), .RECT1_WIDTH(rectangle1_widths[1928]), .RECT1_HEIGHT(rectangle1_heights[1928]), .RECT1_WEIGHT(rectangle1_weights[1928]), .RECT2_X(rectangle2_xs[1928]), .RECT2_Y(rectangle2_ys[1928]), .RECT2_WIDTH(rectangle2_widths[1928]), .RECT2_HEIGHT(rectangle2_heights[1928]), .RECT2_WEIGHT(rectangle2_weights[1928]), .RECT3_X(rectangle3_xs[1928]), .RECT3_Y(rectangle3_ys[1928]), .RECT3_WIDTH(rectangle3_widths[1928]), .RECT3_HEIGHT(rectangle3_heights[1928]), .RECT3_WEIGHT(rectangle3_weights[1928]), .FEAT_THRES(feature_thresholds[1928]), .FEAT_ABOVE(feature_aboves[1928]), .FEAT_BELOW(feature_belows[1928])) ac1928(.scan_win(scan_win1928), .scan_win_std_dev(scan_win_std_dev[1928]), .feature_accum(feature_accums[1928]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1929]), .RECT1_Y(rectangle1_ys[1929]), .RECT1_WIDTH(rectangle1_widths[1929]), .RECT1_HEIGHT(rectangle1_heights[1929]), .RECT1_WEIGHT(rectangle1_weights[1929]), .RECT2_X(rectangle2_xs[1929]), .RECT2_Y(rectangle2_ys[1929]), .RECT2_WIDTH(rectangle2_widths[1929]), .RECT2_HEIGHT(rectangle2_heights[1929]), .RECT2_WEIGHT(rectangle2_weights[1929]), .RECT3_X(rectangle3_xs[1929]), .RECT3_Y(rectangle3_ys[1929]), .RECT3_WIDTH(rectangle3_widths[1929]), .RECT3_HEIGHT(rectangle3_heights[1929]), .RECT3_WEIGHT(rectangle3_weights[1929]), .FEAT_THRES(feature_thresholds[1929]), .FEAT_ABOVE(feature_aboves[1929]), .FEAT_BELOW(feature_belows[1929])) ac1929(.scan_win(scan_win1929), .scan_win_std_dev(scan_win_std_dev[1929]), .feature_accum(feature_accums[1929]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1930]), .RECT1_Y(rectangle1_ys[1930]), .RECT1_WIDTH(rectangle1_widths[1930]), .RECT1_HEIGHT(rectangle1_heights[1930]), .RECT1_WEIGHT(rectangle1_weights[1930]), .RECT2_X(rectangle2_xs[1930]), .RECT2_Y(rectangle2_ys[1930]), .RECT2_WIDTH(rectangle2_widths[1930]), .RECT2_HEIGHT(rectangle2_heights[1930]), .RECT2_WEIGHT(rectangle2_weights[1930]), .RECT3_X(rectangle3_xs[1930]), .RECT3_Y(rectangle3_ys[1930]), .RECT3_WIDTH(rectangle3_widths[1930]), .RECT3_HEIGHT(rectangle3_heights[1930]), .RECT3_WEIGHT(rectangle3_weights[1930]), .FEAT_THRES(feature_thresholds[1930]), .FEAT_ABOVE(feature_aboves[1930]), .FEAT_BELOW(feature_belows[1930])) ac1930(.scan_win(scan_win1930), .scan_win_std_dev(scan_win_std_dev[1930]), .feature_accum(feature_accums[1930]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1931]), .RECT1_Y(rectangle1_ys[1931]), .RECT1_WIDTH(rectangle1_widths[1931]), .RECT1_HEIGHT(rectangle1_heights[1931]), .RECT1_WEIGHT(rectangle1_weights[1931]), .RECT2_X(rectangle2_xs[1931]), .RECT2_Y(rectangle2_ys[1931]), .RECT2_WIDTH(rectangle2_widths[1931]), .RECT2_HEIGHT(rectangle2_heights[1931]), .RECT2_WEIGHT(rectangle2_weights[1931]), .RECT3_X(rectangle3_xs[1931]), .RECT3_Y(rectangle3_ys[1931]), .RECT3_WIDTH(rectangle3_widths[1931]), .RECT3_HEIGHT(rectangle3_heights[1931]), .RECT3_WEIGHT(rectangle3_weights[1931]), .FEAT_THRES(feature_thresholds[1931]), .FEAT_ABOVE(feature_aboves[1931]), .FEAT_BELOW(feature_belows[1931])) ac1931(.scan_win(scan_win1931), .scan_win_std_dev(scan_win_std_dev[1931]), .feature_accum(feature_accums[1931]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1932]), .RECT1_Y(rectangle1_ys[1932]), .RECT1_WIDTH(rectangle1_widths[1932]), .RECT1_HEIGHT(rectangle1_heights[1932]), .RECT1_WEIGHT(rectangle1_weights[1932]), .RECT2_X(rectangle2_xs[1932]), .RECT2_Y(rectangle2_ys[1932]), .RECT2_WIDTH(rectangle2_widths[1932]), .RECT2_HEIGHT(rectangle2_heights[1932]), .RECT2_WEIGHT(rectangle2_weights[1932]), .RECT3_X(rectangle3_xs[1932]), .RECT3_Y(rectangle3_ys[1932]), .RECT3_WIDTH(rectangle3_widths[1932]), .RECT3_HEIGHT(rectangle3_heights[1932]), .RECT3_WEIGHT(rectangle3_weights[1932]), .FEAT_THRES(feature_thresholds[1932]), .FEAT_ABOVE(feature_aboves[1932]), .FEAT_BELOW(feature_belows[1932])) ac1932(.scan_win(scan_win1932), .scan_win_std_dev(scan_win_std_dev[1932]), .feature_accum(feature_accums[1932]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1933]), .RECT1_Y(rectangle1_ys[1933]), .RECT1_WIDTH(rectangle1_widths[1933]), .RECT1_HEIGHT(rectangle1_heights[1933]), .RECT1_WEIGHT(rectangle1_weights[1933]), .RECT2_X(rectangle2_xs[1933]), .RECT2_Y(rectangle2_ys[1933]), .RECT2_WIDTH(rectangle2_widths[1933]), .RECT2_HEIGHT(rectangle2_heights[1933]), .RECT2_WEIGHT(rectangle2_weights[1933]), .RECT3_X(rectangle3_xs[1933]), .RECT3_Y(rectangle3_ys[1933]), .RECT3_WIDTH(rectangle3_widths[1933]), .RECT3_HEIGHT(rectangle3_heights[1933]), .RECT3_WEIGHT(rectangle3_weights[1933]), .FEAT_THRES(feature_thresholds[1933]), .FEAT_ABOVE(feature_aboves[1933]), .FEAT_BELOW(feature_belows[1933])) ac1933(.scan_win(scan_win1933), .scan_win_std_dev(scan_win_std_dev[1933]), .feature_accum(feature_accums[1933]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1934]), .RECT1_Y(rectangle1_ys[1934]), .RECT1_WIDTH(rectangle1_widths[1934]), .RECT1_HEIGHT(rectangle1_heights[1934]), .RECT1_WEIGHT(rectangle1_weights[1934]), .RECT2_X(rectangle2_xs[1934]), .RECT2_Y(rectangle2_ys[1934]), .RECT2_WIDTH(rectangle2_widths[1934]), .RECT2_HEIGHT(rectangle2_heights[1934]), .RECT2_WEIGHT(rectangle2_weights[1934]), .RECT3_X(rectangle3_xs[1934]), .RECT3_Y(rectangle3_ys[1934]), .RECT3_WIDTH(rectangle3_widths[1934]), .RECT3_HEIGHT(rectangle3_heights[1934]), .RECT3_WEIGHT(rectangle3_weights[1934]), .FEAT_THRES(feature_thresholds[1934]), .FEAT_ABOVE(feature_aboves[1934]), .FEAT_BELOW(feature_belows[1934])) ac1934(.scan_win(scan_win1934), .scan_win_std_dev(scan_win_std_dev[1934]), .feature_accum(feature_accums[1934]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1935]), .RECT1_Y(rectangle1_ys[1935]), .RECT1_WIDTH(rectangle1_widths[1935]), .RECT1_HEIGHT(rectangle1_heights[1935]), .RECT1_WEIGHT(rectangle1_weights[1935]), .RECT2_X(rectangle2_xs[1935]), .RECT2_Y(rectangle2_ys[1935]), .RECT2_WIDTH(rectangle2_widths[1935]), .RECT2_HEIGHT(rectangle2_heights[1935]), .RECT2_WEIGHT(rectangle2_weights[1935]), .RECT3_X(rectangle3_xs[1935]), .RECT3_Y(rectangle3_ys[1935]), .RECT3_WIDTH(rectangle3_widths[1935]), .RECT3_HEIGHT(rectangle3_heights[1935]), .RECT3_WEIGHT(rectangle3_weights[1935]), .FEAT_THRES(feature_thresholds[1935]), .FEAT_ABOVE(feature_aboves[1935]), .FEAT_BELOW(feature_belows[1935])) ac1935(.scan_win(scan_win1935), .scan_win_std_dev(scan_win_std_dev[1935]), .feature_accum(feature_accums[1935]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1936]), .RECT1_Y(rectangle1_ys[1936]), .RECT1_WIDTH(rectangle1_widths[1936]), .RECT1_HEIGHT(rectangle1_heights[1936]), .RECT1_WEIGHT(rectangle1_weights[1936]), .RECT2_X(rectangle2_xs[1936]), .RECT2_Y(rectangle2_ys[1936]), .RECT2_WIDTH(rectangle2_widths[1936]), .RECT2_HEIGHT(rectangle2_heights[1936]), .RECT2_WEIGHT(rectangle2_weights[1936]), .RECT3_X(rectangle3_xs[1936]), .RECT3_Y(rectangle3_ys[1936]), .RECT3_WIDTH(rectangle3_widths[1936]), .RECT3_HEIGHT(rectangle3_heights[1936]), .RECT3_WEIGHT(rectangle3_weights[1936]), .FEAT_THRES(feature_thresholds[1936]), .FEAT_ABOVE(feature_aboves[1936]), .FEAT_BELOW(feature_belows[1936])) ac1936(.scan_win(scan_win1936), .scan_win_std_dev(scan_win_std_dev[1936]), .feature_accum(feature_accums[1936]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1937]), .RECT1_Y(rectangle1_ys[1937]), .RECT1_WIDTH(rectangle1_widths[1937]), .RECT1_HEIGHT(rectangle1_heights[1937]), .RECT1_WEIGHT(rectangle1_weights[1937]), .RECT2_X(rectangle2_xs[1937]), .RECT2_Y(rectangle2_ys[1937]), .RECT2_WIDTH(rectangle2_widths[1937]), .RECT2_HEIGHT(rectangle2_heights[1937]), .RECT2_WEIGHT(rectangle2_weights[1937]), .RECT3_X(rectangle3_xs[1937]), .RECT3_Y(rectangle3_ys[1937]), .RECT3_WIDTH(rectangle3_widths[1937]), .RECT3_HEIGHT(rectangle3_heights[1937]), .RECT3_WEIGHT(rectangle3_weights[1937]), .FEAT_THRES(feature_thresholds[1937]), .FEAT_ABOVE(feature_aboves[1937]), .FEAT_BELOW(feature_belows[1937])) ac1937(.scan_win(scan_win1937), .scan_win_std_dev(scan_win_std_dev[1937]), .feature_accum(feature_accums[1937]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1938]), .RECT1_Y(rectangle1_ys[1938]), .RECT1_WIDTH(rectangle1_widths[1938]), .RECT1_HEIGHT(rectangle1_heights[1938]), .RECT1_WEIGHT(rectangle1_weights[1938]), .RECT2_X(rectangle2_xs[1938]), .RECT2_Y(rectangle2_ys[1938]), .RECT2_WIDTH(rectangle2_widths[1938]), .RECT2_HEIGHT(rectangle2_heights[1938]), .RECT2_WEIGHT(rectangle2_weights[1938]), .RECT3_X(rectangle3_xs[1938]), .RECT3_Y(rectangle3_ys[1938]), .RECT3_WIDTH(rectangle3_widths[1938]), .RECT3_HEIGHT(rectangle3_heights[1938]), .RECT3_WEIGHT(rectangle3_weights[1938]), .FEAT_THRES(feature_thresholds[1938]), .FEAT_ABOVE(feature_aboves[1938]), .FEAT_BELOW(feature_belows[1938])) ac1938(.scan_win(scan_win1938), .scan_win_std_dev(scan_win_std_dev[1938]), .feature_accum(feature_accums[1938]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1939]), .RECT1_Y(rectangle1_ys[1939]), .RECT1_WIDTH(rectangle1_widths[1939]), .RECT1_HEIGHT(rectangle1_heights[1939]), .RECT1_WEIGHT(rectangle1_weights[1939]), .RECT2_X(rectangle2_xs[1939]), .RECT2_Y(rectangle2_ys[1939]), .RECT2_WIDTH(rectangle2_widths[1939]), .RECT2_HEIGHT(rectangle2_heights[1939]), .RECT2_WEIGHT(rectangle2_weights[1939]), .RECT3_X(rectangle3_xs[1939]), .RECT3_Y(rectangle3_ys[1939]), .RECT3_WIDTH(rectangle3_widths[1939]), .RECT3_HEIGHT(rectangle3_heights[1939]), .RECT3_WEIGHT(rectangle3_weights[1939]), .FEAT_THRES(feature_thresholds[1939]), .FEAT_ABOVE(feature_aboves[1939]), .FEAT_BELOW(feature_belows[1939])) ac1939(.scan_win(scan_win1939), .scan_win_std_dev(scan_win_std_dev[1939]), .feature_accum(feature_accums[1939]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1940]), .RECT1_Y(rectangle1_ys[1940]), .RECT1_WIDTH(rectangle1_widths[1940]), .RECT1_HEIGHT(rectangle1_heights[1940]), .RECT1_WEIGHT(rectangle1_weights[1940]), .RECT2_X(rectangle2_xs[1940]), .RECT2_Y(rectangle2_ys[1940]), .RECT2_WIDTH(rectangle2_widths[1940]), .RECT2_HEIGHT(rectangle2_heights[1940]), .RECT2_WEIGHT(rectangle2_weights[1940]), .RECT3_X(rectangle3_xs[1940]), .RECT3_Y(rectangle3_ys[1940]), .RECT3_WIDTH(rectangle3_widths[1940]), .RECT3_HEIGHT(rectangle3_heights[1940]), .RECT3_WEIGHT(rectangle3_weights[1940]), .FEAT_THRES(feature_thresholds[1940]), .FEAT_ABOVE(feature_aboves[1940]), .FEAT_BELOW(feature_belows[1940])) ac1940(.scan_win(scan_win1940), .scan_win_std_dev(scan_win_std_dev[1940]), .feature_accum(feature_accums[1940]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1941]), .RECT1_Y(rectangle1_ys[1941]), .RECT1_WIDTH(rectangle1_widths[1941]), .RECT1_HEIGHT(rectangle1_heights[1941]), .RECT1_WEIGHT(rectangle1_weights[1941]), .RECT2_X(rectangle2_xs[1941]), .RECT2_Y(rectangle2_ys[1941]), .RECT2_WIDTH(rectangle2_widths[1941]), .RECT2_HEIGHT(rectangle2_heights[1941]), .RECT2_WEIGHT(rectangle2_weights[1941]), .RECT3_X(rectangle3_xs[1941]), .RECT3_Y(rectangle3_ys[1941]), .RECT3_WIDTH(rectangle3_widths[1941]), .RECT3_HEIGHT(rectangle3_heights[1941]), .RECT3_WEIGHT(rectangle3_weights[1941]), .FEAT_THRES(feature_thresholds[1941]), .FEAT_ABOVE(feature_aboves[1941]), .FEAT_BELOW(feature_belows[1941])) ac1941(.scan_win(scan_win1941), .scan_win_std_dev(scan_win_std_dev[1941]), .feature_accum(feature_accums[1941]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1942]), .RECT1_Y(rectangle1_ys[1942]), .RECT1_WIDTH(rectangle1_widths[1942]), .RECT1_HEIGHT(rectangle1_heights[1942]), .RECT1_WEIGHT(rectangle1_weights[1942]), .RECT2_X(rectangle2_xs[1942]), .RECT2_Y(rectangle2_ys[1942]), .RECT2_WIDTH(rectangle2_widths[1942]), .RECT2_HEIGHT(rectangle2_heights[1942]), .RECT2_WEIGHT(rectangle2_weights[1942]), .RECT3_X(rectangle3_xs[1942]), .RECT3_Y(rectangle3_ys[1942]), .RECT3_WIDTH(rectangle3_widths[1942]), .RECT3_HEIGHT(rectangle3_heights[1942]), .RECT3_WEIGHT(rectangle3_weights[1942]), .FEAT_THRES(feature_thresholds[1942]), .FEAT_ABOVE(feature_aboves[1942]), .FEAT_BELOW(feature_belows[1942])) ac1942(.scan_win(scan_win1942), .scan_win_std_dev(scan_win_std_dev[1942]), .feature_accum(feature_accums[1942]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1943]), .RECT1_Y(rectangle1_ys[1943]), .RECT1_WIDTH(rectangle1_widths[1943]), .RECT1_HEIGHT(rectangle1_heights[1943]), .RECT1_WEIGHT(rectangle1_weights[1943]), .RECT2_X(rectangle2_xs[1943]), .RECT2_Y(rectangle2_ys[1943]), .RECT2_WIDTH(rectangle2_widths[1943]), .RECT2_HEIGHT(rectangle2_heights[1943]), .RECT2_WEIGHT(rectangle2_weights[1943]), .RECT3_X(rectangle3_xs[1943]), .RECT3_Y(rectangle3_ys[1943]), .RECT3_WIDTH(rectangle3_widths[1943]), .RECT3_HEIGHT(rectangle3_heights[1943]), .RECT3_WEIGHT(rectangle3_weights[1943]), .FEAT_THRES(feature_thresholds[1943]), .FEAT_ABOVE(feature_aboves[1943]), .FEAT_BELOW(feature_belows[1943])) ac1943(.scan_win(scan_win1943), .scan_win_std_dev(scan_win_std_dev[1943]), .feature_accum(feature_accums[1943]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1944]), .RECT1_Y(rectangle1_ys[1944]), .RECT1_WIDTH(rectangle1_widths[1944]), .RECT1_HEIGHT(rectangle1_heights[1944]), .RECT1_WEIGHT(rectangle1_weights[1944]), .RECT2_X(rectangle2_xs[1944]), .RECT2_Y(rectangle2_ys[1944]), .RECT2_WIDTH(rectangle2_widths[1944]), .RECT2_HEIGHT(rectangle2_heights[1944]), .RECT2_WEIGHT(rectangle2_weights[1944]), .RECT3_X(rectangle3_xs[1944]), .RECT3_Y(rectangle3_ys[1944]), .RECT3_WIDTH(rectangle3_widths[1944]), .RECT3_HEIGHT(rectangle3_heights[1944]), .RECT3_WEIGHT(rectangle3_weights[1944]), .FEAT_THRES(feature_thresholds[1944]), .FEAT_ABOVE(feature_aboves[1944]), .FEAT_BELOW(feature_belows[1944])) ac1944(.scan_win(scan_win1944), .scan_win_std_dev(scan_win_std_dev[1944]), .feature_accum(feature_accums[1944]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1945]), .RECT1_Y(rectangle1_ys[1945]), .RECT1_WIDTH(rectangle1_widths[1945]), .RECT1_HEIGHT(rectangle1_heights[1945]), .RECT1_WEIGHT(rectangle1_weights[1945]), .RECT2_X(rectangle2_xs[1945]), .RECT2_Y(rectangle2_ys[1945]), .RECT2_WIDTH(rectangle2_widths[1945]), .RECT2_HEIGHT(rectangle2_heights[1945]), .RECT2_WEIGHT(rectangle2_weights[1945]), .RECT3_X(rectangle3_xs[1945]), .RECT3_Y(rectangle3_ys[1945]), .RECT3_WIDTH(rectangle3_widths[1945]), .RECT3_HEIGHT(rectangle3_heights[1945]), .RECT3_WEIGHT(rectangle3_weights[1945]), .FEAT_THRES(feature_thresholds[1945]), .FEAT_ABOVE(feature_aboves[1945]), .FEAT_BELOW(feature_belows[1945])) ac1945(.scan_win(scan_win1945), .scan_win_std_dev(scan_win_std_dev[1945]), .feature_accum(feature_accums[1945]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1946]), .RECT1_Y(rectangle1_ys[1946]), .RECT1_WIDTH(rectangle1_widths[1946]), .RECT1_HEIGHT(rectangle1_heights[1946]), .RECT1_WEIGHT(rectangle1_weights[1946]), .RECT2_X(rectangle2_xs[1946]), .RECT2_Y(rectangle2_ys[1946]), .RECT2_WIDTH(rectangle2_widths[1946]), .RECT2_HEIGHT(rectangle2_heights[1946]), .RECT2_WEIGHT(rectangle2_weights[1946]), .RECT3_X(rectangle3_xs[1946]), .RECT3_Y(rectangle3_ys[1946]), .RECT3_WIDTH(rectangle3_widths[1946]), .RECT3_HEIGHT(rectangle3_heights[1946]), .RECT3_WEIGHT(rectangle3_weights[1946]), .FEAT_THRES(feature_thresholds[1946]), .FEAT_ABOVE(feature_aboves[1946]), .FEAT_BELOW(feature_belows[1946])) ac1946(.scan_win(scan_win1946), .scan_win_std_dev(scan_win_std_dev[1946]), .feature_accum(feature_accums[1946]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1947]), .RECT1_Y(rectangle1_ys[1947]), .RECT1_WIDTH(rectangle1_widths[1947]), .RECT1_HEIGHT(rectangle1_heights[1947]), .RECT1_WEIGHT(rectangle1_weights[1947]), .RECT2_X(rectangle2_xs[1947]), .RECT2_Y(rectangle2_ys[1947]), .RECT2_WIDTH(rectangle2_widths[1947]), .RECT2_HEIGHT(rectangle2_heights[1947]), .RECT2_WEIGHT(rectangle2_weights[1947]), .RECT3_X(rectangle3_xs[1947]), .RECT3_Y(rectangle3_ys[1947]), .RECT3_WIDTH(rectangle3_widths[1947]), .RECT3_HEIGHT(rectangle3_heights[1947]), .RECT3_WEIGHT(rectangle3_weights[1947]), .FEAT_THRES(feature_thresholds[1947]), .FEAT_ABOVE(feature_aboves[1947]), .FEAT_BELOW(feature_belows[1947])) ac1947(.scan_win(scan_win1947), .scan_win_std_dev(scan_win_std_dev[1947]), .feature_accum(feature_accums[1947]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1948]), .RECT1_Y(rectangle1_ys[1948]), .RECT1_WIDTH(rectangle1_widths[1948]), .RECT1_HEIGHT(rectangle1_heights[1948]), .RECT1_WEIGHT(rectangle1_weights[1948]), .RECT2_X(rectangle2_xs[1948]), .RECT2_Y(rectangle2_ys[1948]), .RECT2_WIDTH(rectangle2_widths[1948]), .RECT2_HEIGHT(rectangle2_heights[1948]), .RECT2_WEIGHT(rectangle2_weights[1948]), .RECT3_X(rectangle3_xs[1948]), .RECT3_Y(rectangle3_ys[1948]), .RECT3_WIDTH(rectangle3_widths[1948]), .RECT3_HEIGHT(rectangle3_heights[1948]), .RECT3_WEIGHT(rectangle3_weights[1948]), .FEAT_THRES(feature_thresholds[1948]), .FEAT_ABOVE(feature_aboves[1948]), .FEAT_BELOW(feature_belows[1948])) ac1948(.scan_win(scan_win1948), .scan_win_std_dev(scan_win_std_dev[1948]), .feature_accum(feature_accums[1948]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1949]), .RECT1_Y(rectangle1_ys[1949]), .RECT1_WIDTH(rectangle1_widths[1949]), .RECT1_HEIGHT(rectangle1_heights[1949]), .RECT1_WEIGHT(rectangle1_weights[1949]), .RECT2_X(rectangle2_xs[1949]), .RECT2_Y(rectangle2_ys[1949]), .RECT2_WIDTH(rectangle2_widths[1949]), .RECT2_HEIGHT(rectangle2_heights[1949]), .RECT2_WEIGHT(rectangle2_weights[1949]), .RECT3_X(rectangle3_xs[1949]), .RECT3_Y(rectangle3_ys[1949]), .RECT3_WIDTH(rectangle3_widths[1949]), .RECT3_HEIGHT(rectangle3_heights[1949]), .RECT3_WEIGHT(rectangle3_weights[1949]), .FEAT_THRES(feature_thresholds[1949]), .FEAT_ABOVE(feature_aboves[1949]), .FEAT_BELOW(feature_belows[1949])) ac1949(.scan_win(scan_win1949), .scan_win_std_dev(scan_win_std_dev[1949]), .feature_accum(feature_accums[1949]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1950]), .RECT1_Y(rectangle1_ys[1950]), .RECT1_WIDTH(rectangle1_widths[1950]), .RECT1_HEIGHT(rectangle1_heights[1950]), .RECT1_WEIGHT(rectangle1_weights[1950]), .RECT2_X(rectangle2_xs[1950]), .RECT2_Y(rectangle2_ys[1950]), .RECT2_WIDTH(rectangle2_widths[1950]), .RECT2_HEIGHT(rectangle2_heights[1950]), .RECT2_WEIGHT(rectangle2_weights[1950]), .RECT3_X(rectangle3_xs[1950]), .RECT3_Y(rectangle3_ys[1950]), .RECT3_WIDTH(rectangle3_widths[1950]), .RECT3_HEIGHT(rectangle3_heights[1950]), .RECT3_WEIGHT(rectangle3_weights[1950]), .FEAT_THRES(feature_thresholds[1950]), .FEAT_ABOVE(feature_aboves[1950]), .FEAT_BELOW(feature_belows[1950])) ac1950(.scan_win(scan_win1950), .scan_win_std_dev(scan_win_std_dev[1950]), .feature_accum(feature_accums[1950]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1951]), .RECT1_Y(rectangle1_ys[1951]), .RECT1_WIDTH(rectangle1_widths[1951]), .RECT1_HEIGHT(rectangle1_heights[1951]), .RECT1_WEIGHT(rectangle1_weights[1951]), .RECT2_X(rectangle2_xs[1951]), .RECT2_Y(rectangle2_ys[1951]), .RECT2_WIDTH(rectangle2_widths[1951]), .RECT2_HEIGHT(rectangle2_heights[1951]), .RECT2_WEIGHT(rectangle2_weights[1951]), .RECT3_X(rectangle3_xs[1951]), .RECT3_Y(rectangle3_ys[1951]), .RECT3_WIDTH(rectangle3_widths[1951]), .RECT3_HEIGHT(rectangle3_heights[1951]), .RECT3_WEIGHT(rectangle3_weights[1951]), .FEAT_THRES(feature_thresholds[1951]), .FEAT_ABOVE(feature_aboves[1951]), .FEAT_BELOW(feature_belows[1951])) ac1951(.scan_win(scan_win1951), .scan_win_std_dev(scan_win_std_dev[1951]), .feature_accum(feature_accums[1951]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1952]), .RECT1_Y(rectangle1_ys[1952]), .RECT1_WIDTH(rectangle1_widths[1952]), .RECT1_HEIGHT(rectangle1_heights[1952]), .RECT1_WEIGHT(rectangle1_weights[1952]), .RECT2_X(rectangle2_xs[1952]), .RECT2_Y(rectangle2_ys[1952]), .RECT2_WIDTH(rectangle2_widths[1952]), .RECT2_HEIGHT(rectangle2_heights[1952]), .RECT2_WEIGHT(rectangle2_weights[1952]), .RECT3_X(rectangle3_xs[1952]), .RECT3_Y(rectangle3_ys[1952]), .RECT3_WIDTH(rectangle3_widths[1952]), .RECT3_HEIGHT(rectangle3_heights[1952]), .RECT3_WEIGHT(rectangle3_weights[1952]), .FEAT_THRES(feature_thresholds[1952]), .FEAT_ABOVE(feature_aboves[1952]), .FEAT_BELOW(feature_belows[1952])) ac1952(.scan_win(scan_win1952), .scan_win_std_dev(scan_win_std_dev[1952]), .feature_accum(feature_accums[1952]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1953]), .RECT1_Y(rectangle1_ys[1953]), .RECT1_WIDTH(rectangle1_widths[1953]), .RECT1_HEIGHT(rectangle1_heights[1953]), .RECT1_WEIGHT(rectangle1_weights[1953]), .RECT2_X(rectangle2_xs[1953]), .RECT2_Y(rectangle2_ys[1953]), .RECT2_WIDTH(rectangle2_widths[1953]), .RECT2_HEIGHT(rectangle2_heights[1953]), .RECT2_WEIGHT(rectangle2_weights[1953]), .RECT3_X(rectangle3_xs[1953]), .RECT3_Y(rectangle3_ys[1953]), .RECT3_WIDTH(rectangle3_widths[1953]), .RECT3_HEIGHT(rectangle3_heights[1953]), .RECT3_WEIGHT(rectangle3_weights[1953]), .FEAT_THRES(feature_thresholds[1953]), .FEAT_ABOVE(feature_aboves[1953]), .FEAT_BELOW(feature_belows[1953])) ac1953(.scan_win(scan_win1953), .scan_win_std_dev(scan_win_std_dev[1953]), .feature_accum(feature_accums[1953]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1954]), .RECT1_Y(rectangle1_ys[1954]), .RECT1_WIDTH(rectangle1_widths[1954]), .RECT1_HEIGHT(rectangle1_heights[1954]), .RECT1_WEIGHT(rectangle1_weights[1954]), .RECT2_X(rectangle2_xs[1954]), .RECT2_Y(rectangle2_ys[1954]), .RECT2_WIDTH(rectangle2_widths[1954]), .RECT2_HEIGHT(rectangle2_heights[1954]), .RECT2_WEIGHT(rectangle2_weights[1954]), .RECT3_X(rectangle3_xs[1954]), .RECT3_Y(rectangle3_ys[1954]), .RECT3_WIDTH(rectangle3_widths[1954]), .RECT3_HEIGHT(rectangle3_heights[1954]), .RECT3_WEIGHT(rectangle3_weights[1954]), .FEAT_THRES(feature_thresholds[1954]), .FEAT_ABOVE(feature_aboves[1954]), .FEAT_BELOW(feature_belows[1954])) ac1954(.scan_win(scan_win1954), .scan_win_std_dev(scan_win_std_dev[1954]), .feature_accum(feature_accums[1954]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1955]), .RECT1_Y(rectangle1_ys[1955]), .RECT1_WIDTH(rectangle1_widths[1955]), .RECT1_HEIGHT(rectangle1_heights[1955]), .RECT1_WEIGHT(rectangle1_weights[1955]), .RECT2_X(rectangle2_xs[1955]), .RECT2_Y(rectangle2_ys[1955]), .RECT2_WIDTH(rectangle2_widths[1955]), .RECT2_HEIGHT(rectangle2_heights[1955]), .RECT2_WEIGHT(rectangle2_weights[1955]), .RECT3_X(rectangle3_xs[1955]), .RECT3_Y(rectangle3_ys[1955]), .RECT3_WIDTH(rectangle3_widths[1955]), .RECT3_HEIGHT(rectangle3_heights[1955]), .RECT3_WEIGHT(rectangle3_weights[1955]), .FEAT_THRES(feature_thresholds[1955]), .FEAT_ABOVE(feature_aboves[1955]), .FEAT_BELOW(feature_belows[1955])) ac1955(.scan_win(scan_win1955), .scan_win_std_dev(scan_win_std_dev[1955]), .feature_accum(feature_accums[1955]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1956]), .RECT1_Y(rectangle1_ys[1956]), .RECT1_WIDTH(rectangle1_widths[1956]), .RECT1_HEIGHT(rectangle1_heights[1956]), .RECT1_WEIGHT(rectangle1_weights[1956]), .RECT2_X(rectangle2_xs[1956]), .RECT2_Y(rectangle2_ys[1956]), .RECT2_WIDTH(rectangle2_widths[1956]), .RECT2_HEIGHT(rectangle2_heights[1956]), .RECT2_WEIGHT(rectangle2_weights[1956]), .RECT3_X(rectangle3_xs[1956]), .RECT3_Y(rectangle3_ys[1956]), .RECT3_WIDTH(rectangle3_widths[1956]), .RECT3_HEIGHT(rectangle3_heights[1956]), .RECT3_WEIGHT(rectangle3_weights[1956]), .FEAT_THRES(feature_thresholds[1956]), .FEAT_ABOVE(feature_aboves[1956]), .FEAT_BELOW(feature_belows[1956])) ac1956(.scan_win(scan_win1956), .scan_win_std_dev(scan_win_std_dev[1956]), .feature_accum(feature_accums[1956]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1957]), .RECT1_Y(rectangle1_ys[1957]), .RECT1_WIDTH(rectangle1_widths[1957]), .RECT1_HEIGHT(rectangle1_heights[1957]), .RECT1_WEIGHT(rectangle1_weights[1957]), .RECT2_X(rectangle2_xs[1957]), .RECT2_Y(rectangle2_ys[1957]), .RECT2_WIDTH(rectangle2_widths[1957]), .RECT2_HEIGHT(rectangle2_heights[1957]), .RECT2_WEIGHT(rectangle2_weights[1957]), .RECT3_X(rectangle3_xs[1957]), .RECT3_Y(rectangle3_ys[1957]), .RECT3_WIDTH(rectangle3_widths[1957]), .RECT3_HEIGHT(rectangle3_heights[1957]), .RECT3_WEIGHT(rectangle3_weights[1957]), .FEAT_THRES(feature_thresholds[1957]), .FEAT_ABOVE(feature_aboves[1957]), .FEAT_BELOW(feature_belows[1957])) ac1957(.scan_win(scan_win1957), .scan_win_std_dev(scan_win_std_dev[1957]), .feature_accum(feature_accums[1957]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1958]), .RECT1_Y(rectangle1_ys[1958]), .RECT1_WIDTH(rectangle1_widths[1958]), .RECT1_HEIGHT(rectangle1_heights[1958]), .RECT1_WEIGHT(rectangle1_weights[1958]), .RECT2_X(rectangle2_xs[1958]), .RECT2_Y(rectangle2_ys[1958]), .RECT2_WIDTH(rectangle2_widths[1958]), .RECT2_HEIGHT(rectangle2_heights[1958]), .RECT2_WEIGHT(rectangle2_weights[1958]), .RECT3_X(rectangle3_xs[1958]), .RECT3_Y(rectangle3_ys[1958]), .RECT3_WIDTH(rectangle3_widths[1958]), .RECT3_HEIGHT(rectangle3_heights[1958]), .RECT3_WEIGHT(rectangle3_weights[1958]), .FEAT_THRES(feature_thresholds[1958]), .FEAT_ABOVE(feature_aboves[1958]), .FEAT_BELOW(feature_belows[1958])) ac1958(.scan_win(scan_win1958), .scan_win_std_dev(scan_win_std_dev[1958]), .feature_accum(feature_accums[1958]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1959]), .RECT1_Y(rectangle1_ys[1959]), .RECT1_WIDTH(rectangle1_widths[1959]), .RECT1_HEIGHT(rectangle1_heights[1959]), .RECT1_WEIGHT(rectangle1_weights[1959]), .RECT2_X(rectangle2_xs[1959]), .RECT2_Y(rectangle2_ys[1959]), .RECT2_WIDTH(rectangle2_widths[1959]), .RECT2_HEIGHT(rectangle2_heights[1959]), .RECT2_WEIGHT(rectangle2_weights[1959]), .RECT3_X(rectangle3_xs[1959]), .RECT3_Y(rectangle3_ys[1959]), .RECT3_WIDTH(rectangle3_widths[1959]), .RECT3_HEIGHT(rectangle3_heights[1959]), .RECT3_WEIGHT(rectangle3_weights[1959]), .FEAT_THRES(feature_thresholds[1959]), .FEAT_ABOVE(feature_aboves[1959]), .FEAT_BELOW(feature_belows[1959])) ac1959(.scan_win(scan_win1959), .scan_win_std_dev(scan_win_std_dev[1959]), .feature_accum(feature_accums[1959]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1960]), .RECT1_Y(rectangle1_ys[1960]), .RECT1_WIDTH(rectangle1_widths[1960]), .RECT1_HEIGHT(rectangle1_heights[1960]), .RECT1_WEIGHT(rectangle1_weights[1960]), .RECT2_X(rectangle2_xs[1960]), .RECT2_Y(rectangle2_ys[1960]), .RECT2_WIDTH(rectangle2_widths[1960]), .RECT2_HEIGHT(rectangle2_heights[1960]), .RECT2_WEIGHT(rectangle2_weights[1960]), .RECT3_X(rectangle3_xs[1960]), .RECT3_Y(rectangle3_ys[1960]), .RECT3_WIDTH(rectangle3_widths[1960]), .RECT3_HEIGHT(rectangle3_heights[1960]), .RECT3_WEIGHT(rectangle3_weights[1960]), .FEAT_THRES(feature_thresholds[1960]), .FEAT_ABOVE(feature_aboves[1960]), .FEAT_BELOW(feature_belows[1960])) ac1960(.scan_win(scan_win1960), .scan_win_std_dev(scan_win_std_dev[1960]), .feature_accum(feature_accums[1960]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1961]), .RECT1_Y(rectangle1_ys[1961]), .RECT1_WIDTH(rectangle1_widths[1961]), .RECT1_HEIGHT(rectangle1_heights[1961]), .RECT1_WEIGHT(rectangle1_weights[1961]), .RECT2_X(rectangle2_xs[1961]), .RECT2_Y(rectangle2_ys[1961]), .RECT2_WIDTH(rectangle2_widths[1961]), .RECT2_HEIGHT(rectangle2_heights[1961]), .RECT2_WEIGHT(rectangle2_weights[1961]), .RECT3_X(rectangle3_xs[1961]), .RECT3_Y(rectangle3_ys[1961]), .RECT3_WIDTH(rectangle3_widths[1961]), .RECT3_HEIGHT(rectangle3_heights[1961]), .RECT3_WEIGHT(rectangle3_weights[1961]), .FEAT_THRES(feature_thresholds[1961]), .FEAT_ABOVE(feature_aboves[1961]), .FEAT_BELOW(feature_belows[1961])) ac1961(.scan_win(scan_win1961), .scan_win_std_dev(scan_win_std_dev[1961]), .feature_accum(feature_accums[1961]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1962]), .RECT1_Y(rectangle1_ys[1962]), .RECT1_WIDTH(rectangle1_widths[1962]), .RECT1_HEIGHT(rectangle1_heights[1962]), .RECT1_WEIGHT(rectangle1_weights[1962]), .RECT2_X(rectangle2_xs[1962]), .RECT2_Y(rectangle2_ys[1962]), .RECT2_WIDTH(rectangle2_widths[1962]), .RECT2_HEIGHT(rectangle2_heights[1962]), .RECT2_WEIGHT(rectangle2_weights[1962]), .RECT3_X(rectangle3_xs[1962]), .RECT3_Y(rectangle3_ys[1962]), .RECT3_WIDTH(rectangle3_widths[1962]), .RECT3_HEIGHT(rectangle3_heights[1962]), .RECT3_WEIGHT(rectangle3_weights[1962]), .FEAT_THRES(feature_thresholds[1962]), .FEAT_ABOVE(feature_aboves[1962]), .FEAT_BELOW(feature_belows[1962])) ac1962(.scan_win(scan_win1962), .scan_win_std_dev(scan_win_std_dev[1962]), .feature_accum(feature_accums[1962]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1963]), .RECT1_Y(rectangle1_ys[1963]), .RECT1_WIDTH(rectangle1_widths[1963]), .RECT1_HEIGHT(rectangle1_heights[1963]), .RECT1_WEIGHT(rectangle1_weights[1963]), .RECT2_X(rectangle2_xs[1963]), .RECT2_Y(rectangle2_ys[1963]), .RECT2_WIDTH(rectangle2_widths[1963]), .RECT2_HEIGHT(rectangle2_heights[1963]), .RECT2_WEIGHT(rectangle2_weights[1963]), .RECT3_X(rectangle3_xs[1963]), .RECT3_Y(rectangle3_ys[1963]), .RECT3_WIDTH(rectangle3_widths[1963]), .RECT3_HEIGHT(rectangle3_heights[1963]), .RECT3_WEIGHT(rectangle3_weights[1963]), .FEAT_THRES(feature_thresholds[1963]), .FEAT_ABOVE(feature_aboves[1963]), .FEAT_BELOW(feature_belows[1963])) ac1963(.scan_win(scan_win1963), .scan_win_std_dev(scan_win_std_dev[1963]), .feature_accum(feature_accums[1963]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1964]), .RECT1_Y(rectangle1_ys[1964]), .RECT1_WIDTH(rectangle1_widths[1964]), .RECT1_HEIGHT(rectangle1_heights[1964]), .RECT1_WEIGHT(rectangle1_weights[1964]), .RECT2_X(rectangle2_xs[1964]), .RECT2_Y(rectangle2_ys[1964]), .RECT2_WIDTH(rectangle2_widths[1964]), .RECT2_HEIGHT(rectangle2_heights[1964]), .RECT2_WEIGHT(rectangle2_weights[1964]), .RECT3_X(rectangle3_xs[1964]), .RECT3_Y(rectangle3_ys[1964]), .RECT3_WIDTH(rectangle3_widths[1964]), .RECT3_HEIGHT(rectangle3_heights[1964]), .RECT3_WEIGHT(rectangle3_weights[1964]), .FEAT_THRES(feature_thresholds[1964]), .FEAT_ABOVE(feature_aboves[1964]), .FEAT_BELOW(feature_belows[1964])) ac1964(.scan_win(scan_win1964), .scan_win_std_dev(scan_win_std_dev[1964]), .feature_accum(feature_accums[1964]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1965]), .RECT1_Y(rectangle1_ys[1965]), .RECT1_WIDTH(rectangle1_widths[1965]), .RECT1_HEIGHT(rectangle1_heights[1965]), .RECT1_WEIGHT(rectangle1_weights[1965]), .RECT2_X(rectangle2_xs[1965]), .RECT2_Y(rectangle2_ys[1965]), .RECT2_WIDTH(rectangle2_widths[1965]), .RECT2_HEIGHT(rectangle2_heights[1965]), .RECT2_WEIGHT(rectangle2_weights[1965]), .RECT3_X(rectangle3_xs[1965]), .RECT3_Y(rectangle3_ys[1965]), .RECT3_WIDTH(rectangle3_widths[1965]), .RECT3_HEIGHT(rectangle3_heights[1965]), .RECT3_WEIGHT(rectangle3_weights[1965]), .FEAT_THRES(feature_thresholds[1965]), .FEAT_ABOVE(feature_aboves[1965]), .FEAT_BELOW(feature_belows[1965])) ac1965(.scan_win(scan_win1965), .scan_win_std_dev(scan_win_std_dev[1965]), .feature_accum(feature_accums[1965]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1966]), .RECT1_Y(rectangle1_ys[1966]), .RECT1_WIDTH(rectangle1_widths[1966]), .RECT1_HEIGHT(rectangle1_heights[1966]), .RECT1_WEIGHT(rectangle1_weights[1966]), .RECT2_X(rectangle2_xs[1966]), .RECT2_Y(rectangle2_ys[1966]), .RECT2_WIDTH(rectangle2_widths[1966]), .RECT2_HEIGHT(rectangle2_heights[1966]), .RECT2_WEIGHT(rectangle2_weights[1966]), .RECT3_X(rectangle3_xs[1966]), .RECT3_Y(rectangle3_ys[1966]), .RECT3_WIDTH(rectangle3_widths[1966]), .RECT3_HEIGHT(rectangle3_heights[1966]), .RECT3_WEIGHT(rectangle3_weights[1966]), .FEAT_THRES(feature_thresholds[1966]), .FEAT_ABOVE(feature_aboves[1966]), .FEAT_BELOW(feature_belows[1966])) ac1966(.scan_win(scan_win1966), .scan_win_std_dev(scan_win_std_dev[1966]), .feature_accum(feature_accums[1966]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1967]), .RECT1_Y(rectangle1_ys[1967]), .RECT1_WIDTH(rectangle1_widths[1967]), .RECT1_HEIGHT(rectangle1_heights[1967]), .RECT1_WEIGHT(rectangle1_weights[1967]), .RECT2_X(rectangle2_xs[1967]), .RECT2_Y(rectangle2_ys[1967]), .RECT2_WIDTH(rectangle2_widths[1967]), .RECT2_HEIGHT(rectangle2_heights[1967]), .RECT2_WEIGHT(rectangle2_weights[1967]), .RECT3_X(rectangle3_xs[1967]), .RECT3_Y(rectangle3_ys[1967]), .RECT3_WIDTH(rectangle3_widths[1967]), .RECT3_HEIGHT(rectangle3_heights[1967]), .RECT3_WEIGHT(rectangle3_weights[1967]), .FEAT_THRES(feature_thresholds[1967]), .FEAT_ABOVE(feature_aboves[1967]), .FEAT_BELOW(feature_belows[1967])) ac1967(.scan_win(scan_win1967), .scan_win_std_dev(scan_win_std_dev[1967]), .feature_accum(feature_accums[1967]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1968]), .RECT1_Y(rectangle1_ys[1968]), .RECT1_WIDTH(rectangle1_widths[1968]), .RECT1_HEIGHT(rectangle1_heights[1968]), .RECT1_WEIGHT(rectangle1_weights[1968]), .RECT2_X(rectangle2_xs[1968]), .RECT2_Y(rectangle2_ys[1968]), .RECT2_WIDTH(rectangle2_widths[1968]), .RECT2_HEIGHT(rectangle2_heights[1968]), .RECT2_WEIGHT(rectangle2_weights[1968]), .RECT3_X(rectangle3_xs[1968]), .RECT3_Y(rectangle3_ys[1968]), .RECT3_WIDTH(rectangle3_widths[1968]), .RECT3_HEIGHT(rectangle3_heights[1968]), .RECT3_WEIGHT(rectangle3_weights[1968]), .FEAT_THRES(feature_thresholds[1968]), .FEAT_ABOVE(feature_aboves[1968]), .FEAT_BELOW(feature_belows[1968])) ac1968(.scan_win(scan_win1968), .scan_win_std_dev(scan_win_std_dev[1968]), .feature_accum(feature_accums[1968]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1969]), .RECT1_Y(rectangle1_ys[1969]), .RECT1_WIDTH(rectangle1_widths[1969]), .RECT1_HEIGHT(rectangle1_heights[1969]), .RECT1_WEIGHT(rectangle1_weights[1969]), .RECT2_X(rectangle2_xs[1969]), .RECT2_Y(rectangle2_ys[1969]), .RECT2_WIDTH(rectangle2_widths[1969]), .RECT2_HEIGHT(rectangle2_heights[1969]), .RECT2_WEIGHT(rectangle2_weights[1969]), .RECT3_X(rectangle3_xs[1969]), .RECT3_Y(rectangle3_ys[1969]), .RECT3_WIDTH(rectangle3_widths[1969]), .RECT3_HEIGHT(rectangle3_heights[1969]), .RECT3_WEIGHT(rectangle3_weights[1969]), .FEAT_THRES(feature_thresholds[1969]), .FEAT_ABOVE(feature_aboves[1969]), .FEAT_BELOW(feature_belows[1969])) ac1969(.scan_win(scan_win1969), .scan_win_std_dev(scan_win_std_dev[1969]), .feature_accum(feature_accums[1969]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1970]), .RECT1_Y(rectangle1_ys[1970]), .RECT1_WIDTH(rectangle1_widths[1970]), .RECT1_HEIGHT(rectangle1_heights[1970]), .RECT1_WEIGHT(rectangle1_weights[1970]), .RECT2_X(rectangle2_xs[1970]), .RECT2_Y(rectangle2_ys[1970]), .RECT2_WIDTH(rectangle2_widths[1970]), .RECT2_HEIGHT(rectangle2_heights[1970]), .RECT2_WEIGHT(rectangle2_weights[1970]), .RECT3_X(rectangle3_xs[1970]), .RECT3_Y(rectangle3_ys[1970]), .RECT3_WIDTH(rectangle3_widths[1970]), .RECT3_HEIGHT(rectangle3_heights[1970]), .RECT3_WEIGHT(rectangle3_weights[1970]), .FEAT_THRES(feature_thresholds[1970]), .FEAT_ABOVE(feature_aboves[1970]), .FEAT_BELOW(feature_belows[1970])) ac1970(.scan_win(scan_win1970), .scan_win_std_dev(scan_win_std_dev[1970]), .feature_accum(feature_accums[1970]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1971]), .RECT1_Y(rectangle1_ys[1971]), .RECT1_WIDTH(rectangle1_widths[1971]), .RECT1_HEIGHT(rectangle1_heights[1971]), .RECT1_WEIGHT(rectangle1_weights[1971]), .RECT2_X(rectangle2_xs[1971]), .RECT2_Y(rectangle2_ys[1971]), .RECT2_WIDTH(rectangle2_widths[1971]), .RECT2_HEIGHT(rectangle2_heights[1971]), .RECT2_WEIGHT(rectangle2_weights[1971]), .RECT3_X(rectangle3_xs[1971]), .RECT3_Y(rectangle3_ys[1971]), .RECT3_WIDTH(rectangle3_widths[1971]), .RECT3_HEIGHT(rectangle3_heights[1971]), .RECT3_WEIGHT(rectangle3_weights[1971]), .FEAT_THRES(feature_thresholds[1971]), .FEAT_ABOVE(feature_aboves[1971]), .FEAT_BELOW(feature_belows[1971])) ac1971(.scan_win(scan_win1971), .scan_win_std_dev(scan_win_std_dev[1971]), .feature_accum(feature_accums[1971]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1972]), .RECT1_Y(rectangle1_ys[1972]), .RECT1_WIDTH(rectangle1_widths[1972]), .RECT1_HEIGHT(rectangle1_heights[1972]), .RECT1_WEIGHT(rectangle1_weights[1972]), .RECT2_X(rectangle2_xs[1972]), .RECT2_Y(rectangle2_ys[1972]), .RECT2_WIDTH(rectangle2_widths[1972]), .RECT2_HEIGHT(rectangle2_heights[1972]), .RECT2_WEIGHT(rectangle2_weights[1972]), .RECT3_X(rectangle3_xs[1972]), .RECT3_Y(rectangle3_ys[1972]), .RECT3_WIDTH(rectangle3_widths[1972]), .RECT3_HEIGHT(rectangle3_heights[1972]), .RECT3_WEIGHT(rectangle3_weights[1972]), .FEAT_THRES(feature_thresholds[1972]), .FEAT_ABOVE(feature_aboves[1972]), .FEAT_BELOW(feature_belows[1972])) ac1972(.scan_win(scan_win1972), .scan_win_std_dev(scan_win_std_dev[1972]), .feature_accum(feature_accums[1972]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1973]), .RECT1_Y(rectangle1_ys[1973]), .RECT1_WIDTH(rectangle1_widths[1973]), .RECT1_HEIGHT(rectangle1_heights[1973]), .RECT1_WEIGHT(rectangle1_weights[1973]), .RECT2_X(rectangle2_xs[1973]), .RECT2_Y(rectangle2_ys[1973]), .RECT2_WIDTH(rectangle2_widths[1973]), .RECT2_HEIGHT(rectangle2_heights[1973]), .RECT2_WEIGHT(rectangle2_weights[1973]), .RECT3_X(rectangle3_xs[1973]), .RECT3_Y(rectangle3_ys[1973]), .RECT3_WIDTH(rectangle3_widths[1973]), .RECT3_HEIGHT(rectangle3_heights[1973]), .RECT3_WEIGHT(rectangle3_weights[1973]), .FEAT_THRES(feature_thresholds[1973]), .FEAT_ABOVE(feature_aboves[1973]), .FEAT_BELOW(feature_belows[1973])) ac1973(.scan_win(scan_win1973), .scan_win_std_dev(scan_win_std_dev[1973]), .feature_accum(feature_accums[1973]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1974]), .RECT1_Y(rectangle1_ys[1974]), .RECT1_WIDTH(rectangle1_widths[1974]), .RECT1_HEIGHT(rectangle1_heights[1974]), .RECT1_WEIGHT(rectangle1_weights[1974]), .RECT2_X(rectangle2_xs[1974]), .RECT2_Y(rectangle2_ys[1974]), .RECT2_WIDTH(rectangle2_widths[1974]), .RECT2_HEIGHT(rectangle2_heights[1974]), .RECT2_WEIGHT(rectangle2_weights[1974]), .RECT3_X(rectangle3_xs[1974]), .RECT3_Y(rectangle3_ys[1974]), .RECT3_WIDTH(rectangle3_widths[1974]), .RECT3_HEIGHT(rectangle3_heights[1974]), .RECT3_WEIGHT(rectangle3_weights[1974]), .FEAT_THRES(feature_thresholds[1974]), .FEAT_ABOVE(feature_aboves[1974]), .FEAT_BELOW(feature_belows[1974])) ac1974(.scan_win(scan_win1974), .scan_win_std_dev(scan_win_std_dev[1974]), .feature_accum(feature_accums[1974]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1975]), .RECT1_Y(rectangle1_ys[1975]), .RECT1_WIDTH(rectangle1_widths[1975]), .RECT1_HEIGHT(rectangle1_heights[1975]), .RECT1_WEIGHT(rectangle1_weights[1975]), .RECT2_X(rectangle2_xs[1975]), .RECT2_Y(rectangle2_ys[1975]), .RECT2_WIDTH(rectangle2_widths[1975]), .RECT2_HEIGHT(rectangle2_heights[1975]), .RECT2_WEIGHT(rectangle2_weights[1975]), .RECT3_X(rectangle3_xs[1975]), .RECT3_Y(rectangle3_ys[1975]), .RECT3_WIDTH(rectangle3_widths[1975]), .RECT3_HEIGHT(rectangle3_heights[1975]), .RECT3_WEIGHT(rectangle3_weights[1975]), .FEAT_THRES(feature_thresholds[1975]), .FEAT_ABOVE(feature_aboves[1975]), .FEAT_BELOW(feature_belows[1975])) ac1975(.scan_win(scan_win1975), .scan_win_std_dev(scan_win_std_dev[1975]), .feature_accum(feature_accums[1975]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1976]), .RECT1_Y(rectangle1_ys[1976]), .RECT1_WIDTH(rectangle1_widths[1976]), .RECT1_HEIGHT(rectangle1_heights[1976]), .RECT1_WEIGHT(rectangle1_weights[1976]), .RECT2_X(rectangle2_xs[1976]), .RECT2_Y(rectangle2_ys[1976]), .RECT2_WIDTH(rectangle2_widths[1976]), .RECT2_HEIGHT(rectangle2_heights[1976]), .RECT2_WEIGHT(rectangle2_weights[1976]), .RECT3_X(rectangle3_xs[1976]), .RECT3_Y(rectangle3_ys[1976]), .RECT3_WIDTH(rectangle3_widths[1976]), .RECT3_HEIGHT(rectangle3_heights[1976]), .RECT3_WEIGHT(rectangle3_weights[1976]), .FEAT_THRES(feature_thresholds[1976]), .FEAT_ABOVE(feature_aboves[1976]), .FEAT_BELOW(feature_belows[1976])) ac1976(.scan_win(scan_win1976), .scan_win_std_dev(scan_win_std_dev[1976]), .feature_accum(feature_accums[1976]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1977]), .RECT1_Y(rectangle1_ys[1977]), .RECT1_WIDTH(rectangle1_widths[1977]), .RECT1_HEIGHT(rectangle1_heights[1977]), .RECT1_WEIGHT(rectangle1_weights[1977]), .RECT2_X(rectangle2_xs[1977]), .RECT2_Y(rectangle2_ys[1977]), .RECT2_WIDTH(rectangle2_widths[1977]), .RECT2_HEIGHT(rectangle2_heights[1977]), .RECT2_WEIGHT(rectangle2_weights[1977]), .RECT3_X(rectangle3_xs[1977]), .RECT3_Y(rectangle3_ys[1977]), .RECT3_WIDTH(rectangle3_widths[1977]), .RECT3_HEIGHT(rectangle3_heights[1977]), .RECT3_WEIGHT(rectangle3_weights[1977]), .FEAT_THRES(feature_thresholds[1977]), .FEAT_ABOVE(feature_aboves[1977]), .FEAT_BELOW(feature_belows[1977])) ac1977(.scan_win(scan_win1977), .scan_win_std_dev(scan_win_std_dev[1977]), .feature_accum(feature_accums[1977]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1978]), .RECT1_Y(rectangle1_ys[1978]), .RECT1_WIDTH(rectangle1_widths[1978]), .RECT1_HEIGHT(rectangle1_heights[1978]), .RECT1_WEIGHT(rectangle1_weights[1978]), .RECT2_X(rectangle2_xs[1978]), .RECT2_Y(rectangle2_ys[1978]), .RECT2_WIDTH(rectangle2_widths[1978]), .RECT2_HEIGHT(rectangle2_heights[1978]), .RECT2_WEIGHT(rectangle2_weights[1978]), .RECT3_X(rectangle3_xs[1978]), .RECT3_Y(rectangle3_ys[1978]), .RECT3_WIDTH(rectangle3_widths[1978]), .RECT3_HEIGHT(rectangle3_heights[1978]), .RECT3_WEIGHT(rectangle3_weights[1978]), .FEAT_THRES(feature_thresholds[1978]), .FEAT_ABOVE(feature_aboves[1978]), .FEAT_BELOW(feature_belows[1978])) ac1978(.scan_win(scan_win1978), .scan_win_std_dev(scan_win_std_dev[1978]), .feature_accum(feature_accums[1978]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1979]), .RECT1_Y(rectangle1_ys[1979]), .RECT1_WIDTH(rectangle1_widths[1979]), .RECT1_HEIGHT(rectangle1_heights[1979]), .RECT1_WEIGHT(rectangle1_weights[1979]), .RECT2_X(rectangle2_xs[1979]), .RECT2_Y(rectangle2_ys[1979]), .RECT2_WIDTH(rectangle2_widths[1979]), .RECT2_HEIGHT(rectangle2_heights[1979]), .RECT2_WEIGHT(rectangle2_weights[1979]), .RECT3_X(rectangle3_xs[1979]), .RECT3_Y(rectangle3_ys[1979]), .RECT3_WIDTH(rectangle3_widths[1979]), .RECT3_HEIGHT(rectangle3_heights[1979]), .RECT3_WEIGHT(rectangle3_weights[1979]), .FEAT_THRES(feature_thresholds[1979]), .FEAT_ABOVE(feature_aboves[1979]), .FEAT_BELOW(feature_belows[1979])) ac1979(.scan_win(scan_win1979), .scan_win_std_dev(scan_win_std_dev[1979]), .feature_accum(feature_accums[1979]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1980]), .RECT1_Y(rectangle1_ys[1980]), .RECT1_WIDTH(rectangle1_widths[1980]), .RECT1_HEIGHT(rectangle1_heights[1980]), .RECT1_WEIGHT(rectangle1_weights[1980]), .RECT2_X(rectangle2_xs[1980]), .RECT2_Y(rectangle2_ys[1980]), .RECT2_WIDTH(rectangle2_widths[1980]), .RECT2_HEIGHT(rectangle2_heights[1980]), .RECT2_WEIGHT(rectangle2_weights[1980]), .RECT3_X(rectangle3_xs[1980]), .RECT3_Y(rectangle3_ys[1980]), .RECT3_WIDTH(rectangle3_widths[1980]), .RECT3_HEIGHT(rectangle3_heights[1980]), .RECT3_WEIGHT(rectangle3_weights[1980]), .FEAT_THRES(feature_thresholds[1980]), .FEAT_ABOVE(feature_aboves[1980]), .FEAT_BELOW(feature_belows[1980])) ac1980(.scan_win(scan_win1980), .scan_win_std_dev(scan_win_std_dev[1980]), .feature_accum(feature_accums[1980]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1981]), .RECT1_Y(rectangle1_ys[1981]), .RECT1_WIDTH(rectangle1_widths[1981]), .RECT1_HEIGHT(rectangle1_heights[1981]), .RECT1_WEIGHT(rectangle1_weights[1981]), .RECT2_X(rectangle2_xs[1981]), .RECT2_Y(rectangle2_ys[1981]), .RECT2_WIDTH(rectangle2_widths[1981]), .RECT2_HEIGHT(rectangle2_heights[1981]), .RECT2_WEIGHT(rectangle2_weights[1981]), .RECT3_X(rectangle3_xs[1981]), .RECT3_Y(rectangle3_ys[1981]), .RECT3_WIDTH(rectangle3_widths[1981]), .RECT3_HEIGHT(rectangle3_heights[1981]), .RECT3_WEIGHT(rectangle3_weights[1981]), .FEAT_THRES(feature_thresholds[1981]), .FEAT_ABOVE(feature_aboves[1981]), .FEAT_BELOW(feature_belows[1981])) ac1981(.scan_win(scan_win1981), .scan_win_std_dev(scan_win_std_dev[1981]), .feature_accum(feature_accums[1981]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1982]), .RECT1_Y(rectangle1_ys[1982]), .RECT1_WIDTH(rectangle1_widths[1982]), .RECT1_HEIGHT(rectangle1_heights[1982]), .RECT1_WEIGHT(rectangle1_weights[1982]), .RECT2_X(rectangle2_xs[1982]), .RECT2_Y(rectangle2_ys[1982]), .RECT2_WIDTH(rectangle2_widths[1982]), .RECT2_HEIGHT(rectangle2_heights[1982]), .RECT2_WEIGHT(rectangle2_weights[1982]), .RECT3_X(rectangle3_xs[1982]), .RECT3_Y(rectangle3_ys[1982]), .RECT3_WIDTH(rectangle3_widths[1982]), .RECT3_HEIGHT(rectangle3_heights[1982]), .RECT3_WEIGHT(rectangle3_weights[1982]), .FEAT_THRES(feature_thresholds[1982]), .FEAT_ABOVE(feature_aboves[1982]), .FEAT_BELOW(feature_belows[1982])) ac1982(.scan_win(scan_win1982), .scan_win_std_dev(scan_win_std_dev[1982]), .feature_accum(feature_accums[1982]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1983]), .RECT1_Y(rectangle1_ys[1983]), .RECT1_WIDTH(rectangle1_widths[1983]), .RECT1_HEIGHT(rectangle1_heights[1983]), .RECT1_WEIGHT(rectangle1_weights[1983]), .RECT2_X(rectangle2_xs[1983]), .RECT2_Y(rectangle2_ys[1983]), .RECT2_WIDTH(rectangle2_widths[1983]), .RECT2_HEIGHT(rectangle2_heights[1983]), .RECT2_WEIGHT(rectangle2_weights[1983]), .RECT3_X(rectangle3_xs[1983]), .RECT3_Y(rectangle3_ys[1983]), .RECT3_WIDTH(rectangle3_widths[1983]), .RECT3_HEIGHT(rectangle3_heights[1983]), .RECT3_WEIGHT(rectangle3_weights[1983]), .FEAT_THRES(feature_thresholds[1983]), .FEAT_ABOVE(feature_aboves[1983]), .FEAT_BELOW(feature_belows[1983])) ac1983(.scan_win(scan_win1983), .scan_win_std_dev(scan_win_std_dev[1983]), .feature_accum(feature_accums[1983]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1984]), .RECT1_Y(rectangle1_ys[1984]), .RECT1_WIDTH(rectangle1_widths[1984]), .RECT1_HEIGHT(rectangle1_heights[1984]), .RECT1_WEIGHT(rectangle1_weights[1984]), .RECT2_X(rectangle2_xs[1984]), .RECT2_Y(rectangle2_ys[1984]), .RECT2_WIDTH(rectangle2_widths[1984]), .RECT2_HEIGHT(rectangle2_heights[1984]), .RECT2_WEIGHT(rectangle2_weights[1984]), .RECT3_X(rectangle3_xs[1984]), .RECT3_Y(rectangle3_ys[1984]), .RECT3_WIDTH(rectangle3_widths[1984]), .RECT3_HEIGHT(rectangle3_heights[1984]), .RECT3_WEIGHT(rectangle3_weights[1984]), .FEAT_THRES(feature_thresholds[1984]), .FEAT_ABOVE(feature_aboves[1984]), .FEAT_BELOW(feature_belows[1984])) ac1984(.scan_win(scan_win1984), .scan_win_std_dev(scan_win_std_dev[1984]), .feature_accum(feature_accums[1984]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1985]), .RECT1_Y(rectangle1_ys[1985]), .RECT1_WIDTH(rectangle1_widths[1985]), .RECT1_HEIGHT(rectangle1_heights[1985]), .RECT1_WEIGHT(rectangle1_weights[1985]), .RECT2_X(rectangle2_xs[1985]), .RECT2_Y(rectangle2_ys[1985]), .RECT2_WIDTH(rectangle2_widths[1985]), .RECT2_HEIGHT(rectangle2_heights[1985]), .RECT2_WEIGHT(rectangle2_weights[1985]), .RECT3_X(rectangle3_xs[1985]), .RECT3_Y(rectangle3_ys[1985]), .RECT3_WIDTH(rectangle3_widths[1985]), .RECT3_HEIGHT(rectangle3_heights[1985]), .RECT3_WEIGHT(rectangle3_weights[1985]), .FEAT_THRES(feature_thresholds[1985]), .FEAT_ABOVE(feature_aboves[1985]), .FEAT_BELOW(feature_belows[1985])) ac1985(.scan_win(scan_win1985), .scan_win_std_dev(scan_win_std_dev[1985]), .feature_accum(feature_accums[1985]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1986]), .RECT1_Y(rectangle1_ys[1986]), .RECT1_WIDTH(rectangle1_widths[1986]), .RECT1_HEIGHT(rectangle1_heights[1986]), .RECT1_WEIGHT(rectangle1_weights[1986]), .RECT2_X(rectangle2_xs[1986]), .RECT2_Y(rectangle2_ys[1986]), .RECT2_WIDTH(rectangle2_widths[1986]), .RECT2_HEIGHT(rectangle2_heights[1986]), .RECT2_WEIGHT(rectangle2_weights[1986]), .RECT3_X(rectangle3_xs[1986]), .RECT3_Y(rectangle3_ys[1986]), .RECT3_WIDTH(rectangle3_widths[1986]), .RECT3_HEIGHT(rectangle3_heights[1986]), .RECT3_WEIGHT(rectangle3_weights[1986]), .FEAT_THRES(feature_thresholds[1986]), .FEAT_ABOVE(feature_aboves[1986]), .FEAT_BELOW(feature_belows[1986])) ac1986(.scan_win(scan_win1986), .scan_win_std_dev(scan_win_std_dev[1986]), .feature_accum(feature_accums[1986]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1987]), .RECT1_Y(rectangle1_ys[1987]), .RECT1_WIDTH(rectangle1_widths[1987]), .RECT1_HEIGHT(rectangle1_heights[1987]), .RECT1_WEIGHT(rectangle1_weights[1987]), .RECT2_X(rectangle2_xs[1987]), .RECT2_Y(rectangle2_ys[1987]), .RECT2_WIDTH(rectangle2_widths[1987]), .RECT2_HEIGHT(rectangle2_heights[1987]), .RECT2_WEIGHT(rectangle2_weights[1987]), .RECT3_X(rectangle3_xs[1987]), .RECT3_Y(rectangle3_ys[1987]), .RECT3_WIDTH(rectangle3_widths[1987]), .RECT3_HEIGHT(rectangle3_heights[1987]), .RECT3_WEIGHT(rectangle3_weights[1987]), .FEAT_THRES(feature_thresholds[1987]), .FEAT_ABOVE(feature_aboves[1987]), .FEAT_BELOW(feature_belows[1987])) ac1987(.scan_win(scan_win1987), .scan_win_std_dev(scan_win_std_dev[1987]), .feature_accum(feature_accums[1987]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1988]), .RECT1_Y(rectangle1_ys[1988]), .RECT1_WIDTH(rectangle1_widths[1988]), .RECT1_HEIGHT(rectangle1_heights[1988]), .RECT1_WEIGHT(rectangle1_weights[1988]), .RECT2_X(rectangle2_xs[1988]), .RECT2_Y(rectangle2_ys[1988]), .RECT2_WIDTH(rectangle2_widths[1988]), .RECT2_HEIGHT(rectangle2_heights[1988]), .RECT2_WEIGHT(rectangle2_weights[1988]), .RECT3_X(rectangle3_xs[1988]), .RECT3_Y(rectangle3_ys[1988]), .RECT3_WIDTH(rectangle3_widths[1988]), .RECT3_HEIGHT(rectangle3_heights[1988]), .RECT3_WEIGHT(rectangle3_weights[1988]), .FEAT_THRES(feature_thresholds[1988]), .FEAT_ABOVE(feature_aboves[1988]), .FEAT_BELOW(feature_belows[1988])) ac1988(.scan_win(scan_win1988), .scan_win_std_dev(scan_win_std_dev[1988]), .feature_accum(feature_accums[1988]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1989]), .RECT1_Y(rectangle1_ys[1989]), .RECT1_WIDTH(rectangle1_widths[1989]), .RECT1_HEIGHT(rectangle1_heights[1989]), .RECT1_WEIGHT(rectangle1_weights[1989]), .RECT2_X(rectangle2_xs[1989]), .RECT2_Y(rectangle2_ys[1989]), .RECT2_WIDTH(rectangle2_widths[1989]), .RECT2_HEIGHT(rectangle2_heights[1989]), .RECT2_WEIGHT(rectangle2_weights[1989]), .RECT3_X(rectangle3_xs[1989]), .RECT3_Y(rectangle3_ys[1989]), .RECT3_WIDTH(rectangle3_widths[1989]), .RECT3_HEIGHT(rectangle3_heights[1989]), .RECT3_WEIGHT(rectangle3_weights[1989]), .FEAT_THRES(feature_thresholds[1989]), .FEAT_ABOVE(feature_aboves[1989]), .FEAT_BELOW(feature_belows[1989])) ac1989(.scan_win(scan_win1989), .scan_win_std_dev(scan_win_std_dev[1989]), .feature_accum(feature_accums[1989]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1990]), .RECT1_Y(rectangle1_ys[1990]), .RECT1_WIDTH(rectangle1_widths[1990]), .RECT1_HEIGHT(rectangle1_heights[1990]), .RECT1_WEIGHT(rectangle1_weights[1990]), .RECT2_X(rectangle2_xs[1990]), .RECT2_Y(rectangle2_ys[1990]), .RECT2_WIDTH(rectangle2_widths[1990]), .RECT2_HEIGHT(rectangle2_heights[1990]), .RECT2_WEIGHT(rectangle2_weights[1990]), .RECT3_X(rectangle3_xs[1990]), .RECT3_Y(rectangle3_ys[1990]), .RECT3_WIDTH(rectangle3_widths[1990]), .RECT3_HEIGHT(rectangle3_heights[1990]), .RECT3_WEIGHT(rectangle3_weights[1990]), .FEAT_THRES(feature_thresholds[1990]), .FEAT_ABOVE(feature_aboves[1990]), .FEAT_BELOW(feature_belows[1990])) ac1990(.scan_win(scan_win1990), .scan_win_std_dev(scan_win_std_dev[1990]), .feature_accum(feature_accums[1990]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1991]), .RECT1_Y(rectangle1_ys[1991]), .RECT1_WIDTH(rectangle1_widths[1991]), .RECT1_HEIGHT(rectangle1_heights[1991]), .RECT1_WEIGHT(rectangle1_weights[1991]), .RECT2_X(rectangle2_xs[1991]), .RECT2_Y(rectangle2_ys[1991]), .RECT2_WIDTH(rectangle2_widths[1991]), .RECT2_HEIGHT(rectangle2_heights[1991]), .RECT2_WEIGHT(rectangle2_weights[1991]), .RECT3_X(rectangle3_xs[1991]), .RECT3_Y(rectangle3_ys[1991]), .RECT3_WIDTH(rectangle3_widths[1991]), .RECT3_HEIGHT(rectangle3_heights[1991]), .RECT3_WEIGHT(rectangle3_weights[1991]), .FEAT_THRES(feature_thresholds[1991]), .FEAT_ABOVE(feature_aboves[1991]), .FEAT_BELOW(feature_belows[1991])) ac1991(.scan_win(scan_win1991), .scan_win_std_dev(scan_win_std_dev[1991]), .feature_accum(feature_accums[1991]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1992]), .RECT1_Y(rectangle1_ys[1992]), .RECT1_WIDTH(rectangle1_widths[1992]), .RECT1_HEIGHT(rectangle1_heights[1992]), .RECT1_WEIGHT(rectangle1_weights[1992]), .RECT2_X(rectangle2_xs[1992]), .RECT2_Y(rectangle2_ys[1992]), .RECT2_WIDTH(rectangle2_widths[1992]), .RECT2_HEIGHT(rectangle2_heights[1992]), .RECT2_WEIGHT(rectangle2_weights[1992]), .RECT3_X(rectangle3_xs[1992]), .RECT3_Y(rectangle3_ys[1992]), .RECT3_WIDTH(rectangle3_widths[1992]), .RECT3_HEIGHT(rectangle3_heights[1992]), .RECT3_WEIGHT(rectangle3_weights[1992]), .FEAT_THRES(feature_thresholds[1992]), .FEAT_ABOVE(feature_aboves[1992]), .FEAT_BELOW(feature_belows[1992])) ac1992(.scan_win(scan_win1992), .scan_win_std_dev(scan_win_std_dev[1992]), .feature_accum(feature_accums[1992]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1993]), .RECT1_Y(rectangle1_ys[1993]), .RECT1_WIDTH(rectangle1_widths[1993]), .RECT1_HEIGHT(rectangle1_heights[1993]), .RECT1_WEIGHT(rectangle1_weights[1993]), .RECT2_X(rectangle2_xs[1993]), .RECT2_Y(rectangle2_ys[1993]), .RECT2_WIDTH(rectangle2_widths[1993]), .RECT2_HEIGHT(rectangle2_heights[1993]), .RECT2_WEIGHT(rectangle2_weights[1993]), .RECT3_X(rectangle3_xs[1993]), .RECT3_Y(rectangle3_ys[1993]), .RECT3_WIDTH(rectangle3_widths[1993]), .RECT3_HEIGHT(rectangle3_heights[1993]), .RECT3_WEIGHT(rectangle3_weights[1993]), .FEAT_THRES(feature_thresholds[1993]), .FEAT_ABOVE(feature_aboves[1993]), .FEAT_BELOW(feature_belows[1993])) ac1993(.scan_win(scan_win1993), .scan_win_std_dev(scan_win_std_dev[1993]), .feature_accum(feature_accums[1993]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1994]), .RECT1_Y(rectangle1_ys[1994]), .RECT1_WIDTH(rectangle1_widths[1994]), .RECT1_HEIGHT(rectangle1_heights[1994]), .RECT1_WEIGHT(rectangle1_weights[1994]), .RECT2_X(rectangle2_xs[1994]), .RECT2_Y(rectangle2_ys[1994]), .RECT2_WIDTH(rectangle2_widths[1994]), .RECT2_HEIGHT(rectangle2_heights[1994]), .RECT2_WEIGHT(rectangle2_weights[1994]), .RECT3_X(rectangle3_xs[1994]), .RECT3_Y(rectangle3_ys[1994]), .RECT3_WIDTH(rectangle3_widths[1994]), .RECT3_HEIGHT(rectangle3_heights[1994]), .RECT3_WEIGHT(rectangle3_weights[1994]), .FEAT_THRES(feature_thresholds[1994]), .FEAT_ABOVE(feature_aboves[1994]), .FEAT_BELOW(feature_belows[1994])) ac1994(.scan_win(scan_win1994), .scan_win_std_dev(scan_win_std_dev[1994]), .feature_accum(feature_accums[1994]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1995]), .RECT1_Y(rectangle1_ys[1995]), .RECT1_WIDTH(rectangle1_widths[1995]), .RECT1_HEIGHT(rectangle1_heights[1995]), .RECT1_WEIGHT(rectangle1_weights[1995]), .RECT2_X(rectangle2_xs[1995]), .RECT2_Y(rectangle2_ys[1995]), .RECT2_WIDTH(rectangle2_widths[1995]), .RECT2_HEIGHT(rectangle2_heights[1995]), .RECT2_WEIGHT(rectangle2_weights[1995]), .RECT3_X(rectangle3_xs[1995]), .RECT3_Y(rectangle3_ys[1995]), .RECT3_WIDTH(rectangle3_widths[1995]), .RECT3_HEIGHT(rectangle3_heights[1995]), .RECT3_WEIGHT(rectangle3_weights[1995]), .FEAT_THRES(feature_thresholds[1995]), .FEAT_ABOVE(feature_aboves[1995]), .FEAT_BELOW(feature_belows[1995])) ac1995(.scan_win(scan_win1995), .scan_win_std_dev(scan_win_std_dev[1995]), .feature_accum(feature_accums[1995]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1996]), .RECT1_Y(rectangle1_ys[1996]), .RECT1_WIDTH(rectangle1_widths[1996]), .RECT1_HEIGHT(rectangle1_heights[1996]), .RECT1_WEIGHT(rectangle1_weights[1996]), .RECT2_X(rectangle2_xs[1996]), .RECT2_Y(rectangle2_ys[1996]), .RECT2_WIDTH(rectangle2_widths[1996]), .RECT2_HEIGHT(rectangle2_heights[1996]), .RECT2_WEIGHT(rectangle2_weights[1996]), .RECT3_X(rectangle3_xs[1996]), .RECT3_Y(rectangle3_ys[1996]), .RECT3_WIDTH(rectangle3_widths[1996]), .RECT3_HEIGHT(rectangle3_heights[1996]), .RECT3_WEIGHT(rectangle3_weights[1996]), .FEAT_THRES(feature_thresholds[1996]), .FEAT_ABOVE(feature_aboves[1996]), .FEAT_BELOW(feature_belows[1996])) ac1996(.scan_win(scan_win1996), .scan_win_std_dev(scan_win_std_dev[1996]), .feature_accum(feature_accums[1996]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1997]), .RECT1_Y(rectangle1_ys[1997]), .RECT1_WIDTH(rectangle1_widths[1997]), .RECT1_HEIGHT(rectangle1_heights[1997]), .RECT1_WEIGHT(rectangle1_weights[1997]), .RECT2_X(rectangle2_xs[1997]), .RECT2_Y(rectangle2_ys[1997]), .RECT2_WIDTH(rectangle2_widths[1997]), .RECT2_HEIGHT(rectangle2_heights[1997]), .RECT2_WEIGHT(rectangle2_weights[1997]), .RECT3_X(rectangle3_xs[1997]), .RECT3_Y(rectangle3_ys[1997]), .RECT3_WIDTH(rectangle3_widths[1997]), .RECT3_HEIGHT(rectangle3_heights[1997]), .RECT3_WEIGHT(rectangle3_weights[1997]), .FEAT_THRES(feature_thresholds[1997]), .FEAT_ABOVE(feature_aboves[1997]), .FEAT_BELOW(feature_belows[1997])) ac1997(.scan_win(scan_win1997), .scan_win_std_dev(scan_win_std_dev[1997]), .feature_accum(feature_accums[1997]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1998]), .RECT1_Y(rectangle1_ys[1998]), .RECT1_WIDTH(rectangle1_widths[1998]), .RECT1_HEIGHT(rectangle1_heights[1998]), .RECT1_WEIGHT(rectangle1_weights[1998]), .RECT2_X(rectangle2_xs[1998]), .RECT2_Y(rectangle2_ys[1998]), .RECT2_WIDTH(rectangle2_widths[1998]), .RECT2_HEIGHT(rectangle2_heights[1998]), .RECT2_WEIGHT(rectangle2_weights[1998]), .RECT3_X(rectangle3_xs[1998]), .RECT3_Y(rectangle3_ys[1998]), .RECT3_WIDTH(rectangle3_widths[1998]), .RECT3_HEIGHT(rectangle3_heights[1998]), .RECT3_WEIGHT(rectangle3_weights[1998]), .FEAT_THRES(feature_thresholds[1998]), .FEAT_ABOVE(feature_aboves[1998]), .FEAT_BELOW(feature_belows[1998])) ac1998(.scan_win(scan_win1998), .scan_win_std_dev(scan_win_std_dev[1998]), .feature_accum(feature_accums[1998]));
  accum_calculator #(.RECT1_X(rectangle1_xs[1999]), .RECT1_Y(rectangle1_ys[1999]), .RECT1_WIDTH(rectangle1_widths[1999]), .RECT1_HEIGHT(rectangle1_heights[1999]), .RECT1_WEIGHT(rectangle1_weights[1999]), .RECT2_X(rectangle2_xs[1999]), .RECT2_Y(rectangle2_ys[1999]), .RECT2_WIDTH(rectangle2_widths[1999]), .RECT2_HEIGHT(rectangle2_heights[1999]), .RECT2_WEIGHT(rectangle2_weights[1999]), .RECT3_X(rectangle3_xs[1999]), .RECT3_Y(rectangle3_ys[1999]), .RECT3_WIDTH(rectangle3_widths[1999]), .RECT3_HEIGHT(rectangle3_heights[1999]), .RECT3_WEIGHT(rectangle3_weights[1999]), .FEAT_THRES(feature_thresholds[1999]), .FEAT_ABOVE(feature_aboves[1999]), .FEAT_BELOW(feature_belows[1999])) ac1999(.scan_win(scan_win1999), .scan_win_std_dev(scan_win_std_dev[1999]), .feature_accum(feature_accums[1999]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2000]), .RECT1_Y(rectangle1_ys[2000]), .RECT1_WIDTH(rectangle1_widths[2000]), .RECT1_HEIGHT(rectangle1_heights[2000]), .RECT1_WEIGHT(rectangle1_weights[2000]), .RECT2_X(rectangle2_xs[2000]), .RECT2_Y(rectangle2_ys[2000]), .RECT2_WIDTH(rectangle2_widths[2000]), .RECT2_HEIGHT(rectangle2_heights[2000]), .RECT2_WEIGHT(rectangle2_weights[2000]), .RECT3_X(rectangle3_xs[2000]), .RECT3_Y(rectangle3_ys[2000]), .RECT3_WIDTH(rectangle3_widths[2000]), .RECT3_HEIGHT(rectangle3_heights[2000]), .RECT3_WEIGHT(rectangle3_weights[2000]), .FEAT_THRES(feature_thresholds[2000]), .FEAT_ABOVE(feature_aboves[2000]), .FEAT_BELOW(feature_belows[2000])) ac2000(.scan_win(scan_win2000), .scan_win_std_dev(scan_win_std_dev[2000]), .feature_accum(feature_accums[2000]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2001]), .RECT1_Y(rectangle1_ys[2001]), .RECT1_WIDTH(rectangle1_widths[2001]), .RECT1_HEIGHT(rectangle1_heights[2001]), .RECT1_WEIGHT(rectangle1_weights[2001]), .RECT2_X(rectangle2_xs[2001]), .RECT2_Y(rectangle2_ys[2001]), .RECT2_WIDTH(rectangle2_widths[2001]), .RECT2_HEIGHT(rectangle2_heights[2001]), .RECT2_WEIGHT(rectangle2_weights[2001]), .RECT3_X(rectangle3_xs[2001]), .RECT3_Y(rectangle3_ys[2001]), .RECT3_WIDTH(rectangle3_widths[2001]), .RECT3_HEIGHT(rectangle3_heights[2001]), .RECT3_WEIGHT(rectangle3_weights[2001]), .FEAT_THRES(feature_thresholds[2001]), .FEAT_ABOVE(feature_aboves[2001]), .FEAT_BELOW(feature_belows[2001])) ac2001(.scan_win(scan_win2001), .scan_win_std_dev(scan_win_std_dev[2001]), .feature_accum(feature_accums[2001]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2002]), .RECT1_Y(rectangle1_ys[2002]), .RECT1_WIDTH(rectangle1_widths[2002]), .RECT1_HEIGHT(rectangle1_heights[2002]), .RECT1_WEIGHT(rectangle1_weights[2002]), .RECT2_X(rectangle2_xs[2002]), .RECT2_Y(rectangle2_ys[2002]), .RECT2_WIDTH(rectangle2_widths[2002]), .RECT2_HEIGHT(rectangle2_heights[2002]), .RECT2_WEIGHT(rectangle2_weights[2002]), .RECT3_X(rectangle3_xs[2002]), .RECT3_Y(rectangle3_ys[2002]), .RECT3_WIDTH(rectangle3_widths[2002]), .RECT3_HEIGHT(rectangle3_heights[2002]), .RECT3_WEIGHT(rectangle3_weights[2002]), .FEAT_THRES(feature_thresholds[2002]), .FEAT_ABOVE(feature_aboves[2002]), .FEAT_BELOW(feature_belows[2002])) ac2002(.scan_win(scan_win2002), .scan_win_std_dev(scan_win_std_dev[2002]), .feature_accum(feature_accums[2002]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2003]), .RECT1_Y(rectangle1_ys[2003]), .RECT1_WIDTH(rectangle1_widths[2003]), .RECT1_HEIGHT(rectangle1_heights[2003]), .RECT1_WEIGHT(rectangle1_weights[2003]), .RECT2_X(rectangle2_xs[2003]), .RECT2_Y(rectangle2_ys[2003]), .RECT2_WIDTH(rectangle2_widths[2003]), .RECT2_HEIGHT(rectangle2_heights[2003]), .RECT2_WEIGHT(rectangle2_weights[2003]), .RECT3_X(rectangle3_xs[2003]), .RECT3_Y(rectangle3_ys[2003]), .RECT3_WIDTH(rectangle3_widths[2003]), .RECT3_HEIGHT(rectangle3_heights[2003]), .RECT3_WEIGHT(rectangle3_weights[2003]), .FEAT_THRES(feature_thresholds[2003]), .FEAT_ABOVE(feature_aboves[2003]), .FEAT_BELOW(feature_belows[2003])) ac2003(.scan_win(scan_win2003), .scan_win_std_dev(scan_win_std_dev[2003]), .feature_accum(feature_accums[2003]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2004]), .RECT1_Y(rectangle1_ys[2004]), .RECT1_WIDTH(rectangle1_widths[2004]), .RECT1_HEIGHT(rectangle1_heights[2004]), .RECT1_WEIGHT(rectangle1_weights[2004]), .RECT2_X(rectangle2_xs[2004]), .RECT2_Y(rectangle2_ys[2004]), .RECT2_WIDTH(rectangle2_widths[2004]), .RECT2_HEIGHT(rectangle2_heights[2004]), .RECT2_WEIGHT(rectangle2_weights[2004]), .RECT3_X(rectangle3_xs[2004]), .RECT3_Y(rectangle3_ys[2004]), .RECT3_WIDTH(rectangle3_widths[2004]), .RECT3_HEIGHT(rectangle3_heights[2004]), .RECT3_WEIGHT(rectangle3_weights[2004]), .FEAT_THRES(feature_thresholds[2004]), .FEAT_ABOVE(feature_aboves[2004]), .FEAT_BELOW(feature_belows[2004])) ac2004(.scan_win(scan_win2004), .scan_win_std_dev(scan_win_std_dev[2004]), .feature_accum(feature_accums[2004]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2005]), .RECT1_Y(rectangle1_ys[2005]), .RECT1_WIDTH(rectangle1_widths[2005]), .RECT1_HEIGHT(rectangle1_heights[2005]), .RECT1_WEIGHT(rectangle1_weights[2005]), .RECT2_X(rectangle2_xs[2005]), .RECT2_Y(rectangle2_ys[2005]), .RECT2_WIDTH(rectangle2_widths[2005]), .RECT2_HEIGHT(rectangle2_heights[2005]), .RECT2_WEIGHT(rectangle2_weights[2005]), .RECT3_X(rectangle3_xs[2005]), .RECT3_Y(rectangle3_ys[2005]), .RECT3_WIDTH(rectangle3_widths[2005]), .RECT3_HEIGHT(rectangle3_heights[2005]), .RECT3_WEIGHT(rectangle3_weights[2005]), .FEAT_THRES(feature_thresholds[2005]), .FEAT_ABOVE(feature_aboves[2005]), .FEAT_BELOW(feature_belows[2005])) ac2005(.scan_win(scan_win2005), .scan_win_std_dev(scan_win_std_dev[2005]), .feature_accum(feature_accums[2005]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2006]), .RECT1_Y(rectangle1_ys[2006]), .RECT1_WIDTH(rectangle1_widths[2006]), .RECT1_HEIGHT(rectangle1_heights[2006]), .RECT1_WEIGHT(rectangle1_weights[2006]), .RECT2_X(rectangle2_xs[2006]), .RECT2_Y(rectangle2_ys[2006]), .RECT2_WIDTH(rectangle2_widths[2006]), .RECT2_HEIGHT(rectangle2_heights[2006]), .RECT2_WEIGHT(rectangle2_weights[2006]), .RECT3_X(rectangle3_xs[2006]), .RECT3_Y(rectangle3_ys[2006]), .RECT3_WIDTH(rectangle3_widths[2006]), .RECT3_HEIGHT(rectangle3_heights[2006]), .RECT3_WEIGHT(rectangle3_weights[2006]), .FEAT_THRES(feature_thresholds[2006]), .FEAT_ABOVE(feature_aboves[2006]), .FEAT_BELOW(feature_belows[2006])) ac2006(.scan_win(scan_win2006), .scan_win_std_dev(scan_win_std_dev[2006]), .feature_accum(feature_accums[2006]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2007]), .RECT1_Y(rectangle1_ys[2007]), .RECT1_WIDTH(rectangle1_widths[2007]), .RECT1_HEIGHT(rectangle1_heights[2007]), .RECT1_WEIGHT(rectangle1_weights[2007]), .RECT2_X(rectangle2_xs[2007]), .RECT2_Y(rectangle2_ys[2007]), .RECT2_WIDTH(rectangle2_widths[2007]), .RECT2_HEIGHT(rectangle2_heights[2007]), .RECT2_WEIGHT(rectangle2_weights[2007]), .RECT3_X(rectangle3_xs[2007]), .RECT3_Y(rectangle3_ys[2007]), .RECT3_WIDTH(rectangle3_widths[2007]), .RECT3_HEIGHT(rectangle3_heights[2007]), .RECT3_WEIGHT(rectangle3_weights[2007]), .FEAT_THRES(feature_thresholds[2007]), .FEAT_ABOVE(feature_aboves[2007]), .FEAT_BELOW(feature_belows[2007])) ac2007(.scan_win(scan_win2007), .scan_win_std_dev(scan_win_std_dev[2007]), .feature_accum(feature_accums[2007]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2008]), .RECT1_Y(rectangle1_ys[2008]), .RECT1_WIDTH(rectangle1_widths[2008]), .RECT1_HEIGHT(rectangle1_heights[2008]), .RECT1_WEIGHT(rectangle1_weights[2008]), .RECT2_X(rectangle2_xs[2008]), .RECT2_Y(rectangle2_ys[2008]), .RECT2_WIDTH(rectangle2_widths[2008]), .RECT2_HEIGHT(rectangle2_heights[2008]), .RECT2_WEIGHT(rectangle2_weights[2008]), .RECT3_X(rectangle3_xs[2008]), .RECT3_Y(rectangle3_ys[2008]), .RECT3_WIDTH(rectangle3_widths[2008]), .RECT3_HEIGHT(rectangle3_heights[2008]), .RECT3_WEIGHT(rectangle3_weights[2008]), .FEAT_THRES(feature_thresholds[2008]), .FEAT_ABOVE(feature_aboves[2008]), .FEAT_BELOW(feature_belows[2008])) ac2008(.scan_win(scan_win2008), .scan_win_std_dev(scan_win_std_dev[2008]), .feature_accum(feature_accums[2008]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2009]), .RECT1_Y(rectangle1_ys[2009]), .RECT1_WIDTH(rectangle1_widths[2009]), .RECT1_HEIGHT(rectangle1_heights[2009]), .RECT1_WEIGHT(rectangle1_weights[2009]), .RECT2_X(rectangle2_xs[2009]), .RECT2_Y(rectangle2_ys[2009]), .RECT2_WIDTH(rectangle2_widths[2009]), .RECT2_HEIGHT(rectangle2_heights[2009]), .RECT2_WEIGHT(rectangle2_weights[2009]), .RECT3_X(rectangle3_xs[2009]), .RECT3_Y(rectangle3_ys[2009]), .RECT3_WIDTH(rectangle3_widths[2009]), .RECT3_HEIGHT(rectangle3_heights[2009]), .RECT3_WEIGHT(rectangle3_weights[2009]), .FEAT_THRES(feature_thresholds[2009]), .FEAT_ABOVE(feature_aboves[2009]), .FEAT_BELOW(feature_belows[2009])) ac2009(.scan_win(scan_win2009), .scan_win_std_dev(scan_win_std_dev[2009]), .feature_accum(feature_accums[2009]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2010]), .RECT1_Y(rectangle1_ys[2010]), .RECT1_WIDTH(rectangle1_widths[2010]), .RECT1_HEIGHT(rectangle1_heights[2010]), .RECT1_WEIGHT(rectangle1_weights[2010]), .RECT2_X(rectangle2_xs[2010]), .RECT2_Y(rectangle2_ys[2010]), .RECT2_WIDTH(rectangle2_widths[2010]), .RECT2_HEIGHT(rectangle2_heights[2010]), .RECT2_WEIGHT(rectangle2_weights[2010]), .RECT3_X(rectangle3_xs[2010]), .RECT3_Y(rectangle3_ys[2010]), .RECT3_WIDTH(rectangle3_widths[2010]), .RECT3_HEIGHT(rectangle3_heights[2010]), .RECT3_WEIGHT(rectangle3_weights[2010]), .FEAT_THRES(feature_thresholds[2010]), .FEAT_ABOVE(feature_aboves[2010]), .FEAT_BELOW(feature_belows[2010])) ac2010(.scan_win(scan_win2010), .scan_win_std_dev(scan_win_std_dev[2010]), .feature_accum(feature_accums[2010]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2011]), .RECT1_Y(rectangle1_ys[2011]), .RECT1_WIDTH(rectangle1_widths[2011]), .RECT1_HEIGHT(rectangle1_heights[2011]), .RECT1_WEIGHT(rectangle1_weights[2011]), .RECT2_X(rectangle2_xs[2011]), .RECT2_Y(rectangle2_ys[2011]), .RECT2_WIDTH(rectangle2_widths[2011]), .RECT2_HEIGHT(rectangle2_heights[2011]), .RECT2_WEIGHT(rectangle2_weights[2011]), .RECT3_X(rectangle3_xs[2011]), .RECT3_Y(rectangle3_ys[2011]), .RECT3_WIDTH(rectangle3_widths[2011]), .RECT3_HEIGHT(rectangle3_heights[2011]), .RECT3_WEIGHT(rectangle3_weights[2011]), .FEAT_THRES(feature_thresholds[2011]), .FEAT_ABOVE(feature_aboves[2011]), .FEAT_BELOW(feature_belows[2011])) ac2011(.scan_win(scan_win2011), .scan_win_std_dev(scan_win_std_dev[2011]), .feature_accum(feature_accums[2011]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2012]), .RECT1_Y(rectangle1_ys[2012]), .RECT1_WIDTH(rectangle1_widths[2012]), .RECT1_HEIGHT(rectangle1_heights[2012]), .RECT1_WEIGHT(rectangle1_weights[2012]), .RECT2_X(rectangle2_xs[2012]), .RECT2_Y(rectangle2_ys[2012]), .RECT2_WIDTH(rectangle2_widths[2012]), .RECT2_HEIGHT(rectangle2_heights[2012]), .RECT2_WEIGHT(rectangle2_weights[2012]), .RECT3_X(rectangle3_xs[2012]), .RECT3_Y(rectangle3_ys[2012]), .RECT3_WIDTH(rectangle3_widths[2012]), .RECT3_HEIGHT(rectangle3_heights[2012]), .RECT3_WEIGHT(rectangle3_weights[2012]), .FEAT_THRES(feature_thresholds[2012]), .FEAT_ABOVE(feature_aboves[2012]), .FEAT_BELOW(feature_belows[2012])) ac2012(.scan_win(scan_win2012), .scan_win_std_dev(scan_win_std_dev[2012]), .feature_accum(feature_accums[2012]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2013]), .RECT1_Y(rectangle1_ys[2013]), .RECT1_WIDTH(rectangle1_widths[2013]), .RECT1_HEIGHT(rectangle1_heights[2013]), .RECT1_WEIGHT(rectangle1_weights[2013]), .RECT2_X(rectangle2_xs[2013]), .RECT2_Y(rectangle2_ys[2013]), .RECT2_WIDTH(rectangle2_widths[2013]), .RECT2_HEIGHT(rectangle2_heights[2013]), .RECT2_WEIGHT(rectangle2_weights[2013]), .RECT3_X(rectangle3_xs[2013]), .RECT3_Y(rectangle3_ys[2013]), .RECT3_WIDTH(rectangle3_widths[2013]), .RECT3_HEIGHT(rectangle3_heights[2013]), .RECT3_WEIGHT(rectangle3_weights[2013]), .FEAT_THRES(feature_thresholds[2013]), .FEAT_ABOVE(feature_aboves[2013]), .FEAT_BELOW(feature_belows[2013])) ac2013(.scan_win(scan_win2013), .scan_win_std_dev(scan_win_std_dev[2013]), .feature_accum(feature_accums[2013]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2014]), .RECT1_Y(rectangle1_ys[2014]), .RECT1_WIDTH(rectangle1_widths[2014]), .RECT1_HEIGHT(rectangle1_heights[2014]), .RECT1_WEIGHT(rectangle1_weights[2014]), .RECT2_X(rectangle2_xs[2014]), .RECT2_Y(rectangle2_ys[2014]), .RECT2_WIDTH(rectangle2_widths[2014]), .RECT2_HEIGHT(rectangle2_heights[2014]), .RECT2_WEIGHT(rectangle2_weights[2014]), .RECT3_X(rectangle3_xs[2014]), .RECT3_Y(rectangle3_ys[2014]), .RECT3_WIDTH(rectangle3_widths[2014]), .RECT3_HEIGHT(rectangle3_heights[2014]), .RECT3_WEIGHT(rectangle3_weights[2014]), .FEAT_THRES(feature_thresholds[2014]), .FEAT_ABOVE(feature_aboves[2014]), .FEAT_BELOW(feature_belows[2014])) ac2014(.scan_win(scan_win2014), .scan_win_std_dev(scan_win_std_dev[2014]), .feature_accum(feature_accums[2014]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2015]), .RECT1_Y(rectangle1_ys[2015]), .RECT1_WIDTH(rectangle1_widths[2015]), .RECT1_HEIGHT(rectangle1_heights[2015]), .RECT1_WEIGHT(rectangle1_weights[2015]), .RECT2_X(rectangle2_xs[2015]), .RECT2_Y(rectangle2_ys[2015]), .RECT2_WIDTH(rectangle2_widths[2015]), .RECT2_HEIGHT(rectangle2_heights[2015]), .RECT2_WEIGHT(rectangle2_weights[2015]), .RECT3_X(rectangle3_xs[2015]), .RECT3_Y(rectangle3_ys[2015]), .RECT3_WIDTH(rectangle3_widths[2015]), .RECT3_HEIGHT(rectangle3_heights[2015]), .RECT3_WEIGHT(rectangle3_weights[2015]), .FEAT_THRES(feature_thresholds[2015]), .FEAT_ABOVE(feature_aboves[2015]), .FEAT_BELOW(feature_belows[2015])) ac2015(.scan_win(scan_win2015), .scan_win_std_dev(scan_win_std_dev[2015]), .feature_accum(feature_accums[2015]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2016]), .RECT1_Y(rectangle1_ys[2016]), .RECT1_WIDTH(rectangle1_widths[2016]), .RECT1_HEIGHT(rectangle1_heights[2016]), .RECT1_WEIGHT(rectangle1_weights[2016]), .RECT2_X(rectangle2_xs[2016]), .RECT2_Y(rectangle2_ys[2016]), .RECT2_WIDTH(rectangle2_widths[2016]), .RECT2_HEIGHT(rectangle2_heights[2016]), .RECT2_WEIGHT(rectangle2_weights[2016]), .RECT3_X(rectangle3_xs[2016]), .RECT3_Y(rectangle3_ys[2016]), .RECT3_WIDTH(rectangle3_widths[2016]), .RECT3_HEIGHT(rectangle3_heights[2016]), .RECT3_WEIGHT(rectangle3_weights[2016]), .FEAT_THRES(feature_thresholds[2016]), .FEAT_ABOVE(feature_aboves[2016]), .FEAT_BELOW(feature_belows[2016])) ac2016(.scan_win(scan_win2016), .scan_win_std_dev(scan_win_std_dev[2016]), .feature_accum(feature_accums[2016]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2017]), .RECT1_Y(rectangle1_ys[2017]), .RECT1_WIDTH(rectangle1_widths[2017]), .RECT1_HEIGHT(rectangle1_heights[2017]), .RECT1_WEIGHT(rectangle1_weights[2017]), .RECT2_X(rectangle2_xs[2017]), .RECT2_Y(rectangle2_ys[2017]), .RECT2_WIDTH(rectangle2_widths[2017]), .RECT2_HEIGHT(rectangle2_heights[2017]), .RECT2_WEIGHT(rectangle2_weights[2017]), .RECT3_X(rectangle3_xs[2017]), .RECT3_Y(rectangle3_ys[2017]), .RECT3_WIDTH(rectangle3_widths[2017]), .RECT3_HEIGHT(rectangle3_heights[2017]), .RECT3_WEIGHT(rectangle3_weights[2017]), .FEAT_THRES(feature_thresholds[2017]), .FEAT_ABOVE(feature_aboves[2017]), .FEAT_BELOW(feature_belows[2017])) ac2017(.scan_win(scan_win2017), .scan_win_std_dev(scan_win_std_dev[2017]), .feature_accum(feature_accums[2017]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2018]), .RECT1_Y(rectangle1_ys[2018]), .RECT1_WIDTH(rectangle1_widths[2018]), .RECT1_HEIGHT(rectangle1_heights[2018]), .RECT1_WEIGHT(rectangle1_weights[2018]), .RECT2_X(rectangle2_xs[2018]), .RECT2_Y(rectangle2_ys[2018]), .RECT2_WIDTH(rectangle2_widths[2018]), .RECT2_HEIGHT(rectangle2_heights[2018]), .RECT2_WEIGHT(rectangle2_weights[2018]), .RECT3_X(rectangle3_xs[2018]), .RECT3_Y(rectangle3_ys[2018]), .RECT3_WIDTH(rectangle3_widths[2018]), .RECT3_HEIGHT(rectangle3_heights[2018]), .RECT3_WEIGHT(rectangle3_weights[2018]), .FEAT_THRES(feature_thresholds[2018]), .FEAT_ABOVE(feature_aboves[2018]), .FEAT_BELOW(feature_belows[2018])) ac2018(.scan_win(scan_win2018), .scan_win_std_dev(scan_win_std_dev[2018]), .feature_accum(feature_accums[2018]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2019]), .RECT1_Y(rectangle1_ys[2019]), .RECT1_WIDTH(rectangle1_widths[2019]), .RECT1_HEIGHT(rectangle1_heights[2019]), .RECT1_WEIGHT(rectangle1_weights[2019]), .RECT2_X(rectangle2_xs[2019]), .RECT2_Y(rectangle2_ys[2019]), .RECT2_WIDTH(rectangle2_widths[2019]), .RECT2_HEIGHT(rectangle2_heights[2019]), .RECT2_WEIGHT(rectangle2_weights[2019]), .RECT3_X(rectangle3_xs[2019]), .RECT3_Y(rectangle3_ys[2019]), .RECT3_WIDTH(rectangle3_widths[2019]), .RECT3_HEIGHT(rectangle3_heights[2019]), .RECT3_WEIGHT(rectangle3_weights[2019]), .FEAT_THRES(feature_thresholds[2019]), .FEAT_ABOVE(feature_aboves[2019]), .FEAT_BELOW(feature_belows[2019])) ac2019(.scan_win(scan_win2019), .scan_win_std_dev(scan_win_std_dev[2019]), .feature_accum(feature_accums[2019]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2020]), .RECT1_Y(rectangle1_ys[2020]), .RECT1_WIDTH(rectangle1_widths[2020]), .RECT1_HEIGHT(rectangle1_heights[2020]), .RECT1_WEIGHT(rectangle1_weights[2020]), .RECT2_X(rectangle2_xs[2020]), .RECT2_Y(rectangle2_ys[2020]), .RECT2_WIDTH(rectangle2_widths[2020]), .RECT2_HEIGHT(rectangle2_heights[2020]), .RECT2_WEIGHT(rectangle2_weights[2020]), .RECT3_X(rectangle3_xs[2020]), .RECT3_Y(rectangle3_ys[2020]), .RECT3_WIDTH(rectangle3_widths[2020]), .RECT3_HEIGHT(rectangle3_heights[2020]), .RECT3_WEIGHT(rectangle3_weights[2020]), .FEAT_THRES(feature_thresholds[2020]), .FEAT_ABOVE(feature_aboves[2020]), .FEAT_BELOW(feature_belows[2020])) ac2020(.scan_win(scan_win2020), .scan_win_std_dev(scan_win_std_dev[2020]), .feature_accum(feature_accums[2020]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2021]), .RECT1_Y(rectangle1_ys[2021]), .RECT1_WIDTH(rectangle1_widths[2021]), .RECT1_HEIGHT(rectangle1_heights[2021]), .RECT1_WEIGHT(rectangle1_weights[2021]), .RECT2_X(rectangle2_xs[2021]), .RECT2_Y(rectangle2_ys[2021]), .RECT2_WIDTH(rectangle2_widths[2021]), .RECT2_HEIGHT(rectangle2_heights[2021]), .RECT2_WEIGHT(rectangle2_weights[2021]), .RECT3_X(rectangle3_xs[2021]), .RECT3_Y(rectangle3_ys[2021]), .RECT3_WIDTH(rectangle3_widths[2021]), .RECT3_HEIGHT(rectangle3_heights[2021]), .RECT3_WEIGHT(rectangle3_weights[2021]), .FEAT_THRES(feature_thresholds[2021]), .FEAT_ABOVE(feature_aboves[2021]), .FEAT_BELOW(feature_belows[2021])) ac2021(.scan_win(scan_win2021), .scan_win_std_dev(scan_win_std_dev[2021]), .feature_accum(feature_accums[2021]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2022]), .RECT1_Y(rectangle1_ys[2022]), .RECT1_WIDTH(rectangle1_widths[2022]), .RECT1_HEIGHT(rectangle1_heights[2022]), .RECT1_WEIGHT(rectangle1_weights[2022]), .RECT2_X(rectangle2_xs[2022]), .RECT2_Y(rectangle2_ys[2022]), .RECT2_WIDTH(rectangle2_widths[2022]), .RECT2_HEIGHT(rectangle2_heights[2022]), .RECT2_WEIGHT(rectangle2_weights[2022]), .RECT3_X(rectangle3_xs[2022]), .RECT3_Y(rectangle3_ys[2022]), .RECT3_WIDTH(rectangle3_widths[2022]), .RECT3_HEIGHT(rectangle3_heights[2022]), .RECT3_WEIGHT(rectangle3_weights[2022]), .FEAT_THRES(feature_thresholds[2022]), .FEAT_ABOVE(feature_aboves[2022]), .FEAT_BELOW(feature_belows[2022])) ac2022(.scan_win(scan_win2022), .scan_win_std_dev(scan_win_std_dev[2022]), .feature_accum(feature_accums[2022]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2023]), .RECT1_Y(rectangle1_ys[2023]), .RECT1_WIDTH(rectangle1_widths[2023]), .RECT1_HEIGHT(rectangle1_heights[2023]), .RECT1_WEIGHT(rectangle1_weights[2023]), .RECT2_X(rectangle2_xs[2023]), .RECT2_Y(rectangle2_ys[2023]), .RECT2_WIDTH(rectangle2_widths[2023]), .RECT2_HEIGHT(rectangle2_heights[2023]), .RECT2_WEIGHT(rectangle2_weights[2023]), .RECT3_X(rectangle3_xs[2023]), .RECT3_Y(rectangle3_ys[2023]), .RECT3_WIDTH(rectangle3_widths[2023]), .RECT3_HEIGHT(rectangle3_heights[2023]), .RECT3_WEIGHT(rectangle3_weights[2023]), .FEAT_THRES(feature_thresholds[2023]), .FEAT_ABOVE(feature_aboves[2023]), .FEAT_BELOW(feature_belows[2023])) ac2023(.scan_win(scan_win2023), .scan_win_std_dev(scan_win_std_dev[2023]), .feature_accum(feature_accums[2023]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2024]), .RECT1_Y(rectangle1_ys[2024]), .RECT1_WIDTH(rectangle1_widths[2024]), .RECT1_HEIGHT(rectangle1_heights[2024]), .RECT1_WEIGHT(rectangle1_weights[2024]), .RECT2_X(rectangle2_xs[2024]), .RECT2_Y(rectangle2_ys[2024]), .RECT2_WIDTH(rectangle2_widths[2024]), .RECT2_HEIGHT(rectangle2_heights[2024]), .RECT2_WEIGHT(rectangle2_weights[2024]), .RECT3_X(rectangle3_xs[2024]), .RECT3_Y(rectangle3_ys[2024]), .RECT3_WIDTH(rectangle3_widths[2024]), .RECT3_HEIGHT(rectangle3_heights[2024]), .RECT3_WEIGHT(rectangle3_weights[2024]), .FEAT_THRES(feature_thresholds[2024]), .FEAT_ABOVE(feature_aboves[2024]), .FEAT_BELOW(feature_belows[2024])) ac2024(.scan_win(scan_win2024), .scan_win_std_dev(scan_win_std_dev[2024]), .feature_accum(feature_accums[2024]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2025]), .RECT1_Y(rectangle1_ys[2025]), .RECT1_WIDTH(rectangle1_widths[2025]), .RECT1_HEIGHT(rectangle1_heights[2025]), .RECT1_WEIGHT(rectangle1_weights[2025]), .RECT2_X(rectangle2_xs[2025]), .RECT2_Y(rectangle2_ys[2025]), .RECT2_WIDTH(rectangle2_widths[2025]), .RECT2_HEIGHT(rectangle2_heights[2025]), .RECT2_WEIGHT(rectangle2_weights[2025]), .RECT3_X(rectangle3_xs[2025]), .RECT3_Y(rectangle3_ys[2025]), .RECT3_WIDTH(rectangle3_widths[2025]), .RECT3_HEIGHT(rectangle3_heights[2025]), .RECT3_WEIGHT(rectangle3_weights[2025]), .FEAT_THRES(feature_thresholds[2025]), .FEAT_ABOVE(feature_aboves[2025]), .FEAT_BELOW(feature_belows[2025])) ac2025(.scan_win(scan_win2025), .scan_win_std_dev(scan_win_std_dev[2025]), .feature_accum(feature_accums[2025]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2026]), .RECT1_Y(rectangle1_ys[2026]), .RECT1_WIDTH(rectangle1_widths[2026]), .RECT1_HEIGHT(rectangle1_heights[2026]), .RECT1_WEIGHT(rectangle1_weights[2026]), .RECT2_X(rectangle2_xs[2026]), .RECT2_Y(rectangle2_ys[2026]), .RECT2_WIDTH(rectangle2_widths[2026]), .RECT2_HEIGHT(rectangle2_heights[2026]), .RECT2_WEIGHT(rectangle2_weights[2026]), .RECT3_X(rectangle3_xs[2026]), .RECT3_Y(rectangle3_ys[2026]), .RECT3_WIDTH(rectangle3_widths[2026]), .RECT3_HEIGHT(rectangle3_heights[2026]), .RECT3_WEIGHT(rectangle3_weights[2026]), .FEAT_THRES(feature_thresholds[2026]), .FEAT_ABOVE(feature_aboves[2026]), .FEAT_BELOW(feature_belows[2026])) ac2026(.scan_win(scan_win2026), .scan_win_std_dev(scan_win_std_dev[2026]), .feature_accum(feature_accums[2026]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2027]), .RECT1_Y(rectangle1_ys[2027]), .RECT1_WIDTH(rectangle1_widths[2027]), .RECT1_HEIGHT(rectangle1_heights[2027]), .RECT1_WEIGHT(rectangle1_weights[2027]), .RECT2_X(rectangle2_xs[2027]), .RECT2_Y(rectangle2_ys[2027]), .RECT2_WIDTH(rectangle2_widths[2027]), .RECT2_HEIGHT(rectangle2_heights[2027]), .RECT2_WEIGHT(rectangle2_weights[2027]), .RECT3_X(rectangle3_xs[2027]), .RECT3_Y(rectangle3_ys[2027]), .RECT3_WIDTH(rectangle3_widths[2027]), .RECT3_HEIGHT(rectangle3_heights[2027]), .RECT3_WEIGHT(rectangle3_weights[2027]), .FEAT_THRES(feature_thresholds[2027]), .FEAT_ABOVE(feature_aboves[2027]), .FEAT_BELOW(feature_belows[2027])) ac2027(.scan_win(scan_win2027), .scan_win_std_dev(scan_win_std_dev[2027]), .feature_accum(feature_accums[2027]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2028]), .RECT1_Y(rectangle1_ys[2028]), .RECT1_WIDTH(rectangle1_widths[2028]), .RECT1_HEIGHT(rectangle1_heights[2028]), .RECT1_WEIGHT(rectangle1_weights[2028]), .RECT2_X(rectangle2_xs[2028]), .RECT2_Y(rectangle2_ys[2028]), .RECT2_WIDTH(rectangle2_widths[2028]), .RECT2_HEIGHT(rectangle2_heights[2028]), .RECT2_WEIGHT(rectangle2_weights[2028]), .RECT3_X(rectangle3_xs[2028]), .RECT3_Y(rectangle3_ys[2028]), .RECT3_WIDTH(rectangle3_widths[2028]), .RECT3_HEIGHT(rectangle3_heights[2028]), .RECT3_WEIGHT(rectangle3_weights[2028]), .FEAT_THRES(feature_thresholds[2028]), .FEAT_ABOVE(feature_aboves[2028]), .FEAT_BELOW(feature_belows[2028])) ac2028(.scan_win(scan_win2028), .scan_win_std_dev(scan_win_std_dev[2028]), .feature_accum(feature_accums[2028]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2029]), .RECT1_Y(rectangle1_ys[2029]), .RECT1_WIDTH(rectangle1_widths[2029]), .RECT1_HEIGHT(rectangle1_heights[2029]), .RECT1_WEIGHT(rectangle1_weights[2029]), .RECT2_X(rectangle2_xs[2029]), .RECT2_Y(rectangle2_ys[2029]), .RECT2_WIDTH(rectangle2_widths[2029]), .RECT2_HEIGHT(rectangle2_heights[2029]), .RECT2_WEIGHT(rectangle2_weights[2029]), .RECT3_X(rectangle3_xs[2029]), .RECT3_Y(rectangle3_ys[2029]), .RECT3_WIDTH(rectangle3_widths[2029]), .RECT3_HEIGHT(rectangle3_heights[2029]), .RECT3_WEIGHT(rectangle3_weights[2029]), .FEAT_THRES(feature_thresholds[2029]), .FEAT_ABOVE(feature_aboves[2029]), .FEAT_BELOW(feature_belows[2029])) ac2029(.scan_win(scan_win2029), .scan_win_std_dev(scan_win_std_dev[2029]), .feature_accum(feature_accums[2029]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2030]), .RECT1_Y(rectangle1_ys[2030]), .RECT1_WIDTH(rectangle1_widths[2030]), .RECT1_HEIGHT(rectangle1_heights[2030]), .RECT1_WEIGHT(rectangle1_weights[2030]), .RECT2_X(rectangle2_xs[2030]), .RECT2_Y(rectangle2_ys[2030]), .RECT2_WIDTH(rectangle2_widths[2030]), .RECT2_HEIGHT(rectangle2_heights[2030]), .RECT2_WEIGHT(rectangle2_weights[2030]), .RECT3_X(rectangle3_xs[2030]), .RECT3_Y(rectangle3_ys[2030]), .RECT3_WIDTH(rectangle3_widths[2030]), .RECT3_HEIGHT(rectangle3_heights[2030]), .RECT3_WEIGHT(rectangle3_weights[2030]), .FEAT_THRES(feature_thresholds[2030]), .FEAT_ABOVE(feature_aboves[2030]), .FEAT_BELOW(feature_belows[2030])) ac2030(.scan_win(scan_win2030), .scan_win_std_dev(scan_win_std_dev[2030]), .feature_accum(feature_accums[2030]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2031]), .RECT1_Y(rectangle1_ys[2031]), .RECT1_WIDTH(rectangle1_widths[2031]), .RECT1_HEIGHT(rectangle1_heights[2031]), .RECT1_WEIGHT(rectangle1_weights[2031]), .RECT2_X(rectangle2_xs[2031]), .RECT2_Y(rectangle2_ys[2031]), .RECT2_WIDTH(rectangle2_widths[2031]), .RECT2_HEIGHT(rectangle2_heights[2031]), .RECT2_WEIGHT(rectangle2_weights[2031]), .RECT3_X(rectangle3_xs[2031]), .RECT3_Y(rectangle3_ys[2031]), .RECT3_WIDTH(rectangle3_widths[2031]), .RECT3_HEIGHT(rectangle3_heights[2031]), .RECT3_WEIGHT(rectangle3_weights[2031]), .FEAT_THRES(feature_thresholds[2031]), .FEAT_ABOVE(feature_aboves[2031]), .FEAT_BELOW(feature_belows[2031])) ac2031(.scan_win(scan_win2031), .scan_win_std_dev(scan_win_std_dev[2031]), .feature_accum(feature_accums[2031]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2032]), .RECT1_Y(rectangle1_ys[2032]), .RECT1_WIDTH(rectangle1_widths[2032]), .RECT1_HEIGHT(rectangle1_heights[2032]), .RECT1_WEIGHT(rectangle1_weights[2032]), .RECT2_X(rectangle2_xs[2032]), .RECT2_Y(rectangle2_ys[2032]), .RECT2_WIDTH(rectangle2_widths[2032]), .RECT2_HEIGHT(rectangle2_heights[2032]), .RECT2_WEIGHT(rectangle2_weights[2032]), .RECT3_X(rectangle3_xs[2032]), .RECT3_Y(rectangle3_ys[2032]), .RECT3_WIDTH(rectangle3_widths[2032]), .RECT3_HEIGHT(rectangle3_heights[2032]), .RECT3_WEIGHT(rectangle3_weights[2032]), .FEAT_THRES(feature_thresholds[2032]), .FEAT_ABOVE(feature_aboves[2032]), .FEAT_BELOW(feature_belows[2032])) ac2032(.scan_win(scan_win2032), .scan_win_std_dev(scan_win_std_dev[2032]), .feature_accum(feature_accums[2032]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2033]), .RECT1_Y(rectangle1_ys[2033]), .RECT1_WIDTH(rectangle1_widths[2033]), .RECT1_HEIGHT(rectangle1_heights[2033]), .RECT1_WEIGHT(rectangle1_weights[2033]), .RECT2_X(rectangle2_xs[2033]), .RECT2_Y(rectangle2_ys[2033]), .RECT2_WIDTH(rectangle2_widths[2033]), .RECT2_HEIGHT(rectangle2_heights[2033]), .RECT2_WEIGHT(rectangle2_weights[2033]), .RECT3_X(rectangle3_xs[2033]), .RECT3_Y(rectangle3_ys[2033]), .RECT3_WIDTH(rectangle3_widths[2033]), .RECT3_HEIGHT(rectangle3_heights[2033]), .RECT3_WEIGHT(rectangle3_weights[2033]), .FEAT_THRES(feature_thresholds[2033]), .FEAT_ABOVE(feature_aboves[2033]), .FEAT_BELOW(feature_belows[2033])) ac2033(.scan_win(scan_win2033), .scan_win_std_dev(scan_win_std_dev[2033]), .feature_accum(feature_accums[2033]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2034]), .RECT1_Y(rectangle1_ys[2034]), .RECT1_WIDTH(rectangle1_widths[2034]), .RECT1_HEIGHT(rectangle1_heights[2034]), .RECT1_WEIGHT(rectangle1_weights[2034]), .RECT2_X(rectangle2_xs[2034]), .RECT2_Y(rectangle2_ys[2034]), .RECT2_WIDTH(rectangle2_widths[2034]), .RECT2_HEIGHT(rectangle2_heights[2034]), .RECT2_WEIGHT(rectangle2_weights[2034]), .RECT3_X(rectangle3_xs[2034]), .RECT3_Y(rectangle3_ys[2034]), .RECT3_WIDTH(rectangle3_widths[2034]), .RECT3_HEIGHT(rectangle3_heights[2034]), .RECT3_WEIGHT(rectangle3_weights[2034]), .FEAT_THRES(feature_thresholds[2034]), .FEAT_ABOVE(feature_aboves[2034]), .FEAT_BELOW(feature_belows[2034])) ac2034(.scan_win(scan_win2034), .scan_win_std_dev(scan_win_std_dev[2034]), .feature_accum(feature_accums[2034]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2035]), .RECT1_Y(rectangle1_ys[2035]), .RECT1_WIDTH(rectangle1_widths[2035]), .RECT1_HEIGHT(rectangle1_heights[2035]), .RECT1_WEIGHT(rectangle1_weights[2035]), .RECT2_X(rectangle2_xs[2035]), .RECT2_Y(rectangle2_ys[2035]), .RECT2_WIDTH(rectangle2_widths[2035]), .RECT2_HEIGHT(rectangle2_heights[2035]), .RECT2_WEIGHT(rectangle2_weights[2035]), .RECT3_X(rectangle3_xs[2035]), .RECT3_Y(rectangle3_ys[2035]), .RECT3_WIDTH(rectangle3_widths[2035]), .RECT3_HEIGHT(rectangle3_heights[2035]), .RECT3_WEIGHT(rectangle3_weights[2035]), .FEAT_THRES(feature_thresholds[2035]), .FEAT_ABOVE(feature_aboves[2035]), .FEAT_BELOW(feature_belows[2035])) ac2035(.scan_win(scan_win2035), .scan_win_std_dev(scan_win_std_dev[2035]), .feature_accum(feature_accums[2035]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2036]), .RECT1_Y(rectangle1_ys[2036]), .RECT1_WIDTH(rectangle1_widths[2036]), .RECT1_HEIGHT(rectangle1_heights[2036]), .RECT1_WEIGHT(rectangle1_weights[2036]), .RECT2_X(rectangle2_xs[2036]), .RECT2_Y(rectangle2_ys[2036]), .RECT2_WIDTH(rectangle2_widths[2036]), .RECT2_HEIGHT(rectangle2_heights[2036]), .RECT2_WEIGHT(rectangle2_weights[2036]), .RECT3_X(rectangle3_xs[2036]), .RECT3_Y(rectangle3_ys[2036]), .RECT3_WIDTH(rectangle3_widths[2036]), .RECT3_HEIGHT(rectangle3_heights[2036]), .RECT3_WEIGHT(rectangle3_weights[2036]), .FEAT_THRES(feature_thresholds[2036]), .FEAT_ABOVE(feature_aboves[2036]), .FEAT_BELOW(feature_belows[2036])) ac2036(.scan_win(scan_win2036), .scan_win_std_dev(scan_win_std_dev[2036]), .feature_accum(feature_accums[2036]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2037]), .RECT1_Y(rectangle1_ys[2037]), .RECT1_WIDTH(rectangle1_widths[2037]), .RECT1_HEIGHT(rectangle1_heights[2037]), .RECT1_WEIGHT(rectangle1_weights[2037]), .RECT2_X(rectangle2_xs[2037]), .RECT2_Y(rectangle2_ys[2037]), .RECT2_WIDTH(rectangle2_widths[2037]), .RECT2_HEIGHT(rectangle2_heights[2037]), .RECT2_WEIGHT(rectangle2_weights[2037]), .RECT3_X(rectangle3_xs[2037]), .RECT3_Y(rectangle3_ys[2037]), .RECT3_WIDTH(rectangle3_widths[2037]), .RECT3_HEIGHT(rectangle3_heights[2037]), .RECT3_WEIGHT(rectangle3_weights[2037]), .FEAT_THRES(feature_thresholds[2037]), .FEAT_ABOVE(feature_aboves[2037]), .FEAT_BELOW(feature_belows[2037])) ac2037(.scan_win(scan_win2037), .scan_win_std_dev(scan_win_std_dev[2037]), .feature_accum(feature_accums[2037]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2038]), .RECT1_Y(rectangle1_ys[2038]), .RECT1_WIDTH(rectangle1_widths[2038]), .RECT1_HEIGHT(rectangle1_heights[2038]), .RECT1_WEIGHT(rectangle1_weights[2038]), .RECT2_X(rectangle2_xs[2038]), .RECT2_Y(rectangle2_ys[2038]), .RECT2_WIDTH(rectangle2_widths[2038]), .RECT2_HEIGHT(rectangle2_heights[2038]), .RECT2_WEIGHT(rectangle2_weights[2038]), .RECT3_X(rectangle3_xs[2038]), .RECT3_Y(rectangle3_ys[2038]), .RECT3_WIDTH(rectangle3_widths[2038]), .RECT3_HEIGHT(rectangle3_heights[2038]), .RECT3_WEIGHT(rectangle3_weights[2038]), .FEAT_THRES(feature_thresholds[2038]), .FEAT_ABOVE(feature_aboves[2038]), .FEAT_BELOW(feature_belows[2038])) ac2038(.scan_win(scan_win2038), .scan_win_std_dev(scan_win_std_dev[2038]), .feature_accum(feature_accums[2038]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2039]), .RECT1_Y(rectangle1_ys[2039]), .RECT1_WIDTH(rectangle1_widths[2039]), .RECT1_HEIGHT(rectangle1_heights[2039]), .RECT1_WEIGHT(rectangle1_weights[2039]), .RECT2_X(rectangle2_xs[2039]), .RECT2_Y(rectangle2_ys[2039]), .RECT2_WIDTH(rectangle2_widths[2039]), .RECT2_HEIGHT(rectangle2_heights[2039]), .RECT2_WEIGHT(rectangle2_weights[2039]), .RECT3_X(rectangle3_xs[2039]), .RECT3_Y(rectangle3_ys[2039]), .RECT3_WIDTH(rectangle3_widths[2039]), .RECT3_HEIGHT(rectangle3_heights[2039]), .RECT3_WEIGHT(rectangle3_weights[2039]), .FEAT_THRES(feature_thresholds[2039]), .FEAT_ABOVE(feature_aboves[2039]), .FEAT_BELOW(feature_belows[2039])) ac2039(.scan_win(scan_win2039), .scan_win_std_dev(scan_win_std_dev[2039]), .feature_accum(feature_accums[2039]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2040]), .RECT1_Y(rectangle1_ys[2040]), .RECT1_WIDTH(rectangle1_widths[2040]), .RECT1_HEIGHT(rectangle1_heights[2040]), .RECT1_WEIGHT(rectangle1_weights[2040]), .RECT2_X(rectangle2_xs[2040]), .RECT2_Y(rectangle2_ys[2040]), .RECT2_WIDTH(rectangle2_widths[2040]), .RECT2_HEIGHT(rectangle2_heights[2040]), .RECT2_WEIGHT(rectangle2_weights[2040]), .RECT3_X(rectangle3_xs[2040]), .RECT3_Y(rectangle3_ys[2040]), .RECT3_WIDTH(rectangle3_widths[2040]), .RECT3_HEIGHT(rectangle3_heights[2040]), .RECT3_WEIGHT(rectangle3_weights[2040]), .FEAT_THRES(feature_thresholds[2040]), .FEAT_ABOVE(feature_aboves[2040]), .FEAT_BELOW(feature_belows[2040])) ac2040(.scan_win(scan_win2040), .scan_win_std_dev(scan_win_std_dev[2040]), .feature_accum(feature_accums[2040]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2041]), .RECT1_Y(rectangle1_ys[2041]), .RECT1_WIDTH(rectangle1_widths[2041]), .RECT1_HEIGHT(rectangle1_heights[2041]), .RECT1_WEIGHT(rectangle1_weights[2041]), .RECT2_X(rectangle2_xs[2041]), .RECT2_Y(rectangle2_ys[2041]), .RECT2_WIDTH(rectangle2_widths[2041]), .RECT2_HEIGHT(rectangle2_heights[2041]), .RECT2_WEIGHT(rectangle2_weights[2041]), .RECT3_X(rectangle3_xs[2041]), .RECT3_Y(rectangle3_ys[2041]), .RECT3_WIDTH(rectangle3_widths[2041]), .RECT3_HEIGHT(rectangle3_heights[2041]), .RECT3_WEIGHT(rectangle3_weights[2041]), .FEAT_THRES(feature_thresholds[2041]), .FEAT_ABOVE(feature_aboves[2041]), .FEAT_BELOW(feature_belows[2041])) ac2041(.scan_win(scan_win2041), .scan_win_std_dev(scan_win_std_dev[2041]), .feature_accum(feature_accums[2041]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2042]), .RECT1_Y(rectangle1_ys[2042]), .RECT1_WIDTH(rectangle1_widths[2042]), .RECT1_HEIGHT(rectangle1_heights[2042]), .RECT1_WEIGHT(rectangle1_weights[2042]), .RECT2_X(rectangle2_xs[2042]), .RECT2_Y(rectangle2_ys[2042]), .RECT2_WIDTH(rectangle2_widths[2042]), .RECT2_HEIGHT(rectangle2_heights[2042]), .RECT2_WEIGHT(rectangle2_weights[2042]), .RECT3_X(rectangle3_xs[2042]), .RECT3_Y(rectangle3_ys[2042]), .RECT3_WIDTH(rectangle3_widths[2042]), .RECT3_HEIGHT(rectangle3_heights[2042]), .RECT3_WEIGHT(rectangle3_weights[2042]), .FEAT_THRES(feature_thresholds[2042]), .FEAT_ABOVE(feature_aboves[2042]), .FEAT_BELOW(feature_belows[2042])) ac2042(.scan_win(scan_win2042), .scan_win_std_dev(scan_win_std_dev[2042]), .feature_accum(feature_accums[2042]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2043]), .RECT1_Y(rectangle1_ys[2043]), .RECT1_WIDTH(rectangle1_widths[2043]), .RECT1_HEIGHT(rectangle1_heights[2043]), .RECT1_WEIGHT(rectangle1_weights[2043]), .RECT2_X(rectangle2_xs[2043]), .RECT2_Y(rectangle2_ys[2043]), .RECT2_WIDTH(rectangle2_widths[2043]), .RECT2_HEIGHT(rectangle2_heights[2043]), .RECT2_WEIGHT(rectangle2_weights[2043]), .RECT3_X(rectangle3_xs[2043]), .RECT3_Y(rectangle3_ys[2043]), .RECT3_WIDTH(rectangle3_widths[2043]), .RECT3_HEIGHT(rectangle3_heights[2043]), .RECT3_WEIGHT(rectangle3_weights[2043]), .FEAT_THRES(feature_thresholds[2043]), .FEAT_ABOVE(feature_aboves[2043]), .FEAT_BELOW(feature_belows[2043])) ac2043(.scan_win(scan_win2043), .scan_win_std_dev(scan_win_std_dev[2043]), .feature_accum(feature_accums[2043]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2044]), .RECT1_Y(rectangle1_ys[2044]), .RECT1_WIDTH(rectangle1_widths[2044]), .RECT1_HEIGHT(rectangle1_heights[2044]), .RECT1_WEIGHT(rectangle1_weights[2044]), .RECT2_X(rectangle2_xs[2044]), .RECT2_Y(rectangle2_ys[2044]), .RECT2_WIDTH(rectangle2_widths[2044]), .RECT2_HEIGHT(rectangle2_heights[2044]), .RECT2_WEIGHT(rectangle2_weights[2044]), .RECT3_X(rectangle3_xs[2044]), .RECT3_Y(rectangle3_ys[2044]), .RECT3_WIDTH(rectangle3_widths[2044]), .RECT3_HEIGHT(rectangle3_heights[2044]), .RECT3_WEIGHT(rectangle3_weights[2044]), .FEAT_THRES(feature_thresholds[2044]), .FEAT_ABOVE(feature_aboves[2044]), .FEAT_BELOW(feature_belows[2044])) ac2044(.scan_win(scan_win2044), .scan_win_std_dev(scan_win_std_dev[2044]), .feature_accum(feature_accums[2044]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2045]), .RECT1_Y(rectangle1_ys[2045]), .RECT1_WIDTH(rectangle1_widths[2045]), .RECT1_HEIGHT(rectangle1_heights[2045]), .RECT1_WEIGHT(rectangle1_weights[2045]), .RECT2_X(rectangle2_xs[2045]), .RECT2_Y(rectangle2_ys[2045]), .RECT2_WIDTH(rectangle2_widths[2045]), .RECT2_HEIGHT(rectangle2_heights[2045]), .RECT2_WEIGHT(rectangle2_weights[2045]), .RECT3_X(rectangle3_xs[2045]), .RECT3_Y(rectangle3_ys[2045]), .RECT3_WIDTH(rectangle3_widths[2045]), .RECT3_HEIGHT(rectangle3_heights[2045]), .RECT3_WEIGHT(rectangle3_weights[2045]), .FEAT_THRES(feature_thresholds[2045]), .FEAT_ABOVE(feature_aboves[2045]), .FEAT_BELOW(feature_belows[2045])) ac2045(.scan_win(scan_win2045), .scan_win_std_dev(scan_win_std_dev[2045]), .feature_accum(feature_accums[2045]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2046]), .RECT1_Y(rectangle1_ys[2046]), .RECT1_WIDTH(rectangle1_widths[2046]), .RECT1_HEIGHT(rectangle1_heights[2046]), .RECT1_WEIGHT(rectangle1_weights[2046]), .RECT2_X(rectangle2_xs[2046]), .RECT2_Y(rectangle2_ys[2046]), .RECT2_WIDTH(rectangle2_widths[2046]), .RECT2_HEIGHT(rectangle2_heights[2046]), .RECT2_WEIGHT(rectangle2_weights[2046]), .RECT3_X(rectangle3_xs[2046]), .RECT3_Y(rectangle3_ys[2046]), .RECT3_WIDTH(rectangle3_widths[2046]), .RECT3_HEIGHT(rectangle3_heights[2046]), .RECT3_WEIGHT(rectangle3_weights[2046]), .FEAT_THRES(feature_thresholds[2046]), .FEAT_ABOVE(feature_aboves[2046]), .FEAT_BELOW(feature_belows[2046])) ac2046(.scan_win(scan_win2046), .scan_win_std_dev(scan_win_std_dev[2046]), .feature_accum(feature_accums[2046]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2047]), .RECT1_Y(rectangle1_ys[2047]), .RECT1_WIDTH(rectangle1_widths[2047]), .RECT1_HEIGHT(rectangle1_heights[2047]), .RECT1_WEIGHT(rectangle1_weights[2047]), .RECT2_X(rectangle2_xs[2047]), .RECT2_Y(rectangle2_ys[2047]), .RECT2_WIDTH(rectangle2_widths[2047]), .RECT2_HEIGHT(rectangle2_heights[2047]), .RECT2_WEIGHT(rectangle2_weights[2047]), .RECT3_X(rectangle3_xs[2047]), .RECT3_Y(rectangle3_ys[2047]), .RECT3_WIDTH(rectangle3_widths[2047]), .RECT3_HEIGHT(rectangle3_heights[2047]), .RECT3_WEIGHT(rectangle3_weights[2047]), .FEAT_THRES(feature_thresholds[2047]), .FEAT_ABOVE(feature_aboves[2047]), .FEAT_BELOW(feature_belows[2047])) ac2047(.scan_win(scan_win2047), .scan_win_std_dev(scan_win_std_dev[2047]), .feature_accum(feature_accums[2047]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2048]), .RECT1_Y(rectangle1_ys[2048]), .RECT1_WIDTH(rectangle1_widths[2048]), .RECT1_HEIGHT(rectangle1_heights[2048]), .RECT1_WEIGHT(rectangle1_weights[2048]), .RECT2_X(rectangle2_xs[2048]), .RECT2_Y(rectangle2_ys[2048]), .RECT2_WIDTH(rectangle2_widths[2048]), .RECT2_HEIGHT(rectangle2_heights[2048]), .RECT2_WEIGHT(rectangle2_weights[2048]), .RECT3_X(rectangle3_xs[2048]), .RECT3_Y(rectangle3_ys[2048]), .RECT3_WIDTH(rectangle3_widths[2048]), .RECT3_HEIGHT(rectangle3_heights[2048]), .RECT3_WEIGHT(rectangle3_weights[2048]), .FEAT_THRES(feature_thresholds[2048]), .FEAT_ABOVE(feature_aboves[2048]), .FEAT_BELOW(feature_belows[2048])) ac2048(.scan_win(scan_win2048), .scan_win_std_dev(scan_win_std_dev[2048]), .feature_accum(feature_accums[2048]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2049]), .RECT1_Y(rectangle1_ys[2049]), .RECT1_WIDTH(rectangle1_widths[2049]), .RECT1_HEIGHT(rectangle1_heights[2049]), .RECT1_WEIGHT(rectangle1_weights[2049]), .RECT2_X(rectangle2_xs[2049]), .RECT2_Y(rectangle2_ys[2049]), .RECT2_WIDTH(rectangle2_widths[2049]), .RECT2_HEIGHT(rectangle2_heights[2049]), .RECT2_WEIGHT(rectangle2_weights[2049]), .RECT3_X(rectangle3_xs[2049]), .RECT3_Y(rectangle3_ys[2049]), .RECT3_WIDTH(rectangle3_widths[2049]), .RECT3_HEIGHT(rectangle3_heights[2049]), .RECT3_WEIGHT(rectangle3_weights[2049]), .FEAT_THRES(feature_thresholds[2049]), .FEAT_ABOVE(feature_aboves[2049]), .FEAT_BELOW(feature_belows[2049])) ac2049(.scan_win(scan_win2049), .scan_win_std_dev(scan_win_std_dev[2049]), .feature_accum(feature_accums[2049]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2050]), .RECT1_Y(rectangle1_ys[2050]), .RECT1_WIDTH(rectangle1_widths[2050]), .RECT1_HEIGHT(rectangle1_heights[2050]), .RECT1_WEIGHT(rectangle1_weights[2050]), .RECT2_X(rectangle2_xs[2050]), .RECT2_Y(rectangle2_ys[2050]), .RECT2_WIDTH(rectangle2_widths[2050]), .RECT2_HEIGHT(rectangle2_heights[2050]), .RECT2_WEIGHT(rectangle2_weights[2050]), .RECT3_X(rectangle3_xs[2050]), .RECT3_Y(rectangle3_ys[2050]), .RECT3_WIDTH(rectangle3_widths[2050]), .RECT3_HEIGHT(rectangle3_heights[2050]), .RECT3_WEIGHT(rectangle3_weights[2050]), .FEAT_THRES(feature_thresholds[2050]), .FEAT_ABOVE(feature_aboves[2050]), .FEAT_BELOW(feature_belows[2050])) ac2050(.scan_win(scan_win2050), .scan_win_std_dev(scan_win_std_dev[2050]), .feature_accum(feature_accums[2050]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2051]), .RECT1_Y(rectangle1_ys[2051]), .RECT1_WIDTH(rectangle1_widths[2051]), .RECT1_HEIGHT(rectangle1_heights[2051]), .RECT1_WEIGHT(rectangle1_weights[2051]), .RECT2_X(rectangle2_xs[2051]), .RECT2_Y(rectangle2_ys[2051]), .RECT2_WIDTH(rectangle2_widths[2051]), .RECT2_HEIGHT(rectangle2_heights[2051]), .RECT2_WEIGHT(rectangle2_weights[2051]), .RECT3_X(rectangle3_xs[2051]), .RECT3_Y(rectangle3_ys[2051]), .RECT3_WIDTH(rectangle3_widths[2051]), .RECT3_HEIGHT(rectangle3_heights[2051]), .RECT3_WEIGHT(rectangle3_weights[2051]), .FEAT_THRES(feature_thresholds[2051]), .FEAT_ABOVE(feature_aboves[2051]), .FEAT_BELOW(feature_belows[2051])) ac2051(.scan_win(scan_win2051), .scan_win_std_dev(scan_win_std_dev[2051]), .feature_accum(feature_accums[2051]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2052]), .RECT1_Y(rectangle1_ys[2052]), .RECT1_WIDTH(rectangle1_widths[2052]), .RECT1_HEIGHT(rectangle1_heights[2052]), .RECT1_WEIGHT(rectangle1_weights[2052]), .RECT2_X(rectangle2_xs[2052]), .RECT2_Y(rectangle2_ys[2052]), .RECT2_WIDTH(rectangle2_widths[2052]), .RECT2_HEIGHT(rectangle2_heights[2052]), .RECT2_WEIGHT(rectangle2_weights[2052]), .RECT3_X(rectangle3_xs[2052]), .RECT3_Y(rectangle3_ys[2052]), .RECT3_WIDTH(rectangle3_widths[2052]), .RECT3_HEIGHT(rectangle3_heights[2052]), .RECT3_WEIGHT(rectangle3_weights[2052]), .FEAT_THRES(feature_thresholds[2052]), .FEAT_ABOVE(feature_aboves[2052]), .FEAT_BELOW(feature_belows[2052])) ac2052(.scan_win(scan_win2052), .scan_win_std_dev(scan_win_std_dev[2052]), .feature_accum(feature_accums[2052]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2053]), .RECT1_Y(rectangle1_ys[2053]), .RECT1_WIDTH(rectangle1_widths[2053]), .RECT1_HEIGHT(rectangle1_heights[2053]), .RECT1_WEIGHT(rectangle1_weights[2053]), .RECT2_X(rectangle2_xs[2053]), .RECT2_Y(rectangle2_ys[2053]), .RECT2_WIDTH(rectangle2_widths[2053]), .RECT2_HEIGHT(rectangle2_heights[2053]), .RECT2_WEIGHT(rectangle2_weights[2053]), .RECT3_X(rectangle3_xs[2053]), .RECT3_Y(rectangle3_ys[2053]), .RECT3_WIDTH(rectangle3_widths[2053]), .RECT3_HEIGHT(rectangle3_heights[2053]), .RECT3_WEIGHT(rectangle3_weights[2053]), .FEAT_THRES(feature_thresholds[2053]), .FEAT_ABOVE(feature_aboves[2053]), .FEAT_BELOW(feature_belows[2053])) ac2053(.scan_win(scan_win2053), .scan_win_std_dev(scan_win_std_dev[2053]), .feature_accum(feature_accums[2053]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2054]), .RECT1_Y(rectangle1_ys[2054]), .RECT1_WIDTH(rectangle1_widths[2054]), .RECT1_HEIGHT(rectangle1_heights[2054]), .RECT1_WEIGHT(rectangle1_weights[2054]), .RECT2_X(rectangle2_xs[2054]), .RECT2_Y(rectangle2_ys[2054]), .RECT2_WIDTH(rectangle2_widths[2054]), .RECT2_HEIGHT(rectangle2_heights[2054]), .RECT2_WEIGHT(rectangle2_weights[2054]), .RECT3_X(rectangle3_xs[2054]), .RECT3_Y(rectangle3_ys[2054]), .RECT3_WIDTH(rectangle3_widths[2054]), .RECT3_HEIGHT(rectangle3_heights[2054]), .RECT3_WEIGHT(rectangle3_weights[2054]), .FEAT_THRES(feature_thresholds[2054]), .FEAT_ABOVE(feature_aboves[2054]), .FEAT_BELOW(feature_belows[2054])) ac2054(.scan_win(scan_win2054), .scan_win_std_dev(scan_win_std_dev[2054]), .feature_accum(feature_accums[2054]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2055]), .RECT1_Y(rectangle1_ys[2055]), .RECT1_WIDTH(rectangle1_widths[2055]), .RECT1_HEIGHT(rectangle1_heights[2055]), .RECT1_WEIGHT(rectangle1_weights[2055]), .RECT2_X(rectangle2_xs[2055]), .RECT2_Y(rectangle2_ys[2055]), .RECT2_WIDTH(rectangle2_widths[2055]), .RECT2_HEIGHT(rectangle2_heights[2055]), .RECT2_WEIGHT(rectangle2_weights[2055]), .RECT3_X(rectangle3_xs[2055]), .RECT3_Y(rectangle3_ys[2055]), .RECT3_WIDTH(rectangle3_widths[2055]), .RECT3_HEIGHT(rectangle3_heights[2055]), .RECT3_WEIGHT(rectangle3_weights[2055]), .FEAT_THRES(feature_thresholds[2055]), .FEAT_ABOVE(feature_aboves[2055]), .FEAT_BELOW(feature_belows[2055])) ac2055(.scan_win(scan_win2055), .scan_win_std_dev(scan_win_std_dev[2055]), .feature_accum(feature_accums[2055]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2056]), .RECT1_Y(rectangle1_ys[2056]), .RECT1_WIDTH(rectangle1_widths[2056]), .RECT1_HEIGHT(rectangle1_heights[2056]), .RECT1_WEIGHT(rectangle1_weights[2056]), .RECT2_X(rectangle2_xs[2056]), .RECT2_Y(rectangle2_ys[2056]), .RECT2_WIDTH(rectangle2_widths[2056]), .RECT2_HEIGHT(rectangle2_heights[2056]), .RECT2_WEIGHT(rectangle2_weights[2056]), .RECT3_X(rectangle3_xs[2056]), .RECT3_Y(rectangle3_ys[2056]), .RECT3_WIDTH(rectangle3_widths[2056]), .RECT3_HEIGHT(rectangle3_heights[2056]), .RECT3_WEIGHT(rectangle3_weights[2056]), .FEAT_THRES(feature_thresholds[2056]), .FEAT_ABOVE(feature_aboves[2056]), .FEAT_BELOW(feature_belows[2056])) ac2056(.scan_win(scan_win2056), .scan_win_std_dev(scan_win_std_dev[2056]), .feature_accum(feature_accums[2056]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2057]), .RECT1_Y(rectangle1_ys[2057]), .RECT1_WIDTH(rectangle1_widths[2057]), .RECT1_HEIGHT(rectangle1_heights[2057]), .RECT1_WEIGHT(rectangle1_weights[2057]), .RECT2_X(rectangle2_xs[2057]), .RECT2_Y(rectangle2_ys[2057]), .RECT2_WIDTH(rectangle2_widths[2057]), .RECT2_HEIGHT(rectangle2_heights[2057]), .RECT2_WEIGHT(rectangle2_weights[2057]), .RECT3_X(rectangle3_xs[2057]), .RECT3_Y(rectangle3_ys[2057]), .RECT3_WIDTH(rectangle3_widths[2057]), .RECT3_HEIGHT(rectangle3_heights[2057]), .RECT3_WEIGHT(rectangle3_weights[2057]), .FEAT_THRES(feature_thresholds[2057]), .FEAT_ABOVE(feature_aboves[2057]), .FEAT_BELOW(feature_belows[2057])) ac2057(.scan_win(scan_win2057), .scan_win_std_dev(scan_win_std_dev[2057]), .feature_accum(feature_accums[2057]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2058]), .RECT1_Y(rectangle1_ys[2058]), .RECT1_WIDTH(rectangle1_widths[2058]), .RECT1_HEIGHT(rectangle1_heights[2058]), .RECT1_WEIGHT(rectangle1_weights[2058]), .RECT2_X(rectangle2_xs[2058]), .RECT2_Y(rectangle2_ys[2058]), .RECT2_WIDTH(rectangle2_widths[2058]), .RECT2_HEIGHT(rectangle2_heights[2058]), .RECT2_WEIGHT(rectangle2_weights[2058]), .RECT3_X(rectangle3_xs[2058]), .RECT3_Y(rectangle3_ys[2058]), .RECT3_WIDTH(rectangle3_widths[2058]), .RECT3_HEIGHT(rectangle3_heights[2058]), .RECT3_WEIGHT(rectangle3_weights[2058]), .FEAT_THRES(feature_thresholds[2058]), .FEAT_ABOVE(feature_aboves[2058]), .FEAT_BELOW(feature_belows[2058])) ac2058(.scan_win(scan_win2058), .scan_win_std_dev(scan_win_std_dev[2058]), .feature_accum(feature_accums[2058]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2059]), .RECT1_Y(rectangle1_ys[2059]), .RECT1_WIDTH(rectangle1_widths[2059]), .RECT1_HEIGHT(rectangle1_heights[2059]), .RECT1_WEIGHT(rectangle1_weights[2059]), .RECT2_X(rectangle2_xs[2059]), .RECT2_Y(rectangle2_ys[2059]), .RECT2_WIDTH(rectangle2_widths[2059]), .RECT2_HEIGHT(rectangle2_heights[2059]), .RECT2_WEIGHT(rectangle2_weights[2059]), .RECT3_X(rectangle3_xs[2059]), .RECT3_Y(rectangle3_ys[2059]), .RECT3_WIDTH(rectangle3_widths[2059]), .RECT3_HEIGHT(rectangle3_heights[2059]), .RECT3_WEIGHT(rectangle3_weights[2059]), .FEAT_THRES(feature_thresholds[2059]), .FEAT_ABOVE(feature_aboves[2059]), .FEAT_BELOW(feature_belows[2059])) ac2059(.scan_win(scan_win2059), .scan_win_std_dev(scan_win_std_dev[2059]), .feature_accum(feature_accums[2059]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2060]), .RECT1_Y(rectangle1_ys[2060]), .RECT1_WIDTH(rectangle1_widths[2060]), .RECT1_HEIGHT(rectangle1_heights[2060]), .RECT1_WEIGHT(rectangle1_weights[2060]), .RECT2_X(rectangle2_xs[2060]), .RECT2_Y(rectangle2_ys[2060]), .RECT2_WIDTH(rectangle2_widths[2060]), .RECT2_HEIGHT(rectangle2_heights[2060]), .RECT2_WEIGHT(rectangle2_weights[2060]), .RECT3_X(rectangle3_xs[2060]), .RECT3_Y(rectangle3_ys[2060]), .RECT3_WIDTH(rectangle3_widths[2060]), .RECT3_HEIGHT(rectangle3_heights[2060]), .RECT3_WEIGHT(rectangle3_weights[2060]), .FEAT_THRES(feature_thresholds[2060]), .FEAT_ABOVE(feature_aboves[2060]), .FEAT_BELOW(feature_belows[2060])) ac2060(.scan_win(scan_win2060), .scan_win_std_dev(scan_win_std_dev[2060]), .feature_accum(feature_accums[2060]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2061]), .RECT1_Y(rectangle1_ys[2061]), .RECT1_WIDTH(rectangle1_widths[2061]), .RECT1_HEIGHT(rectangle1_heights[2061]), .RECT1_WEIGHT(rectangle1_weights[2061]), .RECT2_X(rectangle2_xs[2061]), .RECT2_Y(rectangle2_ys[2061]), .RECT2_WIDTH(rectangle2_widths[2061]), .RECT2_HEIGHT(rectangle2_heights[2061]), .RECT2_WEIGHT(rectangle2_weights[2061]), .RECT3_X(rectangle3_xs[2061]), .RECT3_Y(rectangle3_ys[2061]), .RECT3_WIDTH(rectangle3_widths[2061]), .RECT3_HEIGHT(rectangle3_heights[2061]), .RECT3_WEIGHT(rectangle3_weights[2061]), .FEAT_THRES(feature_thresholds[2061]), .FEAT_ABOVE(feature_aboves[2061]), .FEAT_BELOW(feature_belows[2061])) ac2061(.scan_win(scan_win2061), .scan_win_std_dev(scan_win_std_dev[2061]), .feature_accum(feature_accums[2061]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2062]), .RECT1_Y(rectangle1_ys[2062]), .RECT1_WIDTH(rectangle1_widths[2062]), .RECT1_HEIGHT(rectangle1_heights[2062]), .RECT1_WEIGHT(rectangle1_weights[2062]), .RECT2_X(rectangle2_xs[2062]), .RECT2_Y(rectangle2_ys[2062]), .RECT2_WIDTH(rectangle2_widths[2062]), .RECT2_HEIGHT(rectangle2_heights[2062]), .RECT2_WEIGHT(rectangle2_weights[2062]), .RECT3_X(rectangle3_xs[2062]), .RECT3_Y(rectangle3_ys[2062]), .RECT3_WIDTH(rectangle3_widths[2062]), .RECT3_HEIGHT(rectangle3_heights[2062]), .RECT3_WEIGHT(rectangle3_weights[2062]), .FEAT_THRES(feature_thresholds[2062]), .FEAT_ABOVE(feature_aboves[2062]), .FEAT_BELOW(feature_belows[2062])) ac2062(.scan_win(scan_win2062), .scan_win_std_dev(scan_win_std_dev[2062]), .feature_accum(feature_accums[2062]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2063]), .RECT1_Y(rectangle1_ys[2063]), .RECT1_WIDTH(rectangle1_widths[2063]), .RECT1_HEIGHT(rectangle1_heights[2063]), .RECT1_WEIGHT(rectangle1_weights[2063]), .RECT2_X(rectangle2_xs[2063]), .RECT2_Y(rectangle2_ys[2063]), .RECT2_WIDTH(rectangle2_widths[2063]), .RECT2_HEIGHT(rectangle2_heights[2063]), .RECT2_WEIGHT(rectangle2_weights[2063]), .RECT3_X(rectangle3_xs[2063]), .RECT3_Y(rectangle3_ys[2063]), .RECT3_WIDTH(rectangle3_widths[2063]), .RECT3_HEIGHT(rectangle3_heights[2063]), .RECT3_WEIGHT(rectangle3_weights[2063]), .FEAT_THRES(feature_thresholds[2063]), .FEAT_ABOVE(feature_aboves[2063]), .FEAT_BELOW(feature_belows[2063])) ac2063(.scan_win(scan_win2063), .scan_win_std_dev(scan_win_std_dev[2063]), .feature_accum(feature_accums[2063]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2064]), .RECT1_Y(rectangle1_ys[2064]), .RECT1_WIDTH(rectangle1_widths[2064]), .RECT1_HEIGHT(rectangle1_heights[2064]), .RECT1_WEIGHT(rectangle1_weights[2064]), .RECT2_X(rectangle2_xs[2064]), .RECT2_Y(rectangle2_ys[2064]), .RECT2_WIDTH(rectangle2_widths[2064]), .RECT2_HEIGHT(rectangle2_heights[2064]), .RECT2_WEIGHT(rectangle2_weights[2064]), .RECT3_X(rectangle3_xs[2064]), .RECT3_Y(rectangle3_ys[2064]), .RECT3_WIDTH(rectangle3_widths[2064]), .RECT3_HEIGHT(rectangle3_heights[2064]), .RECT3_WEIGHT(rectangle3_weights[2064]), .FEAT_THRES(feature_thresholds[2064]), .FEAT_ABOVE(feature_aboves[2064]), .FEAT_BELOW(feature_belows[2064])) ac2064(.scan_win(scan_win2064), .scan_win_std_dev(scan_win_std_dev[2064]), .feature_accum(feature_accums[2064]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2065]), .RECT1_Y(rectangle1_ys[2065]), .RECT1_WIDTH(rectangle1_widths[2065]), .RECT1_HEIGHT(rectangle1_heights[2065]), .RECT1_WEIGHT(rectangle1_weights[2065]), .RECT2_X(rectangle2_xs[2065]), .RECT2_Y(rectangle2_ys[2065]), .RECT2_WIDTH(rectangle2_widths[2065]), .RECT2_HEIGHT(rectangle2_heights[2065]), .RECT2_WEIGHT(rectangle2_weights[2065]), .RECT3_X(rectangle3_xs[2065]), .RECT3_Y(rectangle3_ys[2065]), .RECT3_WIDTH(rectangle3_widths[2065]), .RECT3_HEIGHT(rectangle3_heights[2065]), .RECT3_WEIGHT(rectangle3_weights[2065]), .FEAT_THRES(feature_thresholds[2065]), .FEAT_ABOVE(feature_aboves[2065]), .FEAT_BELOW(feature_belows[2065])) ac2065(.scan_win(scan_win2065), .scan_win_std_dev(scan_win_std_dev[2065]), .feature_accum(feature_accums[2065]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2066]), .RECT1_Y(rectangle1_ys[2066]), .RECT1_WIDTH(rectangle1_widths[2066]), .RECT1_HEIGHT(rectangle1_heights[2066]), .RECT1_WEIGHT(rectangle1_weights[2066]), .RECT2_X(rectangle2_xs[2066]), .RECT2_Y(rectangle2_ys[2066]), .RECT2_WIDTH(rectangle2_widths[2066]), .RECT2_HEIGHT(rectangle2_heights[2066]), .RECT2_WEIGHT(rectangle2_weights[2066]), .RECT3_X(rectangle3_xs[2066]), .RECT3_Y(rectangle3_ys[2066]), .RECT3_WIDTH(rectangle3_widths[2066]), .RECT3_HEIGHT(rectangle3_heights[2066]), .RECT3_WEIGHT(rectangle3_weights[2066]), .FEAT_THRES(feature_thresholds[2066]), .FEAT_ABOVE(feature_aboves[2066]), .FEAT_BELOW(feature_belows[2066])) ac2066(.scan_win(scan_win2066), .scan_win_std_dev(scan_win_std_dev[2066]), .feature_accum(feature_accums[2066]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2067]), .RECT1_Y(rectangle1_ys[2067]), .RECT1_WIDTH(rectangle1_widths[2067]), .RECT1_HEIGHT(rectangle1_heights[2067]), .RECT1_WEIGHT(rectangle1_weights[2067]), .RECT2_X(rectangle2_xs[2067]), .RECT2_Y(rectangle2_ys[2067]), .RECT2_WIDTH(rectangle2_widths[2067]), .RECT2_HEIGHT(rectangle2_heights[2067]), .RECT2_WEIGHT(rectangle2_weights[2067]), .RECT3_X(rectangle3_xs[2067]), .RECT3_Y(rectangle3_ys[2067]), .RECT3_WIDTH(rectangle3_widths[2067]), .RECT3_HEIGHT(rectangle3_heights[2067]), .RECT3_WEIGHT(rectangle3_weights[2067]), .FEAT_THRES(feature_thresholds[2067]), .FEAT_ABOVE(feature_aboves[2067]), .FEAT_BELOW(feature_belows[2067])) ac2067(.scan_win(scan_win2067), .scan_win_std_dev(scan_win_std_dev[2067]), .feature_accum(feature_accums[2067]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2068]), .RECT1_Y(rectangle1_ys[2068]), .RECT1_WIDTH(rectangle1_widths[2068]), .RECT1_HEIGHT(rectangle1_heights[2068]), .RECT1_WEIGHT(rectangle1_weights[2068]), .RECT2_X(rectangle2_xs[2068]), .RECT2_Y(rectangle2_ys[2068]), .RECT2_WIDTH(rectangle2_widths[2068]), .RECT2_HEIGHT(rectangle2_heights[2068]), .RECT2_WEIGHT(rectangle2_weights[2068]), .RECT3_X(rectangle3_xs[2068]), .RECT3_Y(rectangle3_ys[2068]), .RECT3_WIDTH(rectangle3_widths[2068]), .RECT3_HEIGHT(rectangle3_heights[2068]), .RECT3_WEIGHT(rectangle3_weights[2068]), .FEAT_THRES(feature_thresholds[2068]), .FEAT_ABOVE(feature_aboves[2068]), .FEAT_BELOW(feature_belows[2068])) ac2068(.scan_win(scan_win2068), .scan_win_std_dev(scan_win_std_dev[2068]), .feature_accum(feature_accums[2068]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2069]), .RECT1_Y(rectangle1_ys[2069]), .RECT1_WIDTH(rectangle1_widths[2069]), .RECT1_HEIGHT(rectangle1_heights[2069]), .RECT1_WEIGHT(rectangle1_weights[2069]), .RECT2_X(rectangle2_xs[2069]), .RECT2_Y(rectangle2_ys[2069]), .RECT2_WIDTH(rectangle2_widths[2069]), .RECT2_HEIGHT(rectangle2_heights[2069]), .RECT2_WEIGHT(rectangle2_weights[2069]), .RECT3_X(rectangle3_xs[2069]), .RECT3_Y(rectangle3_ys[2069]), .RECT3_WIDTH(rectangle3_widths[2069]), .RECT3_HEIGHT(rectangle3_heights[2069]), .RECT3_WEIGHT(rectangle3_weights[2069]), .FEAT_THRES(feature_thresholds[2069]), .FEAT_ABOVE(feature_aboves[2069]), .FEAT_BELOW(feature_belows[2069])) ac2069(.scan_win(scan_win2069), .scan_win_std_dev(scan_win_std_dev[2069]), .feature_accum(feature_accums[2069]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2070]), .RECT1_Y(rectangle1_ys[2070]), .RECT1_WIDTH(rectangle1_widths[2070]), .RECT1_HEIGHT(rectangle1_heights[2070]), .RECT1_WEIGHT(rectangle1_weights[2070]), .RECT2_X(rectangle2_xs[2070]), .RECT2_Y(rectangle2_ys[2070]), .RECT2_WIDTH(rectangle2_widths[2070]), .RECT2_HEIGHT(rectangle2_heights[2070]), .RECT2_WEIGHT(rectangle2_weights[2070]), .RECT3_X(rectangle3_xs[2070]), .RECT3_Y(rectangle3_ys[2070]), .RECT3_WIDTH(rectangle3_widths[2070]), .RECT3_HEIGHT(rectangle3_heights[2070]), .RECT3_WEIGHT(rectangle3_weights[2070]), .FEAT_THRES(feature_thresholds[2070]), .FEAT_ABOVE(feature_aboves[2070]), .FEAT_BELOW(feature_belows[2070])) ac2070(.scan_win(scan_win2070), .scan_win_std_dev(scan_win_std_dev[2070]), .feature_accum(feature_accums[2070]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2071]), .RECT1_Y(rectangle1_ys[2071]), .RECT1_WIDTH(rectangle1_widths[2071]), .RECT1_HEIGHT(rectangle1_heights[2071]), .RECT1_WEIGHT(rectangle1_weights[2071]), .RECT2_X(rectangle2_xs[2071]), .RECT2_Y(rectangle2_ys[2071]), .RECT2_WIDTH(rectangle2_widths[2071]), .RECT2_HEIGHT(rectangle2_heights[2071]), .RECT2_WEIGHT(rectangle2_weights[2071]), .RECT3_X(rectangle3_xs[2071]), .RECT3_Y(rectangle3_ys[2071]), .RECT3_WIDTH(rectangle3_widths[2071]), .RECT3_HEIGHT(rectangle3_heights[2071]), .RECT3_WEIGHT(rectangle3_weights[2071]), .FEAT_THRES(feature_thresholds[2071]), .FEAT_ABOVE(feature_aboves[2071]), .FEAT_BELOW(feature_belows[2071])) ac2071(.scan_win(scan_win2071), .scan_win_std_dev(scan_win_std_dev[2071]), .feature_accum(feature_accums[2071]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2072]), .RECT1_Y(rectangle1_ys[2072]), .RECT1_WIDTH(rectangle1_widths[2072]), .RECT1_HEIGHT(rectangle1_heights[2072]), .RECT1_WEIGHT(rectangle1_weights[2072]), .RECT2_X(rectangle2_xs[2072]), .RECT2_Y(rectangle2_ys[2072]), .RECT2_WIDTH(rectangle2_widths[2072]), .RECT2_HEIGHT(rectangle2_heights[2072]), .RECT2_WEIGHT(rectangle2_weights[2072]), .RECT3_X(rectangle3_xs[2072]), .RECT3_Y(rectangle3_ys[2072]), .RECT3_WIDTH(rectangle3_widths[2072]), .RECT3_HEIGHT(rectangle3_heights[2072]), .RECT3_WEIGHT(rectangle3_weights[2072]), .FEAT_THRES(feature_thresholds[2072]), .FEAT_ABOVE(feature_aboves[2072]), .FEAT_BELOW(feature_belows[2072])) ac2072(.scan_win(scan_win2072), .scan_win_std_dev(scan_win_std_dev[2072]), .feature_accum(feature_accums[2072]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2073]), .RECT1_Y(rectangle1_ys[2073]), .RECT1_WIDTH(rectangle1_widths[2073]), .RECT1_HEIGHT(rectangle1_heights[2073]), .RECT1_WEIGHT(rectangle1_weights[2073]), .RECT2_X(rectangle2_xs[2073]), .RECT2_Y(rectangle2_ys[2073]), .RECT2_WIDTH(rectangle2_widths[2073]), .RECT2_HEIGHT(rectangle2_heights[2073]), .RECT2_WEIGHT(rectangle2_weights[2073]), .RECT3_X(rectangle3_xs[2073]), .RECT3_Y(rectangle3_ys[2073]), .RECT3_WIDTH(rectangle3_widths[2073]), .RECT3_HEIGHT(rectangle3_heights[2073]), .RECT3_WEIGHT(rectangle3_weights[2073]), .FEAT_THRES(feature_thresholds[2073]), .FEAT_ABOVE(feature_aboves[2073]), .FEAT_BELOW(feature_belows[2073])) ac2073(.scan_win(scan_win2073), .scan_win_std_dev(scan_win_std_dev[2073]), .feature_accum(feature_accums[2073]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2074]), .RECT1_Y(rectangle1_ys[2074]), .RECT1_WIDTH(rectangle1_widths[2074]), .RECT1_HEIGHT(rectangle1_heights[2074]), .RECT1_WEIGHT(rectangle1_weights[2074]), .RECT2_X(rectangle2_xs[2074]), .RECT2_Y(rectangle2_ys[2074]), .RECT2_WIDTH(rectangle2_widths[2074]), .RECT2_HEIGHT(rectangle2_heights[2074]), .RECT2_WEIGHT(rectangle2_weights[2074]), .RECT3_X(rectangle3_xs[2074]), .RECT3_Y(rectangle3_ys[2074]), .RECT3_WIDTH(rectangle3_widths[2074]), .RECT3_HEIGHT(rectangle3_heights[2074]), .RECT3_WEIGHT(rectangle3_weights[2074]), .FEAT_THRES(feature_thresholds[2074]), .FEAT_ABOVE(feature_aboves[2074]), .FEAT_BELOW(feature_belows[2074])) ac2074(.scan_win(scan_win2074), .scan_win_std_dev(scan_win_std_dev[2074]), .feature_accum(feature_accums[2074]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2075]), .RECT1_Y(rectangle1_ys[2075]), .RECT1_WIDTH(rectangle1_widths[2075]), .RECT1_HEIGHT(rectangle1_heights[2075]), .RECT1_WEIGHT(rectangle1_weights[2075]), .RECT2_X(rectangle2_xs[2075]), .RECT2_Y(rectangle2_ys[2075]), .RECT2_WIDTH(rectangle2_widths[2075]), .RECT2_HEIGHT(rectangle2_heights[2075]), .RECT2_WEIGHT(rectangle2_weights[2075]), .RECT3_X(rectangle3_xs[2075]), .RECT3_Y(rectangle3_ys[2075]), .RECT3_WIDTH(rectangle3_widths[2075]), .RECT3_HEIGHT(rectangle3_heights[2075]), .RECT3_WEIGHT(rectangle3_weights[2075]), .FEAT_THRES(feature_thresholds[2075]), .FEAT_ABOVE(feature_aboves[2075]), .FEAT_BELOW(feature_belows[2075])) ac2075(.scan_win(scan_win2075), .scan_win_std_dev(scan_win_std_dev[2075]), .feature_accum(feature_accums[2075]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2076]), .RECT1_Y(rectangle1_ys[2076]), .RECT1_WIDTH(rectangle1_widths[2076]), .RECT1_HEIGHT(rectangle1_heights[2076]), .RECT1_WEIGHT(rectangle1_weights[2076]), .RECT2_X(rectangle2_xs[2076]), .RECT2_Y(rectangle2_ys[2076]), .RECT2_WIDTH(rectangle2_widths[2076]), .RECT2_HEIGHT(rectangle2_heights[2076]), .RECT2_WEIGHT(rectangle2_weights[2076]), .RECT3_X(rectangle3_xs[2076]), .RECT3_Y(rectangle3_ys[2076]), .RECT3_WIDTH(rectangle3_widths[2076]), .RECT3_HEIGHT(rectangle3_heights[2076]), .RECT3_WEIGHT(rectangle3_weights[2076]), .FEAT_THRES(feature_thresholds[2076]), .FEAT_ABOVE(feature_aboves[2076]), .FEAT_BELOW(feature_belows[2076])) ac2076(.scan_win(scan_win2076), .scan_win_std_dev(scan_win_std_dev[2076]), .feature_accum(feature_accums[2076]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2077]), .RECT1_Y(rectangle1_ys[2077]), .RECT1_WIDTH(rectangle1_widths[2077]), .RECT1_HEIGHT(rectangle1_heights[2077]), .RECT1_WEIGHT(rectangle1_weights[2077]), .RECT2_X(rectangle2_xs[2077]), .RECT2_Y(rectangle2_ys[2077]), .RECT2_WIDTH(rectangle2_widths[2077]), .RECT2_HEIGHT(rectangle2_heights[2077]), .RECT2_WEIGHT(rectangle2_weights[2077]), .RECT3_X(rectangle3_xs[2077]), .RECT3_Y(rectangle3_ys[2077]), .RECT3_WIDTH(rectangle3_widths[2077]), .RECT3_HEIGHT(rectangle3_heights[2077]), .RECT3_WEIGHT(rectangle3_weights[2077]), .FEAT_THRES(feature_thresholds[2077]), .FEAT_ABOVE(feature_aboves[2077]), .FEAT_BELOW(feature_belows[2077])) ac2077(.scan_win(scan_win2077), .scan_win_std_dev(scan_win_std_dev[2077]), .feature_accum(feature_accums[2077]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2078]), .RECT1_Y(rectangle1_ys[2078]), .RECT1_WIDTH(rectangle1_widths[2078]), .RECT1_HEIGHT(rectangle1_heights[2078]), .RECT1_WEIGHT(rectangle1_weights[2078]), .RECT2_X(rectangle2_xs[2078]), .RECT2_Y(rectangle2_ys[2078]), .RECT2_WIDTH(rectangle2_widths[2078]), .RECT2_HEIGHT(rectangle2_heights[2078]), .RECT2_WEIGHT(rectangle2_weights[2078]), .RECT3_X(rectangle3_xs[2078]), .RECT3_Y(rectangle3_ys[2078]), .RECT3_WIDTH(rectangle3_widths[2078]), .RECT3_HEIGHT(rectangle3_heights[2078]), .RECT3_WEIGHT(rectangle3_weights[2078]), .FEAT_THRES(feature_thresholds[2078]), .FEAT_ABOVE(feature_aboves[2078]), .FEAT_BELOW(feature_belows[2078])) ac2078(.scan_win(scan_win2078), .scan_win_std_dev(scan_win_std_dev[2078]), .feature_accum(feature_accums[2078]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2079]), .RECT1_Y(rectangle1_ys[2079]), .RECT1_WIDTH(rectangle1_widths[2079]), .RECT1_HEIGHT(rectangle1_heights[2079]), .RECT1_WEIGHT(rectangle1_weights[2079]), .RECT2_X(rectangle2_xs[2079]), .RECT2_Y(rectangle2_ys[2079]), .RECT2_WIDTH(rectangle2_widths[2079]), .RECT2_HEIGHT(rectangle2_heights[2079]), .RECT2_WEIGHT(rectangle2_weights[2079]), .RECT3_X(rectangle3_xs[2079]), .RECT3_Y(rectangle3_ys[2079]), .RECT3_WIDTH(rectangle3_widths[2079]), .RECT3_HEIGHT(rectangle3_heights[2079]), .RECT3_WEIGHT(rectangle3_weights[2079]), .FEAT_THRES(feature_thresholds[2079]), .FEAT_ABOVE(feature_aboves[2079]), .FEAT_BELOW(feature_belows[2079])) ac2079(.scan_win(scan_win2079), .scan_win_std_dev(scan_win_std_dev[2079]), .feature_accum(feature_accums[2079]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2080]), .RECT1_Y(rectangle1_ys[2080]), .RECT1_WIDTH(rectangle1_widths[2080]), .RECT1_HEIGHT(rectangle1_heights[2080]), .RECT1_WEIGHT(rectangle1_weights[2080]), .RECT2_X(rectangle2_xs[2080]), .RECT2_Y(rectangle2_ys[2080]), .RECT2_WIDTH(rectangle2_widths[2080]), .RECT2_HEIGHT(rectangle2_heights[2080]), .RECT2_WEIGHT(rectangle2_weights[2080]), .RECT3_X(rectangle3_xs[2080]), .RECT3_Y(rectangle3_ys[2080]), .RECT3_WIDTH(rectangle3_widths[2080]), .RECT3_HEIGHT(rectangle3_heights[2080]), .RECT3_WEIGHT(rectangle3_weights[2080]), .FEAT_THRES(feature_thresholds[2080]), .FEAT_ABOVE(feature_aboves[2080]), .FEAT_BELOW(feature_belows[2080])) ac2080(.scan_win(scan_win2080), .scan_win_std_dev(scan_win_std_dev[2080]), .feature_accum(feature_accums[2080]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2081]), .RECT1_Y(rectangle1_ys[2081]), .RECT1_WIDTH(rectangle1_widths[2081]), .RECT1_HEIGHT(rectangle1_heights[2081]), .RECT1_WEIGHT(rectangle1_weights[2081]), .RECT2_X(rectangle2_xs[2081]), .RECT2_Y(rectangle2_ys[2081]), .RECT2_WIDTH(rectangle2_widths[2081]), .RECT2_HEIGHT(rectangle2_heights[2081]), .RECT2_WEIGHT(rectangle2_weights[2081]), .RECT3_X(rectangle3_xs[2081]), .RECT3_Y(rectangle3_ys[2081]), .RECT3_WIDTH(rectangle3_widths[2081]), .RECT3_HEIGHT(rectangle3_heights[2081]), .RECT3_WEIGHT(rectangle3_weights[2081]), .FEAT_THRES(feature_thresholds[2081]), .FEAT_ABOVE(feature_aboves[2081]), .FEAT_BELOW(feature_belows[2081])) ac2081(.scan_win(scan_win2081), .scan_win_std_dev(scan_win_std_dev[2081]), .feature_accum(feature_accums[2081]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2082]), .RECT1_Y(rectangle1_ys[2082]), .RECT1_WIDTH(rectangle1_widths[2082]), .RECT1_HEIGHT(rectangle1_heights[2082]), .RECT1_WEIGHT(rectangle1_weights[2082]), .RECT2_X(rectangle2_xs[2082]), .RECT2_Y(rectangle2_ys[2082]), .RECT2_WIDTH(rectangle2_widths[2082]), .RECT2_HEIGHT(rectangle2_heights[2082]), .RECT2_WEIGHT(rectangle2_weights[2082]), .RECT3_X(rectangle3_xs[2082]), .RECT3_Y(rectangle3_ys[2082]), .RECT3_WIDTH(rectangle3_widths[2082]), .RECT3_HEIGHT(rectangle3_heights[2082]), .RECT3_WEIGHT(rectangle3_weights[2082]), .FEAT_THRES(feature_thresholds[2082]), .FEAT_ABOVE(feature_aboves[2082]), .FEAT_BELOW(feature_belows[2082])) ac2082(.scan_win(scan_win2082), .scan_win_std_dev(scan_win_std_dev[2082]), .feature_accum(feature_accums[2082]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2083]), .RECT1_Y(rectangle1_ys[2083]), .RECT1_WIDTH(rectangle1_widths[2083]), .RECT1_HEIGHT(rectangle1_heights[2083]), .RECT1_WEIGHT(rectangle1_weights[2083]), .RECT2_X(rectangle2_xs[2083]), .RECT2_Y(rectangle2_ys[2083]), .RECT2_WIDTH(rectangle2_widths[2083]), .RECT2_HEIGHT(rectangle2_heights[2083]), .RECT2_WEIGHT(rectangle2_weights[2083]), .RECT3_X(rectangle3_xs[2083]), .RECT3_Y(rectangle3_ys[2083]), .RECT3_WIDTH(rectangle3_widths[2083]), .RECT3_HEIGHT(rectangle3_heights[2083]), .RECT3_WEIGHT(rectangle3_weights[2083]), .FEAT_THRES(feature_thresholds[2083]), .FEAT_ABOVE(feature_aboves[2083]), .FEAT_BELOW(feature_belows[2083])) ac2083(.scan_win(scan_win2083), .scan_win_std_dev(scan_win_std_dev[2083]), .feature_accum(feature_accums[2083]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2084]), .RECT1_Y(rectangle1_ys[2084]), .RECT1_WIDTH(rectangle1_widths[2084]), .RECT1_HEIGHT(rectangle1_heights[2084]), .RECT1_WEIGHT(rectangle1_weights[2084]), .RECT2_X(rectangle2_xs[2084]), .RECT2_Y(rectangle2_ys[2084]), .RECT2_WIDTH(rectangle2_widths[2084]), .RECT2_HEIGHT(rectangle2_heights[2084]), .RECT2_WEIGHT(rectangle2_weights[2084]), .RECT3_X(rectangle3_xs[2084]), .RECT3_Y(rectangle3_ys[2084]), .RECT3_WIDTH(rectangle3_widths[2084]), .RECT3_HEIGHT(rectangle3_heights[2084]), .RECT3_WEIGHT(rectangle3_weights[2084]), .FEAT_THRES(feature_thresholds[2084]), .FEAT_ABOVE(feature_aboves[2084]), .FEAT_BELOW(feature_belows[2084])) ac2084(.scan_win(scan_win2084), .scan_win_std_dev(scan_win_std_dev[2084]), .feature_accum(feature_accums[2084]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2085]), .RECT1_Y(rectangle1_ys[2085]), .RECT1_WIDTH(rectangle1_widths[2085]), .RECT1_HEIGHT(rectangle1_heights[2085]), .RECT1_WEIGHT(rectangle1_weights[2085]), .RECT2_X(rectangle2_xs[2085]), .RECT2_Y(rectangle2_ys[2085]), .RECT2_WIDTH(rectangle2_widths[2085]), .RECT2_HEIGHT(rectangle2_heights[2085]), .RECT2_WEIGHT(rectangle2_weights[2085]), .RECT3_X(rectangle3_xs[2085]), .RECT3_Y(rectangle3_ys[2085]), .RECT3_WIDTH(rectangle3_widths[2085]), .RECT3_HEIGHT(rectangle3_heights[2085]), .RECT3_WEIGHT(rectangle3_weights[2085]), .FEAT_THRES(feature_thresholds[2085]), .FEAT_ABOVE(feature_aboves[2085]), .FEAT_BELOW(feature_belows[2085])) ac2085(.scan_win(scan_win2085), .scan_win_std_dev(scan_win_std_dev[2085]), .feature_accum(feature_accums[2085]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2086]), .RECT1_Y(rectangle1_ys[2086]), .RECT1_WIDTH(rectangle1_widths[2086]), .RECT1_HEIGHT(rectangle1_heights[2086]), .RECT1_WEIGHT(rectangle1_weights[2086]), .RECT2_X(rectangle2_xs[2086]), .RECT2_Y(rectangle2_ys[2086]), .RECT2_WIDTH(rectangle2_widths[2086]), .RECT2_HEIGHT(rectangle2_heights[2086]), .RECT2_WEIGHT(rectangle2_weights[2086]), .RECT3_X(rectangle3_xs[2086]), .RECT3_Y(rectangle3_ys[2086]), .RECT3_WIDTH(rectangle3_widths[2086]), .RECT3_HEIGHT(rectangle3_heights[2086]), .RECT3_WEIGHT(rectangle3_weights[2086]), .FEAT_THRES(feature_thresholds[2086]), .FEAT_ABOVE(feature_aboves[2086]), .FEAT_BELOW(feature_belows[2086])) ac2086(.scan_win(scan_win2086), .scan_win_std_dev(scan_win_std_dev[2086]), .feature_accum(feature_accums[2086]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2087]), .RECT1_Y(rectangle1_ys[2087]), .RECT1_WIDTH(rectangle1_widths[2087]), .RECT1_HEIGHT(rectangle1_heights[2087]), .RECT1_WEIGHT(rectangle1_weights[2087]), .RECT2_X(rectangle2_xs[2087]), .RECT2_Y(rectangle2_ys[2087]), .RECT2_WIDTH(rectangle2_widths[2087]), .RECT2_HEIGHT(rectangle2_heights[2087]), .RECT2_WEIGHT(rectangle2_weights[2087]), .RECT3_X(rectangle3_xs[2087]), .RECT3_Y(rectangle3_ys[2087]), .RECT3_WIDTH(rectangle3_widths[2087]), .RECT3_HEIGHT(rectangle3_heights[2087]), .RECT3_WEIGHT(rectangle3_weights[2087]), .FEAT_THRES(feature_thresholds[2087]), .FEAT_ABOVE(feature_aboves[2087]), .FEAT_BELOW(feature_belows[2087])) ac2087(.scan_win(scan_win2087), .scan_win_std_dev(scan_win_std_dev[2087]), .feature_accum(feature_accums[2087]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2088]), .RECT1_Y(rectangle1_ys[2088]), .RECT1_WIDTH(rectangle1_widths[2088]), .RECT1_HEIGHT(rectangle1_heights[2088]), .RECT1_WEIGHT(rectangle1_weights[2088]), .RECT2_X(rectangle2_xs[2088]), .RECT2_Y(rectangle2_ys[2088]), .RECT2_WIDTH(rectangle2_widths[2088]), .RECT2_HEIGHT(rectangle2_heights[2088]), .RECT2_WEIGHT(rectangle2_weights[2088]), .RECT3_X(rectangle3_xs[2088]), .RECT3_Y(rectangle3_ys[2088]), .RECT3_WIDTH(rectangle3_widths[2088]), .RECT3_HEIGHT(rectangle3_heights[2088]), .RECT3_WEIGHT(rectangle3_weights[2088]), .FEAT_THRES(feature_thresholds[2088]), .FEAT_ABOVE(feature_aboves[2088]), .FEAT_BELOW(feature_belows[2088])) ac2088(.scan_win(scan_win2088), .scan_win_std_dev(scan_win_std_dev[2088]), .feature_accum(feature_accums[2088]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2089]), .RECT1_Y(rectangle1_ys[2089]), .RECT1_WIDTH(rectangle1_widths[2089]), .RECT1_HEIGHT(rectangle1_heights[2089]), .RECT1_WEIGHT(rectangle1_weights[2089]), .RECT2_X(rectangle2_xs[2089]), .RECT2_Y(rectangle2_ys[2089]), .RECT2_WIDTH(rectangle2_widths[2089]), .RECT2_HEIGHT(rectangle2_heights[2089]), .RECT2_WEIGHT(rectangle2_weights[2089]), .RECT3_X(rectangle3_xs[2089]), .RECT3_Y(rectangle3_ys[2089]), .RECT3_WIDTH(rectangle3_widths[2089]), .RECT3_HEIGHT(rectangle3_heights[2089]), .RECT3_WEIGHT(rectangle3_weights[2089]), .FEAT_THRES(feature_thresholds[2089]), .FEAT_ABOVE(feature_aboves[2089]), .FEAT_BELOW(feature_belows[2089])) ac2089(.scan_win(scan_win2089), .scan_win_std_dev(scan_win_std_dev[2089]), .feature_accum(feature_accums[2089]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2090]), .RECT1_Y(rectangle1_ys[2090]), .RECT1_WIDTH(rectangle1_widths[2090]), .RECT1_HEIGHT(rectangle1_heights[2090]), .RECT1_WEIGHT(rectangle1_weights[2090]), .RECT2_X(rectangle2_xs[2090]), .RECT2_Y(rectangle2_ys[2090]), .RECT2_WIDTH(rectangle2_widths[2090]), .RECT2_HEIGHT(rectangle2_heights[2090]), .RECT2_WEIGHT(rectangle2_weights[2090]), .RECT3_X(rectangle3_xs[2090]), .RECT3_Y(rectangle3_ys[2090]), .RECT3_WIDTH(rectangle3_widths[2090]), .RECT3_HEIGHT(rectangle3_heights[2090]), .RECT3_WEIGHT(rectangle3_weights[2090]), .FEAT_THRES(feature_thresholds[2090]), .FEAT_ABOVE(feature_aboves[2090]), .FEAT_BELOW(feature_belows[2090])) ac2090(.scan_win(scan_win2090), .scan_win_std_dev(scan_win_std_dev[2090]), .feature_accum(feature_accums[2090]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2091]), .RECT1_Y(rectangle1_ys[2091]), .RECT1_WIDTH(rectangle1_widths[2091]), .RECT1_HEIGHT(rectangle1_heights[2091]), .RECT1_WEIGHT(rectangle1_weights[2091]), .RECT2_X(rectangle2_xs[2091]), .RECT2_Y(rectangle2_ys[2091]), .RECT2_WIDTH(rectangle2_widths[2091]), .RECT2_HEIGHT(rectangle2_heights[2091]), .RECT2_WEIGHT(rectangle2_weights[2091]), .RECT3_X(rectangle3_xs[2091]), .RECT3_Y(rectangle3_ys[2091]), .RECT3_WIDTH(rectangle3_widths[2091]), .RECT3_HEIGHT(rectangle3_heights[2091]), .RECT3_WEIGHT(rectangle3_weights[2091]), .FEAT_THRES(feature_thresholds[2091]), .FEAT_ABOVE(feature_aboves[2091]), .FEAT_BELOW(feature_belows[2091])) ac2091(.scan_win(scan_win2091), .scan_win_std_dev(scan_win_std_dev[2091]), .feature_accum(feature_accums[2091]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2092]), .RECT1_Y(rectangle1_ys[2092]), .RECT1_WIDTH(rectangle1_widths[2092]), .RECT1_HEIGHT(rectangle1_heights[2092]), .RECT1_WEIGHT(rectangle1_weights[2092]), .RECT2_X(rectangle2_xs[2092]), .RECT2_Y(rectangle2_ys[2092]), .RECT2_WIDTH(rectangle2_widths[2092]), .RECT2_HEIGHT(rectangle2_heights[2092]), .RECT2_WEIGHT(rectangle2_weights[2092]), .RECT3_X(rectangle3_xs[2092]), .RECT3_Y(rectangle3_ys[2092]), .RECT3_WIDTH(rectangle3_widths[2092]), .RECT3_HEIGHT(rectangle3_heights[2092]), .RECT3_WEIGHT(rectangle3_weights[2092]), .FEAT_THRES(feature_thresholds[2092]), .FEAT_ABOVE(feature_aboves[2092]), .FEAT_BELOW(feature_belows[2092])) ac2092(.scan_win(scan_win2092), .scan_win_std_dev(scan_win_std_dev[2092]), .feature_accum(feature_accums[2092]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2093]), .RECT1_Y(rectangle1_ys[2093]), .RECT1_WIDTH(rectangle1_widths[2093]), .RECT1_HEIGHT(rectangle1_heights[2093]), .RECT1_WEIGHT(rectangle1_weights[2093]), .RECT2_X(rectangle2_xs[2093]), .RECT2_Y(rectangle2_ys[2093]), .RECT2_WIDTH(rectangle2_widths[2093]), .RECT2_HEIGHT(rectangle2_heights[2093]), .RECT2_WEIGHT(rectangle2_weights[2093]), .RECT3_X(rectangle3_xs[2093]), .RECT3_Y(rectangle3_ys[2093]), .RECT3_WIDTH(rectangle3_widths[2093]), .RECT3_HEIGHT(rectangle3_heights[2093]), .RECT3_WEIGHT(rectangle3_weights[2093]), .FEAT_THRES(feature_thresholds[2093]), .FEAT_ABOVE(feature_aboves[2093]), .FEAT_BELOW(feature_belows[2093])) ac2093(.scan_win(scan_win2093), .scan_win_std_dev(scan_win_std_dev[2093]), .feature_accum(feature_accums[2093]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2094]), .RECT1_Y(rectangle1_ys[2094]), .RECT1_WIDTH(rectangle1_widths[2094]), .RECT1_HEIGHT(rectangle1_heights[2094]), .RECT1_WEIGHT(rectangle1_weights[2094]), .RECT2_X(rectangle2_xs[2094]), .RECT2_Y(rectangle2_ys[2094]), .RECT2_WIDTH(rectangle2_widths[2094]), .RECT2_HEIGHT(rectangle2_heights[2094]), .RECT2_WEIGHT(rectangle2_weights[2094]), .RECT3_X(rectangle3_xs[2094]), .RECT3_Y(rectangle3_ys[2094]), .RECT3_WIDTH(rectangle3_widths[2094]), .RECT3_HEIGHT(rectangle3_heights[2094]), .RECT3_WEIGHT(rectangle3_weights[2094]), .FEAT_THRES(feature_thresholds[2094]), .FEAT_ABOVE(feature_aboves[2094]), .FEAT_BELOW(feature_belows[2094])) ac2094(.scan_win(scan_win2094), .scan_win_std_dev(scan_win_std_dev[2094]), .feature_accum(feature_accums[2094]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2095]), .RECT1_Y(rectangle1_ys[2095]), .RECT1_WIDTH(rectangle1_widths[2095]), .RECT1_HEIGHT(rectangle1_heights[2095]), .RECT1_WEIGHT(rectangle1_weights[2095]), .RECT2_X(rectangle2_xs[2095]), .RECT2_Y(rectangle2_ys[2095]), .RECT2_WIDTH(rectangle2_widths[2095]), .RECT2_HEIGHT(rectangle2_heights[2095]), .RECT2_WEIGHT(rectangle2_weights[2095]), .RECT3_X(rectangle3_xs[2095]), .RECT3_Y(rectangle3_ys[2095]), .RECT3_WIDTH(rectangle3_widths[2095]), .RECT3_HEIGHT(rectangle3_heights[2095]), .RECT3_WEIGHT(rectangle3_weights[2095]), .FEAT_THRES(feature_thresholds[2095]), .FEAT_ABOVE(feature_aboves[2095]), .FEAT_BELOW(feature_belows[2095])) ac2095(.scan_win(scan_win2095), .scan_win_std_dev(scan_win_std_dev[2095]), .feature_accum(feature_accums[2095]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2096]), .RECT1_Y(rectangle1_ys[2096]), .RECT1_WIDTH(rectangle1_widths[2096]), .RECT1_HEIGHT(rectangle1_heights[2096]), .RECT1_WEIGHT(rectangle1_weights[2096]), .RECT2_X(rectangle2_xs[2096]), .RECT2_Y(rectangle2_ys[2096]), .RECT2_WIDTH(rectangle2_widths[2096]), .RECT2_HEIGHT(rectangle2_heights[2096]), .RECT2_WEIGHT(rectangle2_weights[2096]), .RECT3_X(rectangle3_xs[2096]), .RECT3_Y(rectangle3_ys[2096]), .RECT3_WIDTH(rectangle3_widths[2096]), .RECT3_HEIGHT(rectangle3_heights[2096]), .RECT3_WEIGHT(rectangle3_weights[2096]), .FEAT_THRES(feature_thresholds[2096]), .FEAT_ABOVE(feature_aboves[2096]), .FEAT_BELOW(feature_belows[2096])) ac2096(.scan_win(scan_win2096), .scan_win_std_dev(scan_win_std_dev[2096]), .feature_accum(feature_accums[2096]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2097]), .RECT1_Y(rectangle1_ys[2097]), .RECT1_WIDTH(rectangle1_widths[2097]), .RECT1_HEIGHT(rectangle1_heights[2097]), .RECT1_WEIGHT(rectangle1_weights[2097]), .RECT2_X(rectangle2_xs[2097]), .RECT2_Y(rectangle2_ys[2097]), .RECT2_WIDTH(rectangle2_widths[2097]), .RECT2_HEIGHT(rectangle2_heights[2097]), .RECT2_WEIGHT(rectangle2_weights[2097]), .RECT3_X(rectangle3_xs[2097]), .RECT3_Y(rectangle3_ys[2097]), .RECT3_WIDTH(rectangle3_widths[2097]), .RECT3_HEIGHT(rectangle3_heights[2097]), .RECT3_WEIGHT(rectangle3_weights[2097]), .FEAT_THRES(feature_thresholds[2097]), .FEAT_ABOVE(feature_aboves[2097]), .FEAT_BELOW(feature_belows[2097])) ac2097(.scan_win(scan_win2097), .scan_win_std_dev(scan_win_std_dev[2097]), .feature_accum(feature_accums[2097]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2098]), .RECT1_Y(rectangle1_ys[2098]), .RECT1_WIDTH(rectangle1_widths[2098]), .RECT1_HEIGHT(rectangle1_heights[2098]), .RECT1_WEIGHT(rectangle1_weights[2098]), .RECT2_X(rectangle2_xs[2098]), .RECT2_Y(rectangle2_ys[2098]), .RECT2_WIDTH(rectangle2_widths[2098]), .RECT2_HEIGHT(rectangle2_heights[2098]), .RECT2_WEIGHT(rectangle2_weights[2098]), .RECT3_X(rectangle3_xs[2098]), .RECT3_Y(rectangle3_ys[2098]), .RECT3_WIDTH(rectangle3_widths[2098]), .RECT3_HEIGHT(rectangle3_heights[2098]), .RECT3_WEIGHT(rectangle3_weights[2098]), .FEAT_THRES(feature_thresholds[2098]), .FEAT_ABOVE(feature_aboves[2098]), .FEAT_BELOW(feature_belows[2098])) ac2098(.scan_win(scan_win2098), .scan_win_std_dev(scan_win_std_dev[2098]), .feature_accum(feature_accums[2098]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2099]), .RECT1_Y(rectangle1_ys[2099]), .RECT1_WIDTH(rectangle1_widths[2099]), .RECT1_HEIGHT(rectangle1_heights[2099]), .RECT1_WEIGHT(rectangle1_weights[2099]), .RECT2_X(rectangle2_xs[2099]), .RECT2_Y(rectangle2_ys[2099]), .RECT2_WIDTH(rectangle2_widths[2099]), .RECT2_HEIGHT(rectangle2_heights[2099]), .RECT2_WEIGHT(rectangle2_weights[2099]), .RECT3_X(rectangle3_xs[2099]), .RECT3_Y(rectangle3_ys[2099]), .RECT3_WIDTH(rectangle3_widths[2099]), .RECT3_HEIGHT(rectangle3_heights[2099]), .RECT3_WEIGHT(rectangle3_weights[2099]), .FEAT_THRES(feature_thresholds[2099]), .FEAT_ABOVE(feature_aboves[2099]), .FEAT_BELOW(feature_belows[2099])) ac2099(.scan_win(scan_win2099), .scan_win_std_dev(scan_win_std_dev[2099]), .feature_accum(feature_accums[2099]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2100]), .RECT1_Y(rectangle1_ys[2100]), .RECT1_WIDTH(rectangle1_widths[2100]), .RECT1_HEIGHT(rectangle1_heights[2100]), .RECT1_WEIGHT(rectangle1_weights[2100]), .RECT2_X(rectangle2_xs[2100]), .RECT2_Y(rectangle2_ys[2100]), .RECT2_WIDTH(rectangle2_widths[2100]), .RECT2_HEIGHT(rectangle2_heights[2100]), .RECT2_WEIGHT(rectangle2_weights[2100]), .RECT3_X(rectangle3_xs[2100]), .RECT3_Y(rectangle3_ys[2100]), .RECT3_WIDTH(rectangle3_widths[2100]), .RECT3_HEIGHT(rectangle3_heights[2100]), .RECT3_WEIGHT(rectangle3_weights[2100]), .FEAT_THRES(feature_thresholds[2100]), .FEAT_ABOVE(feature_aboves[2100]), .FEAT_BELOW(feature_belows[2100])) ac2100(.scan_win(scan_win2100), .scan_win_std_dev(scan_win_std_dev[2100]), .feature_accum(feature_accums[2100]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2101]), .RECT1_Y(rectangle1_ys[2101]), .RECT1_WIDTH(rectangle1_widths[2101]), .RECT1_HEIGHT(rectangle1_heights[2101]), .RECT1_WEIGHT(rectangle1_weights[2101]), .RECT2_X(rectangle2_xs[2101]), .RECT2_Y(rectangle2_ys[2101]), .RECT2_WIDTH(rectangle2_widths[2101]), .RECT2_HEIGHT(rectangle2_heights[2101]), .RECT2_WEIGHT(rectangle2_weights[2101]), .RECT3_X(rectangle3_xs[2101]), .RECT3_Y(rectangle3_ys[2101]), .RECT3_WIDTH(rectangle3_widths[2101]), .RECT3_HEIGHT(rectangle3_heights[2101]), .RECT3_WEIGHT(rectangle3_weights[2101]), .FEAT_THRES(feature_thresholds[2101]), .FEAT_ABOVE(feature_aboves[2101]), .FEAT_BELOW(feature_belows[2101])) ac2101(.scan_win(scan_win2101), .scan_win_std_dev(scan_win_std_dev[2101]), .feature_accum(feature_accums[2101]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2102]), .RECT1_Y(rectangle1_ys[2102]), .RECT1_WIDTH(rectangle1_widths[2102]), .RECT1_HEIGHT(rectangle1_heights[2102]), .RECT1_WEIGHT(rectangle1_weights[2102]), .RECT2_X(rectangle2_xs[2102]), .RECT2_Y(rectangle2_ys[2102]), .RECT2_WIDTH(rectangle2_widths[2102]), .RECT2_HEIGHT(rectangle2_heights[2102]), .RECT2_WEIGHT(rectangle2_weights[2102]), .RECT3_X(rectangle3_xs[2102]), .RECT3_Y(rectangle3_ys[2102]), .RECT3_WIDTH(rectangle3_widths[2102]), .RECT3_HEIGHT(rectangle3_heights[2102]), .RECT3_WEIGHT(rectangle3_weights[2102]), .FEAT_THRES(feature_thresholds[2102]), .FEAT_ABOVE(feature_aboves[2102]), .FEAT_BELOW(feature_belows[2102])) ac2102(.scan_win(scan_win2102), .scan_win_std_dev(scan_win_std_dev[2102]), .feature_accum(feature_accums[2102]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2103]), .RECT1_Y(rectangle1_ys[2103]), .RECT1_WIDTH(rectangle1_widths[2103]), .RECT1_HEIGHT(rectangle1_heights[2103]), .RECT1_WEIGHT(rectangle1_weights[2103]), .RECT2_X(rectangle2_xs[2103]), .RECT2_Y(rectangle2_ys[2103]), .RECT2_WIDTH(rectangle2_widths[2103]), .RECT2_HEIGHT(rectangle2_heights[2103]), .RECT2_WEIGHT(rectangle2_weights[2103]), .RECT3_X(rectangle3_xs[2103]), .RECT3_Y(rectangle3_ys[2103]), .RECT3_WIDTH(rectangle3_widths[2103]), .RECT3_HEIGHT(rectangle3_heights[2103]), .RECT3_WEIGHT(rectangle3_weights[2103]), .FEAT_THRES(feature_thresholds[2103]), .FEAT_ABOVE(feature_aboves[2103]), .FEAT_BELOW(feature_belows[2103])) ac2103(.scan_win(scan_win2103), .scan_win_std_dev(scan_win_std_dev[2103]), .feature_accum(feature_accums[2103]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2104]), .RECT1_Y(rectangle1_ys[2104]), .RECT1_WIDTH(rectangle1_widths[2104]), .RECT1_HEIGHT(rectangle1_heights[2104]), .RECT1_WEIGHT(rectangle1_weights[2104]), .RECT2_X(rectangle2_xs[2104]), .RECT2_Y(rectangle2_ys[2104]), .RECT2_WIDTH(rectangle2_widths[2104]), .RECT2_HEIGHT(rectangle2_heights[2104]), .RECT2_WEIGHT(rectangle2_weights[2104]), .RECT3_X(rectangle3_xs[2104]), .RECT3_Y(rectangle3_ys[2104]), .RECT3_WIDTH(rectangle3_widths[2104]), .RECT3_HEIGHT(rectangle3_heights[2104]), .RECT3_WEIGHT(rectangle3_weights[2104]), .FEAT_THRES(feature_thresholds[2104]), .FEAT_ABOVE(feature_aboves[2104]), .FEAT_BELOW(feature_belows[2104])) ac2104(.scan_win(scan_win2104), .scan_win_std_dev(scan_win_std_dev[2104]), .feature_accum(feature_accums[2104]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2105]), .RECT1_Y(rectangle1_ys[2105]), .RECT1_WIDTH(rectangle1_widths[2105]), .RECT1_HEIGHT(rectangle1_heights[2105]), .RECT1_WEIGHT(rectangle1_weights[2105]), .RECT2_X(rectangle2_xs[2105]), .RECT2_Y(rectangle2_ys[2105]), .RECT2_WIDTH(rectangle2_widths[2105]), .RECT2_HEIGHT(rectangle2_heights[2105]), .RECT2_WEIGHT(rectangle2_weights[2105]), .RECT3_X(rectangle3_xs[2105]), .RECT3_Y(rectangle3_ys[2105]), .RECT3_WIDTH(rectangle3_widths[2105]), .RECT3_HEIGHT(rectangle3_heights[2105]), .RECT3_WEIGHT(rectangle3_weights[2105]), .FEAT_THRES(feature_thresholds[2105]), .FEAT_ABOVE(feature_aboves[2105]), .FEAT_BELOW(feature_belows[2105])) ac2105(.scan_win(scan_win2105), .scan_win_std_dev(scan_win_std_dev[2105]), .feature_accum(feature_accums[2105]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2106]), .RECT1_Y(rectangle1_ys[2106]), .RECT1_WIDTH(rectangle1_widths[2106]), .RECT1_HEIGHT(rectangle1_heights[2106]), .RECT1_WEIGHT(rectangle1_weights[2106]), .RECT2_X(rectangle2_xs[2106]), .RECT2_Y(rectangle2_ys[2106]), .RECT2_WIDTH(rectangle2_widths[2106]), .RECT2_HEIGHT(rectangle2_heights[2106]), .RECT2_WEIGHT(rectangle2_weights[2106]), .RECT3_X(rectangle3_xs[2106]), .RECT3_Y(rectangle3_ys[2106]), .RECT3_WIDTH(rectangle3_widths[2106]), .RECT3_HEIGHT(rectangle3_heights[2106]), .RECT3_WEIGHT(rectangle3_weights[2106]), .FEAT_THRES(feature_thresholds[2106]), .FEAT_ABOVE(feature_aboves[2106]), .FEAT_BELOW(feature_belows[2106])) ac2106(.scan_win(scan_win2106), .scan_win_std_dev(scan_win_std_dev[2106]), .feature_accum(feature_accums[2106]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2107]), .RECT1_Y(rectangle1_ys[2107]), .RECT1_WIDTH(rectangle1_widths[2107]), .RECT1_HEIGHT(rectangle1_heights[2107]), .RECT1_WEIGHT(rectangle1_weights[2107]), .RECT2_X(rectangle2_xs[2107]), .RECT2_Y(rectangle2_ys[2107]), .RECT2_WIDTH(rectangle2_widths[2107]), .RECT2_HEIGHT(rectangle2_heights[2107]), .RECT2_WEIGHT(rectangle2_weights[2107]), .RECT3_X(rectangle3_xs[2107]), .RECT3_Y(rectangle3_ys[2107]), .RECT3_WIDTH(rectangle3_widths[2107]), .RECT3_HEIGHT(rectangle3_heights[2107]), .RECT3_WEIGHT(rectangle3_weights[2107]), .FEAT_THRES(feature_thresholds[2107]), .FEAT_ABOVE(feature_aboves[2107]), .FEAT_BELOW(feature_belows[2107])) ac2107(.scan_win(scan_win2107), .scan_win_std_dev(scan_win_std_dev[2107]), .feature_accum(feature_accums[2107]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2108]), .RECT1_Y(rectangle1_ys[2108]), .RECT1_WIDTH(rectangle1_widths[2108]), .RECT1_HEIGHT(rectangle1_heights[2108]), .RECT1_WEIGHT(rectangle1_weights[2108]), .RECT2_X(rectangle2_xs[2108]), .RECT2_Y(rectangle2_ys[2108]), .RECT2_WIDTH(rectangle2_widths[2108]), .RECT2_HEIGHT(rectangle2_heights[2108]), .RECT2_WEIGHT(rectangle2_weights[2108]), .RECT3_X(rectangle3_xs[2108]), .RECT3_Y(rectangle3_ys[2108]), .RECT3_WIDTH(rectangle3_widths[2108]), .RECT3_HEIGHT(rectangle3_heights[2108]), .RECT3_WEIGHT(rectangle3_weights[2108]), .FEAT_THRES(feature_thresholds[2108]), .FEAT_ABOVE(feature_aboves[2108]), .FEAT_BELOW(feature_belows[2108])) ac2108(.scan_win(scan_win2108), .scan_win_std_dev(scan_win_std_dev[2108]), .feature_accum(feature_accums[2108]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2109]), .RECT1_Y(rectangle1_ys[2109]), .RECT1_WIDTH(rectangle1_widths[2109]), .RECT1_HEIGHT(rectangle1_heights[2109]), .RECT1_WEIGHT(rectangle1_weights[2109]), .RECT2_X(rectangle2_xs[2109]), .RECT2_Y(rectangle2_ys[2109]), .RECT2_WIDTH(rectangle2_widths[2109]), .RECT2_HEIGHT(rectangle2_heights[2109]), .RECT2_WEIGHT(rectangle2_weights[2109]), .RECT3_X(rectangle3_xs[2109]), .RECT3_Y(rectangle3_ys[2109]), .RECT3_WIDTH(rectangle3_widths[2109]), .RECT3_HEIGHT(rectangle3_heights[2109]), .RECT3_WEIGHT(rectangle3_weights[2109]), .FEAT_THRES(feature_thresholds[2109]), .FEAT_ABOVE(feature_aboves[2109]), .FEAT_BELOW(feature_belows[2109])) ac2109(.scan_win(scan_win2109), .scan_win_std_dev(scan_win_std_dev[2109]), .feature_accum(feature_accums[2109]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2110]), .RECT1_Y(rectangle1_ys[2110]), .RECT1_WIDTH(rectangle1_widths[2110]), .RECT1_HEIGHT(rectangle1_heights[2110]), .RECT1_WEIGHT(rectangle1_weights[2110]), .RECT2_X(rectangle2_xs[2110]), .RECT2_Y(rectangle2_ys[2110]), .RECT2_WIDTH(rectangle2_widths[2110]), .RECT2_HEIGHT(rectangle2_heights[2110]), .RECT2_WEIGHT(rectangle2_weights[2110]), .RECT3_X(rectangle3_xs[2110]), .RECT3_Y(rectangle3_ys[2110]), .RECT3_WIDTH(rectangle3_widths[2110]), .RECT3_HEIGHT(rectangle3_heights[2110]), .RECT3_WEIGHT(rectangle3_weights[2110]), .FEAT_THRES(feature_thresholds[2110]), .FEAT_ABOVE(feature_aboves[2110]), .FEAT_BELOW(feature_belows[2110])) ac2110(.scan_win(scan_win2110), .scan_win_std_dev(scan_win_std_dev[2110]), .feature_accum(feature_accums[2110]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2111]), .RECT1_Y(rectangle1_ys[2111]), .RECT1_WIDTH(rectangle1_widths[2111]), .RECT1_HEIGHT(rectangle1_heights[2111]), .RECT1_WEIGHT(rectangle1_weights[2111]), .RECT2_X(rectangle2_xs[2111]), .RECT2_Y(rectangle2_ys[2111]), .RECT2_WIDTH(rectangle2_widths[2111]), .RECT2_HEIGHT(rectangle2_heights[2111]), .RECT2_WEIGHT(rectangle2_weights[2111]), .RECT3_X(rectangle3_xs[2111]), .RECT3_Y(rectangle3_ys[2111]), .RECT3_WIDTH(rectangle3_widths[2111]), .RECT3_HEIGHT(rectangle3_heights[2111]), .RECT3_WEIGHT(rectangle3_weights[2111]), .FEAT_THRES(feature_thresholds[2111]), .FEAT_ABOVE(feature_aboves[2111]), .FEAT_BELOW(feature_belows[2111])) ac2111(.scan_win(scan_win2111), .scan_win_std_dev(scan_win_std_dev[2111]), .feature_accum(feature_accums[2111]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2112]), .RECT1_Y(rectangle1_ys[2112]), .RECT1_WIDTH(rectangle1_widths[2112]), .RECT1_HEIGHT(rectangle1_heights[2112]), .RECT1_WEIGHT(rectangle1_weights[2112]), .RECT2_X(rectangle2_xs[2112]), .RECT2_Y(rectangle2_ys[2112]), .RECT2_WIDTH(rectangle2_widths[2112]), .RECT2_HEIGHT(rectangle2_heights[2112]), .RECT2_WEIGHT(rectangle2_weights[2112]), .RECT3_X(rectangle3_xs[2112]), .RECT3_Y(rectangle3_ys[2112]), .RECT3_WIDTH(rectangle3_widths[2112]), .RECT3_HEIGHT(rectangle3_heights[2112]), .RECT3_WEIGHT(rectangle3_weights[2112]), .FEAT_THRES(feature_thresholds[2112]), .FEAT_ABOVE(feature_aboves[2112]), .FEAT_BELOW(feature_belows[2112])) ac2112(.scan_win(scan_win2112), .scan_win_std_dev(scan_win_std_dev[2112]), .feature_accum(feature_accums[2112]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2113]), .RECT1_Y(rectangle1_ys[2113]), .RECT1_WIDTH(rectangle1_widths[2113]), .RECT1_HEIGHT(rectangle1_heights[2113]), .RECT1_WEIGHT(rectangle1_weights[2113]), .RECT2_X(rectangle2_xs[2113]), .RECT2_Y(rectangle2_ys[2113]), .RECT2_WIDTH(rectangle2_widths[2113]), .RECT2_HEIGHT(rectangle2_heights[2113]), .RECT2_WEIGHT(rectangle2_weights[2113]), .RECT3_X(rectangle3_xs[2113]), .RECT3_Y(rectangle3_ys[2113]), .RECT3_WIDTH(rectangle3_widths[2113]), .RECT3_HEIGHT(rectangle3_heights[2113]), .RECT3_WEIGHT(rectangle3_weights[2113]), .FEAT_THRES(feature_thresholds[2113]), .FEAT_ABOVE(feature_aboves[2113]), .FEAT_BELOW(feature_belows[2113])) ac2113(.scan_win(scan_win2113), .scan_win_std_dev(scan_win_std_dev[2113]), .feature_accum(feature_accums[2113]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2114]), .RECT1_Y(rectangle1_ys[2114]), .RECT1_WIDTH(rectangle1_widths[2114]), .RECT1_HEIGHT(rectangle1_heights[2114]), .RECT1_WEIGHT(rectangle1_weights[2114]), .RECT2_X(rectangle2_xs[2114]), .RECT2_Y(rectangle2_ys[2114]), .RECT2_WIDTH(rectangle2_widths[2114]), .RECT2_HEIGHT(rectangle2_heights[2114]), .RECT2_WEIGHT(rectangle2_weights[2114]), .RECT3_X(rectangle3_xs[2114]), .RECT3_Y(rectangle3_ys[2114]), .RECT3_WIDTH(rectangle3_widths[2114]), .RECT3_HEIGHT(rectangle3_heights[2114]), .RECT3_WEIGHT(rectangle3_weights[2114]), .FEAT_THRES(feature_thresholds[2114]), .FEAT_ABOVE(feature_aboves[2114]), .FEAT_BELOW(feature_belows[2114])) ac2114(.scan_win(scan_win2114), .scan_win_std_dev(scan_win_std_dev[2114]), .feature_accum(feature_accums[2114]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2115]), .RECT1_Y(rectangle1_ys[2115]), .RECT1_WIDTH(rectangle1_widths[2115]), .RECT1_HEIGHT(rectangle1_heights[2115]), .RECT1_WEIGHT(rectangle1_weights[2115]), .RECT2_X(rectangle2_xs[2115]), .RECT2_Y(rectangle2_ys[2115]), .RECT2_WIDTH(rectangle2_widths[2115]), .RECT2_HEIGHT(rectangle2_heights[2115]), .RECT2_WEIGHT(rectangle2_weights[2115]), .RECT3_X(rectangle3_xs[2115]), .RECT3_Y(rectangle3_ys[2115]), .RECT3_WIDTH(rectangle3_widths[2115]), .RECT3_HEIGHT(rectangle3_heights[2115]), .RECT3_WEIGHT(rectangle3_weights[2115]), .FEAT_THRES(feature_thresholds[2115]), .FEAT_ABOVE(feature_aboves[2115]), .FEAT_BELOW(feature_belows[2115])) ac2115(.scan_win(scan_win2115), .scan_win_std_dev(scan_win_std_dev[2115]), .feature_accum(feature_accums[2115]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2116]), .RECT1_Y(rectangle1_ys[2116]), .RECT1_WIDTH(rectangle1_widths[2116]), .RECT1_HEIGHT(rectangle1_heights[2116]), .RECT1_WEIGHT(rectangle1_weights[2116]), .RECT2_X(rectangle2_xs[2116]), .RECT2_Y(rectangle2_ys[2116]), .RECT2_WIDTH(rectangle2_widths[2116]), .RECT2_HEIGHT(rectangle2_heights[2116]), .RECT2_WEIGHT(rectangle2_weights[2116]), .RECT3_X(rectangle3_xs[2116]), .RECT3_Y(rectangle3_ys[2116]), .RECT3_WIDTH(rectangle3_widths[2116]), .RECT3_HEIGHT(rectangle3_heights[2116]), .RECT3_WEIGHT(rectangle3_weights[2116]), .FEAT_THRES(feature_thresholds[2116]), .FEAT_ABOVE(feature_aboves[2116]), .FEAT_BELOW(feature_belows[2116])) ac2116(.scan_win(scan_win2116), .scan_win_std_dev(scan_win_std_dev[2116]), .feature_accum(feature_accums[2116]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2117]), .RECT1_Y(rectangle1_ys[2117]), .RECT1_WIDTH(rectangle1_widths[2117]), .RECT1_HEIGHT(rectangle1_heights[2117]), .RECT1_WEIGHT(rectangle1_weights[2117]), .RECT2_X(rectangle2_xs[2117]), .RECT2_Y(rectangle2_ys[2117]), .RECT2_WIDTH(rectangle2_widths[2117]), .RECT2_HEIGHT(rectangle2_heights[2117]), .RECT2_WEIGHT(rectangle2_weights[2117]), .RECT3_X(rectangle3_xs[2117]), .RECT3_Y(rectangle3_ys[2117]), .RECT3_WIDTH(rectangle3_widths[2117]), .RECT3_HEIGHT(rectangle3_heights[2117]), .RECT3_WEIGHT(rectangle3_weights[2117]), .FEAT_THRES(feature_thresholds[2117]), .FEAT_ABOVE(feature_aboves[2117]), .FEAT_BELOW(feature_belows[2117])) ac2117(.scan_win(scan_win2117), .scan_win_std_dev(scan_win_std_dev[2117]), .feature_accum(feature_accums[2117]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2118]), .RECT1_Y(rectangle1_ys[2118]), .RECT1_WIDTH(rectangle1_widths[2118]), .RECT1_HEIGHT(rectangle1_heights[2118]), .RECT1_WEIGHT(rectangle1_weights[2118]), .RECT2_X(rectangle2_xs[2118]), .RECT2_Y(rectangle2_ys[2118]), .RECT2_WIDTH(rectangle2_widths[2118]), .RECT2_HEIGHT(rectangle2_heights[2118]), .RECT2_WEIGHT(rectangle2_weights[2118]), .RECT3_X(rectangle3_xs[2118]), .RECT3_Y(rectangle3_ys[2118]), .RECT3_WIDTH(rectangle3_widths[2118]), .RECT3_HEIGHT(rectangle3_heights[2118]), .RECT3_WEIGHT(rectangle3_weights[2118]), .FEAT_THRES(feature_thresholds[2118]), .FEAT_ABOVE(feature_aboves[2118]), .FEAT_BELOW(feature_belows[2118])) ac2118(.scan_win(scan_win2118), .scan_win_std_dev(scan_win_std_dev[2118]), .feature_accum(feature_accums[2118]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2119]), .RECT1_Y(rectangle1_ys[2119]), .RECT1_WIDTH(rectangle1_widths[2119]), .RECT1_HEIGHT(rectangle1_heights[2119]), .RECT1_WEIGHT(rectangle1_weights[2119]), .RECT2_X(rectangle2_xs[2119]), .RECT2_Y(rectangle2_ys[2119]), .RECT2_WIDTH(rectangle2_widths[2119]), .RECT2_HEIGHT(rectangle2_heights[2119]), .RECT2_WEIGHT(rectangle2_weights[2119]), .RECT3_X(rectangle3_xs[2119]), .RECT3_Y(rectangle3_ys[2119]), .RECT3_WIDTH(rectangle3_widths[2119]), .RECT3_HEIGHT(rectangle3_heights[2119]), .RECT3_WEIGHT(rectangle3_weights[2119]), .FEAT_THRES(feature_thresholds[2119]), .FEAT_ABOVE(feature_aboves[2119]), .FEAT_BELOW(feature_belows[2119])) ac2119(.scan_win(scan_win2119), .scan_win_std_dev(scan_win_std_dev[2119]), .feature_accum(feature_accums[2119]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2120]), .RECT1_Y(rectangle1_ys[2120]), .RECT1_WIDTH(rectangle1_widths[2120]), .RECT1_HEIGHT(rectangle1_heights[2120]), .RECT1_WEIGHT(rectangle1_weights[2120]), .RECT2_X(rectangle2_xs[2120]), .RECT2_Y(rectangle2_ys[2120]), .RECT2_WIDTH(rectangle2_widths[2120]), .RECT2_HEIGHT(rectangle2_heights[2120]), .RECT2_WEIGHT(rectangle2_weights[2120]), .RECT3_X(rectangle3_xs[2120]), .RECT3_Y(rectangle3_ys[2120]), .RECT3_WIDTH(rectangle3_widths[2120]), .RECT3_HEIGHT(rectangle3_heights[2120]), .RECT3_WEIGHT(rectangle3_weights[2120]), .FEAT_THRES(feature_thresholds[2120]), .FEAT_ABOVE(feature_aboves[2120]), .FEAT_BELOW(feature_belows[2120])) ac2120(.scan_win(scan_win2120), .scan_win_std_dev(scan_win_std_dev[2120]), .feature_accum(feature_accums[2120]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2121]), .RECT1_Y(rectangle1_ys[2121]), .RECT1_WIDTH(rectangle1_widths[2121]), .RECT1_HEIGHT(rectangle1_heights[2121]), .RECT1_WEIGHT(rectangle1_weights[2121]), .RECT2_X(rectangle2_xs[2121]), .RECT2_Y(rectangle2_ys[2121]), .RECT2_WIDTH(rectangle2_widths[2121]), .RECT2_HEIGHT(rectangle2_heights[2121]), .RECT2_WEIGHT(rectangle2_weights[2121]), .RECT3_X(rectangle3_xs[2121]), .RECT3_Y(rectangle3_ys[2121]), .RECT3_WIDTH(rectangle3_widths[2121]), .RECT3_HEIGHT(rectangle3_heights[2121]), .RECT3_WEIGHT(rectangle3_weights[2121]), .FEAT_THRES(feature_thresholds[2121]), .FEAT_ABOVE(feature_aboves[2121]), .FEAT_BELOW(feature_belows[2121])) ac2121(.scan_win(scan_win2121), .scan_win_std_dev(scan_win_std_dev[2121]), .feature_accum(feature_accums[2121]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2122]), .RECT1_Y(rectangle1_ys[2122]), .RECT1_WIDTH(rectangle1_widths[2122]), .RECT1_HEIGHT(rectangle1_heights[2122]), .RECT1_WEIGHT(rectangle1_weights[2122]), .RECT2_X(rectangle2_xs[2122]), .RECT2_Y(rectangle2_ys[2122]), .RECT2_WIDTH(rectangle2_widths[2122]), .RECT2_HEIGHT(rectangle2_heights[2122]), .RECT2_WEIGHT(rectangle2_weights[2122]), .RECT3_X(rectangle3_xs[2122]), .RECT3_Y(rectangle3_ys[2122]), .RECT3_WIDTH(rectangle3_widths[2122]), .RECT3_HEIGHT(rectangle3_heights[2122]), .RECT3_WEIGHT(rectangle3_weights[2122]), .FEAT_THRES(feature_thresholds[2122]), .FEAT_ABOVE(feature_aboves[2122]), .FEAT_BELOW(feature_belows[2122])) ac2122(.scan_win(scan_win2122), .scan_win_std_dev(scan_win_std_dev[2122]), .feature_accum(feature_accums[2122]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2123]), .RECT1_Y(rectangle1_ys[2123]), .RECT1_WIDTH(rectangle1_widths[2123]), .RECT1_HEIGHT(rectangle1_heights[2123]), .RECT1_WEIGHT(rectangle1_weights[2123]), .RECT2_X(rectangle2_xs[2123]), .RECT2_Y(rectangle2_ys[2123]), .RECT2_WIDTH(rectangle2_widths[2123]), .RECT2_HEIGHT(rectangle2_heights[2123]), .RECT2_WEIGHT(rectangle2_weights[2123]), .RECT3_X(rectangle3_xs[2123]), .RECT3_Y(rectangle3_ys[2123]), .RECT3_WIDTH(rectangle3_widths[2123]), .RECT3_HEIGHT(rectangle3_heights[2123]), .RECT3_WEIGHT(rectangle3_weights[2123]), .FEAT_THRES(feature_thresholds[2123]), .FEAT_ABOVE(feature_aboves[2123]), .FEAT_BELOW(feature_belows[2123])) ac2123(.scan_win(scan_win2123), .scan_win_std_dev(scan_win_std_dev[2123]), .feature_accum(feature_accums[2123]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2124]), .RECT1_Y(rectangle1_ys[2124]), .RECT1_WIDTH(rectangle1_widths[2124]), .RECT1_HEIGHT(rectangle1_heights[2124]), .RECT1_WEIGHT(rectangle1_weights[2124]), .RECT2_X(rectangle2_xs[2124]), .RECT2_Y(rectangle2_ys[2124]), .RECT2_WIDTH(rectangle2_widths[2124]), .RECT2_HEIGHT(rectangle2_heights[2124]), .RECT2_WEIGHT(rectangle2_weights[2124]), .RECT3_X(rectangle3_xs[2124]), .RECT3_Y(rectangle3_ys[2124]), .RECT3_WIDTH(rectangle3_widths[2124]), .RECT3_HEIGHT(rectangle3_heights[2124]), .RECT3_WEIGHT(rectangle3_weights[2124]), .FEAT_THRES(feature_thresholds[2124]), .FEAT_ABOVE(feature_aboves[2124]), .FEAT_BELOW(feature_belows[2124])) ac2124(.scan_win(scan_win2124), .scan_win_std_dev(scan_win_std_dev[2124]), .feature_accum(feature_accums[2124]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2125]), .RECT1_Y(rectangle1_ys[2125]), .RECT1_WIDTH(rectangle1_widths[2125]), .RECT1_HEIGHT(rectangle1_heights[2125]), .RECT1_WEIGHT(rectangle1_weights[2125]), .RECT2_X(rectangle2_xs[2125]), .RECT2_Y(rectangle2_ys[2125]), .RECT2_WIDTH(rectangle2_widths[2125]), .RECT2_HEIGHT(rectangle2_heights[2125]), .RECT2_WEIGHT(rectangle2_weights[2125]), .RECT3_X(rectangle3_xs[2125]), .RECT3_Y(rectangle3_ys[2125]), .RECT3_WIDTH(rectangle3_widths[2125]), .RECT3_HEIGHT(rectangle3_heights[2125]), .RECT3_WEIGHT(rectangle3_weights[2125]), .FEAT_THRES(feature_thresholds[2125]), .FEAT_ABOVE(feature_aboves[2125]), .FEAT_BELOW(feature_belows[2125])) ac2125(.scan_win(scan_win2125), .scan_win_std_dev(scan_win_std_dev[2125]), .feature_accum(feature_accums[2125]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2126]), .RECT1_Y(rectangle1_ys[2126]), .RECT1_WIDTH(rectangle1_widths[2126]), .RECT1_HEIGHT(rectangle1_heights[2126]), .RECT1_WEIGHT(rectangle1_weights[2126]), .RECT2_X(rectangle2_xs[2126]), .RECT2_Y(rectangle2_ys[2126]), .RECT2_WIDTH(rectangle2_widths[2126]), .RECT2_HEIGHT(rectangle2_heights[2126]), .RECT2_WEIGHT(rectangle2_weights[2126]), .RECT3_X(rectangle3_xs[2126]), .RECT3_Y(rectangle3_ys[2126]), .RECT3_WIDTH(rectangle3_widths[2126]), .RECT3_HEIGHT(rectangle3_heights[2126]), .RECT3_WEIGHT(rectangle3_weights[2126]), .FEAT_THRES(feature_thresholds[2126]), .FEAT_ABOVE(feature_aboves[2126]), .FEAT_BELOW(feature_belows[2126])) ac2126(.scan_win(scan_win2126), .scan_win_std_dev(scan_win_std_dev[2126]), .feature_accum(feature_accums[2126]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2127]), .RECT1_Y(rectangle1_ys[2127]), .RECT1_WIDTH(rectangle1_widths[2127]), .RECT1_HEIGHT(rectangle1_heights[2127]), .RECT1_WEIGHT(rectangle1_weights[2127]), .RECT2_X(rectangle2_xs[2127]), .RECT2_Y(rectangle2_ys[2127]), .RECT2_WIDTH(rectangle2_widths[2127]), .RECT2_HEIGHT(rectangle2_heights[2127]), .RECT2_WEIGHT(rectangle2_weights[2127]), .RECT3_X(rectangle3_xs[2127]), .RECT3_Y(rectangle3_ys[2127]), .RECT3_WIDTH(rectangle3_widths[2127]), .RECT3_HEIGHT(rectangle3_heights[2127]), .RECT3_WEIGHT(rectangle3_weights[2127]), .FEAT_THRES(feature_thresholds[2127]), .FEAT_ABOVE(feature_aboves[2127]), .FEAT_BELOW(feature_belows[2127])) ac2127(.scan_win(scan_win2127), .scan_win_std_dev(scan_win_std_dev[2127]), .feature_accum(feature_accums[2127]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2128]), .RECT1_Y(rectangle1_ys[2128]), .RECT1_WIDTH(rectangle1_widths[2128]), .RECT1_HEIGHT(rectangle1_heights[2128]), .RECT1_WEIGHT(rectangle1_weights[2128]), .RECT2_X(rectangle2_xs[2128]), .RECT2_Y(rectangle2_ys[2128]), .RECT2_WIDTH(rectangle2_widths[2128]), .RECT2_HEIGHT(rectangle2_heights[2128]), .RECT2_WEIGHT(rectangle2_weights[2128]), .RECT3_X(rectangle3_xs[2128]), .RECT3_Y(rectangle3_ys[2128]), .RECT3_WIDTH(rectangle3_widths[2128]), .RECT3_HEIGHT(rectangle3_heights[2128]), .RECT3_WEIGHT(rectangle3_weights[2128]), .FEAT_THRES(feature_thresholds[2128]), .FEAT_ABOVE(feature_aboves[2128]), .FEAT_BELOW(feature_belows[2128])) ac2128(.scan_win(scan_win2128), .scan_win_std_dev(scan_win_std_dev[2128]), .feature_accum(feature_accums[2128]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2129]), .RECT1_Y(rectangle1_ys[2129]), .RECT1_WIDTH(rectangle1_widths[2129]), .RECT1_HEIGHT(rectangle1_heights[2129]), .RECT1_WEIGHT(rectangle1_weights[2129]), .RECT2_X(rectangle2_xs[2129]), .RECT2_Y(rectangle2_ys[2129]), .RECT2_WIDTH(rectangle2_widths[2129]), .RECT2_HEIGHT(rectangle2_heights[2129]), .RECT2_WEIGHT(rectangle2_weights[2129]), .RECT3_X(rectangle3_xs[2129]), .RECT3_Y(rectangle3_ys[2129]), .RECT3_WIDTH(rectangle3_widths[2129]), .RECT3_HEIGHT(rectangle3_heights[2129]), .RECT3_WEIGHT(rectangle3_weights[2129]), .FEAT_THRES(feature_thresholds[2129]), .FEAT_ABOVE(feature_aboves[2129]), .FEAT_BELOW(feature_belows[2129])) ac2129(.scan_win(scan_win2129), .scan_win_std_dev(scan_win_std_dev[2129]), .feature_accum(feature_accums[2129]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2130]), .RECT1_Y(rectangle1_ys[2130]), .RECT1_WIDTH(rectangle1_widths[2130]), .RECT1_HEIGHT(rectangle1_heights[2130]), .RECT1_WEIGHT(rectangle1_weights[2130]), .RECT2_X(rectangle2_xs[2130]), .RECT2_Y(rectangle2_ys[2130]), .RECT2_WIDTH(rectangle2_widths[2130]), .RECT2_HEIGHT(rectangle2_heights[2130]), .RECT2_WEIGHT(rectangle2_weights[2130]), .RECT3_X(rectangle3_xs[2130]), .RECT3_Y(rectangle3_ys[2130]), .RECT3_WIDTH(rectangle3_widths[2130]), .RECT3_HEIGHT(rectangle3_heights[2130]), .RECT3_WEIGHT(rectangle3_weights[2130]), .FEAT_THRES(feature_thresholds[2130]), .FEAT_ABOVE(feature_aboves[2130]), .FEAT_BELOW(feature_belows[2130])) ac2130(.scan_win(scan_win2130), .scan_win_std_dev(scan_win_std_dev[2130]), .feature_accum(feature_accums[2130]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2131]), .RECT1_Y(rectangle1_ys[2131]), .RECT1_WIDTH(rectangle1_widths[2131]), .RECT1_HEIGHT(rectangle1_heights[2131]), .RECT1_WEIGHT(rectangle1_weights[2131]), .RECT2_X(rectangle2_xs[2131]), .RECT2_Y(rectangle2_ys[2131]), .RECT2_WIDTH(rectangle2_widths[2131]), .RECT2_HEIGHT(rectangle2_heights[2131]), .RECT2_WEIGHT(rectangle2_weights[2131]), .RECT3_X(rectangle3_xs[2131]), .RECT3_Y(rectangle3_ys[2131]), .RECT3_WIDTH(rectangle3_widths[2131]), .RECT3_HEIGHT(rectangle3_heights[2131]), .RECT3_WEIGHT(rectangle3_weights[2131]), .FEAT_THRES(feature_thresholds[2131]), .FEAT_ABOVE(feature_aboves[2131]), .FEAT_BELOW(feature_belows[2131])) ac2131(.scan_win(scan_win2131), .scan_win_std_dev(scan_win_std_dev[2131]), .feature_accum(feature_accums[2131]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2132]), .RECT1_Y(rectangle1_ys[2132]), .RECT1_WIDTH(rectangle1_widths[2132]), .RECT1_HEIGHT(rectangle1_heights[2132]), .RECT1_WEIGHT(rectangle1_weights[2132]), .RECT2_X(rectangle2_xs[2132]), .RECT2_Y(rectangle2_ys[2132]), .RECT2_WIDTH(rectangle2_widths[2132]), .RECT2_HEIGHT(rectangle2_heights[2132]), .RECT2_WEIGHT(rectangle2_weights[2132]), .RECT3_X(rectangle3_xs[2132]), .RECT3_Y(rectangle3_ys[2132]), .RECT3_WIDTH(rectangle3_widths[2132]), .RECT3_HEIGHT(rectangle3_heights[2132]), .RECT3_WEIGHT(rectangle3_weights[2132]), .FEAT_THRES(feature_thresholds[2132]), .FEAT_ABOVE(feature_aboves[2132]), .FEAT_BELOW(feature_belows[2132])) ac2132(.scan_win(scan_win2132), .scan_win_std_dev(scan_win_std_dev[2132]), .feature_accum(feature_accums[2132]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2133]), .RECT1_Y(rectangle1_ys[2133]), .RECT1_WIDTH(rectangle1_widths[2133]), .RECT1_HEIGHT(rectangle1_heights[2133]), .RECT1_WEIGHT(rectangle1_weights[2133]), .RECT2_X(rectangle2_xs[2133]), .RECT2_Y(rectangle2_ys[2133]), .RECT2_WIDTH(rectangle2_widths[2133]), .RECT2_HEIGHT(rectangle2_heights[2133]), .RECT2_WEIGHT(rectangle2_weights[2133]), .RECT3_X(rectangle3_xs[2133]), .RECT3_Y(rectangle3_ys[2133]), .RECT3_WIDTH(rectangle3_widths[2133]), .RECT3_HEIGHT(rectangle3_heights[2133]), .RECT3_WEIGHT(rectangle3_weights[2133]), .FEAT_THRES(feature_thresholds[2133]), .FEAT_ABOVE(feature_aboves[2133]), .FEAT_BELOW(feature_belows[2133])) ac2133(.scan_win(scan_win2133), .scan_win_std_dev(scan_win_std_dev[2133]), .feature_accum(feature_accums[2133]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2134]), .RECT1_Y(rectangle1_ys[2134]), .RECT1_WIDTH(rectangle1_widths[2134]), .RECT1_HEIGHT(rectangle1_heights[2134]), .RECT1_WEIGHT(rectangle1_weights[2134]), .RECT2_X(rectangle2_xs[2134]), .RECT2_Y(rectangle2_ys[2134]), .RECT2_WIDTH(rectangle2_widths[2134]), .RECT2_HEIGHT(rectangle2_heights[2134]), .RECT2_WEIGHT(rectangle2_weights[2134]), .RECT3_X(rectangle3_xs[2134]), .RECT3_Y(rectangle3_ys[2134]), .RECT3_WIDTH(rectangle3_widths[2134]), .RECT3_HEIGHT(rectangle3_heights[2134]), .RECT3_WEIGHT(rectangle3_weights[2134]), .FEAT_THRES(feature_thresholds[2134]), .FEAT_ABOVE(feature_aboves[2134]), .FEAT_BELOW(feature_belows[2134])) ac2134(.scan_win(scan_win2134), .scan_win_std_dev(scan_win_std_dev[2134]), .feature_accum(feature_accums[2134]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2135]), .RECT1_Y(rectangle1_ys[2135]), .RECT1_WIDTH(rectangle1_widths[2135]), .RECT1_HEIGHT(rectangle1_heights[2135]), .RECT1_WEIGHT(rectangle1_weights[2135]), .RECT2_X(rectangle2_xs[2135]), .RECT2_Y(rectangle2_ys[2135]), .RECT2_WIDTH(rectangle2_widths[2135]), .RECT2_HEIGHT(rectangle2_heights[2135]), .RECT2_WEIGHT(rectangle2_weights[2135]), .RECT3_X(rectangle3_xs[2135]), .RECT3_Y(rectangle3_ys[2135]), .RECT3_WIDTH(rectangle3_widths[2135]), .RECT3_HEIGHT(rectangle3_heights[2135]), .RECT3_WEIGHT(rectangle3_weights[2135]), .FEAT_THRES(feature_thresholds[2135]), .FEAT_ABOVE(feature_aboves[2135]), .FEAT_BELOW(feature_belows[2135])) ac2135(.scan_win(scan_win2135), .scan_win_std_dev(scan_win_std_dev[2135]), .feature_accum(feature_accums[2135]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2136]), .RECT1_Y(rectangle1_ys[2136]), .RECT1_WIDTH(rectangle1_widths[2136]), .RECT1_HEIGHT(rectangle1_heights[2136]), .RECT1_WEIGHT(rectangle1_weights[2136]), .RECT2_X(rectangle2_xs[2136]), .RECT2_Y(rectangle2_ys[2136]), .RECT2_WIDTH(rectangle2_widths[2136]), .RECT2_HEIGHT(rectangle2_heights[2136]), .RECT2_WEIGHT(rectangle2_weights[2136]), .RECT3_X(rectangle3_xs[2136]), .RECT3_Y(rectangle3_ys[2136]), .RECT3_WIDTH(rectangle3_widths[2136]), .RECT3_HEIGHT(rectangle3_heights[2136]), .RECT3_WEIGHT(rectangle3_weights[2136]), .FEAT_THRES(feature_thresholds[2136]), .FEAT_ABOVE(feature_aboves[2136]), .FEAT_BELOW(feature_belows[2136])) ac2136(.scan_win(scan_win2136), .scan_win_std_dev(scan_win_std_dev[2136]), .feature_accum(feature_accums[2136]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2137]), .RECT1_Y(rectangle1_ys[2137]), .RECT1_WIDTH(rectangle1_widths[2137]), .RECT1_HEIGHT(rectangle1_heights[2137]), .RECT1_WEIGHT(rectangle1_weights[2137]), .RECT2_X(rectangle2_xs[2137]), .RECT2_Y(rectangle2_ys[2137]), .RECT2_WIDTH(rectangle2_widths[2137]), .RECT2_HEIGHT(rectangle2_heights[2137]), .RECT2_WEIGHT(rectangle2_weights[2137]), .RECT3_X(rectangle3_xs[2137]), .RECT3_Y(rectangle3_ys[2137]), .RECT3_WIDTH(rectangle3_widths[2137]), .RECT3_HEIGHT(rectangle3_heights[2137]), .RECT3_WEIGHT(rectangle3_weights[2137]), .FEAT_THRES(feature_thresholds[2137]), .FEAT_ABOVE(feature_aboves[2137]), .FEAT_BELOW(feature_belows[2137])) ac2137(.scan_win(scan_win2137), .scan_win_std_dev(scan_win_std_dev[2137]), .feature_accum(feature_accums[2137]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2138]), .RECT1_Y(rectangle1_ys[2138]), .RECT1_WIDTH(rectangle1_widths[2138]), .RECT1_HEIGHT(rectangle1_heights[2138]), .RECT1_WEIGHT(rectangle1_weights[2138]), .RECT2_X(rectangle2_xs[2138]), .RECT2_Y(rectangle2_ys[2138]), .RECT2_WIDTH(rectangle2_widths[2138]), .RECT2_HEIGHT(rectangle2_heights[2138]), .RECT2_WEIGHT(rectangle2_weights[2138]), .RECT3_X(rectangle3_xs[2138]), .RECT3_Y(rectangle3_ys[2138]), .RECT3_WIDTH(rectangle3_widths[2138]), .RECT3_HEIGHT(rectangle3_heights[2138]), .RECT3_WEIGHT(rectangle3_weights[2138]), .FEAT_THRES(feature_thresholds[2138]), .FEAT_ABOVE(feature_aboves[2138]), .FEAT_BELOW(feature_belows[2138])) ac2138(.scan_win(scan_win2138), .scan_win_std_dev(scan_win_std_dev[2138]), .feature_accum(feature_accums[2138]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2139]), .RECT1_Y(rectangle1_ys[2139]), .RECT1_WIDTH(rectangle1_widths[2139]), .RECT1_HEIGHT(rectangle1_heights[2139]), .RECT1_WEIGHT(rectangle1_weights[2139]), .RECT2_X(rectangle2_xs[2139]), .RECT2_Y(rectangle2_ys[2139]), .RECT2_WIDTH(rectangle2_widths[2139]), .RECT2_HEIGHT(rectangle2_heights[2139]), .RECT2_WEIGHT(rectangle2_weights[2139]), .RECT3_X(rectangle3_xs[2139]), .RECT3_Y(rectangle3_ys[2139]), .RECT3_WIDTH(rectangle3_widths[2139]), .RECT3_HEIGHT(rectangle3_heights[2139]), .RECT3_WEIGHT(rectangle3_weights[2139]), .FEAT_THRES(feature_thresholds[2139]), .FEAT_ABOVE(feature_aboves[2139]), .FEAT_BELOW(feature_belows[2139])) ac2139(.scan_win(scan_win2139), .scan_win_std_dev(scan_win_std_dev[2139]), .feature_accum(feature_accums[2139]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2140]), .RECT1_Y(rectangle1_ys[2140]), .RECT1_WIDTH(rectangle1_widths[2140]), .RECT1_HEIGHT(rectangle1_heights[2140]), .RECT1_WEIGHT(rectangle1_weights[2140]), .RECT2_X(rectangle2_xs[2140]), .RECT2_Y(rectangle2_ys[2140]), .RECT2_WIDTH(rectangle2_widths[2140]), .RECT2_HEIGHT(rectangle2_heights[2140]), .RECT2_WEIGHT(rectangle2_weights[2140]), .RECT3_X(rectangle3_xs[2140]), .RECT3_Y(rectangle3_ys[2140]), .RECT3_WIDTH(rectangle3_widths[2140]), .RECT3_HEIGHT(rectangle3_heights[2140]), .RECT3_WEIGHT(rectangle3_weights[2140]), .FEAT_THRES(feature_thresholds[2140]), .FEAT_ABOVE(feature_aboves[2140]), .FEAT_BELOW(feature_belows[2140])) ac2140(.scan_win(scan_win2140), .scan_win_std_dev(scan_win_std_dev[2140]), .feature_accum(feature_accums[2140]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2141]), .RECT1_Y(rectangle1_ys[2141]), .RECT1_WIDTH(rectangle1_widths[2141]), .RECT1_HEIGHT(rectangle1_heights[2141]), .RECT1_WEIGHT(rectangle1_weights[2141]), .RECT2_X(rectangle2_xs[2141]), .RECT2_Y(rectangle2_ys[2141]), .RECT2_WIDTH(rectangle2_widths[2141]), .RECT2_HEIGHT(rectangle2_heights[2141]), .RECT2_WEIGHT(rectangle2_weights[2141]), .RECT3_X(rectangle3_xs[2141]), .RECT3_Y(rectangle3_ys[2141]), .RECT3_WIDTH(rectangle3_widths[2141]), .RECT3_HEIGHT(rectangle3_heights[2141]), .RECT3_WEIGHT(rectangle3_weights[2141]), .FEAT_THRES(feature_thresholds[2141]), .FEAT_ABOVE(feature_aboves[2141]), .FEAT_BELOW(feature_belows[2141])) ac2141(.scan_win(scan_win2141), .scan_win_std_dev(scan_win_std_dev[2141]), .feature_accum(feature_accums[2141]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2142]), .RECT1_Y(rectangle1_ys[2142]), .RECT1_WIDTH(rectangle1_widths[2142]), .RECT1_HEIGHT(rectangle1_heights[2142]), .RECT1_WEIGHT(rectangle1_weights[2142]), .RECT2_X(rectangle2_xs[2142]), .RECT2_Y(rectangle2_ys[2142]), .RECT2_WIDTH(rectangle2_widths[2142]), .RECT2_HEIGHT(rectangle2_heights[2142]), .RECT2_WEIGHT(rectangle2_weights[2142]), .RECT3_X(rectangle3_xs[2142]), .RECT3_Y(rectangle3_ys[2142]), .RECT3_WIDTH(rectangle3_widths[2142]), .RECT3_HEIGHT(rectangle3_heights[2142]), .RECT3_WEIGHT(rectangle3_weights[2142]), .FEAT_THRES(feature_thresholds[2142]), .FEAT_ABOVE(feature_aboves[2142]), .FEAT_BELOW(feature_belows[2142])) ac2142(.scan_win(scan_win2142), .scan_win_std_dev(scan_win_std_dev[2142]), .feature_accum(feature_accums[2142]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2143]), .RECT1_Y(rectangle1_ys[2143]), .RECT1_WIDTH(rectangle1_widths[2143]), .RECT1_HEIGHT(rectangle1_heights[2143]), .RECT1_WEIGHT(rectangle1_weights[2143]), .RECT2_X(rectangle2_xs[2143]), .RECT2_Y(rectangle2_ys[2143]), .RECT2_WIDTH(rectangle2_widths[2143]), .RECT2_HEIGHT(rectangle2_heights[2143]), .RECT2_WEIGHT(rectangle2_weights[2143]), .RECT3_X(rectangle3_xs[2143]), .RECT3_Y(rectangle3_ys[2143]), .RECT3_WIDTH(rectangle3_widths[2143]), .RECT3_HEIGHT(rectangle3_heights[2143]), .RECT3_WEIGHT(rectangle3_weights[2143]), .FEAT_THRES(feature_thresholds[2143]), .FEAT_ABOVE(feature_aboves[2143]), .FEAT_BELOW(feature_belows[2143])) ac2143(.scan_win(scan_win2143), .scan_win_std_dev(scan_win_std_dev[2143]), .feature_accum(feature_accums[2143]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2144]), .RECT1_Y(rectangle1_ys[2144]), .RECT1_WIDTH(rectangle1_widths[2144]), .RECT1_HEIGHT(rectangle1_heights[2144]), .RECT1_WEIGHT(rectangle1_weights[2144]), .RECT2_X(rectangle2_xs[2144]), .RECT2_Y(rectangle2_ys[2144]), .RECT2_WIDTH(rectangle2_widths[2144]), .RECT2_HEIGHT(rectangle2_heights[2144]), .RECT2_WEIGHT(rectangle2_weights[2144]), .RECT3_X(rectangle3_xs[2144]), .RECT3_Y(rectangle3_ys[2144]), .RECT3_WIDTH(rectangle3_widths[2144]), .RECT3_HEIGHT(rectangle3_heights[2144]), .RECT3_WEIGHT(rectangle3_weights[2144]), .FEAT_THRES(feature_thresholds[2144]), .FEAT_ABOVE(feature_aboves[2144]), .FEAT_BELOW(feature_belows[2144])) ac2144(.scan_win(scan_win2144), .scan_win_std_dev(scan_win_std_dev[2144]), .feature_accum(feature_accums[2144]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2145]), .RECT1_Y(rectangle1_ys[2145]), .RECT1_WIDTH(rectangle1_widths[2145]), .RECT1_HEIGHT(rectangle1_heights[2145]), .RECT1_WEIGHT(rectangle1_weights[2145]), .RECT2_X(rectangle2_xs[2145]), .RECT2_Y(rectangle2_ys[2145]), .RECT2_WIDTH(rectangle2_widths[2145]), .RECT2_HEIGHT(rectangle2_heights[2145]), .RECT2_WEIGHT(rectangle2_weights[2145]), .RECT3_X(rectangle3_xs[2145]), .RECT3_Y(rectangle3_ys[2145]), .RECT3_WIDTH(rectangle3_widths[2145]), .RECT3_HEIGHT(rectangle3_heights[2145]), .RECT3_WEIGHT(rectangle3_weights[2145]), .FEAT_THRES(feature_thresholds[2145]), .FEAT_ABOVE(feature_aboves[2145]), .FEAT_BELOW(feature_belows[2145])) ac2145(.scan_win(scan_win2145), .scan_win_std_dev(scan_win_std_dev[2145]), .feature_accum(feature_accums[2145]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2146]), .RECT1_Y(rectangle1_ys[2146]), .RECT1_WIDTH(rectangle1_widths[2146]), .RECT1_HEIGHT(rectangle1_heights[2146]), .RECT1_WEIGHT(rectangle1_weights[2146]), .RECT2_X(rectangle2_xs[2146]), .RECT2_Y(rectangle2_ys[2146]), .RECT2_WIDTH(rectangle2_widths[2146]), .RECT2_HEIGHT(rectangle2_heights[2146]), .RECT2_WEIGHT(rectangle2_weights[2146]), .RECT3_X(rectangle3_xs[2146]), .RECT3_Y(rectangle3_ys[2146]), .RECT3_WIDTH(rectangle3_widths[2146]), .RECT3_HEIGHT(rectangle3_heights[2146]), .RECT3_WEIGHT(rectangle3_weights[2146]), .FEAT_THRES(feature_thresholds[2146]), .FEAT_ABOVE(feature_aboves[2146]), .FEAT_BELOW(feature_belows[2146])) ac2146(.scan_win(scan_win2146), .scan_win_std_dev(scan_win_std_dev[2146]), .feature_accum(feature_accums[2146]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2147]), .RECT1_Y(rectangle1_ys[2147]), .RECT1_WIDTH(rectangle1_widths[2147]), .RECT1_HEIGHT(rectangle1_heights[2147]), .RECT1_WEIGHT(rectangle1_weights[2147]), .RECT2_X(rectangle2_xs[2147]), .RECT2_Y(rectangle2_ys[2147]), .RECT2_WIDTH(rectangle2_widths[2147]), .RECT2_HEIGHT(rectangle2_heights[2147]), .RECT2_WEIGHT(rectangle2_weights[2147]), .RECT3_X(rectangle3_xs[2147]), .RECT3_Y(rectangle3_ys[2147]), .RECT3_WIDTH(rectangle3_widths[2147]), .RECT3_HEIGHT(rectangle3_heights[2147]), .RECT3_WEIGHT(rectangle3_weights[2147]), .FEAT_THRES(feature_thresholds[2147]), .FEAT_ABOVE(feature_aboves[2147]), .FEAT_BELOW(feature_belows[2147])) ac2147(.scan_win(scan_win2147), .scan_win_std_dev(scan_win_std_dev[2147]), .feature_accum(feature_accums[2147]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2148]), .RECT1_Y(rectangle1_ys[2148]), .RECT1_WIDTH(rectangle1_widths[2148]), .RECT1_HEIGHT(rectangle1_heights[2148]), .RECT1_WEIGHT(rectangle1_weights[2148]), .RECT2_X(rectangle2_xs[2148]), .RECT2_Y(rectangle2_ys[2148]), .RECT2_WIDTH(rectangle2_widths[2148]), .RECT2_HEIGHT(rectangle2_heights[2148]), .RECT2_WEIGHT(rectangle2_weights[2148]), .RECT3_X(rectangle3_xs[2148]), .RECT3_Y(rectangle3_ys[2148]), .RECT3_WIDTH(rectangle3_widths[2148]), .RECT3_HEIGHT(rectangle3_heights[2148]), .RECT3_WEIGHT(rectangle3_weights[2148]), .FEAT_THRES(feature_thresholds[2148]), .FEAT_ABOVE(feature_aboves[2148]), .FEAT_BELOW(feature_belows[2148])) ac2148(.scan_win(scan_win2148), .scan_win_std_dev(scan_win_std_dev[2148]), .feature_accum(feature_accums[2148]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2149]), .RECT1_Y(rectangle1_ys[2149]), .RECT1_WIDTH(rectangle1_widths[2149]), .RECT1_HEIGHT(rectangle1_heights[2149]), .RECT1_WEIGHT(rectangle1_weights[2149]), .RECT2_X(rectangle2_xs[2149]), .RECT2_Y(rectangle2_ys[2149]), .RECT2_WIDTH(rectangle2_widths[2149]), .RECT2_HEIGHT(rectangle2_heights[2149]), .RECT2_WEIGHT(rectangle2_weights[2149]), .RECT3_X(rectangle3_xs[2149]), .RECT3_Y(rectangle3_ys[2149]), .RECT3_WIDTH(rectangle3_widths[2149]), .RECT3_HEIGHT(rectangle3_heights[2149]), .RECT3_WEIGHT(rectangle3_weights[2149]), .FEAT_THRES(feature_thresholds[2149]), .FEAT_ABOVE(feature_aboves[2149]), .FEAT_BELOW(feature_belows[2149])) ac2149(.scan_win(scan_win2149), .scan_win_std_dev(scan_win_std_dev[2149]), .feature_accum(feature_accums[2149]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2150]), .RECT1_Y(rectangle1_ys[2150]), .RECT1_WIDTH(rectangle1_widths[2150]), .RECT1_HEIGHT(rectangle1_heights[2150]), .RECT1_WEIGHT(rectangle1_weights[2150]), .RECT2_X(rectangle2_xs[2150]), .RECT2_Y(rectangle2_ys[2150]), .RECT2_WIDTH(rectangle2_widths[2150]), .RECT2_HEIGHT(rectangle2_heights[2150]), .RECT2_WEIGHT(rectangle2_weights[2150]), .RECT3_X(rectangle3_xs[2150]), .RECT3_Y(rectangle3_ys[2150]), .RECT3_WIDTH(rectangle3_widths[2150]), .RECT3_HEIGHT(rectangle3_heights[2150]), .RECT3_WEIGHT(rectangle3_weights[2150]), .FEAT_THRES(feature_thresholds[2150]), .FEAT_ABOVE(feature_aboves[2150]), .FEAT_BELOW(feature_belows[2150])) ac2150(.scan_win(scan_win2150), .scan_win_std_dev(scan_win_std_dev[2150]), .feature_accum(feature_accums[2150]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2151]), .RECT1_Y(rectangle1_ys[2151]), .RECT1_WIDTH(rectangle1_widths[2151]), .RECT1_HEIGHT(rectangle1_heights[2151]), .RECT1_WEIGHT(rectangle1_weights[2151]), .RECT2_X(rectangle2_xs[2151]), .RECT2_Y(rectangle2_ys[2151]), .RECT2_WIDTH(rectangle2_widths[2151]), .RECT2_HEIGHT(rectangle2_heights[2151]), .RECT2_WEIGHT(rectangle2_weights[2151]), .RECT3_X(rectangle3_xs[2151]), .RECT3_Y(rectangle3_ys[2151]), .RECT3_WIDTH(rectangle3_widths[2151]), .RECT3_HEIGHT(rectangle3_heights[2151]), .RECT3_WEIGHT(rectangle3_weights[2151]), .FEAT_THRES(feature_thresholds[2151]), .FEAT_ABOVE(feature_aboves[2151]), .FEAT_BELOW(feature_belows[2151])) ac2151(.scan_win(scan_win2151), .scan_win_std_dev(scan_win_std_dev[2151]), .feature_accum(feature_accums[2151]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2152]), .RECT1_Y(rectangle1_ys[2152]), .RECT1_WIDTH(rectangle1_widths[2152]), .RECT1_HEIGHT(rectangle1_heights[2152]), .RECT1_WEIGHT(rectangle1_weights[2152]), .RECT2_X(rectangle2_xs[2152]), .RECT2_Y(rectangle2_ys[2152]), .RECT2_WIDTH(rectangle2_widths[2152]), .RECT2_HEIGHT(rectangle2_heights[2152]), .RECT2_WEIGHT(rectangle2_weights[2152]), .RECT3_X(rectangle3_xs[2152]), .RECT3_Y(rectangle3_ys[2152]), .RECT3_WIDTH(rectangle3_widths[2152]), .RECT3_HEIGHT(rectangle3_heights[2152]), .RECT3_WEIGHT(rectangle3_weights[2152]), .FEAT_THRES(feature_thresholds[2152]), .FEAT_ABOVE(feature_aboves[2152]), .FEAT_BELOW(feature_belows[2152])) ac2152(.scan_win(scan_win2152), .scan_win_std_dev(scan_win_std_dev[2152]), .feature_accum(feature_accums[2152]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2153]), .RECT1_Y(rectangle1_ys[2153]), .RECT1_WIDTH(rectangle1_widths[2153]), .RECT1_HEIGHT(rectangle1_heights[2153]), .RECT1_WEIGHT(rectangle1_weights[2153]), .RECT2_X(rectangle2_xs[2153]), .RECT2_Y(rectangle2_ys[2153]), .RECT2_WIDTH(rectangle2_widths[2153]), .RECT2_HEIGHT(rectangle2_heights[2153]), .RECT2_WEIGHT(rectangle2_weights[2153]), .RECT3_X(rectangle3_xs[2153]), .RECT3_Y(rectangle3_ys[2153]), .RECT3_WIDTH(rectangle3_widths[2153]), .RECT3_HEIGHT(rectangle3_heights[2153]), .RECT3_WEIGHT(rectangle3_weights[2153]), .FEAT_THRES(feature_thresholds[2153]), .FEAT_ABOVE(feature_aboves[2153]), .FEAT_BELOW(feature_belows[2153])) ac2153(.scan_win(scan_win2153), .scan_win_std_dev(scan_win_std_dev[2153]), .feature_accum(feature_accums[2153]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2154]), .RECT1_Y(rectangle1_ys[2154]), .RECT1_WIDTH(rectangle1_widths[2154]), .RECT1_HEIGHT(rectangle1_heights[2154]), .RECT1_WEIGHT(rectangle1_weights[2154]), .RECT2_X(rectangle2_xs[2154]), .RECT2_Y(rectangle2_ys[2154]), .RECT2_WIDTH(rectangle2_widths[2154]), .RECT2_HEIGHT(rectangle2_heights[2154]), .RECT2_WEIGHT(rectangle2_weights[2154]), .RECT3_X(rectangle3_xs[2154]), .RECT3_Y(rectangle3_ys[2154]), .RECT3_WIDTH(rectangle3_widths[2154]), .RECT3_HEIGHT(rectangle3_heights[2154]), .RECT3_WEIGHT(rectangle3_weights[2154]), .FEAT_THRES(feature_thresholds[2154]), .FEAT_ABOVE(feature_aboves[2154]), .FEAT_BELOW(feature_belows[2154])) ac2154(.scan_win(scan_win2154), .scan_win_std_dev(scan_win_std_dev[2154]), .feature_accum(feature_accums[2154]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2155]), .RECT1_Y(rectangle1_ys[2155]), .RECT1_WIDTH(rectangle1_widths[2155]), .RECT1_HEIGHT(rectangle1_heights[2155]), .RECT1_WEIGHT(rectangle1_weights[2155]), .RECT2_X(rectangle2_xs[2155]), .RECT2_Y(rectangle2_ys[2155]), .RECT2_WIDTH(rectangle2_widths[2155]), .RECT2_HEIGHT(rectangle2_heights[2155]), .RECT2_WEIGHT(rectangle2_weights[2155]), .RECT3_X(rectangle3_xs[2155]), .RECT3_Y(rectangle3_ys[2155]), .RECT3_WIDTH(rectangle3_widths[2155]), .RECT3_HEIGHT(rectangle3_heights[2155]), .RECT3_WEIGHT(rectangle3_weights[2155]), .FEAT_THRES(feature_thresholds[2155]), .FEAT_ABOVE(feature_aboves[2155]), .FEAT_BELOW(feature_belows[2155])) ac2155(.scan_win(scan_win2155), .scan_win_std_dev(scan_win_std_dev[2155]), .feature_accum(feature_accums[2155]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2156]), .RECT1_Y(rectangle1_ys[2156]), .RECT1_WIDTH(rectangle1_widths[2156]), .RECT1_HEIGHT(rectangle1_heights[2156]), .RECT1_WEIGHT(rectangle1_weights[2156]), .RECT2_X(rectangle2_xs[2156]), .RECT2_Y(rectangle2_ys[2156]), .RECT2_WIDTH(rectangle2_widths[2156]), .RECT2_HEIGHT(rectangle2_heights[2156]), .RECT2_WEIGHT(rectangle2_weights[2156]), .RECT3_X(rectangle3_xs[2156]), .RECT3_Y(rectangle3_ys[2156]), .RECT3_WIDTH(rectangle3_widths[2156]), .RECT3_HEIGHT(rectangle3_heights[2156]), .RECT3_WEIGHT(rectangle3_weights[2156]), .FEAT_THRES(feature_thresholds[2156]), .FEAT_ABOVE(feature_aboves[2156]), .FEAT_BELOW(feature_belows[2156])) ac2156(.scan_win(scan_win2156), .scan_win_std_dev(scan_win_std_dev[2156]), .feature_accum(feature_accums[2156]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2157]), .RECT1_Y(rectangle1_ys[2157]), .RECT1_WIDTH(rectangle1_widths[2157]), .RECT1_HEIGHT(rectangle1_heights[2157]), .RECT1_WEIGHT(rectangle1_weights[2157]), .RECT2_X(rectangle2_xs[2157]), .RECT2_Y(rectangle2_ys[2157]), .RECT2_WIDTH(rectangle2_widths[2157]), .RECT2_HEIGHT(rectangle2_heights[2157]), .RECT2_WEIGHT(rectangle2_weights[2157]), .RECT3_X(rectangle3_xs[2157]), .RECT3_Y(rectangle3_ys[2157]), .RECT3_WIDTH(rectangle3_widths[2157]), .RECT3_HEIGHT(rectangle3_heights[2157]), .RECT3_WEIGHT(rectangle3_weights[2157]), .FEAT_THRES(feature_thresholds[2157]), .FEAT_ABOVE(feature_aboves[2157]), .FEAT_BELOW(feature_belows[2157])) ac2157(.scan_win(scan_win2157), .scan_win_std_dev(scan_win_std_dev[2157]), .feature_accum(feature_accums[2157]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2158]), .RECT1_Y(rectangle1_ys[2158]), .RECT1_WIDTH(rectangle1_widths[2158]), .RECT1_HEIGHT(rectangle1_heights[2158]), .RECT1_WEIGHT(rectangle1_weights[2158]), .RECT2_X(rectangle2_xs[2158]), .RECT2_Y(rectangle2_ys[2158]), .RECT2_WIDTH(rectangle2_widths[2158]), .RECT2_HEIGHT(rectangle2_heights[2158]), .RECT2_WEIGHT(rectangle2_weights[2158]), .RECT3_X(rectangle3_xs[2158]), .RECT3_Y(rectangle3_ys[2158]), .RECT3_WIDTH(rectangle3_widths[2158]), .RECT3_HEIGHT(rectangle3_heights[2158]), .RECT3_WEIGHT(rectangle3_weights[2158]), .FEAT_THRES(feature_thresholds[2158]), .FEAT_ABOVE(feature_aboves[2158]), .FEAT_BELOW(feature_belows[2158])) ac2158(.scan_win(scan_win2158), .scan_win_std_dev(scan_win_std_dev[2158]), .feature_accum(feature_accums[2158]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2159]), .RECT1_Y(rectangle1_ys[2159]), .RECT1_WIDTH(rectangle1_widths[2159]), .RECT1_HEIGHT(rectangle1_heights[2159]), .RECT1_WEIGHT(rectangle1_weights[2159]), .RECT2_X(rectangle2_xs[2159]), .RECT2_Y(rectangle2_ys[2159]), .RECT2_WIDTH(rectangle2_widths[2159]), .RECT2_HEIGHT(rectangle2_heights[2159]), .RECT2_WEIGHT(rectangle2_weights[2159]), .RECT3_X(rectangle3_xs[2159]), .RECT3_Y(rectangle3_ys[2159]), .RECT3_WIDTH(rectangle3_widths[2159]), .RECT3_HEIGHT(rectangle3_heights[2159]), .RECT3_WEIGHT(rectangle3_weights[2159]), .FEAT_THRES(feature_thresholds[2159]), .FEAT_ABOVE(feature_aboves[2159]), .FEAT_BELOW(feature_belows[2159])) ac2159(.scan_win(scan_win2159), .scan_win_std_dev(scan_win_std_dev[2159]), .feature_accum(feature_accums[2159]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2160]), .RECT1_Y(rectangle1_ys[2160]), .RECT1_WIDTH(rectangle1_widths[2160]), .RECT1_HEIGHT(rectangle1_heights[2160]), .RECT1_WEIGHT(rectangle1_weights[2160]), .RECT2_X(rectangle2_xs[2160]), .RECT2_Y(rectangle2_ys[2160]), .RECT2_WIDTH(rectangle2_widths[2160]), .RECT2_HEIGHT(rectangle2_heights[2160]), .RECT2_WEIGHT(rectangle2_weights[2160]), .RECT3_X(rectangle3_xs[2160]), .RECT3_Y(rectangle3_ys[2160]), .RECT3_WIDTH(rectangle3_widths[2160]), .RECT3_HEIGHT(rectangle3_heights[2160]), .RECT3_WEIGHT(rectangle3_weights[2160]), .FEAT_THRES(feature_thresholds[2160]), .FEAT_ABOVE(feature_aboves[2160]), .FEAT_BELOW(feature_belows[2160])) ac2160(.scan_win(scan_win2160), .scan_win_std_dev(scan_win_std_dev[2160]), .feature_accum(feature_accums[2160]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2161]), .RECT1_Y(rectangle1_ys[2161]), .RECT1_WIDTH(rectangle1_widths[2161]), .RECT1_HEIGHT(rectangle1_heights[2161]), .RECT1_WEIGHT(rectangle1_weights[2161]), .RECT2_X(rectangle2_xs[2161]), .RECT2_Y(rectangle2_ys[2161]), .RECT2_WIDTH(rectangle2_widths[2161]), .RECT2_HEIGHT(rectangle2_heights[2161]), .RECT2_WEIGHT(rectangle2_weights[2161]), .RECT3_X(rectangle3_xs[2161]), .RECT3_Y(rectangle3_ys[2161]), .RECT3_WIDTH(rectangle3_widths[2161]), .RECT3_HEIGHT(rectangle3_heights[2161]), .RECT3_WEIGHT(rectangle3_weights[2161]), .FEAT_THRES(feature_thresholds[2161]), .FEAT_ABOVE(feature_aboves[2161]), .FEAT_BELOW(feature_belows[2161])) ac2161(.scan_win(scan_win2161), .scan_win_std_dev(scan_win_std_dev[2161]), .feature_accum(feature_accums[2161]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2162]), .RECT1_Y(rectangle1_ys[2162]), .RECT1_WIDTH(rectangle1_widths[2162]), .RECT1_HEIGHT(rectangle1_heights[2162]), .RECT1_WEIGHT(rectangle1_weights[2162]), .RECT2_X(rectangle2_xs[2162]), .RECT2_Y(rectangle2_ys[2162]), .RECT2_WIDTH(rectangle2_widths[2162]), .RECT2_HEIGHT(rectangle2_heights[2162]), .RECT2_WEIGHT(rectangle2_weights[2162]), .RECT3_X(rectangle3_xs[2162]), .RECT3_Y(rectangle3_ys[2162]), .RECT3_WIDTH(rectangle3_widths[2162]), .RECT3_HEIGHT(rectangle3_heights[2162]), .RECT3_WEIGHT(rectangle3_weights[2162]), .FEAT_THRES(feature_thresholds[2162]), .FEAT_ABOVE(feature_aboves[2162]), .FEAT_BELOW(feature_belows[2162])) ac2162(.scan_win(scan_win2162), .scan_win_std_dev(scan_win_std_dev[2162]), .feature_accum(feature_accums[2162]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2163]), .RECT1_Y(rectangle1_ys[2163]), .RECT1_WIDTH(rectangle1_widths[2163]), .RECT1_HEIGHT(rectangle1_heights[2163]), .RECT1_WEIGHT(rectangle1_weights[2163]), .RECT2_X(rectangle2_xs[2163]), .RECT2_Y(rectangle2_ys[2163]), .RECT2_WIDTH(rectangle2_widths[2163]), .RECT2_HEIGHT(rectangle2_heights[2163]), .RECT2_WEIGHT(rectangle2_weights[2163]), .RECT3_X(rectangle3_xs[2163]), .RECT3_Y(rectangle3_ys[2163]), .RECT3_WIDTH(rectangle3_widths[2163]), .RECT3_HEIGHT(rectangle3_heights[2163]), .RECT3_WEIGHT(rectangle3_weights[2163]), .FEAT_THRES(feature_thresholds[2163]), .FEAT_ABOVE(feature_aboves[2163]), .FEAT_BELOW(feature_belows[2163])) ac2163(.scan_win(scan_win2163), .scan_win_std_dev(scan_win_std_dev[2163]), .feature_accum(feature_accums[2163]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2164]), .RECT1_Y(rectangle1_ys[2164]), .RECT1_WIDTH(rectangle1_widths[2164]), .RECT1_HEIGHT(rectangle1_heights[2164]), .RECT1_WEIGHT(rectangle1_weights[2164]), .RECT2_X(rectangle2_xs[2164]), .RECT2_Y(rectangle2_ys[2164]), .RECT2_WIDTH(rectangle2_widths[2164]), .RECT2_HEIGHT(rectangle2_heights[2164]), .RECT2_WEIGHT(rectangle2_weights[2164]), .RECT3_X(rectangle3_xs[2164]), .RECT3_Y(rectangle3_ys[2164]), .RECT3_WIDTH(rectangle3_widths[2164]), .RECT3_HEIGHT(rectangle3_heights[2164]), .RECT3_WEIGHT(rectangle3_weights[2164]), .FEAT_THRES(feature_thresholds[2164]), .FEAT_ABOVE(feature_aboves[2164]), .FEAT_BELOW(feature_belows[2164])) ac2164(.scan_win(scan_win2164), .scan_win_std_dev(scan_win_std_dev[2164]), .feature_accum(feature_accums[2164]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2165]), .RECT1_Y(rectangle1_ys[2165]), .RECT1_WIDTH(rectangle1_widths[2165]), .RECT1_HEIGHT(rectangle1_heights[2165]), .RECT1_WEIGHT(rectangle1_weights[2165]), .RECT2_X(rectangle2_xs[2165]), .RECT2_Y(rectangle2_ys[2165]), .RECT2_WIDTH(rectangle2_widths[2165]), .RECT2_HEIGHT(rectangle2_heights[2165]), .RECT2_WEIGHT(rectangle2_weights[2165]), .RECT3_X(rectangle3_xs[2165]), .RECT3_Y(rectangle3_ys[2165]), .RECT3_WIDTH(rectangle3_widths[2165]), .RECT3_HEIGHT(rectangle3_heights[2165]), .RECT3_WEIGHT(rectangle3_weights[2165]), .FEAT_THRES(feature_thresholds[2165]), .FEAT_ABOVE(feature_aboves[2165]), .FEAT_BELOW(feature_belows[2165])) ac2165(.scan_win(scan_win2165), .scan_win_std_dev(scan_win_std_dev[2165]), .feature_accum(feature_accums[2165]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2166]), .RECT1_Y(rectangle1_ys[2166]), .RECT1_WIDTH(rectangle1_widths[2166]), .RECT1_HEIGHT(rectangle1_heights[2166]), .RECT1_WEIGHT(rectangle1_weights[2166]), .RECT2_X(rectangle2_xs[2166]), .RECT2_Y(rectangle2_ys[2166]), .RECT2_WIDTH(rectangle2_widths[2166]), .RECT2_HEIGHT(rectangle2_heights[2166]), .RECT2_WEIGHT(rectangle2_weights[2166]), .RECT3_X(rectangle3_xs[2166]), .RECT3_Y(rectangle3_ys[2166]), .RECT3_WIDTH(rectangle3_widths[2166]), .RECT3_HEIGHT(rectangle3_heights[2166]), .RECT3_WEIGHT(rectangle3_weights[2166]), .FEAT_THRES(feature_thresholds[2166]), .FEAT_ABOVE(feature_aboves[2166]), .FEAT_BELOW(feature_belows[2166])) ac2166(.scan_win(scan_win2166), .scan_win_std_dev(scan_win_std_dev[2166]), .feature_accum(feature_accums[2166]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2167]), .RECT1_Y(rectangle1_ys[2167]), .RECT1_WIDTH(rectangle1_widths[2167]), .RECT1_HEIGHT(rectangle1_heights[2167]), .RECT1_WEIGHT(rectangle1_weights[2167]), .RECT2_X(rectangle2_xs[2167]), .RECT2_Y(rectangle2_ys[2167]), .RECT2_WIDTH(rectangle2_widths[2167]), .RECT2_HEIGHT(rectangle2_heights[2167]), .RECT2_WEIGHT(rectangle2_weights[2167]), .RECT3_X(rectangle3_xs[2167]), .RECT3_Y(rectangle3_ys[2167]), .RECT3_WIDTH(rectangle3_widths[2167]), .RECT3_HEIGHT(rectangle3_heights[2167]), .RECT3_WEIGHT(rectangle3_weights[2167]), .FEAT_THRES(feature_thresholds[2167]), .FEAT_ABOVE(feature_aboves[2167]), .FEAT_BELOW(feature_belows[2167])) ac2167(.scan_win(scan_win2167), .scan_win_std_dev(scan_win_std_dev[2167]), .feature_accum(feature_accums[2167]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2168]), .RECT1_Y(rectangle1_ys[2168]), .RECT1_WIDTH(rectangle1_widths[2168]), .RECT1_HEIGHT(rectangle1_heights[2168]), .RECT1_WEIGHT(rectangle1_weights[2168]), .RECT2_X(rectangle2_xs[2168]), .RECT2_Y(rectangle2_ys[2168]), .RECT2_WIDTH(rectangle2_widths[2168]), .RECT2_HEIGHT(rectangle2_heights[2168]), .RECT2_WEIGHT(rectangle2_weights[2168]), .RECT3_X(rectangle3_xs[2168]), .RECT3_Y(rectangle3_ys[2168]), .RECT3_WIDTH(rectangle3_widths[2168]), .RECT3_HEIGHT(rectangle3_heights[2168]), .RECT3_WEIGHT(rectangle3_weights[2168]), .FEAT_THRES(feature_thresholds[2168]), .FEAT_ABOVE(feature_aboves[2168]), .FEAT_BELOW(feature_belows[2168])) ac2168(.scan_win(scan_win2168), .scan_win_std_dev(scan_win_std_dev[2168]), .feature_accum(feature_accums[2168]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2169]), .RECT1_Y(rectangle1_ys[2169]), .RECT1_WIDTH(rectangle1_widths[2169]), .RECT1_HEIGHT(rectangle1_heights[2169]), .RECT1_WEIGHT(rectangle1_weights[2169]), .RECT2_X(rectangle2_xs[2169]), .RECT2_Y(rectangle2_ys[2169]), .RECT2_WIDTH(rectangle2_widths[2169]), .RECT2_HEIGHT(rectangle2_heights[2169]), .RECT2_WEIGHT(rectangle2_weights[2169]), .RECT3_X(rectangle3_xs[2169]), .RECT3_Y(rectangle3_ys[2169]), .RECT3_WIDTH(rectangle3_widths[2169]), .RECT3_HEIGHT(rectangle3_heights[2169]), .RECT3_WEIGHT(rectangle3_weights[2169]), .FEAT_THRES(feature_thresholds[2169]), .FEAT_ABOVE(feature_aboves[2169]), .FEAT_BELOW(feature_belows[2169])) ac2169(.scan_win(scan_win2169), .scan_win_std_dev(scan_win_std_dev[2169]), .feature_accum(feature_accums[2169]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2170]), .RECT1_Y(rectangle1_ys[2170]), .RECT1_WIDTH(rectangle1_widths[2170]), .RECT1_HEIGHT(rectangle1_heights[2170]), .RECT1_WEIGHT(rectangle1_weights[2170]), .RECT2_X(rectangle2_xs[2170]), .RECT2_Y(rectangle2_ys[2170]), .RECT2_WIDTH(rectangle2_widths[2170]), .RECT2_HEIGHT(rectangle2_heights[2170]), .RECT2_WEIGHT(rectangle2_weights[2170]), .RECT3_X(rectangle3_xs[2170]), .RECT3_Y(rectangle3_ys[2170]), .RECT3_WIDTH(rectangle3_widths[2170]), .RECT3_HEIGHT(rectangle3_heights[2170]), .RECT3_WEIGHT(rectangle3_weights[2170]), .FEAT_THRES(feature_thresholds[2170]), .FEAT_ABOVE(feature_aboves[2170]), .FEAT_BELOW(feature_belows[2170])) ac2170(.scan_win(scan_win2170), .scan_win_std_dev(scan_win_std_dev[2170]), .feature_accum(feature_accums[2170]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2171]), .RECT1_Y(rectangle1_ys[2171]), .RECT1_WIDTH(rectangle1_widths[2171]), .RECT1_HEIGHT(rectangle1_heights[2171]), .RECT1_WEIGHT(rectangle1_weights[2171]), .RECT2_X(rectangle2_xs[2171]), .RECT2_Y(rectangle2_ys[2171]), .RECT2_WIDTH(rectangle2_widths[2171]), .RECT2_HEIGHT(rectangle2_heights[2171]), .RECT2_WEIGHT(rectangle2_weights[2171]), .RECT3_X(rectangle3_xs[2171]), .RECT3_Y(rectangle3_ys[2171]), .RECT3_WIDTH(rectangle3_widths[2171]), .RECT3_HEIGHT(rectangle3_heights[2171]), .RECT3_WEIGHT(rectangle3_weights[2171]), .FEAT_THRES(feature_thresholds[2171]), .FEAT_ABOVE(feature_aboves[2171]), .FEAT_BELOW(feature_belows[2171])) ac2171(.scan_win(scan_win2171), .scan_win_std_dev(scan_win_std_dev[2171]), .feature_accum(feature_accums[2171]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2172]), .RECT1_Y(rectangle1_ys[2172]), .RECT1_WIDTH(rectangle1_widths[2172]), .RECT1_HEIGHT(rectangle1_heights[2172]), .RECT1_WEIGHT(rectangle1_weights[2172]), .RECT2_X(rectangle2_xs[2172]), .RECT2_Y(rectangle2_ys[2172]), .RECT2_WIDTH(rectangle2_widths[2172]), .RECT2_HEIGHT(rectangle2_heights[2172]), .RECT2_WEIGHT(rectangle2_weights[2172]), .RECT3_X(rectangle3_xs[2172]), .RECT3_Y(rectangle3_ys[2172]), .RECT3_WIDTH(rectangle3_widths[2172]), .RECT3_HEIGHT(rectangle3_heights[2172]), .RECT3_WEIGHT(rectangle3_weights[2172]), .FEAT_THRES(feature_thresholds[2172]), .FEAT_ABOVE(feature_aboves[2172]), .FEAT_BELOW(feature_belows[2172])) ac2172(.scan_win(scan_win2172), .scan_win_std_dev(scan_win_std_dev[2172]), .feature_accum(feature_accums[2172]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2173]), .RECT1_Y(rectangle1_ys[2173]), .RECT1_WIDTH(rectangle1_widths[2173]), .RECT1_HEIGHT(rectangle1_heights[2173]), .RECT1_WEIGHT(rectangle1_weights[2173]), .RECT2_X(rectangle2_xs[2173]), .RECT2_Y(rectangle2_ys[2173]), .RECT2_WIDTH(rectangle2_widths[2173]), .RECT2_HEIGHT(rectangle2_heights[2173]), .RECT2_WEIGHT(rectangle2_weights[2173]), .RECT3_X(rectangle3_xs[2173]), .RECT3_Y(rectangle3_ys[2173]), .RECT3_WIDTH(rectangle3_widths[2173]), .RECT3_HEIGHT(rectangle3_heights[2173]), .RECT3_WEIGHT(rectangle3_weights[2173]), .FEAT_THRES(feature_thresholds[2173]), .FEAT_ABOVE(feature_aboves[2173]), .FEAT_BELOW(feature_belows[2173])) ac2173(.scan_win(scan_win2173), .scan_win_std_dev(scan_win_std_dev[2173]), .feature_accum(feature_accums[2173]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2174]), .RECT1_Y(rectangle1_ys[2174]), .RECT1_WIDTH(rectangle1_widths[2174]), .RECT1_HEIGHT(rectangle1_heights[2174]), .RECT1_WEIGHT(rectangle1_weights[2174]), .RECT2_X(rectangle2_xs[2174]), .RECT2_Y(rectangle2_ys[2174]), .RECT2_WIDTH(rectangle2_widths[2174]), .RECT2_HEIGHT(rectangle2_heights[2174]), .RECT2_WEIGHT(rectangle2_weights[2174]), .RECT3_X(rectangle3_xs[2174]), .RECT3_Y(rectangle3_ys[2174]), .RECT3_WIDTH(rectangle3_widths[2174]), .RECT3_HEIGHT(rectangle3_heights[2174]), .RECT3_WEIGHT(rectangle3_weights[2174]), .FEAT_THRES(feature_thresholds[2174]), .FEAT_ABOVE(feature_aboves[2174]), .FEAT_BELOW(feature_belows[2174])) ac2174(.scan_win(scan_win2174), .scan_win_std_dev(scan_win_std_dev[2174]), .feature_accum(feature_accums[2174]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2175]), .RECT1_Y(rectangle1_ys[2175]), .RECT1_WIDTH(rectangle1_widths[2175]), .RECT1_HEIGHT(rectangle1_heights[2175]), .RECT1_WEIGHT(rectangle1_weights[2175]), .RECT2_X(rectangle2_xs[2175]), .RECT2_Y(rectangle2_ys[2175]), .RECT2_WIDTH(rectangle2_widths[2175]), .RECT2_HEIGHT(rectangle2_heights[2175]), .RECT2_WEIGHT(rectangle2_weights[2175]), .RECT3_X(rectangle3_xs[2175]), .RECT3_Y(rectangle3_ys[2175]), .RECT3_WIDTH(rectangle3_widths[2175]), .RECT3_HEIGHT(rectangle3_heights[2175]), .RECT3_WEIGHT(rectangle3_weights[2175]), .FEAT_THRES(feature_thresholds[2175]), .FEAT_ABOVE(feature_aboves[2175]), .FEAT_BELOW(feature_belows[2175])) ac2175(.scan_win(scan_win2175), .scan_win_std_dev(scan_win_std_dev[2175]), .feature_accum(feature_accums[2175]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2176]), .RECT1_Y(rectangle1_ys[2176]), .RECT1_WIDTH(rectangle1_widths[2176]), .RECT1_HEIGHT(rectangle1_heights[2176]), .RECT1_WEIGHT(rectangle1_weights[2176]), .RECT2_X(rectangle2_xs[2176]), .RECT2_Y(rectangle2_ys[2176]), .RECT2_WIDTH(rectangle2_widths[2176]), .RECT2_HEIGHT(rectangle2_heights[2176]), .RECT2_WEIGHT(rectangle2_weights[2176]), .RECT3_X(rectangle3_xs[2176]), .RECT3_Y(rectangle3_ys[2176]), .RECT3_WIDTH(rectangle3_widths[2176]), .RECT3_HEIGHT(rectangle3_heights[2176]), .RECT3_WEIGHT(rectangle3_weights[2176]), .FEAT_THRES(feature_thresholds[2176]), .FEAT_ABOVE(feature_aboves[2176]), .FEAT_BELOW(feature_belows[2176])) ac2176(.scan_win(scan_win2176), .scan_win_std_dev(scan_win_std_dev[2176]), .feature_accum(feature_accums[2176]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2177]), .RECT1_Y(rectangle1_ys[2177]), .RECT1_WIDTH(rectangle1_widths[2177]), .RECT1_HEIGHT(rectangle1_heights[2177]), .RECT1_WEIGHT(rectangle1_weights[2177]), .RECT2_X(rectangle2_xs[2177]), .RECT2_Y(rectangle2_ys[2177]), .RECT2_WIDTH(rectangle2_widths[2177]), .RECT2_HEIGHT(rectangle2_heights[2177]), .RECT2_WEIGHT(rectangle2_weights[2177]), .RECT3_X(rectangle3_xs[2177]), .RECT3_Y(rectangle3_ys[2177]), .RECT3_WIDTH(rectangle3_widths[2177]), .RECT3_HEIGHT(rectangle3_heights[2177]), .RECT3_WEIGHT(rectangle3_weights[2177]), .FEAT_THRES(feature_thresholds[2177]), .FEAT_ABOVE(feature_aboves[2177]), .FEAT_BELOW(feature_belows[2177])) ac2177(.scan_win(scan_win2177), .scan_win_std_dev(scan_win_std_dev[2177]), .feature_accum(feature_accums[2177]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2178]), .RECT1_Y(rectangle1_ys[2178]), .RECT1_WIDTH(rectangle1_widths[2178]), .RECT1_HEIGHT(rectangle1_heights[2178]), .RECT1_WEIGHT(rectangle1_weights[2178]), .RECT2_X(rectangle2_xs[2178]), .RECT2_Y(rectangle2_ys[2178]), .RECT2_WIDTH(rectangle2_widths[2178]), .RECT2_HEIGHT(rectangle2_heights[2178]), .RECT2_WEIGHT(rectangle2_weights[2178]), .RECT3_X(rectangle3_xs[2178]), .RECT3_Y(rectangle3_ys[2178]), .RECT3_WIDTH(rectangle3_widths[2178]), .RECT3_HEIGHT(rectangle3_heights[2178]), .RECT3_WEIGHT(rectangle3_weights[2178]), .FEAT_THRES(feature_thresholds[2178]), .FEAT_ABOVE(feature_aboves[2178]), .FEAT_BELOW(feature_belows[2178])) ac2178(.scan_win(scan_win2178), .scan_win_std_dev(scan_win_std_dev[2178]), .feature_accum(feature_accums[2178]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2179]), .RECT1_Y(rectangle1_ys[2179]), .RECT1_WIDTH(rectangle1_widths[2179]), .RECT1_HEIGHT(rectangle1_heights[2179]), .RECT1_WEIGHT(rectangle1_weights[2179]), .RECT2_X(rectangle2_xs[2179]), .RECT2_Y(rectangle2_ys[2179]), .RECT2_WIDTH(rectangle2_widths[2179]), .RECT2_HEIGHT(rectangle2_heights[2179]), .RECT2_WEIGHT(rectangle2_weights[2179]), .RECT3_X(rectangle3_xs[2179]), .RECT3_Y(rectangle3_ys[2179]), .RECT3_WIDTH(rectangle3_widths[2179]), .RECT3_HEIGHT(rectangle3_heights[2179]), .RECT3_WEIGHT(rectangle3_weights[2179]), .FEAT_THRES(feature_thresholds[2179]), .FEAT_ABOVE(feature_aboves[2179]), .FEAT_BELOW(feature_belows[2179])) ac2179(.scan_win(scan_win2179), .scan_win_std_dev(scan_win_std_dev[2179]), .feature_accum(feature_accums[2179]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2180]), .RECT1_Y(rectangle1_ys[2180]), .RECT1_WIDTH(rectangle1_widths[2180]), .RECT1_HEIGHT(rectangle1_heights[2180]), .RECT1_WEIGHT(rectangle1_weights[2180]), .RECT2_X(rectangle2_xs[2180]), .RECT2_Y(rectangle2_ys[2180]), .RECT2_WIDTH(rectangle2_widths[2180]), .RECT2_HEIGHT(rectangle2_heights[2180]), .RECT2_WEIGHT(rectangle2_weights[2180]), .RECT3_X(rectangle3_xs[2180]), .RECT3_Y(rectangle3_ys[2180]), .RECT3_WIDTH(rectangle3_widths[2180]), .RECT3_HEIGHT(rectangle3_heights[2180]), .RECT3_WEIGHT(rectangle3_weights[2180]), .FEAT_THRES(feature_thresholds[2180]), .FEAT_ABOVE(feature_aboves[2180]), .FEAT_BELOW(feature_belows[2180])) ac2180(.scan_win(scan_win2180), .scan_win_std_dev(scan_win_std_dev[2180]), .feature_accum(feature_accums[2180]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2181]), .RECT1_Y(rectangle1_ys[2181]), .RECT1_WIDTH(rectangle1_widths[2181]), .RECT1_HEIGHT(rectangle1_heights[2181]), .RECT1_WEIGHT(rectangle1_weights[2181]), .RECT2_X(rectangle2_xs[2181]), .RECT2_Y(rectangle2_ys[2181]), .RECT2_WIDTH(rectangle2_widths[2181]), .RECT2_HEIGHT(rectangle2_heights[2181]), .RECT2_WEIGHT(rectangle2_weights[2181]), .RECT3_X(rectangle3_xs[2181]), .RECT3_Y(rectangle3_ys[2181]), .RECT3_WIDTH(rectangle3_widths[2181]), .RECT3_HEIGHT(rectangle3_heights[2181]), .RECT3_WEIGHT(rectangle3_weights[2181]), .FEAT_THRES(feature_thresholds[2181]), .FEAT_ABOVE(feature_aboves[2181]), .FEAT_BELOW(feature_belows[2181])) ac2181(.scan_win(scan_win2181), .scan_win_std_dev(scan_win_std_dev[2181]), .feature_accum(feature_accums[2181]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2182]), .RECT1_Y(rectangle1_ys[2182]), .RECT1_WIDTH(rectangle1_widths[2182]), .RECT1_HEIGHT(rectangle1_heights[2182]), .RECT1_WEIGHT(rectangle1_weights[2182]), .RECT2_X(rectangle2_xs[2182]), .RECT2_Y(rectangle2_ys[2182]), .RECT2_WIDTH(rectangle2_widths[2182]), .RECT2_HEIGHT(rectangle2_heights[2182]), .RECT2_WEIGHT(rectangle2_weights[2182]), .RECT3_X(rectangle3_xs[2182]), .RECT3_Y(rectangle3_ys[2182]), .RECT3_WIDTH(rectangle3_widths[2182]), .RECT3_HEIGHT(rectangle3_heights[2182]), .RECT3_WEIGHT(rectangle3_weights[2182]), .FEAT_THRES(feature_thresholds[2182]), .FEAT_ABOVE(feature_aboves[2182]), .FEAT_BELOW(feature_belows[2182])) ac2182(.scan_win(scan_win2182), .scan_win_std_dev(scan_win_std_dev[2182]), .feature_accum(feature_accums[2182]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2183]), .RECT1_Y(rectangle1_ys[2183]), .RECT1_WIDTH(rectangle1_widths[2183]), .RECT1_HEIGHT(rectangle1_heights[2183]), .RECT1_WEIGHT(rectangle1_weights[2183]), .RECT2_X(rectangle2_xs[2183]), .RECT2_Y(rectangle2_ys[2183]), .RECT2_WIDTH(rectangle2_widths[2183]), .RECT2_HEIGHT(rectangle2_heights[2183]), .RECT2_WEIGHT(rectangle2_weights[2183]), .RECT3_X(rectangle3_xs[2183]), .RECT3_Y(rectangle3_ys[2183]), .RECT3_WIDTH(rectangle3_widths[2183]), .RECT3_HEIGHT(rectangle3_heights[2183]), .RECT3_WEIGHT(rectangle3_weights[2183]), .FEAT_THRES(feature_thresholds[2183]), .FEAT_ABOVE(feature_aboves[2183]), .FEAT_BELOW(feature_belows[2183])) ac2183(.scan_win(scan_win2183), .scan_win_std_dev(scan_win_std_dev[2183]), .feature_accum(feature_accums[2183]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2184]), .RECT1_Y(rectangle1_ys[2184]), .RECT1_WIDTH(rectangle1_widths[2184]), .RECT1_HEIGHT(rectangle1_heights[2184]), .RECT1_WEIGHT(rectangle1_weights[2184]), .RECT2_X(rectangle2_xs[2184]), .RECT2_Y(rectangle2_ys[2184]), .RECT2_WIDTH(rectangle2_widths[2184]), .RECT2_HEIGHT(rectangle2_heights[2184]), .RECT2_WEIGHT(rectangle2_weights[2184]), .RECT3_X(rectangle3_xs[2184]), .RECT3_Y(rectangle3_ys[2184]), .RECT3_WIDTH(rectangle3_widths[2184]), .RECT3_HEIGHT(rectangle3_heights[2184]), .RECT3_WEIGHT(rectangle3_weights[2184]), .FEAT_THRES(feature_thresholds[2184]), .FEAT_ABOVE(feature_aboves[2184]), .FEAT_BELOW(feature_belows[2184])) ac2184(.scan_win(scan_win2184), .scan_win_std_dev(scan_win_std_dev[2184]), .feature_accum(feature_accums[2184]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2185]), .RECT1_Y(rectangle1_ys[2185]), .RECT1_WIDTH(rectangle1_widths[2185]), .RECT1_HEIGHT(rectangle1_heights[2185]), .RECT1_WEIGHT(rectangle1_weights[2185]), .RECT2_X(rectangle2_xs[2185]), .RECT2_Y(rectangle2_ys[2185]), .RECT2_WIDTH(rectangle2_widths[2185]), .RECT2_HEIGHT(rectangle2_heights[2185]), .RECT2_WEIGHT(rectangle2_weights[2185]), .RECT3_X(rectangle3_xs[2185]), .RECT3_Y(rectangle3_ys[2185]), .RECT3_WIDTH(rectangle3_widths[2185]), .RECT3_HEIGHT(rectangle3_heights[2185]), .RECT3_WEIGHT(rectangle3_weights[2185]), .FEAT_THRES(feature_thresholds[2185]), .FEAT_ABOVE(feature_aboves[2185]), .FEAT_BELOW(feature_belows[2185])) ac2185(.scan_win(scan_win2185), .scan_win_std_dev(scan_win_std_dev[2185]), .feature_accum(feature_accums[2185]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2186]), .RECT1_Y(rectangle1_ys[2186]), .RECT1_WIDTH(rectangle1_widths[2186]), .RECT1_HEIGHT(rectangle1_heights[2186]), .RECT1_WEIGHT(rectangle1_weights[2186]), .RECT2_X(rectangle2_xs[2186]), .RECT2_Y(rectangle2_ys[2186]), .RECT2_WIDTH(rectangle2_widths[2186]), .RECT2_HEIGHT(rectangle2_heights[2186]), .RECT2_WEIGHT(rectangle2_weights[2186]), .RECT3_X(rectangle3_xs[2186]), .RECT3_Y(rectangle3_ys[2186]), .RECT3_WIDTH(rectangle3_widths[2186]), .RECT3_HEIGHT(rectangle3_heights[2186]), .RECT3_WEIGHT(rectangle3_weights[2186]), .FEAT_THRES(feature_thresholds[2186]), .FEAT_ABOVE(feature_aboves[2186]), .FEAT_BELOW(feature_belows[2186])) ac2186(.scan_win(scan_win2186), .scan_win_std_dev(scan_win_std_dev[2186]), .feature_accum(feature_accums[2186]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2187]), .RECT1_Y(rectangle1_ys[2187]), .RECT1_WIDTH(rectangle1_widths[2187]), .RECT1_HEIGHT(rectangle1_heights[2187]), .RECT1_WEIGHT(rectangle1_weights[2187]), .RECT2_X(rectangle2_xs[2187]), .RECT2_Y(rectangle2_ys[2187]), .RECT2_WIDTH(rectangle2_widths[2187]), .RECT2_HEIGHT(rectangle2_heights[2187]), .RECT2_WEIGHT(rectangle2_weights[2187]), .RECT3_X(rectangle3_xs[2187]), .RECT3_Y(rectangle3_ys[2187]), .RECT3_WIDTH(rectangle3_widths[2187]), .RECT3_HEIGHT(rectangle3_heights[2187]), .RECT3_WEIGHT(rectangle3_weights[2187]), .FEAT_THRES(feature_thresholds[2187]), .FEAT_ABOVE(feature_aboves[2187]), .FEAT_BELOW(feature_belows[2187])) ac2187(.scan_win(scan_win2187), .scan_win_std_dev(scan_win_std_dev[2187]), .feature_accum(feature_accums[2187]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2188]), .RECT1_Y(rectangle1_ys[2188]), .RECT1_WIDTH(rectangle1_widths[2188]), .RECT1_HEIGHT(rectangle1_heights[2188]), .RECT1_WEIGHT(rectangle1_weights[2188]), .RECT2_X(rectangle2_xs[2188]), .RECT2_Y(rectangle2_ys[2188]), .RECT2_WIDTH(rectangle2_widths[2188]), .RECT2_HEIGHT(rectangle2_heights[2188]), .RECT2_WEIGHT(rectangle2_weights[2188]), .RECT3_X(rectangle3_xs[2188]), .RECT3_Y(rectangle3_ys[2188]), .RECT3_WIDTH(rectangle3_widths[2188]), .RECT3_HEIGHT(rectangle3_heights[2188]), .RECT3_WEIGHT(rectangle3_weights[2188]), .FEAT_THRES(feature_thresholds[2188]), .FEAT_ABOVE(feature_aboves[2188]), .FEAT_BELOW(feature_belows[2188])) ac2188(.scan_win(scan_win2188), .scan_win_std_dev(scan_win_std_dev[2188]), .feature_accum(feature_accums[2188]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2189]), .RECT1_Y(rectangle1_ys[2189]), .RECT1_WIDTH(rectangle1_widths[2189]), .RECT1_HEIGHT(rectangle1_heights[2189]), .RECT1_WEIGHT(rectangle1_weights[2189]), .RECT2_X(rectangle2_xs[2189]), .RECT2_Y(rectangle2_ys[2189]), .RECT2_WIDTH(rectangle2_widths[2189]), .RECT2_HEIGHT(rectangle2_heights[2189]), .RECT2_WEIGHT(rectangle2_weights[2189]), .RECT3_X(rectangle3_xs[2189]), .RECT3_Y(rectangle3_ys[2189]), .RECT3_WIDTH(rectangle3_widths[2189]), .RECT3_HEIGHT(rectangle3_heights[2189]), .RECT3_WEIGHT(rectangle3_weights[2189]), .FEAT_THRES(feature_thresholds[2189]), .FEAT_ABOVE(feature_aboves[2189]), .FEAT_BELOW(feature_belows[2189])) ac2189(.scan_win(scan_win2189), .scan_win_std_dev(scan_win_std_dev[2189]), .feature_accum(feature_accums[2189]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2190]), .RECT1_Y(rectangle1_ys[2190]), .RECT1_WIDTH(rectangle1_widths[2190]), .RECT1_HEIGHT(rectangle1_heights[2190]), .RECT1_WEIGHT(rectangle1_weights[2190]), .RECT2_X(rectangle2_xs[2190]), .RECT2_Y(rectangle2_ys[2190]), .RECT2_WIDTH(rectangle2_widths[2190]), .RECT2_HEIGHT(rectangle2_heights[2190]), .RECT2_WEIGHT(rectangle2_weights[2190]), .RECT3_X(rectangle3_xs[2190]), .RECT3_Y(rectangle3_ys[2190]), .RECT3_WIDTH(rectangle3_widths[2190]), .RECT3_HEIGHT(rectangle3_heights[2190]), .RECT3_WEIGHT(rectangle3_weights[2190]), .FEAT_THRES(feature_thresholds[2190]), .FEAT_ABOVE(feature_aboves[2190]), .FEAT_BELOW(feature_belows[2190])) ac2190(.scan_win(scan_win2190), .scan_win_std_dev(scan_win_std_dev[2190]), .feature_accum(feature_accums[2190]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2191]), .RECT1_Y(rectangle1_ys[2191]), .RECT1_WIDTH(rectangle1_widths[2191]), .RECT1_HEIGHT(rectangle1_heights[2191]), .RECT1_WEIGHT(rectangle1_weights[2191]), .RECT2_X(rectangle2_xs[2191]), .RECT2_Y(rectangle2_ys[2191]), .RECT2_WIDTH(rectangle2_widths[2191]), .RECT2_HEIGHT(rectangle2_heights[2191]), .RECT2_WEIGHT(rectangle2_weights[2191]), .RECT3_X(rectangle3_xs[2191]), .RECT3_Y(rectangle3_ys[2191]), .RECT3_WIDTH(rectangle3_widths[2191]), .RECT3_HEIGHT(rectangle3_heights[2191]), .RECT3_WEIGHT(rectangle3_weights[2191]), .FEAT_THRES(feature_thresholds[2191]), .FEAT_ABOVE(feature_aboves[2191]), .FEAT_BELOW(feature_belows[2191])) ac2191(.scan_win(scan_win2191), .scan_win_std_dev(scan_win_std_dev[2191]), .feature_accum(feature_accums[2191]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2192]), .RECT1_Y(rectangle1_ys[2192]), .RECT1_WIDTH(rectangle1_widths[2192]), .RECT1_HEIGHT(rectangle1_heights[2192]), .RECT1_WEIGHT(rectangle1_weights[2192]), .RECT2_X(rectangle2_xs[2192]), .RECT2_Y(rectangle2_ys[2192]), .RECT2_WIDTH(rectangle2_widths[2192]), .RECT2_HEIGHT(rectangle2_heights[2192]), .RECT2_WEIGHT(rectangle2_weights[2192]), .RECT3_X(rectangle3_xs[2192]), .RECT3_Y(rectangle3_ys[2192]), .RECT3_WIDTH(rectangle3_widths[2192]), .RECT3_HEIGHT(rectangle3_heights[2192]), .RECT3_WEIGHT(rectangle3_weights[2192]), .FEAT_THRES(feature_thresholds[2192]), .FEAT_ABOVE(feature_aboves[2192]), .FEAT_BELOW(feature_belows[2192])) ac2192(.scan_win(scan_win2192), .scan_win_std_dev(scan_win_std_dev[2192]), .feature_accum(feature_accums[2192]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2193]), .RECT1_Y(rectangle1_ys[2193]), .RECT1_WIDTH(rectangle1_widths[2193]), .RECT1_HEIGHT(rectangle1_heights[2193]), .RECT1_WEIGHT(rectangle1_weights[2193]), .RECT2_X(rectangle2_xs[2193]), .RECT2_Y(rectangle2_ys[2193]), .RECT2_WIDTH(rectangle2_widths[2193]), .RECT2_HEIGHT(rectangle2_heights[2193]), .RECT2_WEIGHT(rectangle2_weights[2193]), .RECT3_X(rectangle3_xs[2193]), .RECT3_Y(rectangle3_ys[2193]), .RECT3_WIDTH(rectangle3_widths[2193]), .RECT3_HEIGHT(rectangle3_heights[2193]), .RECT3_WEIGHT(rectangle3_weights[2193]), .FEAT_THRES(feature_thresholds[2193]), .FEAT_ABOVE(feature_aboves[2193]), .FEAT_BELOW(feature_belows[2193])) ac2193(.scan_win(scan_win2193), .scan_win_std_dev(scan_win_std_dev[2193]), .feature_accum(feature_accums[2193]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2194]), .RECT1_Y(rectangle1_ys[2194]), .RECT1_WIDTH(rectangle1_widths[2194]), .RECT1_HEIGHT(rectangle1_heights[2194]), .RECT1_WEIGHT(rectangle1_weights[2194]), .RECT2_X(rectangle2_xs[2194]), .RECT2_Y(rectangle2_ys[2194]), .RECT2_WIDTH(rectangle2_widths[2194]), .RECT2_HEIGHT(rectangle2_heights[2194]), .RECT2_WEIGHT(rectangle2_weights[2194]), .RECT3_X(rectangle3_xs[2194]), .RECT3_Y(rectangle3_ys[2194]), .RECT3_WIDTH(rectangle3_widths[2194]), .RECT3_HEIGHT(rectangle3_heights[2194]), .RECT3_WEIGHT(rectangle3_weights[2194]), .FEAT_THRES(feature_thresholds[2194]), .FEAT_ABOVE(feature_aboves[2194]), .FEAT_BELOW(feature_belows[2194])) ac2194(.scan_win(scan_win2194), .scan_win_std_dev(scan_win_std_dev[2194]), .feature_accum(feature_accums[2194]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2195]), .RECT1_Y(rectangle1_ys[2195]), .RECT1_WIDTH(rectangle1_widths[2195]), .RECT1_HEIGHT(rectangle1_heights[2195]), .RECT1_WEIGHT(rectangle1_weights[2195]), .RECT2_X(rectangle2_xs[2195]), .RECT2_Y(rectangle2_ys[2195]), .RECT2_WIDTH(rectangle2_widths[2195]), .RECT2_HEIGHT(rectangle2_heights[2195]), .RECT2_WEIGHT(rectangle2_weights[2195]), .RECT3_X(rectangle3_xs[2195]), .RECT3_Y(rectangle3_ys[2195]), .RECT3_WIDTH(rectangle3_widths[2195]), .RECT3_HEIGHT(rectangle3_heights[2195]), .RECT3_WEIGHT(rectangle3_weights[2195]), .FEAT_THRES(feature_thresholds[2195]), .FEAT_ABOVE(feature_aboves[2195]), .FEAT_BELOW(feature_belows[2195])) ac2195(.scan_win(scan_win2195), .scan_win_std_dev(scan_win_std_dev[2195]), .feature_accum(feature_accums[2195]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2196]), .RECT1_Y(rectangle1_ys[2196]), .RECT1_WIDTH(rectangle1_widths[2196]), .RECT1_HEIGHT(rectangle1_heights[2196]), .RECT1_WEIGHT(rectangle1_weights[2196]), .RECT2_X(rectangle2_xs[2196]), .RECT2_Y(rectangle2_ys[2196]), .RECT2_WIDTH(rectangle2_widths[2196]), .RECT2_HEIGHT(rectangle2_heights[2196]), .RECT2_WEIGHT(rectangle2_weights[2196]), .RECT3_X(rectangle3_xs[2196]), .RECT3_Y(rectangle3_ys[2196]), .RECT3_WIDTH(rectangle3_widths[2196]), .RECT3_HEIGHT(rectangle3_heights[2196]), .RECT3_WEIGHT(rectangle3_weights[2196]), .FEAT_THRES(feature_thresholds[2196]), .FEAT_ABOVE(feature_aboves[2196]), .FEAT_BELOW(feature_belows[2196])) ac2196(.scan_win(scan_win2196), .scan_win_std_dev(scan_win_std_dev[2196]), .feature_accum(feature_accums[2196]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2197]), .RECT1_Y(rectangle1_ys[2197]), .RECT1_WIDTH(rectangle1_widths[2197]), .RECT1_HEIGHT(rectangle1_heights[2197]), .RECT1_WEIGHT(rectangle1_weights[2197]), .RECT2_X(rectangle2_xs[2197]), .RECT2_Y(rectangle2_ys[2197]), .RECT2_WIDTH(rectangle2_widths[2197]), .RECT2_HEIGHT(rectangle2_heights[2197]), .RECT2_WEIGHT(rectangle2_weights[2197]), .RECT3_X(rectangle3_xs[2197]), .RECT3_Y(rectangle3_ys[2197]), .RECT3_WIDTH(rectangle3_widths[2197]), .RECT3_HEIGHT(rectangle3_heights[2197]), .RECT3_WEIGHT(rectangle3_weights[2197]), .FEAT_THRES(feature_thresholds[2197]), .FEAT_ABOVE(feature_aboves[2197]), .FEAT_BELOW(feature_belows[2197])) ac2197(.scan_win(scan_win2197), .scan_win_std_dev(scan_win_std_dev[2197]), .feature_accum(feature_accums[2197]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2198]), .RECT1_Y(rectangle1_ys[2198]), .RECT1_WIDTH(rectangle1_widths[2198]), .RECT1_HEIGHT(rectangle1_heights[2198]), .RECT1_WEIGHT(rectangle1_weights[2198]), .RECT2_X(rectangle2_xs[2198]), .RECT2_Y(rectangle2_ys[2198]), .RECT2_WIDTH(rectangle2_widths[2198]), .RECT2_HEIGHT(rectangle2_heights[2198]), .RECT2_WEIGHT(rectangle2_weights[2198]), .RECT3_X(rectangle3_xs[2198]), .RECT3_Y(rectangle3_ys[2198]), .RECT3_WIDTH(rectangle3_widths[2198]), .RECT3_HEIGHT(rectangle3_heights[2198]), .RECT3_WEIGHT(rectangle3_weights[2198]), .FEAT_THRES(feature_thresholds[2198]), .FEAT_ABOVE(feature_aboves[2198]), .FEAT_BELOW(feature_belows[2198])) ac2198(.scan_win(scan_win2198), .scan_win_std_dev(scan_win_std_dev[2198]), .feature_accum(feature_accums[2198]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2199]), .RECT1_Y(rectangle1_ys[2199]), .RECT1_WIDTH(rectangle1_widths[2199]), .RECT1_HEIGHT(rectangle1_heights[2199]), .RECT1_WEIGHT(rectangle1_weights[2199]), .RECT2_X(rectangle2_xs[2199]), .RECT2_Y(rectangle2_ys[2199]), .RECT2_WIDTH(rectangle2_widths[2199]), .RECT2_HEIGHT(rectangle2_heights[2199]), .RECT2_WEIGHT(rectangle2_weights[2199]), .RECT3_X(rectangle3_xs[2199]), .RECT3_Y(rectangle3_ys[2199]), .RECT3_WIDTH(rectangle3_widths[2199]), .RECT3_HEIGHT(rectangle3_heights[2199]), .RECT3_WEIGHT(rectangle3_weights[2199]), .FEAT_THRES(feature_thresholds[2199]), .FEAT_ABOVE(feature_aboves[2199]), .FEAT_BELOW(feature_belows[2199])) ac2199(.scan_win(scan_win2199), .scan_win_std_dev(scan_win_std_dev[2199]), .feature_accum(feature_accums[2199]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2200]), .RECT1_Y(rectangle1_ys[2200]), .RECT1_WIDTH(rectangle1_widths[2200]), .RECT1_HEIGHT(rectangle1_heights[2200]), .RECT1_WEIGHT(rectangle1_weights[2200]), .RECT2_X(rectangle2_xs[2200]), .RECT2_Y(rectangle2_ys[2200]), .RECT2_WIDTH(rectangle2_widths[2200]), .RECT2_HEIGHT(rectangle2_heights[2200]), .RECT2_WEIGHT(rectangle2_weights[2200]), .RECT3_X(rectangle3_xs[2200]), .RECT3_Y(rectangle3_ys[2200]), .RECT3_WIDTH(rectangle3_widths[2200]), .RECT3_HEIGHT(rectangle3_heights[2200]), .RECT3_WEIGHT(rectangle3_weights[2200]), .FEAT_THRES(feature_thresholds[2200]), .FEAT_ABOVE(feature_aboves[2200]), .FEAT_BELOW(feature_belows[2200])) ac2200(.scan_win(scan_win2200), .scan_win_std_dev(scan_win_std_dev[2200]), .feature_accum(feature_accums[2200]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2201]), .RECT1_Y(rectangle1_ys[2201]), .RECT1_WIDTH(rectangle1_widths[2201]), .RECT1_HEIGHT(rectangle1_heights[2201]), .RECT1_WEIGHT(rectangle1_weights[2201]), .RECT2_X(rectangle2_xs[2201]), .RECT2_Y(rectangle2_ys[2201]), .RECT2_WIDTH(rectangle2_widths[2201]), .RECT2_HEIGHT(rectangle2_heights[2201]), .RECT2_WEIGHT(rectangle2_weights[2201]), .RECT3_X(rectangle3_xs[2201]), .RECT3_Y(rectangle3_ys[2201]), .RECT3_WIDTH(rectangle3_widths[2201]), .RECT3_HEIGHT(rectangle3_heights[2201]), .RECT3_WEIGHT(rectangle3_weights[2201]), .FEAT_THRES(feature_thresholds[2201]), .FEAT_ABOVE(feature_aboves[2201]), .FEAT_BELOW(feature_belows[2201])) ac2201(.scan_win(scan_win2201), .scan_win_std_dev(scan_win_std_dev[2201]), .feature_accum(feature_accums[2201]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2202]), .RECT1_Y(rectangle1_ys[2202]), .RECT1_WIDTH(rectangle1_widths[2202]), .RECT1_HEIGHT(rectangle1_heights[2202]), .RECT1_WEIGHT(rectangle1_weights[2202]), .RECT2_X(rectangle2_xs[2202]), .RECT2_Y(rectangle2_ys[2202]), .RECT2_WIDTH(rectangle2_widths[2202]), .RECT2_HEIGHT(rectangle2_heights[2202]), .RECT2_WEIGHT(rectangle2_weights[2202]), .RECT3_X(rectangle3_xs[2202]), .RECT3_Y(rectangle3_ys[2202]), .RECT3_WIDTH(rectangle3_widths[2202]), .RECT3_HEIGHT(rectangle3_heights[2202]), .RECT3_WEIGHT(rectangle3_weights[2202]), .FEAT_THRES(feature_thresholds[2202]), .FEAT_ABOVE(feature_aboves[2202]), .FEAT_BELOW(feature_belows[2202])) ac2202(.scan_win(scan_win2202), .scan_win_std_dev(scan_win_std_dev[2202]), .feature_accum(feature_accums[2202]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2203]), .RECT1_Y(rectangle1_ys[2203]), .RECT1_WIDTH(rectangle1_widths[2203]), .RECT1_HEIGHT(rectangle1_heights[2203]), .RECT1_WEIGHT(rectangle1_weights[2203]), .RECT2_X(rectangle2_xs[2203]), .RECT2_Y(rectangle2_ys[2203]), .RECT2_WIDTH(rectangle2_widths[2203]), .RECT2_HEIGHT(rectangle2_heights[2203]), .RECT2_WEIGHT(rectangle2_weights[2203]), .RECT3_X(rectangle3_xs[2203]), .RECT3_Y(rectangle3_ys[2203]), .RECT3_WIDTH(rectangle3_widths[2203]), .RECT3_HEIGHT(rectangle3_heights[2203]), .RECT3_WEIGHT(rectangle3_weights[2203]), .FEAT_THRES(feature_thresholds[2203]), .FEAT_ABOVE(feature_aboves[2203]), .FEAT_BELOW(feature_belows[2203])) ac2203(.scan_win(scan_win2203), .scan_win_std_dev(scan_win_std_dev[2203]), .feature_accum(feature_accums[2203]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2204]), .RECT1_Y(rectangle1_ys[2204]), .RECT1_WIDTH(rectangle1_widths[2204]), .RECT1_HEIGHT(rectangle1_heights[2204]), .RECT1_WEIGHT(rectangle1_weights[2204]), .RECT2_X(rectangle2_xs[2204]), .RECT2_Y(rectangle2_ys[2204]), .RECT2_WIDTH(rectangle2_widths[2204]), .RECT2_HEIGHT(rectangle2_heights[2204]), .RECT2_WEIGHT(rectangle2_weights[2204]), .RECT3_X(rectangle3_xs[2204]), .RECT3_Y(rectangle3_ys[2204]), .RECT3_WIDTH(rectangle3_widths[2204]), .RECT3_HEIGHT(rectangle3_heights[2204]), .RECT3_WEIGHT(rectangle3_weights[2204]), .FEAT_THRES(feature_thresholds[2204]), .FEAT_ABOVE(feature_aboves[2204]), .FEAT_BELOW(feature_belows[2204])) ac2204(.scan_win(scan_win2204), .scan_win_std_dev(scan_win_std_dev[2204]), .feature_accum(feature_accums[2204]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2205]), .RECT1_Y(rectangle1_ys[2205]), .RECT1_WIDTH(rectangle1_widths[2205]), .RECT1_HEIGHT(rectangle1_heights[2205]), .RECT1_WEIGHT(rectangle1_weights[2205]), .RECT2_X(rectangle2_xs[2205]), .RECT2_Y(rectangle2_ys[2205]), .RECT2_WIDTH(rectangle2_widths[2205]), .RECT2_HEIGHT(rectangle2_heights[2205]), .RECT2_WEIGHT(rectangle2_weights[2205]), .RECT3_X(rectangle3_xs[2205]), .RECT3_Y(rectangle3_ys[2205]), .RECT3_WIDTH(rectangle3_widths[2205]), .RECT3_HEIGHT(rectangle3_heights[2205]), .RECT3_WEIGHT(rectangle3_weights[2205]), .FEAT_THRES(feature_thresholds[2205]), .FEAT_ABOVE(feature_aboves[2205]), .FEAT_BELOW(feature_belows[2205])) ac2205(.scan_win(scan_win2205), .scan_win_std_dev(scan_win_std_dev[2205]), .feature_accum(feature_accums[2205]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2206]), .RECT1_Y(rectangle1_ys[2206]), .RECT1_WIDTH(rectangle1_widths[2206]), .RECT1_HEIGHT(rectangle1_heights[2206]), .RECT1_WEIGHT(rectangle1_weights[2206]), .RECT2_X(rectangle2_xs[2206]), .RECT2_Y(rectangle2_ys[2206]), .RECT2_WIDTH(rectangle2_widths[2206]), .RECT2_HEIGHT(rectangle2_heights[2206]), .RECT2_WEIGHT(rectangle2_weights[2206]), .RECT3_X(rectangle3_xs[2206]), .RECT3_Y(rectangle3_ys[2206]), .RECT3_WIDTH(rectangle3_widths[2206]), .RECT3_HEIGHT(rectangle3_heights[2206]), .RECT3_WEIGHT(rectangle3_weights[2206]), .FEAT_THRES(feature_thresholds[2206]), .FEAT_ABOVE(feature_aboves[2206]), .FEAT_BELOW(feature_belows[2206])) ac2206(.scan_win(scan_win2206), .scan_win_std_dev(scan_win_std_dev[2206]), .feature_accum(feature_accums[2206]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2207]), .RECT1_Y(rectangle1_ys[2207]), .RECT1_WIDTH(rectangle1_widths[2207]), .RECT1_HEIGHT(rectangle1_heights[2207]), .RECT1_WEIGHT(rectangle1_weights[2207]), .RECT2_X(rectangle2_xs[2207]), .RECT2_Y(rectangle2_ys[2207]), .RECT2_WIDTH(rectangle2_widths[2207]), .RECT2_HEIGHT(rectangle2_heights[2207]), .RECT2_WEIGHT(rectangle2_weights[2207]), .RECT3_X(rectangle3_xs[2207]), .RECT3_Y(rectangle3_ys[2207]), .RECT3_WIDTH(rectangle3_widths[2207]), .RECT3_HEIGHT(rectangle3_heights[2207]), .RECT3_WEIGHT(rectangle3_weights[2207]), .FEAT_THRES(feature_thresholds[2207]), .FEAT_ABOVE(feature_aboves[2207]), .FEAT_BELOW(feature_belows[2207])) ac2207(.scan_win(scan_win2207), .scan_win_std_dev(scan_win_std_dev[2207]), .feature_accum(feature_accums[2207]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2208]), .RECT1_Y(rectangle1_ys[2208]), .RECT1_WIDTH(rectangle1_widths[2208]), .RECT1_HEIGHT(rectangle1_heights[2208]), .RECT1_WEIGHT(rectangle1_weights[2208]), .RECT2_X(rectangle2_xs[2208]), .RECT2_Y(rectangle2_ys[2208]), .RECT2_WIDTH(rectangle2_widths[2208]), .RECT2_HEIGHT(rectangle2_heights[2208]), .RECT2_WEIGHT(rectangle2_weights[2208]), .RECT3_X(rectangle3_xs[2208]), .RECT3_Y(rectangle3_ys[2208]), .RECT3_WIDTH(rectangle3_widths[2208]), .RECT3_HEIGHT(rectangle3_heights[2208]), .RECT3_WEIGHT(rectangle3_weights[2208]), .FEAT_THRES(feature_thresholds[2208]), .FEAT_ABOVE(feature_aboves[2208]), .FEAT_BELOW(feature_belows[2208])) ac2208(.scan_win(scan_win2208), .scan_win_std_dev(scan_win_std_dev[2208]), .feature_accum(feature_accums[2208]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2209]), .RECT1_Y(rectangle1_ys[2209]), .RECT1_WIDTH(rectangle1_widths[2209]), .RECT1_HEIGHT(rectangle1_heights[2209]), .RECT1_WEIGHT(rectangle1_weights[2209]), .RECT2_X(rectangle2_xs[2209]), .RECT2_Y(rectangle2_ys[2209]), .RECT2_WIDTH(rectangle2_widths[2209]), .RECT2_HEIGHT(rectangle2_heights[2209]), .RECT2_WEIGHT(rectangle2_weights[2209]), .RECT3_X(rectangle3_xs[2209]), .RECT3_Y(rectangle3_ys[2209]), .RECT3_WIDTH(rectangle3_widths[2209]), .RECT3_HEIGHT(rectangle3_heights[2209]), .RECT3_WEIGHT(rectangle3_weights[2209]), .FEAT_THRES(feature_thresholds[2209]), .FEAT_ABOVE(feature_aboves[2209]), .FEAT_BELOW(feature_belows[2209])) ac2209(.scan_win(scan_win2209), .scan_win_std_dev(scan_win_std_dev[2209]), .feature_accum(feature_accums[2209]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2210]), .RECT1_Y(rectangle1_ys[2210]), .RECT1_WIDTH(rectangle1_widths[2210]), .RECT1_HEIGHT(rectangle1_heights[2210]), .RECT1_WEIGHT(rectangle1_weights[2210]), .RECT2_X(rectangle2_xs[2210]), .RECT2_Y(rectangle2_ys[2210]), .RECT2_WIDTH(rectangle2_widths[2210]), .RECT2_HEIGHT(rectangle2_heights[2210]), .RECT2_WEIGHT(rectangle2_weights[2210]), .RECT3_X(rectangle3_xs[2210]), .RECT3_Y(rectangle3_ys[2210]), .RECT3_WIDTH(rectangle3_widths[2210]), .RECT3_HEIGHT(rectangle3_heights[2210]), .RECT3_WEIGHT(rectangle3_weights[2210]), .FEAT_THRES(feature_thresholds[2210]), .FEAT_ABOVE(feature_aboves[2210]), .FEAT_BELOW(feature_belows[2210])) ac2210(.scan_win(scan_win2210), .scan_win_std_dev(scan_win_std_dev[2210]), .feature_accum(feature_accums[2210]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2211]), .RECT1_Y(rectangle1_ys[2211]), .RECT1_WIDTH(rectangle1_widths[2211]), .RECT1_HEIGHT(rectangle1_heights[2211]), .RECT1_WEIGHT(rectangle1_weights[2211]), .RECT2_X(rectangle2_xs[2211]), .RECT2_Y(rectangle2_ys[2211]), .RECT2_WIDTH(rectangle2_widths[2211]), .RECT2_HEIGHT(rectangle2_heights[2211]), .RECT2_WEIGHT(rectangle2_weights[2211]), .RECT3_X(rectangle3_xs[2211]), .RECT3_Y(rectangle3_ys[2211]), .RECT3_WIDTH(rectangle3_widths[2211]), .RECT3_HEIGHT(rectangle3_heights[2211]), .RECT3_WEIGHT(rectangle3_weights[2211]), .FEAT_THRES(feature_thresholds[2211]), .FEAT_ABOVE(feature_aboves[2211]), .FEAT_BELOW(feature_belows[2211])) ac2211(.scan_win(scan_win2211), .scan_win_std_dev(scan_win_std_dev[2211]), .feature_accum(feature_accums[2211]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2212]), .RECT1_Y(rectangle1_ys[2212]), .RECT1_WIDTH(rectangle1_widths[2212]), .RECT1_HEIGHT(rectangle1_heights[2212]), .RECT1_WEIGHT(rectangle1_weights[2212]), .RECT2_X(rectangle2_xs[2212]), .RECT2_Y(rectangle2_ys[2212]), .RECT2_WIDTH(rectangle2_widths[2212]), .RECT2_HEIGHT(rectangle2_heights[2212]), .RECT2_WEIGHT(rectangle2_weights[2212]), .RECT3_X(rectangle3_xs[2212]), .RECT3_Y(rectangle3_ys[2212]), .RECT3_WIDTH(rectangle3_widths[2212]), .RECT3_HEIGHT(rectangle3_heights[2212]), .RECT3_WEIGHT(rectangle3_weights[2212]), .FEAT_THRES(feature_thresholds[2212]), .FEAT_ABOVE(feature_aboves[2212]), .FEAT_BELOW(feature_belows[2212])) ac2212(.scan_win(scan_win2212), .scan_win_std_dev(scan_win_std_dev[2212]), .feature_accum(feature_accums[2212]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2213]), .RECT1_Y(rectangle1_ys[2213]), .RECT1_WIDTH(rectangle1_widths[2213]), .RECT1_HEIGHT(rectangle1_heights[2213]), .RECT1_WEIGHT(rectangle1_weights[2213]), .RECT2_X(rectangle2_xs[2213]), .RECT2_Y(rectangle2_ys[2213]), .RECT2_WIDTH(rectangle2_widths[2213]), .RECT2_HEIGHT(rectangle2_heights[2213]), .RECT2_WEIGHT(rectangle2_weights[2213]), .RECT3_X(rectangle3_xs[2213]), .RECT3_Y(rectangle3_ys[2213]), .RECT3_WIDTH(rectangle3_widths[2213]), .RECT3_HEIGHT(rectangle3_heights[2213]), .RECT3_WEIGHT(rectangle3_weights[2213]), .FEAT_THRES(feature_thresholds[2213]), .FEAT_ABOVE(feature_aboves[2213]), .FEAT_BELOW(feature_belows[2213])) ac2213(.scan_win(scan_win2213), .scan_win_std_dev(scan_win_std_dev[2213]), .feature_accum(feature_accums[2213]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2214]), .RECT1_Y(rectangle1_ys[2214]), .RECT1_WIDTH(rectangle1_widths[2214]), .RECT1_HEIGHT(rectangle1_heights[2214]), .RECT1_WEIGHT(rectangle1_weights[2214]), .RECT2_X(rectangle2_xs[2214]), .RECT2_Y(rectangle2_ys[2214]), .RECT2_WIDTH(rectangle2_widths[2214]), .RECT2_HEIGHT(rectangle2_heights[2214]), .RECT2_WEIGHT(rectangle2_weights[2214]), .RECT3_X(rectangle3_xs[2214]), .RECT3_Y(rectangle3_ys[2214]), .RECT3_WIDTH(rectangle3_widths[2214]), .RECT3_HEIGHT(rectangle3_heights[2214]), .RECT3_WEIGHT(rectangle3_weights[2214]), .FEAT_THRES(feature_thresholds[2214]), .FEAT_ABOVE(feature_aboves[2214]), .FEAT_BELOW(feature_belows[2214])) ac2214(.scan_win(scan_win2214), .scan_win_std_dev(scan_win_std_dev[2214]), .feature_accum(feature_accums[2214]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2215]), .RECT1_Y(rectangle1_ys[2215]), .RECT1_WIDTH(rectangle1_widths[2215]), .RECT1_HEIGHT(rectangle1_heights[2215]), .RECT1_WEIGHT(rectangle1_weights[2215]), .RECT2_X(rectangle2_xs[2215]), .RECT2_Y(rectangle2_ys[2215]), .RECT2_WIDTH(rectangle2_widths[2215]), .RECT2_HEIGHT(rectangle2_heights[2215]), .RECT2_WEIGHT(rectangle2_weights[2215]), .RECT3_X(rectangle3_xs[2215]), .RECT3_Y(rectangle3_ys[2215]), .RECT3_WIDTH(rectangle3_widths[2215]), .RECT3_HEIGHT(rectangle3_heights[2215]), .RECT3_WEIGHT(rectangle3_weights[2215]), .FEAT_THRES(feature_thresholds[2215]), .FEAT_ABOVE(feature_aboves[2215]), .FEAT_BELOW(feature_belows[2215])) ac2215(.scan_win(scan_win2215), .scan_win_std_dev(scan_win_std_dev[2215]), .feature_accum(feature_accums[2215]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2216]), .RECT1_Y(rectangle1_ys[2216]), .RECT1_WIDTH(rectangle1_widths[2216]), .RECT1_HEIGHT(rectangle1_heights[2216]), .RECT1_WEIGHT(rectangle1_weights[2216]), .RECT2_X(rectangle2_xs[2216]), .RECT2_Y(rectangle2_ys[2216]), .RECT2_WIDTH(rectangle2_widths[2216]), .RECT2_HEIGHT(rectangle2_heights[2216]), .RECT2_WEIGHT(rectangle2_weights[2216]), .RECT3_X(rectangle3_xs[2216]), .RECT3_Y(rectangle3_ys[2216]), .RECT3_WIDTH(rectangle3_widths[2216]), .RECT3_HEIGHT(rectangle3_heights[2216]), .RECT3_WEIGHT(rectangle3_weights[2216]), .FEAT_THRES(feature_thresholds[2216]), .FEAT_ABOVE(feature_aboves[2216]), .FEAT_BELOW(feature_belows[2216])) ac2216(.scan_win(scan_win2216), .scan_win_std_dev(scan_win_std_dev[2216]), .feature_accum(feature_accums[2216]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2217]), .RECT1_Y(rectangle1_ys[2217]), .RECT1_WIDTH(rectangle1_widths[2217]), .RECT1_HEIGHT(rectangle1_heights[2217]), .RECT1_WEIGHT(rectangle1_weights[2217]), .RECT2_X(rectangle2_xs[2217]), .RECT2_Y(rectangle2_ys[2217]), .RECT2_WIDTH(rectangle2_widths[2217]), .RECT2_HEIGHT(rectangle2_heights[2217]), .RECT2_WEIGHT(rectangle2_weights[2217]), .RECT3_X(rectangle3_xs[2217]), .RECT3_Y(rectangle3_ys[2217]), .RECT3_WIDTH(rectangle3_widths[2217]), .RECT3_HEIGHT(rectangle3_heights[2217]), .RECT3_WEIGHT(rectangle3_weights[2217]), .FEAT_THRES(feature_thresholds[2217]), .FEAT_ABOVE(feature_aboves[2217]), .FEAT_BELOW(feature_belows[2217])) ac2217(.scan_win(scan_win2217), .scan_win_std_dev(scan_win_std_dev[2217]), .feature_accum(feature_accums[2217]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2218]), .RECT1_Y(rectangle1_ys[2218]), .RECT1_WIDTH(rectangle1_widths[2218]), .RECT1_HEIGHT(rectangle1_heights[2218]), .RECT1_WEIGHT(rectangle1_weights[2218]), .RECT2_X(rectangle2_xs[2218]), .RECT2_Y(rectangle2_ys[2218]), .RECT2_WIDTH(rectangle2_widths[2218]), .RECT2_HEIGHT(rectangle2_heights[2218]), .RECT2_WEIGHT(rectangle2_weights[2218]), .RECT3_X(rectangle3_xs[2218]), .RECT3_Y(rectangle3_ys[2218]), .RECT3_WIDTH(rectangle3_widths[2218]), .RECT3_HEIGHT(rectangle3_heights[2218]), .RECT3_WEIGHT(rectangle3_weights[2218]), .FEAT_THRES(feature_thresholds[2218]), .FEAT_ABOVE(feature_aboves[2218]), .FEAT_BELOW(feature_belows[2218])) ac2218(.scan_win(scan_win2218), .scan_win_std_dev(scan_win_std_dev[2218]), .feature_accum(feature_accums[2218]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2219]), .RECT1_Y(rectangle1_ys[2219]), .RECT1_WIDTH(rectangle1_widths[2219]), .RECT1_HEIGHT(rectangle1_heights[2219]), .RECT1_WEIGHT(rectangle1_weights[2219]), .RECT2_X(rectangle2_xs[2219]), .RECT2_Y(rectangle2_ys[2219]), .RECT2_WIDTH(rectangle2_widths[2219]), .RECT2_HEIGHT(rectangle2_heights[2219]), .RECT2_WEIGHT(rectangle2_weights[2219]), .RECT3_X(rectangle3_xs[2219]), .RECT3_Y(rectangle3_ys[2219]), .RECT3_WIDTH(rectangle3_widths[2219]), .RECT3_HEIGHT(rectangle3_heights[2219]), .RECT3_WEIGHT(rectangle3_weights[2219]), .FEAT_THRES(feature_thresholds[2219]), .FEAT_ABOVE(feature_aboves[2219]), .FEAT_BELOW(feature_belows[2219])) ac2219(.scan_win(scan_win2219), .scan_win_std_dev(scan_win_std_dev[2219]), .feature_accum(feature_accums[2219]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2220]), .RECT1_Y(rectangle1_ys[2220]), .RECT1_WIDTH(rectangle1_widths[2220]), .RECT1_HEIGHT(rectangle1_heights[2220]), .RECT1_WEIGHT(rectangle1_weights[2220]), .RECT2_X(rectangle2_xs[2220]), .RECT2_Y(rectangle2_ys[2220]), .RECT2_WIDTH(rectangle2_widths[2220]), .RECT2_HEIGHT(rectangle2_heights[2220]), .RECT2_WEIGHT(rectangle2_weights[2220]), .RECT3_X(rectangle3_xs[2220]), .RECT3_Y(rectangle3_ys[2220]), .RECT3_WIDTH(rectangle3_widths[2220]), .RECT3_HEIGHT(rectangle3_heights[2220]), .RECT3_WEIGHT(rectangle3_weights[2220]), .FEAT_THRES(feature_thresholds[2220]), .FEAT_ABOVE(feature_aboves[2220]), .FEAT_BELOW(feature_belows[2220])) ac2220(.scan_win(scan_win2220), .scan_win_std_dev(scan_win_std_dev[2220]), .feature_accum(feature_accums[2220]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2221]), .RECT1_Y(rectangle1_ys[2221]), .RECT1_WIDTH(rectangle1_widths[2221]), .RECT1_HEIGHT(rectangle1_heights[2221]), .RECT1_WEIGHT(rectangle1_weights[2221]), .RECT2_X(rectangle2_xs[2221]), .RECT2_Y(rectangle2_ys[2221]), .RECT2_WIDTH(rectangle2_widths[2221]), .RECT2_HEIGHT(rectangle2_heights[2221]), .RECT2_WEIGHT(rectangle2_weights[2221]), .RECT3_X(rectangle3_xs[2221]), .RECT3_Y(rectangle3_ys[2221]), .RECT3_WIDTH(rectangle3_widths[2221]), .RECT3_HEIGHT(rectangle3_heights[2221]), .RECT3_WEIGHT(rectangle3_weights[2221]), .FEAT_THRES(feature_thresholds[2221]), .FEAT_ABOVE(feature_aboves[2221]), .FEAT_BELOW(feature_belows[2221])) ac2221(.scan_win(scan_win2221), .scan_win_std_dev(scan_win_std_dev[2221]), .feature_accum(feature_accums[2221]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2222]), .RECT1_Y(rectangle1_ys[2222]), .RECT1_WIDTH(rectangle1_widths[2222]), .RECT1_HEIGHT(rectangle1_heights[2222]), .RECT1_WEIGHT(rectangle1_weights[2222]), .RECT2_X(rectangle2_xs[2222]), .RECT2_Y(rectangle2_ys[2222]), .RECT2_WIDTH(rectangle2_widths[2222]), .RECT2_HEIGHT(rectangle2_heights[2222]), .RECT2_WEIGHT(rectangle2_weights[2222]), .RECT3_X(rectangle3_xs[2222]), .RECT3_Y(rectangle3_ys[2222]), .RECT3_WIDTH(rectangle3_widths[2222]), .RECT3_HEIGHT(rectangle3_heights[2222]), .RECT3_WEIGHT(rectangle3_weights[2222]), .FEAT_THRES(feature_thresholds[2222]), .FEAT_ABOVE(feature_aboves[2222]), .FEAT_BELOW(feature_belows[2222])) ac2222(.scan_win(scan_win2222), .scan_win_std_dev(scan_win_std_dev[2222]), .feature_accum(feature_accums[2222]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2223]), .RECT1_Y(rectangle1_ys[2223]), .RECT1_WIDTH(rectangle1_widths[2223]), .RECT1_HEIGHT(rectangle1_heights[2223]), .RECT1_WEIGHT(rectangle1_weights[2223]), .RECT2_X(rectangle2_xs[2223]), .RECT2_Y(rectangle2_ys[2223]), .RECT2_WIDTH(rectangle2_widths[2223]), .RECT2_HEIGHT(rectangle2_heights[2223]), .RECT2_WEIGHT(rectangle2_weights[2223]), .RECT3_X(rectangle3_xs[2223]), .RECT3_Y(rectangle3_ys[2223]), .RECT3_WIDTH(rectangle3_widths[2223]), .RECT3_HEIGHT(rectangle3_heights[2223]), .RECT3_WEIGHT(rectangle3_weights[2223]), .FEAT_THRES(feature_thresholds[2223]), .FEAT_ABOVE(feature_aboves[2223]), .FEAT_BELOW(feature_belows[2223])) ac2223(.scan_win(scan_win2223), .scan_win_std_dev(scan_win_std_dev[2223]), .feature_accum(feature_accums[2223]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2224]), .RECT1_Y(rectangle1_ys[2224]), .RECT1_WIDTH(rectangle1_widths[2224]), .RECT1_HEIGHT(rectangle1_heights[2224]), .RECT1_WEIGHT(rectangle1_weights[2224]), .RECT2_X(rectangle2_xs[2224]), .RECT2_Y(rectangle2_ys[2224]), .RECT2_WIDTH(rectangle2_widths[2224]), .RECT2_HEIGHT(rectangle2_heights[2224]), .RECT2_WEIGHT(rectangle2_weights[2224]), .RECT3_X(rectangle3_xs[2224]), .RECT3_Y(rectangle3_ys[2224]), .RECT3_WIDTH(rectangle3_widths[2224]), .RECT3_HEIGHT(rectangle3_heights[2224]), .RECT3_WEIGHT(rectangle3_weights[2224]), .FEAT_THRES(feature_thresholds[2224]), .FEAT_ABOVE(feature_aboves[2224]), .FEAT_BELOW(feature_belows[2224])) ac2224(.scan_win(scan_win2224), .scan_win_std_dev(scan_win_std_dev[2224]), .feature_accum(feature_accums[2224]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2225]), .RECT1_Y(rectangle1_ys[2225]), .RECT1_WIDTH(rectangle1_widths[2225]), .RECT1_HEIGHT(rectangle1_heights[2225]), .RECT1_WEIGHT(rectangle1_weights[2225]), .RECT2_X(rectangle2_xs[2225]), .RECT2_Y(rectangle2_ys[2225]), .RECT2_WIDTH(rectangle2_widths[2225]), .RECT2_HEIGHT(rectangle2_heights[2225]), .RECT2_WEIGHT(rectangle2_weights[2225]), .RECT3_X(rectangle3_xs[2225]), .RECT3_Y(rectangle3_ys[2225]), .RECT3_WIDTH(rectangle3_widths[2225]), .RECT3_HEIGHT(rectangle3_heights[2225]), .RECT3_WEIGHT(rectangle3_weights[2225]), .FEAT_THRES(feature_thresholds[2225]), .FEAT_ABOVE(feature_aboves[2225]), .FEAT_BELOW(feature_belows[2225])) ac2225(.scan_win(scan_win2225), .scan_win_std_dev(scan_win_std_dev[2225]), .feature_accum(feature_accums[2225]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2226]), .RECT1_Y(rectangle1_ys[2226]), .RECT1_WIDTH(rectangle1_widths[2226]), .RECT1_HEIGHT(rectangle1_heights[2226]), .RECT1_WEIGHT(rectangle1_weights[2226]), .RECT2_X(rectangle2_xs[2226]), .RECT2_Y(rectangle2_ys[2226]), .RECT2_WIDTH(rectangle2_widths[2226]), .RECT2_HEIGHT(rectangle2_heights[2226]), .RECT2_WEIGHT(rectangle2_weights[2226]), .RECT3_X(rectangle3_xs[2226]), .RECT3_Y(rectangle3_ys[2226]), .RECT3_WIDTH(rectangle3_widths[2226]), .RECT3_HEIGHT(rectangle3_heights[2226]), .RECT3_WEIGHT(rectangle3_weights[2226]), .FEAT_THRES(feature_thresholds[2226]), .FEAT_ABOVE(feature_aboves[2226]), .FEAT_BELOW(feature_belows[2226])) ac2226(.scan_win(scan_win2226), .scan_win_std_dev(scan_win_std_dev[2226]), .feature_accum(feature_accums[2226]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2227]), .RECT1_Y(rectangle1_ys[2227]), .RECT1_WIDTH(rectangle1_widths[2227]), .RECT1_HEIGHT(rectangle1_heights[2227]), .RECT1_WEIGHT(rectangle1_weights[2227]), .RECT2_X(rectangle2_xs[2227]), .RECT2_Y(rectangle2_ys[2227]), .RECT2_WIDTH(rectangle2_widths[2227]), .RECT2_HEIGHT(rectangle2_heights[2227]), .RECT2_WEIGHT(rectangle2_weights[2227]), .RECT3_X(rectangle3_xs[2227]), .RECT3_Y(rectangle3_ys[2227]), .RECT3_WIDTH(rectangle3_widths[2227]), .RECT3_HEIGHT(rectangle3_heights[2227]), .RECT3_WEIGHT(rectangle3_weights[2227]), .FEAT_THRES(feature_thresholds[2227]), .FEAT_ABOVE(feature_aboves[2227]), .FEAT_BELOW(feature_belows[2227])) ac2227(.scan_win(scan_win2227), .scan_win_std_dev(scan_win_std_dev[2227]), .feature_accum(feature_accums[2227]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2228]), .RECT1_Y(rectangle1_ys[2228]), .RECT1_WIDTH(rectangle1_widths[2228]), .RECT1_HEIGHT(rectangle1_heights[2228]), .RECT1_WEIGHT(rectangle1_weights[2228]), .RECT2_X(rectangle2_xs[2228]), .RECT2_Y(rectangle2_ys[2228]), .RECT2_WIDTH(rectangle2_widths[2228]), .RECT2_HEIGHT(rectangle2_heights[2228]), .RECT2_WEIGHT(rectangle2_weights[2228]), .RECT3_X(rectangle3_xs[2228]), .RECT3_Y(rectangle3_ys[2228]), .RECT3_WIDTH(rectangle3_widths[2228]), .RECT3_HEIGHT(rectangle3_heights[2228]), .RECT3_WEIGHT(rectangle3_weights[2228]), .FEAT_THRES(feature_thresholds[2228]), .FEAT_ABOVE(feature_aboves[2228]), .FEAT_BELOW(feature_belows[2228])) ac2228(.scan_win(scan_win2228), .scan_win_std_dev(scan_win_std_dev[2228]), .feature_accum(feature_accums[2228]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2229]), .RECT1_Y(rectangle1_ys[2229]), .RECT1_WIDTH(rectangle1_widths[2229]), .RECT1_HEIGHT(rectangle1_heights[2229]), .RECT1_WEIGHT(rectangle1_weights[2229]), .RECT2_X(rectangle2_xs[2229]), .RECT2_Y(rectangle2_ys[2229]), .RECT2_WIDTH(rectangle2_widths[2229]), .RECT2_HEIGHT(rectangle2_heights[2229]), .RECT2_WEIGHT(rectangle2_weights[2229]), .RECT3_X(rectangle3_xs[2229]), .RECT3_Y(rectangle3_ys[2229]), .RECT3_WIDTH(rectangle3_widths[2229]), .RECT3_HEIGHT(rectangle3_heights[2229]), .RECT3_WEIGHT(rectangle3_weights[2229]), .FEAT_THRES(feature_thresholds[2229]), .FEAT_ABOVE(feature_aboves[2229]), .FEAT_BELOW(feature_belows[2229])) ac2229(.scan_win(scan_win2229), .scan_win_std_dev(scan_win_std_dev[2229]), .feature_accum(feature_accums[2229]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2230]), .RECT1_Y(rectangle1_ys[2230]), .RECT1_WIDTH(rectangle1_widths[2230]), .RECT1_HEIGHT(rectangle1_heights[2230]), .RECT1_WEIGHT(rectangle1_weights[2230]), .RECT2_X(rectangle2_xs[2230]), .RECT2_Y(rectangle2_ys[2230]), .RECT2_WIDTH(rectangle2_widths[2230]), .RECT2_HEIGHT(rectangle2_heights[2230]), .RECT2_WEIGHT(rectangle2_weights[2230]), .RECT3_X(rectangle3_xs[2230]), .RECT3_Y(rectangle3_ys[2230]), .RECT3_WIDTH(rectangle3_widths[2230]), .RECT3_HEIGHT(rectangle3_heights[2230]), .RECT3_WEIGHT(rectangle3_weights[2230]), .FEAT_THRES(feature_thresholds[2230]), .FEAT_ABOVE(feature_aboves[2230]), .FEAT_BELOW(feature_belows[2230])) ac2230(.scan_win(scan_win2230), .scan_win_std_dev(scan_win_std_dev[2230]), .feature_accum(feature_accums[2230]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2231]), .RECT1_Y(rectangle1_ys[2231]), .RECT1_WIDTH(rectangle1_widths[2231]), .RECT1_HEIGHT(rectangle1_heights[2231]), .RECT1_WEIGHT(rectangle1_weights[2231]), .RECT2_X(rectangle2_xs[2231]), .RECT2_Y(rectangle2_ys[2231]), .RECT2_WIDTH(rectangle2_widths[2231]), .RECT2_HEIGHT(rectangle2_heights[2231]), .RECT2_WEIGHT(rectangle2_weights[2231]), .RECT3_X(rectangle3_xs[2231]), .RECT3_Y(rectangle3_ys[2231]), .RECT3_WIDTH(rectangle3_widths[2231]), .RECT3_HEIGHT(rectangle3_heights[2231]), .RECT3_WEIGHT(rectangle3_weights[2231]), .FEAT_THRES(feature_thresholds[2231]), .FEAT_ABOVE(feature_aboves[2231]), .FEAT_BELOW(feature_belows[2231])) ac2231(.scan_win(scan_win2231), .scan_win_std_dev(scan_win_std_dev[2231]), .feature_accum(feature_accums[2231]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2232]), .RECT1_Y(rectangle1_ys[2232]), .RECT1_WIDTH(rectangle1_widths[2232]), .RECT1_HEIGHT(rectangle1_heights[2232]), .RECT1_WEIGHT(rectangle1_weights[2232]), .RECT2_X(rectangle2_xs[2232]), .RECT2_Y(rectangle2_ys[2232]), .RECT2_WIDTH(rectangle2_widths[2232]), .RECT2_HEIGHT(rectangle2_heights[2232]), .RECT2_WEIGHT(rectangle2_weights[2232]), .RECT3_X(rectangle3_xs[2232]), .RECT3_Y(rectangle3_ys[2232]), .RECT3_WIDTH(rectangle3_widths[2232]), .RECT3_HEIGHT(rectangle3_heights[2232]), .RECT3_WEIGHT(rectangle3_weights[2232]), .FEAT_THRES(feature_thresholds[2232]), .FEAT_ABOVE(feature_aboves[2232]), .FEAT_BELOW(feature_belows[2232])) ac2232(.scan_win(scan_win2232), .scan_win_std_dev(scan_win_std_dev[2232]), .feature_accum(feature_accums[2232]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2233]), .RECT1_Y(rectangle1_ys[2233]), .RECT1_WIDTH(rectangle1_widths[2233]), .RECT1_HEIGHT(rectangle1_heights[2233]), .RECT1_WEIGHT(rectangle1_weights[2233]), .RECT2_X(rectangle2_xs[2233]), .RECT2_Y(rectangle2_ys[2233]), .RECT2_WIDTH(rectangle2_widths[2233]), .RECT2_HEIGHT(rectangle2_heights[2233]), .RECT2_WEIGHT(rectangle2_weights[2233]), .RECT3_X(rectangle3_xs[2233]), .RECT3_Y(rectangle3_ys[2233]), .RECT3_WIDTH(rectangle3_widths[2233]), .RECT3_HEIGHT(rectangle3_heights[2233]), .RECT3_WEIGHT(rectangle3_weights[2233]), .FEAT_THRES(feature_thresholds[2233]), .FEAT_ABOVE(feature_aboves[2233]), .FEAT_BELOW(feature_belows[2233])) ac2233(.scan_win(scan_win2233), .scan_win_std_dev(scan_win_std_dev[2233]), .feature_accum(feature_accums[2233]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2234]), .RECT1_Y(rectangle1_ys[2234]), .RECT1_WIDTH(rectangle1_widths[2234]), .RECT1_HEIGHT(rectangle1_heights[2234]), .RECT1_WEIGHT(rectangle1_weights[2234]), .RECT2_X(rectangle2_xs[2234]), .RECT2_Y(rectangle2_ys[2234]), .RECT2_WIDTH(rectangle2_widths[2234]), .RECT2_HEIGHT(rectangle2_heights[2234]), .RECT2_WEIGHT(rectangle2_weights[2234]), .RECT3_X(rectangle3_xs[2234]), .RECT3_Y(rectangle3_ys[2234]), .RECT3_WIDTH(rectangle3_widths[2234]), .RECT3_HEIGHT(rectangle3_heights[2234]), .RECT3_WEIGHT(rectangle3_weights[2234]), .FEAT_THRES(feature_thresholds[2234]), .FEAT_ABOVE(feature_aboves[2234]), .FEAT_BELOW(feature_belows[2234])) ac2234(.scan_win(scan_win2234), .scan_win_std_dev(scan_win_std_dev[2234]), .feature_accum(feature_accums[2234]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2235]), .RECT1_Y(rectangle1_ys[2235]), .RECT1_WIDTH(rectangle1_widths[2235]), .RECT1_HEIGHT(rectangle1_heights[2235]), .RECT1_WEIGHT(rectangle1_weights[2235]), .RECT2_X(rectangle2_xs[2235]), .RECT2_Y(rectangle2_ys[2235]), .RECT2_WIDTH(rectangle2_widths[2235]), .RECT2_HEIGHT(rectangle2_heights[2235]), .RECT2_WEIGHT(rectangle2_weights[2235]), .RECT3_X(rectangle3_xs[2235]), .RECT3_Y(rectangle3_ys[2235]), .RECT3_WIDTH(rectangle3_widths[2235]), .RECT3_HEIGHT(rectangle3_heights[2235]), .RECT3_WEIGHT(rectangle3_weights[2235]), .FEAT_THRES(feature_thresholds[2235]), .FEAT_ABOVE(feature_aboves[2235]), .FEAT_BELOW(feature_belows[2235])) ac2235(.scan_win(scan_win2235), .scan_win_std_dev(scan_win_std_dev[2235]), .feature_accum(feature_accums[2235]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2236]), .RECT1_Y(rectangle1_ys[2236]), .RECT1_WIDTH(rectangle1_widths[2236]), .RECT1_HEIGHT(rectangle1_heights[2236]), .RECT1_WEIGHT(rectangle1_weights[2236]), .RECT2_X(rectangle2_xs[2236]), .RECT2_Y(rectangle2_ys[2236]), .RECT2_WIDTH(rectangle2_widths[2236]), .RECT2_HEIGHT(rectangle2_heights[2236]), .RECT2_WEIGHT(rectangle2_weights[2236]), .RECT3_X(rectangle3_xs[2236]), .RECT3_Y(rectangle3_ys[2236]), .RECT3_WIDTH(rectangle3_widths[2236]), .RECT3_HEIGHT(rectangle3_heights[2236]), .RECT3_WEIGHT(rectangle3_weights[2236]), .FEAT_THRES(feature_thresholds[2236]), .FEAT_ABOVE(feature_aboves[2236]), .FEAT_BELOW(feature_belows[2236])) ac2236(.scan_win(scan_win2236), .scan_win_std_dev(scan_win_std_dev[2236]), .feature_accum(feature_accums[2236]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2237]), .RECT1_Y(rectangle1_ys[2237]), .RECT1_WIDTH(rectangle1_widths[2237]), .RECT1_HEIGHT(rectangle1_heights[2237]), .RECT1_WEIGHT(rectangle1_weights[2237]), .RECT2_X(rectangle2_xs[2237]), .RECT2_Y(rectangle2_ys[2237]), .RECT2_WIDTH(rectangle2_widths[2237]), .RECT2_HEIGHT(rectangle2_heights[2237]), .RECT2_WEIGHT(rectangle2_weights[2237]), .RECT3_X(rectangle3_xs[2237]), .RECT3_Y(rectangle3_ys[2237]), .RECT3_WIDTH(rectangle3_widths[2237]), .RECT3_HEIGHT(rectangle3_heights[2237]), .RECT3_WEIGHT(rectangle3_weights[2237]), .FEAT_THRES(feature_thresholds[2237]), .FEAT_ABOVE(feature_aboves[2237]), .FEAT_BELOW(feature_belows[2237])) ac2237(.scan_win(scan_win2237), .scan_win_std_dev(scan_win_std_dev[2237]), .feature_accum(feature_accums[2237]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2238]), .RECT1_Y(rectangle1_ys[2238]), .RECT1_WIDTH(rectangle1_widths[2238]), .RECT1_HEIGHT(rectangle1_heights[2238]), .RECT1_WEIGHT(rectangle1_weights[2238]), .RECT2_X(rectangle2_xs[2238]), .RECT2_Y(rectangle2_ys[2238]), .RECT2_WIDTH(rectangle2_widths[2238]), .RECT2_HEIGHT(rectangle2_heights[2238]), .RECT2_WEIGHT(rectangle2_weights[2238]), .RECT3_X(rectangle3_xs[2238]), .RECT3_Y(rectangle3_ys[2238]), .RECT3_WIDTH(rectangle3_widths[2238]), .RECT3_HEIGHT(rectangle3_heights[2238]), .RECT3_WEIGHT(rectangle3_weights[2238]), .FEAT_THRES(feature_thresholds[2238]), .FEAT_ABOVE(feature_aboves[2238]), .FEAT_BELOW(feature_belows[2238])) ac2238(.scan_win(scan_win2238), .scan_win_std_dev(scan_win_std_dev[2238]), .feature_accum(feature_accums[2238]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2239]), .RECT1_Y(rectangle1_ys[2239]), .RECT1_WIDTH(rectangle1_widths[2239]), .RECT1_HEIGHT(rectangle1_heights[2239]), .RECT1_WEIGHT(rectangle1_weights[2239]), .RECT2_X(rectangle2_xs[2239]), .RECT2_Y(rectangle2_ys[2239]), .RECT2_WIDTH(rectangle2_widths[2239]), .RECT2_HEIGHT(rectangle2_heights[2239]), .RECT2_WEIGHT(rectangle2_weights[2239]), .RECT3_X(rectangle3_xs[2239]), .RECT3_Y(rectangle3_ys[2239]), .RECT3_WIDTH(rectangle3_widths[2239]), .RECT3_HEIGHT(rectangle3_heights[2239]), .RECT3_WEIGHT(rectangle3_weights[2239]), .FEAT_THRES(feature_thresholds[2239]), .FEAT_ABOVE(feature_aboves[2239]), .FEAT_BELOW(feature_belows[2239])) ac2239(.scan_win(scan_win2239), .scan_win_std_dev(scan_win_std_dev[2239]), .feature_accum(feature_accums[2239]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2240]), .RECT1_Y(rectangle1_ys[2240]), .RECT1_WIDTH(rectangle1_widths[2240]), .RECT1_HEIGHT(rectangle1_heights[2240]), .RECT1_WEIGHT(rectangle1_weights[2240]), .RECT2_X(rectangle2_xs[2240]), .RECT2_Y(rectangle2_ys[2240]), .RECT2_WIDTH(rectangle2_widths[2240]), .RECT2_HEIGHT(rectangle2_heights[2240]), .RECT2_WEIGHT(rectangle2_weights[2240]), .RECT3_X(rectangle3_xs[2240]), .RECT3_Y(rectangle3_ys[2240]), .RECT3_WIDTH(rectangle3_widths[2240]), .RECT3_HEIGHT(rectangle3_heights[2240]), .RECT3_WEIGHT(rectangle3_weights[2240]), .FEAT_THRES(feature_thresholds[2240]), .FEAT_ABOVE(feature_aboves[2240]), .FEAT_BELOW(feature_belows[2240])) ac2240(.scan_win(scan_win2240), .scan_win_std_dev(scan_win_std_dev[2240]), .feature_accum(feature_accums[2240]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2241]), .RECT1_Y(rectangle1_ys[2241]), .RECT1_WIDTH(rectangle1_widths[2241]), .RECT1_HEIGHT(rectangle1_heights[2241]), .RECT1_WEIGHT(rectangle1_weights[2241]), .RECT2_X(rectangle2_xs[2241]), .RECT2_Y(rectangle2_ys[2241]), .RECT2_WIDTH(rectangle2_widths[2241]), .RECT2_HEIGHT(rectangle2_heights[2241]), .RECT2_WEIGHT(rectangle2_weights[2241]), .RECT3_X(rectangle3_xs[2241]), .RECT3_Y(rectangle3_ys[2241]), .RECT3_WIDTH(rectangle3_widths[2241]), .RECT3_HEIGHT(rectangle3_heights[2241]), .RECT3_WEIGHT(rectangle3_weights[2241]), .FEAT_THRES(feature_thresholds[2241]), .FEAT_ABOVE(feature_aboves[2241]), .FEAT_BELOW(feature_belows[2241])) ac2241(.scan_win(scan_win2241), .scan_win_std_dev(scan_win_std_dev[2241]), .feature_accum(feature_accums[2241]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2242]), .RECT1_Y(rectangle1_ys[2242]), .RECT1_WIDTH(rectangle1_widths[2242]), .RECT1_HEIGHT(rectangle1_heights[2242]), .RECT1_WEIGHT(rectangle1_weights[2242]), .RECT2_X(rectangle2_xs[2242]), .RECT2_Y(rectangle2_ys[2242]), .RECT2_WIDTH(rectangle2_widths[2242]), .RECT2_HEIGHT(rectangle2_heights[2242]), .RECT2_WEIGHT(rectangle2_weights[2242]), .RECT3_X(rectangle3_xs[2242]), .RECT3_Y(rectangle3_ys[2242]), .RECT3_WIDTH(rectangle3_widths[2242]), .RECT3_HEIGHT(rectangle3_heights[2242]), .RECT3_WEIGHT(rectangle3_weights[2242]), .FEAT_THRES(feature_thresholds[2242]), .FEAT_ABOVE(feature_aboves[2242]), .FEAT_BELOW(feature_belows[2242])) ac2242(.scan_win(scan_win2242), .scan_win_std_dev(scan_win_std_dev[2242]), .feature_accum(feature_accums[2242]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2243]), .RECT1_Y(rectangle1_ys[2243]), .RECT1_WIDTH(rectangle1_widths[2243]), .RECT1_HEIGHT(rectangle1_heights[2243]), .RECT1_WEIGHT(rectangle1_weights[2243]), .RECT2_X(rectangle2_xs[2243]), .RECT2_Y(rectangle2_ys[2243]), .RECT2_WIDTH(rectangle2_widths[2243]), .RECT2_HEIGHT(rectangle2_heights[2243]), .RECT2_WEIGHT(rectangle2_weights[2243]), .RECT3_X(rectangle3_xs[2243]), .RECT3_Y(rectangle3_ys[2243]), .RECT3_WIDTH(rectangle3_widths[2243]), .RECT3_HEIGHT(rectangle3_heights[2243]), .RECT3_WEIGHT(rectangle3_weights[2243]), .FEAT_THRES(feature_thresholds[2243]), .FEAT_ABOVE(feature_aboves[2243]), .FEAT_BELOW(feature_belows[2243])) ac2243(.scan_win(scan_win2243), .scan_win_std_dev(scan_win_std_dev[2243]), .feature_accum(feature_accums[2243]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2244]), .RECT1_Y(rectangle1_ys[2244]), .RECT1_WIDTH(rectangle1_widths[2244]), .RECT1_HEIGHT(rectangle1_heights[2244]), .RECT1_WEIGHT(rectangle1_weights[2244]), .RECT2_X(rectangle2_xs[2244]), .RECT2_Y(rectangle2_ys[2244]), .RECT2_WIDTH(rectangle2_widths[2244]), .RECT2_HEIGHT(rectangle2_heights[2244]), .RECT2_WEIGHT(rectangle2_weights[2244]), .RECT3_X(rectangle3_xs[2244]), .RECT3_Y(rectangle3_ys[2244]), .RECT3_WIDTH(rectangle3_widths[2244]), .RECT3_HEIGHT(rectangle3_heights[2244]), .RECT3_WEIGHT(rectangle3_weights[2244]), .FEAT_THRES(feature_thresholds[2244]), .FEAT_ABOVE(feature_aboves[2244]), .FEAT_BELOW(feature_belows[2244])) ac2244(.scan_win(scan_win2244), .scan_win_std_dev(scan_win_std_dev[2244]), .feature_accum(feature_accums[2244]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2245]), .RECT1_Y(rectangle1_ys[2245]), .RECT1_WIDTH(rectangle1_widths[2245]), .RECT1_HEIGHT(rectangle1_heights[2245]), .RECT1_WEIGHT(rectangle1_weights[2245]), .RECT2_X(rectangle2_xs[2245]), .RECT2_Y(rectangle2_ys[2245]), .RECT2_WIDTH(rectangle2_widths[2245]), .RECT2_HEIGHT(rectangle2_heights[2245]), .RECT2_WEIGHT(rectangle2_weights[2245]), .RECT3_X(rectangle3_xs[2245]), .RECT3_Y(rectangle3_ys[2245]), .RECT3_WIDTH(rectangle3_widths[2245]), .RECT3_HEIGHT(rectangle3_heights[2245]), .RECT3_WEIGHT(rectangle3_weights[2245]), .FEAT_THRES(feature_thresholds[2245]), .FEAT_ABOVE(feature_aboves[2245]), .FEAT_BELOW(feature_belows[2245])) ac2245(.scan_win(scan_win2245), .scan_win_std_dev(scan_win_std_dev[2245]), .feature_accum(feature_accums[2245]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2246]), .RECT1_Y(rectangle1_ys[2246]), .RECT1_WIDTH(rectangle1_widths[2246]), .RECT1_HEIGHT(rectangle1_heights[2246]), .RECT1_WEIGHT(rectangle1_weights[2246]), .RECT2_X(rectangle2_xs[2246]), .RECT2_Y(rectangle2_ys[2246]), .RECT2_WIDTH(rectangle2_widths[2246]), .RECT2_HEIGHT(rectangle2_heights[2246]), .RECT2_WEIGHT(rectangle2_weights[2246]), .RECT3_X(rectangle3_xs[2246]), .RECT3_Y(rectangle3_ys[2246]), .RECT3_WIDTH(rectangle3_widths[2246]), .RECT3_HEIGHT(rectangle3_heights[2246]), .RECT3_WEIGHT(rectangle3_weights[2246]), .FEAT_THRES(feature_thresholds[2246]), .FEAT_ABOVE(feature_aboves[2246]), .FEAT_BELOW(feature_belows[2246])) ac2246(.scan_win(scan_win2246), .scan_win_std_dev(scan_win_std_dev[2246]), .feature_accum(feature_accums[2246]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2247]), .RECT1_Y(rectangle1_ys[2247]), .RECT1_WIDTH(rectangle1_widths[2247]), .RECT1_HEIGHT(rectangle1_heights[2247]), .RECT1_WEIGHT(rectangle1_weights[2247]), .RECT2_X(rectangle2_xs[2247]), .RECT2_Y(rectangle2_ys[2247]), .RECT2_WIDTH(rectangle2_widths[2247]), .RECT2_HEIGHT(rectangle2_heights[2247]), .RECT2_WEIGHT(rectangle2_weights[2247]), .RECT3_X(rectangle3_xs[2247]), .RECT3_Y(rectangle3_ys[2247]), .RECT3_WIDTH(rectangle3_widths[2247]), .RECT3_HEIGHT(rectangle3_heights[2247]), .RECT3_WEIGHT(rectangle3_weights[2247]), .FEAT_THRES(feature_thresholds[2247]), .FEAT_ABOVE(feature_aboves[2247]), .FEAT_BELOW(feature_belows[2247])) ac2247(.scan_win(scan_win2247), .scan_win_std_dev(scan_win_std_dev[2247]), .feature_accum(feature_accums[2247]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2248]), .RECT1_Y(rectangle1_ys[2248]), .RECT1_WIDTH(rectangle1_widths[2248]), .RECT1_HEIGHT(rectangle1_heights[2248]), .RECT1_WEIGHT(rectangle1_weights[2248]), .RECT2_X(rectangle2_xs[2248]), .RECT2_Y(rectangle2_ys[2248]), .RECT2_WIDTH(rectangle2_widths[2248]), .RECT2_HEIGHT(rectangle2_heights[2248]), .RECT2_WEIGHT(rectangle2_weights[2248]), .RECT3_X(rectangle3_xs[2248]), .RECT3_Y(rectangle3_ys[2248]), .RECT3_WIDTH(rectangle3_widths[2248]), .RECT3_HEIGHT(rectangle3_heights[2248]), .RECT3_WEIGHT(rectangle3_weights[2248]), .FEAT_THRES(feature_thresholds[2248]), .FEAT_ABOVE(feature_aboves[2248]), .FEAT_BELOW(feature_belows[2248])) ac2248(.scan_win(scan_win2248), .scan_win_std_dev(scan_win_std_dev[2248]), .feature_accum(feature_accums[2248]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2249]), .RECT1_Y(rectangle1_ys[2249]), .RECT1_WIDTH(rectangle1_widths[2249]), .RECT1_HEIGHT(rectangle1_heights[2249]), .RECT1_WEIGHT(rectangle1_weights[2249]), .RECT2_X(rectangle2_xs[2249]), .RECT2_Y(rectangle2_ys[2249]), .RECT2_WIDTH(rectangle2_widths[2249]), .RECT2_HEIGHT(rectangle2_heights[2249]), .RECT2_WEIGHT(rectangle2_weights[2249]), .RECT3_X(rectangle3_xs[2249]), .RECT3_Y(rectangle3_ys[2249]), .RECT3_WIDTH(rectangle3_widths[2249]), .RECT3_HEIGHT(rectangle3_heights[2249]), .RECT3_WEIGHT(rectangle3_weights[2249]), .FEAT_THRES(feature_thresholds[2249]), .FEAT_ABOVE(feature_aboves[2249]), .FEAT_BELOW(feature_belows[2249])) ac2249(.scan_win(scan_win2249), .scan_win_std_dev(scan_win_std_dev[2249]), .feature_accum(feature_accums[2249]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2250]), .RECT1_Y(rectangle1_ys[2250]), .RECT1_WIDTH(rectangle1_widths[2250]), .RECT1_HEIGHT(rectangle1_heights[2250]), .RECT1_WEIGHT(rectangle1_weights[2250]), .RECT2_X(rectangle2_xs[2250]), .RECT2_Y(rectangle2_ys[2250]), .RECT2_WIDTH(rectangle2_widths[2250]), .RECT2_HEIGHT(rectangle2_heights[2250]), .RECT2_WEIGHT(rectangle2_weights[2250]), .RECT3_X(rectangle3_xs[2250]), .RECT3_Y(rectangle3_ys[2250]), .RECT3_WIDTH(rectangle3_widths[2250]), .RECT3_HEIGHT(rectangle3_heights[2250]), .RECT3_WEIGHT(rectangle3_weights[2250]), .FEAT_THRES(feature_thresholds[2250]), .FEAT_ABOVE(feature_aboves[2250]), .FEAT_BELOW(feature_belows[2250])) ac2250(.scan_win(scan_win2250), .scan_win_std_dev(scan_win_std_dev[2250]), .feature_accum(feature_accums[2250]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2251]), .RECT1_Y(rectangle1_ys[2251]), .RECT1_WIDTH(rectangle1_widths[2251]), .RECT1_HEIGHT(rectangle1_heights[2251]), .RECT1_WEIGHT(rectangle1_weights[2251]), .RECT2_X(rectangle2_xs[2251]), .RECT2_Y(rectangle2_ys[2251]), .RECT2_WIDTH(rectangle2_widths[2251]), .RECT2_HEIGHT(rectangle2_heights[2251]), .RECT2_WEIGHT(rectangle2_weights[2251]), .RECT3_X(rectangle3_xs[2251]), .RECT3_Y(rectangle3_ys[2251]), .RECT3_WIDTH(rectangle3_widths[2251]), .RECT3_HEIGHT(rectangle3_heights[2251]), .RECT3_WEIGHT(rectangle3_weights[2251]), .FEAT_THRES(feature_thresholds[2251]), .FEAT_ABOVE(feature_aboves[2251]), .FEAT_BELOW(feature_belows[2251])) ac2251(.scan_win(scan_win2251), .scan_win_std_dev(scan_win_std_dev[2251]), .feature_accum(feature_accums[2251]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2252]), .RECT1_Y(rectangle1_ys[2252]), .RECT1_WIDTH(rectangle1_widths[2252]), .RECT1_HEIGHT(rectangle1_heights[2252]), .RECT1_WEIGHT(rectangle1_weights[2252]), .RECT2_X(rectangle2_xs[2252]), .RECT2_Y(rectangle2_ys[2252]), .RECT2_WIDTH(rectangle2_widths[2252]), .RECT2_HEIGHT(rectangle2_heights[2252]), .RECT2_WEIGHT(rectangle2_weights[2252]), .RECT3_X(rectangle3_xs[2252]), .RECT3_Y(rectangle3_ys[2252]), .RECT3_WIDTH(rectangle3_widths[2252]), .RECT3_HEIGHT(rectangle3_heights[2252]), .RECT3_WEIGHT(rectangle3_weights[2252]), .FEAT_THRES(feature_thresholds[2252]), .FEAT_ABOVE(feature_aboves[2252]), .FEAT_BELOW(feature_belows[2252])) ac2252(.scan_win(scan_win2252), .scan_win_std_dev(scan_win_std_dev[2252]), .feature_accum(feature_accums[2252]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2253]), .RECT1_Y(rectangle1_ys[2253]), .RECT1_WIDTH(rectangle1_widths[2253]), .RECT1_HEIGHT(rectangle1_heights[2253]), .RECT1_WEIGHT(rectangle1_weights[2253]), .RECT2_X(rectangle2_xs[2253]), .RECT2_Y(rectangle2_ys[2253]), .RECT2_WIDTH(rectangle2_widths[2253]), .RECT2_HEIGHT(rectangle2_heights[2253]), .RECT2_WEIGHT(rectangle2_weights[2253]), .RECT3_X(rectangle3_xs[2253]), .RECT3_Y(rectangle3_ys[2253]), .RECT3_WIDTH(rectangle3_widths[2253]), .RECT3_HEIGHT(rectangle3_heights[2253]), .RECT3_WEIGHT(rectangle3_weights[2253]), .FEAT_THRES(feature_thresholds[2253]), .FEAT_ABOVE(feature_aboves[2253]), .FEAT_BELOW(feature_belows[2253])) ac2253(.scan_win(scan_win2253), .scan_win_std_dev(scan_win_std_dev[2253]), .feature_accum(feature_accums[2253]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2254]), .RECT1_Y(rectangle1_ys[2254]), .RECT1_WIDTH(rectangle1_widths[2254]), .RECT1_HEIGHT(rectangle1_heights[2254]), .RECT1_WEIGHT(rectangle1_weights[2254]), .RECT2_X(rectangle2_xs[2254]), .RECT2_Y(rectangle2_ys[2254]), .RECT2_WIDTH(rectangle2_widths[2254]), .RECT2_HEIGHT(rectangle2_heights[2254]), .RECT2_WEIGHT(rectangle2_weights[2254]), .RECT3_X(rectangle3_xs[2254]), .RECT3_Y(rectangle3_ys[2254]), .RECT3_WIDTH(rectangle3_widths[2254]), .RECT3_HEIGHT(rectangle3_heights[2254]), .RECT3_WEIGHT(rectangle3_weights[2254]), .FEAT_THRES(feature_thresholds[2254]), .FEAT_ABOVE(feature_aboves[2254]), .FEAT_BELOW(feature_belows[2254])) ac2254(.scan_win(scan_win2254), .scan_win_std_dev(scan_win_std_dev[2254]), .feature_accum(feature_accums[2254]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2255]), .RECT1_Y(rectangle1_ys[2255]), .RECT1_WIDTH(rectangle1_widths[2255]), .RECT1_HEIGHT(rectangle1_heights[2255]), .RECT1_WEIGHT(rectangle1_weights[2255]), .RECT2_X(rectangle2_xs[2255]), .RECT2_Y(rectangle2_ys[2255]), .RECT2_WIDTH(rectangle2_widths[2255]), .RECT2_HEIGHT(rectangle2_heights[2255]), .RECT2_WEIGHT(rectangle2_weights[2255]), .RECT3_X(rectangle3_xs[2255]), .RECT3_Y(rectangle3_ys[2255]), .RECT3_WIDTH(rectangle3_widths[2255]), .RECT3_HEIGHT(rectangle3_heights[2255]), .RECT3_WEIGHT(rectangle3_weights[2255]), .FEAT_THRES(feature_thresholds[2255]), .FEAT_ABOVE(feature_aboves[2255]), .FEAT_BELOW(feature_belows[2255])) ac2255(.scan_win(scan_win2255), .scan_win_std_dev(scan_win_std_dev[2255]), .feature_accum(feature_accums[2255]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2256]), .RECT1_Y(rectangle1_ys[2256]), .RECT1_WIDTH(rectangle1_widths[2256]), .RECT1_HEIGHT(rectangle1_heights[2256]), .RECT1_WEIGHT(rectangle1_weights[2256]), .RECT2_X(rectangle2_xs[2256]), .RECT2_Y(rectangle2_ys[2256]), .RECT2_WIDTH(rectangle2_widths[2256]), .RECT2_HEIGHT(rectangle2_heights[2256]), .RECT2_WEIGHT(rectangle2_weights[2256]), .RECT3_X(rectangle3_xs[2256]), .RECT3_Y(rectangle3_ys[2256]), .RECT3_WIDTH(rectangle3_widths[2256]), .RECT3_HEIGHT(rectangle3_heights[2256]), .RECT3_WEIGHT(rectangle3_weights[2256]), .FEAT_THRES(feature_thresholds[2256]), .FEAT_ABOVE(feature_aboves[2256]), .FEAT_BELOW(feature_belows[2256])) ac2256(.scan_win(scan_win2256), .scan_win_std_dev(scan_win_std_dev[2256]), .feature_accum(feature_accums[2256]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2257]), .RECT1_Y(rectangle1_ys[2257]), .RECT1_WIDTH(rectangle1_widths[2257]), .RECT1_HEIGHT(rectangle1_heights[2257]), .RECT1_WEIGHT(rectangle1_weights[2257]), .RECT2_X(rectangle2_xs[2257]), .RECT2_Y(rectangle2_ys[2257]), .RECT2_WIDTH(rectangle2_widths[2257]), .RECT2_HEIGHT(rectangle2_heights[2257]), .RECT2_WEIGHT(rectangle2_weights[2257]), .RECT3_X(rectangle3_xs[2257]), .RECT3_Y(rectangle3_ys[2257]), .RECT3_WIDTH(rectangle3_widths[2257]), .RECT3_HEIGHT(rectangle3_heights[2257]), .RECT3_WEIGHT(rectangle3_weights[2257]), .FEAT_THRES(feature_thresholds[2257]), .FEAT_ABOVE(feature_aboves[2257]), .FEAT_BELOW(feature_belows[2257])) ac2257(.scan_win(scan_win2257), .scan_win_std_dev(scan_win_std_dev[2257]), .feature_accum(feature_accums[2257]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2258]), .RECT1_Y(rectangle1_ys[2258]), .RECT1_WIDTH(rectangle1_widths[2258]), .RECT1_HEIGHT(rectangle1_heights[2258]), .RECT1_WEIGHT(rectangle1_weights[2258]), .RECT2_X(rectangle2_xs[2258]), .RECT2_Y(rectangle2_ys[2258]), .RECT2_WIDTH(rectangle2_widths[2258]), .RECT2_HEIGHT(rectangle2_heights[2258]), .RECT2_WEIGHT(rectangle2_weights[2258]), .RECT3_X(rectangle3_xs[2258]), .RECT3_Y(rectangle3_ys[2258]), .RECT3_WIDTH(rectangle3_widths[2258]), .RECT3_HEIGHT(rectangle3_heights[2258]), .RECT3_WEIGHT(rectangle3_weights[2258]), .FEAT_THRES(feature_thresholds[2258]), .FEAT_ABOVE(feature_aboves[2258]), .FEAT_BELOW(feature_belows[2258])) ac2258(.scan_win(scan_win2258), .scan_win_std_dev(scan_win_std_dev[2258]), .feature_accum(feature_accums[2258]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2259]), .RECT1_Y(rectangle1_ys[2259]), .RECT1_WIDTH(rectangle1_widths[2259]), .RECT1_HEIGHT(rectangle1_heights[2259]), .RECT1_WEIGHT(rectangle1_weights[2259]), .RECT2_X(rectangle2_xs[2259]), .RECT2_Y(rectangle2_ys[2259]), .RECT2_WIDTH(rectangle2_widths[2259]), .RECT2_HEIGHT(rectangle2_heights[2259]), .RECT2_WEIGHT(rectangle2_weights[2259]), .RECT3_X(rectangle3_xs[2259]), .RECT3_Y(rectangle3_ys[2259]), .RECT3_WIDTH(rectangle3_widths[2259]), .RECT3_HEIGHT(rectangle3_heights[2259]), .RECT3_WEIGHT(rectangle3_weights[2259]), .FEAT_THRES(feature_thresholds[2259]), .FEAT_ABOVE(feature_aboves[2259]), .FEAT_BELOW(feature_belows[2259])) ac2259(.scan_win(scan_win2259), .scan_win_std_dev(scan_win_std_dev[2259]), .feature_accum(feature_accums[2259]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2260]), .RECT1_Y(rectangle1_ys[2260]), .RECT1_WIDTH(rectangle1_widths[2260]), .RECT1_HEIGHT(rectangle1_heights[2260]), .RECT1_WEIGHT(rectangle1_weights[2260]), .RECT2_X(rectangle2_xs[2260]), .RECT2_Y(rectangle2_ys[2260]), .RECT2_WIDTH(rectangle2_widths[2260]), .RECT2_HEIGHT(rectangle2_heights[2260]), .RECT2_WEIGHT(rectangle2_weights[2260]), .RECT3_X(rectangle3_xs[2260]), .RECT3_Y(rectangle3_ys[2260]), .RECT3_WIDTH(rectangle3_widths[2260]), .RECT3_HEIGHT(rectangle3_heights[2260]), .RECT3_WEIGHT(rectangle3_weights[2260]), .FEAT_THRES(feature_thresholds[2260]), .FEAT_ABOVE(feature_aboves[2260]), .FEAT_BELOW(feature_belows[2260])) ac2260(.scan_win(scan_win2260), .scan_win_std_dev(scan_win_std_dev[2260]), .feature_accum(feature_accums[2260]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2261]), .RECT1_Y(rectangle1_ys[2261]), .RECT1_WIDTH(rectangle1_widths[2261]), .RECT1_HEIGHT(rectangle1_heights[2261]), .RECT1_WEIGHT(rectangle1_weights[2261]), .RECT2_X(rectangle2_xs[2261]), .RECT2_Y(rectangle2_ys[2261]), .RECT2_WIDTH(rectangle2_widths[2261]), .RECT2_HEIGHT(rectangle2_heights[2261]), .RECT2_WEIGHT(rectangle2_weights[2261]), .RECT3_X(rectangle3_xs[2261]), .RECT3_Y(rectangle3_ys[2261]), .RECT3_WIDTH(rectangle3_widths[2261]), .RECT3_HEIGHT(rectangle3_heights[2261]), .RECT3_WEIGHT(rectangle3_weights[2261]), .FEAT_THRES(feature_thresholds[2261]), .FEAT_ABOVE(feature_aboves[2261]), .FEAT_BELOW(feature_belows[2261])) ac2261(.scan_win(scan_win2261), .scan_win_std_dev(scan_win_std_dev[2261]), .feature_accum(feature_accums[2261]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2262]), .RECT1_Y(rectangle1_ys[2262]), .RECT1_WIDTH(rectangle1_widths[2262]), .RECT1_HEIGHT(rectangle1_heights[2262]), .RECT1_WEIGHT(rectangle1_weights[2262]), .RECT2_X(rectangle2_xs[2262]), .RECT2_Y(rectangle2_ys[2262]), .RECT2_WIDTH(rectangle2_widths[2262]), .RECT2_HEIGHT(rectangle2_heights[2262]), .RECT2_WEIGHT(rectangle2_weights[2262]), .RECT3_X(rectangle3_xs[2262]), .RECT3_Y(rectangle3_ys[2262]), .RECT3_WIDTH(rectangle3_widths[2262]), .RECT3_HEIGHT(rectangle3_heights[2262]), .RECT3_WEIGHT(rectangle3_weights[2262]), .FEAT_THRES(feature_thresholds[2262]), .FEAT_ABOVE(feature_aboves[2262]), .FEAT_BELOW(feature_belows[2262])) ac2262(.scan_win(scan_win2262), .scan_win_std_dev(scan_win_std_dev[2262]), .feature_accum(feature_accums[2262]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2263]), .RECT1_Y(rectangle1_ys[2263]), .RECT1_WIDTH(rectangle1_widths[2263]), .RECT1_HEIGHT(rectangle1_heights[2263]), .RECT1_WEIGHT(rectangle1_weights[2263]), .RECT2_X(rectangle2_xs[2263]), .RECT2_Y(rectangle2_ys[2263]), .RECT2_WIDTH(rectangle2_widths[2263]), .RECT2_HEIGHT(rectangle2_heights[2263]), .RECT2_WEIGHT(rectangle2_weights[2263]), .RECT3_X(rectangle3_xs[2263]), .RECT3_Y(rectangle3_ys[2263]), .RECT3_WIDTH(rectangle3_widths[2263]), .RECT3_HEIGHT(rectangle3_heights[2263]), .RECT3_WEIGHT(rectangle3_weights[2263]), .FEAT_THRES(feature_thresholds[2263]), .FEAT_ABOVE(feature_aboves[2263]), .FEAT_BELOW(feature_belows[2263])) ac2263(.scan_win(scan_win2263), .scan_win_std_dev(scan_win_std_dev[2263]), .feature_accum(feature_accums[2263]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2264]), .RECT1_Y(rectangle1_ys[2264]), .RECT1_WIDTH(rectangle1_widths[2264]), .RECT1_HEIGHT(rectangle1_heights[2264]), .RECT1_WEIGHT(rectangle1_weights[2264]), .RECT2_X(rectangle2_xs[2264]), .RECT2_Y(rectangle2_ys[2264]), .RECT2_WIDTH(rectangle2_widths[2264]), .RECT2_HEIGHT(rectangle2_heights[2264]), .RECT2_WEIGHT(rectangle2_weights[2264]), .RECT3_X(rectangle3_xs[2264]), .RECT3_Y(rectangle3_ys[2264]), .RECT3_WIDTH(rectangle3_widths[2264]), .RECT3_HEIGHT(rectangle3_heights[2264]), .RECT3_WEIGHT(rectangle3_weights[2264]), .FEAT_THRES(feature_thresholds[2264]), .FEAT_ABOVE(feature_aboves[2264]), .FEAT_BELOW(feature_belows[2264])) ac2264(.scan_win(scan_win2264), .scan_win_std_dev(scan_win_std_dev[2264]), .feature_accum(feature_accums[2264]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2265]), .RECT1_Y(rectangle1_ys[2265]), .RECT1_WIDTH(rectangle1_widths[2265]), .RECT1_HEIGHT(rectangle1_heights[2265]), .RECT1_WEIGHT(rectangle1_weights[2265]), .RECT2_X(rectangle2_xs[2265]), .RECT2_Y(rectangle2_ys[2265]), .RECT2_WIDTH(rectangle2_widths[2265]), .RECT2_HEIGHT(rectangle2_heights[2265]), .RECT2_WEIGHT(rectangle2_weights[2265]), .RECT3_X(rectangle3_xs[2265]), .RECT3_Y(rectangle3_ys[2265]), .RECT3_WIDTH(rectangle3_widths[2265]), .RECT3_HEIGHT(rectangle3_heights[2265]), .RECT3_WEIGHT(rectangle3_weights[2265]), .FEAT_THRES(feature_thresholds[2265]), .FEAT_ABOVE(feature_aboves[2265]), .FEAT_BELOW(feature_belows[2265])) ac2265(.scan_win(scan_win2265), .scan_win_std_dev(scan_win_std_dev[2265]), .feature_accum(feature_accums[2265]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2266]), .RECT1_Y(rectangle1_ys[2266]), .RECT1_WIDTH(rectangle1_widths[2266]), .RECT1_HEIGHT(rectangle1_heights[2266]), .RECT1_WEIGHT(rectangle1_weights[2266]), .RECT2_X(rectangle2_xs[2266]), .RECT2_Y(rectangle2_ys[2266]), .RECT2_WIDTH(rectangle2_widths[2266]), .RECT2_HEIGHT(rectangle2_heights[2266]), .RECT2_WEIGHT(rectangle2_weights[2266]), .RECT3_X(rectangle3_xs[2266]), .RECT3_Y(rectangle3_ys[2266]), .RECT3_WIDTH(rectangle3_widths[2266]), .RECT3_HEIGHT(rectangle3_heights[2266]), .RECT3_WEIGHT(rectangle3_weights[2266]), .FEAT_THRES(feature_thresholds[2266]), .FEAT_ABOVE(feature_aboves[2266]), .FEAT_BELOW(feature_belows[2266])) ac2266(.scan_win(scan_win2266), .scan_win_std_dev(scan_win_std_dev[2266]), .feature_accum(feature_accums[2266]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2267]), .RECT1_Y(rectangle1_ys[2267]), .RECT1_WIDTH(rectangle1_widths[2267]), .RECT1_HEIGHT(rectangle1_heights[2267]), .RECT1_WEIGHT(rectangle1_weights[2267]), .RECT2_X(rectangle2_xs[2267]), .RECT2_Y(rectangle2_ys[2267]), .RECT2_WIDTH(rectangle2_widths[2267]), .RECT2_HEIGHT(rectangle2_heights[2267]), .RECT2_WEIGHT(rectangle2_weights[2267]), .RECT3_X(rectangle3_xs[2267]), .RECT3_Y(rectangle3_ys[2267]), .RECT3_WIDTH(rectangle3_widths[2267]), .RECT3_HEIGHT(rectangle3_heights[2267]), .RECT3_WEIGHT(rectangle3_weights[2267]), .FEAT_THRES(feature_thresholds[2267]), .FEAT_ABOVE(feature_aboves[2267]), .FEAT_BELOW(feature_belows[2267])) ac2267(.scan_win(scan_win2267), .scan_win_std_dev(scan_win_std_dev[2267]), .feature_accum(feature_accums[2267]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2268]), .RECT1_Y(rectangle1_ys[2268]), .RECT1_WIDTH(rectangle1_widths[2268]), .RECT1_HEIGHT(rectangle1_heights[2268]), .RECT1_WEIGHT(rectangle1_weights[2268]), .RECT2_X(rectangle2_xs[2268]), .RECT2_Y(rectangle2_ys[2268]), .RECT2_WIDTH(rectangle2_widths[2268]), .RECT2_HEIGHT(rectangle2_heights[2268]), .RECT2_WEIGHT(rectangle2_weights[2268]), .RECT3_X(rectangle3_xs[2268]), .RECT3_Y(rectangle3_ys[2268]), .RECT3_WIDTH(rectangle3_widths[2268]), .RECT3_HEIGHT(rectangle3_heights[2268]), .RECT3_WEIGHT(rectangle3_weights[2268]), .FEAT_THRES(feature_thresholds[2268]), .FEAT_ABOVE(feature_aboves[2268]), .FEAT_BELOW(feature_belows[2268])) ac2268(.scan_win(scan_win2268), .scan_win_std_dev(scan_win_std_dev[2268]), .feature_accum(feature_accums[2268]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2269]), .RECT1_Y(rectangle1_ys[2269]), .RECT1_WIDTH(rectangle1_widths[2269]), .RECT1_HEIGHT(rectangle1_heights[2269]), .RECT1_WEIGHT(rectangle1_weights[2269]), .RECT2_X(rectangle2_xs[2269]), .RECT2_Y(rectangle2_ys[2269]), .RECT2_WIDTH(rectangle2_widths[2269]), .RECT2_HEIGHT(rectangle2_heights[2269]), .RECT2_WEIGHT(rectangle2_weights[2269]), .RECT3_X(rectangle3_xs[2269]), .RECT3_Y(rectangle3_ys[2269]), .RECT3_WIDTH(rectangle3_widths[2269]), .RECT3_HEIGHT(rectangle3_heights[2269]), .RECT3_WEIGHT(rectangle3_weights[2269]), .FEAT_THRES(feature_thresholds[2269]), .FEAT_ABOVE(feature_aboves[2269]), .FEAT_BELOW(feature_belows[2269])) ac2269(.scan_win(scan_win2269), .scan_win_std_dev(scan_win_std_dev[2269]), .feature_accum(feature_accums[2269]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2270]), .RECT1_Y(rectangle1_ys[2270]), .RECT1_WIDTH(rectangle1_widths[2270]), .RECT1_HEIGHT(rectangle1_heights[2270]), .RECT1_WEIGHT(rectangle1_weights[2270]), .RECT2_X(rectangle2_xs[2270]), .RECT2_Y(rectangle2_ys[2270]), .RECT2_WIDTH(rectangle2_widths[2270]), .RECT2_HEIGHT(rectangle2_heights[2270]), .RECT2_WEIGHT(rectangle2_weights[2270]), .RECT3_X(rectangle3_xs[2270]), .RECT3_Y(rectangle3_ys[2270]), .RECT3_WIDTH(rectangle3_widths[2270]), .RECT3_HEIGHT(rectangle3_heights[2270]), .RECT3_WEIGHT(rectangle3_weights[2270]), .FEAT_THRES(feature_thresholds[2270]), .FEAT_ABOVE(feature_aboves[2270]), .FEAT_BELOW(feature_belows[2270])) ac2270(.scan_win(scan_win2270), .scan_win_std_dev(scan_win_std_dev[2270]), .feature_accum(feature_accums[2270]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2271]), .RECT1_Y(rectangle1_ys[2271]), .RECT1_WIDTH(rectangle1_widths[2271]), .RECT1_HEIGHT(rectangle1_heights[2271]), .RECT1_WEIGHT(rectangle1_weights[2271]), .RECT2_X(rectangle2_xs[2271]), .RECT2_Y(rectangle2_ys[2271]), .RECT2_WIDTH(rectangle2_widths[2271]), .RECT2_HEIGHT(rectangle2_heights[2271]), .RECT2_WEIGHT(rectangle2_weights[2271]), .RECT3_X(rectangle3_xs[2271]), .RECT3_Y(rectangle3_ys[2271]), .RECT3_WIDTH(rectangle3_widths[2271]), .RECT3_HEIGHT(rectangle3_heights[2271]), .RECT3_WEIGHT(rectangle3_weights[2271]), .FEAT_THRES(feature_thresholds[2271]), .FEAT_ABOVE(feature_aboves[2271]), .FEAT_BELOW(feature_belows[2271])) ac2271(.scan_win(scan_win2271), .scan_win_std_dev(scan_win_std_dev[2271]), .feature_accum(feature_accums[2271]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2272]), .RECT1_Y(rectangle1_ys[2272]), .RECT1_WIDTH(rectangle1_widths[2272]), .RECT1_HEIGHT(rectangle1_heights[2272]), .RECT1_WEIGHT(rectangle1_weights[2272]), .RECT2_X(rectangle2_xs[2272]), .RECT2_Y(rectangle2_ys[2272]), .RECT2_WIDTH(rectangle2_widths[2272]), .RECT2_HEIGHT(rectangle2_heights[2272]), .RECT2_WEIGHT(rectangle2_weights[2272]), .RECT3_X(rectangle3_xs[2272]), .RECT3_Y(rectangle3_ys[2272]), .RECT3_WIDTH(rectangle3_widths[2272]), .RECT3_HEIGHT(rectangle3_heights[2272]), .RECT3_WEIGHT(rectangle3_weights[2272]), .FEAT_THRES(feature_thresholds[2272]), .FEAT_ABOVE(feature_aboves[2272]), .FEAT_BELOW(feature_belows[2272])) ac2272(.scan_win(scan_win2272), .scan_win_std_dev(scan_win_std_dev[2272]), .feature_accum(feature_accums[2272]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2273]), .RECT1_Y(rectangle1_ys[2273]), .RECT1_WIDTH(rectangle1_widths[2273]), .RECT1_HEIGHT(rectangle1_heights[2273]), .RECT1_WEIGHT(rectangle1_weights[2273]), .RECT2_X(rectangle2_xs[2273]), .RECT2_Y(rectangle2_ys[2273]), .RECT2_WIDTH(rectangle2_widths[2273]), .RECT2_HEIGHT(rectangle2_heights[2273]), .RECT2_WEIGHT(rectangle2_weights[2273]), .RECT3_X(rectangle3_xs[2273]), .RECT3_Y(rectangle3_ys[2273]), .RECT3_WIDTH(rectangle3_widths[2273]), .RECT3_HEIGHT(rectangle3_heights[2273]), .RECT3_WEIGHT(rectangle3_weights[2273]), .FEAT_THRES(feature_thresholds[2273]), .FEAT_ABOVE(feature_aboves[2273]), .FEAT_BELOW(feature_belows[2273])) ac2273(.scan_win(scan_win2273), .scan_win_std_dev(scan_win_std_dev[2273]), .feature_accum(feature_accums[2273]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2274]), .RECT1_Y(rectangle1_ys[2274]), .RECT1_WIDTH(rectangle1_widths[2274]), .RECT1_HEIGHT(rectangle1_heights[2274]), .RECT1_WEIGHT(rectangle1_weights[2274]), .RECT2_X(rectangle2_xs[2274]), .RECT2_Y(rectangle2_ys[2274]), .RECT2_WIDTH(rectangle2_widths[2274]), .RECT2_HEIGHT(rectangle2_heights[2274]), .RECT2_WEIGHT(rectangle2_weights[2274]), .RECT3_X(rectangle3_xs[2274]), .RECT3_Y(rectangle3_ys[2274]), .RECT3_WIDTH(rectangle3_widths[2274]), .RECT3_HEIGHT(rectangle3_heights[2274]), .RECT3_WEIGHT(rectangle3_weights[2274]), .FEAT_THRES(feature_thresholds[2274]), .FEAT_ABOVE(feature_aboves[2274]), .FEAT_BELOW(feature_belows[2274])) ac2274(.scan_win(scan_win2274), .scan_win_std_dev(scan_win_std_dev[2274]), .feature_accum(feature_accums[2274]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2275]), .RECT1_Y(rectangle1_ys[2275]), .RECT1_WIDTH(rectangle1_widths[2275]), .RECT1_HEIGHT(rectangle1_heights[2275]), .RECT1_WEIGHT(rectangle1_weights[2275]), .RECT2_X(rectangle2_xs[2275]), .RECT2_Y(rectangle2_ys[2275]), .RECT2_WIDTH(rectangle2_widths[2275]), .RECT2_HEIGHT(rectangle2_heights[2275]), .RECT2_WEIGHT(rectangle2_weights[2275]), .RECT3_X(rectangle3_xs[2275]), .RECT3_Y(rectangle3_ys[2275]), .RECT3_WIDTH(rectangle3_widths[2275]), .RECT3_HEIGHT(rectangle3_heights[2275]), .RECT3_WEIGHT(rectangle3_weights[2275]), .FEAT_THRES(feature_thresholds[2275]), .FEAT_ABOVE(feature_aboves[2275]), .FEAT_BELOW(feature_belows[2275])) ac2275(.scan_win(scan_win2275), .scan_win_std_dev(scan_win_std_dev[2275]), .feature_accum(feature_accums[2275]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2276]), .RECT1_Y(rectangle1_ys[2276]), .RECT1_WIDTH(rectangle1_widths[2276]), .RECT1_HEIGHT(rectangle1_heights[2276]), .RECT1_WEIGHT(rectangle1_weights[2276]), .RECT2_X(rectangle2_xs[2276]), .RECT2_Y(rectangle2_ys[2276]), .RECT2_WIDTH(rectangle2_widths[2276]), .RECT2_HEIGHT(rectangle2_heights[2276]), .RECT2_WEIGHT(rectangle2_weights[2276]), .RECT3_X(rectangle3_xs[2276]), .RECT3_Y(rectangle3_ys[2276]), .RECT3_WIDTH(rectangle3_widths[2276]), .RECT3_HEIGHT(rectangle3_heights[2276]), .RECT3_WEIGHT(rectangle3_weights[2276]), .FEAT_THRES(feature_thresholds[2276]), .FEAT_ABOVE(feature_aboves[2276]), .FEAT_BELOW(feature_belows[2276])) ac2276(.scan_win(scan_win2276), .scan_win_std_dev(scan_win_std_dev[2276]), .feature_accum(feature_accums[2276]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2277]), .RECT1_Y(rectangle1_ys[2277]), .RECT1_WIDTH(rectangle1_widths[2277]), .RECT1_HEIGHT(rectangle1_heights[2277]), .RECT1_WEIGHT(rectangle1_weights[2277]), .RECT2_X(rectangle2_xs[2277]), .RECT2_Y(rectangle2_ys[2277]), .RECT2_WIDTH(rectangle2_widths[2277]), .RECT2_HEIGHT(rectangle2_heights[2277]), .RECT2_WEIGHT(rectangle2_weights[2277]), .RECT3_X(rectangle3_xs[2277]), .RECT3_Y(rectangle3_ys[2277]), .RECT3_WIDTH(rectangle3_widths[2277]), .RECT3_HEIGHT(rectangle3_heights[2277]), .RECT3_WEIGHT(rectangle3_weights[2277]), .FEAT_THRES(feature_thresholds[2277]), .FEAT_ABOVE(feature_aboves[2277]), .FEAT_BELOW(feature_belows[2277])) ac2277(.scan_win(scan_win2277), .scan_win_std_dev(scan_win_std_dev[2277]), .feature_accum(feature_accums[2277]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2278]), .RECT1_Y(rectangle1_ys[2278]), .RECT1_WIDTH(rectangle1_widths[2278]), .RECT1_HEIGHT(rectangle1_heights[2278]), .RECT1_WEIGHT(rectangle1_weights[2278]), .RECT2_X(rectangle2_xs[2278]), .RECT2_Y(rectangle2_ys[2278]), .RECT2_WIDTH(rectangle2_widths[2278]), .RECT2_HEIGHT(rectangle2_heights[2278]), .RECT2_WEIGHT(rectangle2_weights[2278]), .RECT3_X(rectangle3_xs[2278]), .RECT3_Y(rectangle3_ys[2278]), .RECT3_WIDTH(rectangle3_widths[2278]), .RECT3_HEIGHT(rectangle3_heights[2278]), .RECT3_WEIGHT(rectangle3_weights[2278]), .FEAT_THRES(feature_thresholds[2278]), .FEAT_ABOVE(feature_aboves[2278]), .FEAT_BELOW(feature_belows[2278])) ac2278(.scan_win(scan_win2278), .scan_win_std_dev(scan_win_std_dev[2278]), .feature_accum(feature_accums[2278]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2279]), .RECT1_Y(rectangle1_ys[2279]), .RECT1_WIDTH(rectangle1_widths[2279]), .RECT1_HEIGHT(rectangle1_heights[2279]), .RECT1_WEIGHT(rectangle1_weights[2279]), .RECT2_X(rectangle2_xs[2279]), .RECT2_Y(rectangle2_ys[2279]), .RECT2_WIDTH(rectangle2_widths[2279]), .RECT2_HEIGHT(rectangle2_heights[2279]), .RECT2_WEIGHT(rectangle2_weights[2279]), .RECT3_X(rectangle3_xs[2279]), .RECT3_Y(rectangle3_ys[2279]), .RECT3_WIDTH(rectangle3_widths[2279]), .RECT3_HEIGHT(rectangle3_heights[2279]), .RECT3_WEIGHT(rectangle3_weights[2279]), .FEAT_THRES(feature_thresholds[2279]), .FEAT_ABOVE(feature_aboves[2279]), .FEAT_BELOW(feature_belows[2279])) ac2279(.scan_win(scan_win2279), .scan_win_std_dev(scan_win_std_dev[2279]), .feature_accum(feature_accums[2279]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2280]), .RECT1_Y(rectangle1_ys[2280]), .RECT1_WIDTH(rectangle1_widths[2280]), .RECT1_HEIGHT(rectangle1_heights[2280]), .RECT1_WEIGHT(rectangle1_weights[2280]), .RECT2_X(rectangle2_xs[2280]), .RECT2_Y(rectangle2_ys[2280]), .RECT2_WIDTH(rectangle2_widths[2280]), .RECT2_HEIGHT(rectangle2_heights[2280]), .RECT2_WEIGHT(rectangle2_weights[2280]), .RECT3_X(rectangle3_xs[2280]), .RECT3_Y(rectangle3_ys[2280]), .RECT3_WIDTH(rectangle3_widths[2280]), .RECT3_HEIGHT(rectangle3_heights[2280]), .RECT3_WEIGHT(rectangle3_weights[2280]), .FEAT_THRES(feature_thresholds[2280]), .FEAT_ABOVE(feature_aboves[2280]), .FEAT_BELOW(feature_belows[2280])) ac2280(.scan_win(scan_win2280), .scan_win_std_dev(scan_win_std_dev[2280]), .feature_accum(feature_accums[2280]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2281]), .RECT1_Y(rectangle1_ys[2281]), .RECT1_WIDTH(rectangle1_widths[2281]), .RECT1_HEIGHT(rectangle1_heights[2281]), .RECT1_WEIGHT(rectangle1_weights[2281]), .RECT2_X(rectangle2_xs[2281]), .RECT2_Y(rectangle2_ys[2281]), .RECT2_WIDTH(rectangle2_widths[2281]), .RECT2_HEIGHT(rectangle2_heights[2281]), .RECT2_WEIGHT(rectangle2_weights[2281]), .RECT3_X(rectangle3_xs[2281]), .RECT3_Y(rectangle3_ys[2281]), .RECT3_WIDTH(rectangle3_widths[2281]), .RECT3_HEIGHT(rectangle3_heights[2281]), .RECT3_WEIGHT(rectangle3_weights[2281]), .FEAT_THRES(feature_thresholds[2281]), .FEAT_ABOVE(feature_aboves[2281]), .FEAT_BELOW(feature_belows[2281])) ac2281(.scan_win(scan_win2281), .scan_win_std_dev(scan_win_std_dev[2281]), .feature_accum(feature_accums[2281]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2282]), .RECT1_Y(rectangle1_ys[2282]), .RECT1_WIDTH(rectangle1_widths[2282]), .RECT1_HEIGHT(rectangle1_heights[2282]), .RECT1_WEIGHT(rectangle1_weights[2282]), .RECT2_X(rectangle2_xs[2282]), .RECT2_Y(rectangle2_ys[2282]), .RECT2_WIDTH(rectangle2_widths[2282]), .RECT2_HEIGHT(rectangle2_heights[2282]), .RECT2_WEIGHT(rectangle2_weights[2282]), .RECT3_X(rectangle3_xs[2282]), .RECT3_Y(rectangle3_ys[2282]), .RECT3_WIDTH(rectangle3_widths[2282]), .RECT3_HEIGHT(rectangle3_heights[2282]), .RECT3_WEIGHT(rectangle3_weights[2282]), .FEAT_THRES(feature_thresholds[2282]), .FEAT_ABOVE(feature_aboves[2282]), .FEAT_BELOW(feature_belows[2282])) ac2282(.scan_win(scan_win2282), .scan_win_std_dev(scan_win_std_dev[2282]), .feature_accum(feature_accums[2282]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2283]), .RECT1_Y(rectangle1_ys[2283]), .RECT1_WIDTH(rectangle1_widths[2283]), .RECT1_HEIGHT(rectangle1_heights[2283]), .RECT1_WEIGHT(rectangle1_weights[2283]), .RECT2_X(rectangle2_xs[2283]), .RECT2_Y(rectangle2_ys[2283]), .RECT2_WIDTH(rectangle2_widths[2283]), .RECT2_HEIGHT(rectangle2_heights[2283]), .RECT2_WEIGHT(rectangle2_weights[2283]), .RECT3_X(rectangle3_xs[2283]), .RECT3_Y(rectangle3_ys[2283]), .RECT3_WIDTH(rectangle3_widths[2283]), .RECT3_HEIGHT(rectangle3_heights[2283]), .RECT3_WEIGHT(rectangle3_weights[2283]), .FEAT_THRES(feature_thresholds[2283]), .FEAT_ABOVE(feature_aboves[2283]), .FEAT_BELOW(feature_belows[2283])) ac2283(.scan_win(scan_win2283), .scan_win_std_dev(scan_win_std_dev[2283]), .feature_accum(feature_accums[2283]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2284]), .RECT1_Y(rectangle1_ys[2284]), .RECT1_WIDTH(rectangle1_widths[2284]), .RECT1_HEIGHT(rectangle1_heights[2284]), .RECT1_WEIGHT(rectangle1_weights[2284]), .RECT2_X(rectangle2_xs[2284]), .RECT2_Y(rectangle2_ys[2284]), .RECT2_WIDTH(rectangle2_widths[2284]), .RECT2_HEIGHT(rectangle2_heights[2284]), .RECT2_WEIGHT(rectangle2_weights[2284]), .RECT3_X(rectangle3_xs[2284]), .RECT3_Y(rectangle3_ys[2284]), .RECT3_WIDTH(rectangle3_widths[2284]), .RECT3_HEIGHT(rectangle3_heights[2284]), .RECT3_WEIGHT(rectangle3_weights[2284]), .FEAT_THRES(feature_thresholds[2284]), .FEAT_ABOVE(feature_aboves[2284]), .FEAT_BELOW(feature_belows[2284])) ac2284(.scan_win(scan_win2284), .scan_win_std_dev(scan_win_std_dev[2284]), .feature_accum(feature_accums[2284]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2285]), .RECT1_Y(rectangle1_ys[2285]), .RECT1_WIDTH(rectangle1_widths[2285]), .RECT1_HEIGHT(rectangle1_heights[2285]), .RECT1_WEIGHT(rectangle1_weights[2285]), .RECT2_X(rectangle2_xs[2285]), .RECT2_Y(rectangle2_ys[2285]), .RECT2_WIDTH(rectangle2_widths[2285]), .RECT2_HEIGHT(rectangle2_heights[2285]), .RECT2_WEIGHT(rectangle2_weights[2285]), .RECT3_X(rectangle3_xs[2285]), .RECT3_Y(rectangle3_ys[2285]), .RECT3_WIDTH(rectangle3_widths[2285]), .RECT3_HEIGHT(rectangle3_heights[2285]), .RECT3_WEIGHT(rectangle3_weights[2285]), .FEAT_THRES(feature_thresholds[2285]), .FEAT_ABOVE(feature_aboves[2285]), .FEAT_BELOW(feature_belows[2285])) ac2285(.scan_win(scan_win2285), .scan_win_std_dev(scan_win_std_dev[2285]), .feature_accum(feature_accums[2285]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2286]), .RECT1_Y(rectangle1_ys[2286]), .RECT1_WIDTH(rectangle1_widths[2286]), .RECT1_HEIGHT(rectangle1_heights[2286]), .RECT1_WEIGHT(rectangle1_weights[2286]), .RECT2_X(rectangle2_xs[2286]), .RECT2_Y(rectangle2_ys[2286]), .RECT2_WIDTH(rectangle2_widths[2286]), .RECT2_HEIGHT(rectangle2_heights[2286]), .RECT2_WEIGHT(rectangle2_weights[2286]), .RECT3_X(rectangle3_xs[2286]), .RECT3_Y(rectangle3_ys[2286]), .RECT3_WIDTH(rectangle3_widths[2286]), .RECT3_HEIGHT(rectangle3_heights[2286]), .RECT3_WEIGHT(rectangle3_weights[2286]), .FEAT_THRES(feature_thresholds[2286]), .FEAT_ABOVE(feature_aboves[2286]), .FEAT_BELOW(feature_belows[2286])) ac2286(.scan_win(scan_win2286), .scan_win_std_dev(scan_win_std_dev[2286]), .feature_accum(feature_accums[2286]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2287]), .RECT1_Y(rectangle1_ys[2287]), .RECT1_WIDTH(rectangle1_widths[2287]), .RECT1_HEIGHT(rectangle1_heights[2287]), .RECT1_WEIGHT(rectangle1_weights[2287]), .RECT2_X(rectangle2_xs[2287]), .RECT2_Y(rectangle2_ys[2287]), .RECT2_WIDTH(rectangle2_widths[2287]), .RECT2_HEIGHT(rectangle2_heights[2287]), .RECT2_WEIGHT(rectangle2_weights[2287]), .RECT3_X(rectangle3_xs[2287]), .RECT3_Y(rectangle3_ys[2287]), .RECT3_WIDTH(rectangle3_widths[2287]), .RECT3_HEIGHT(rectangle3_heights[2287]), .RECT3_WEIGHT(rectangle3_weights[2287]), .FEAT_THRES(feature_thresholds[2287]), .FEAT_ABOVE(feature_aboves[2287]), .FEAT_BELOW(feature_belows[2287])) ac2287(.scan_win(scan_win2287), .scan_win_std_dev(scan_win_std_dev[2287]), .feature_accum(feature_accums[2287]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2288]), .RECT1_Y(rectangle1_ys[2288]), .RECT1_WIDTH(rectangle1_widths[2288]), .RECT1_HEIGHT(rectangle1_heights[2288]), .RECT1_WEIGHT(rectangle1_weights[2288]), .RECT2_X(rectangle2_xs[2288]), .RECT2_Y(rectangle2_ys[2288]), .RECT2_WIDTH(rectangle2_widths[2288]), .RECT2_HEIGHT(rectangle2_heights[2288]), .RECT2_WEIGHT(rectangle2_weights[2288]), .RECT3_X(rectangle3_xs[2288]), .RECT3_Y(rectangle3_ys[2288]), .RECT3_WIDTH(rectangle3_widths[2288]), .RECT3_HEIGHT(rectangle3_heights[2288]), .RECT3_WEIGHT(rectangle3_weights[2288]), .FEAT_THRES(feature_thresholds[2288]), .FEAT_ABOVE(feature_aboves[2288]), .FEAT_BELOW(feature_belows[2288])) ac2288(.scan_win(scan_win2288), .scan_win_std_dev(scan_win_std_dev[2288]), .feature_accum(feature_accums[2288]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2289]), .RECT1_Y(rectangle1_ys[2289]), .RECT1_WIDTH(rectangle1_widths[2289]), .RECT1_HEIGHT(rectangle1_heights[2289]), .RECT1_WEIGHT(rectangle1_weights[2289]), .RECT2_X(rectangle2_xs[2289]), .RECT2_Y(rectangle2_ys[2289]), .RECT2_WIDTH(rectangle2_widths[2289]), .RECT2_HEIGHT(rectangle2_heights[2289]), .RECT2_WEIGHT(rectangle2_weights[2289]), .RECT3_X(rectangle3_xs[2289]), .RECT3_Y(rectangle3_ys[2289]), .RECT3_WIDTH(rectangle3_widths[2289]), .RECT3_HEIGHT(rectangle3_heights[2289]), .RECT3_WEIGHT(rectangle3_weights[2289]), .FEAT_THRES(feature_thresholds[2289]), .FEAT_ABOVE(feature_aboves[2289]), .FEAT_BELOW(feature_belows[2289])) ac2289(.scan_win(scan_win2289), .scan_win_std_dev(scan_win_std_dev[2289]), .feature_accum(feature_accums[2289]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2290]), .RECT1_Y(rectangle1_ys[2290]), .RECT1_WIDTH(rectangle1_widths[2290]), .RECT1_HEIGHT(rectangle1_heights[2290]), .RECT1_WEIGHT(rectangle1_weights[2290]), .RECT2_X(rectangle2_xs[2290]), .RECT2_Y(rectangle2_ys[2290]), .RECT2_WIDTH(rectangle2_widths[2290]), .RECT2_HEIGHT(rectangle2_heights[2290]), .RECT2_WEIGHT(rectangle2_weights[2290]), .RECT3_X(rectangle3_xs[2290]), .RECT3_Y(rectangle3_ys[2290]), .RECT3_WIDTH(rectangle3_widths[2290]), .RECT3_HEIGHT(rectangle3_heights[2290]), .RECT3_WEIGHT(rectangle3_weights[2290]), .FEAT_THRES(feature_thresholds[2290]), .FEAT_ABOVE(feature_aboves[2290]), .FEAT_BELOW(feature_belows[2290])) ac2290(.scan_win(scan_win2290), .scan_win_std_dev(scan_win_std_dev[2290]), .feature_accum(feature_accums[2290]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2291]), .RECT1_Y(rectangle1_ys[2291]), .RECT1_WIDTH(rectangle1_widths[2291]), .RECT1_HEIGHT(rectangle1_heights[2291]), .RECT1_WEIGHT(rectangle1_weights[2291]), .RECT2_X(rectangle2_xs[2291]), .RECT2_Y(rectangle2_ys[2291]), .RECT2_WIDTH(rectangle2_widths[2291]), .RECT2_HEIGHT(rectangle2_heights[2291]), .RECT2_WEIGHT(rectangle2_weights[2291]), .RECT3_X(rectangle3_xs[2291]), .RECT3_Y(rectangle3_ys[2291]), .RECT3_WIDTH(rectangle3_widths[2291]), .RECT3_HEIGHT(rectangle3_heights[2291]), .RECT3_WEIGHT(rectangle3_weights[2291]), .FEAT_THRES(feature_thresholds[2291]), .FEAT_ABOVE(feature_aboves[2291]), .FEAT_BELOW(feature_belows[2291])) ac2291(.scan_win(scan_win2291), .scan_win_std_dev(scan_win_std_dev[2291]), .feature_accum(feature_accums[2291]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2292]), .RECT1_Y(rectangle1_ys[2292]), .RECT1_WIDTH(rectangle1_widths[2292]), .RECT1_HEIGHT(rectangle1_heights[2292]), .RECT1_WEIGHT(rectangle1_weights[2292]), .RECT2_X(rectangle2_xs[2292]), .RECT2_Y(rectangle2_ys[2292]), .RECT2_WIDTH(rectangle2_widths[2292]), .RECT2_HEIGHT(rectangle2_heights[2292]), .RECT2_WEIGHT(rectangle2_weights[2292]), .RECT3_X(rectangle3_xs[2292]), .RECT3_Y(rectangle3_ys[2292]), .RECT3_WIDTH(rectangle3_widths[2292]), .RECT3_HEIGHT(rectangle3_heights[2292]), .RECT3_WEIGHT(rectangle3_weights[2292]), .FEAT_THRES(feature_thresholds[2292]), .FEAT_ABOVE(feature_aboves[2292]), .FEAT_BELOW(feature_belows[2292])) ac2292(.scan_win(scan_win2292), .scan_win_std_dev(scan_win_std_dev[2292]), .feature_accum(feature_accums[2292]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2293]), .RECT1_Y(rectangle1_ys[2293]), .RECT1_WIDTH(rectangle1_widths[2293]), .RECT1_HEIGHT(rectangle1_heights[2293]), .RECT1_WEIGHT(rectangle1_weights[2293]), .RECT2_X(rectangle2_xs[2293]), .RECT2_Y(rectangle2_ys[2293]), .RECT2_WIDTH(rectangle2_widths[2293]), .RECT2_HEIGHT(rectangle2_heights[2293]), .RECT2_WEIGHT(rectangle2_weights[2293]), .RECT3_X(rectangle3_xs[2293]), .RECT3_Y(rectangle3_ys[2293]), .RECT3_WIDTH(rectangle3_widths[2293]), .RECT3_HEIGHT(rectangle3_heights[2293]), .RECT3_WEIGHT(rectangle3_weights[2293]), .FEAT_THRES(feature_thresholds[2293]), .FEAT_ABOVE(feature_aboves[2293]), .FEAT_BELOW(feature_belows[2293])) ac2293(.scan_win(scan_win2293), .scan_win_std_dev(scan_win_std_dev[2293]), .feature_accum(feature_accums[2293]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2294]), .RECT1_Y(rectangle1_ys[2294]), .RECT1_WIDTH(rectangle1_widths[2294]), .RECT1_HEIGHT(rectangle1_heights[2294]), .RECT1_WEIGHT(rectangle1_weights[2294]), .RECT2_X(rectangle2_xs[2294]), .RECT2_Y(rectangle2_ys[2294]), .RECT2_WIDTH(rectangle2_widths[2294]), .RECT2_HEIGHT(rectangle2_heights[2294]), .RECT2_WEIGHT(rectangle2_weights[2294]), .RECT3_X(rectangle3_xs[2294]), .RECT3_Y(rectangle3_ys[2294]), .RECT3_WIDTH(rectangle3_widths[2294]), .RECT3_HEIGHT(rectangle3_heights[2294]), .RECT3_WEIGHT(rectangle3_weights[2294]), .FEAT_THRES(feature_thresholds[2294]), .FEAT_ABOVE(feature_aboves[2294]), .FEAT_BELOW(feature_belows[2294])) ac2294(.scan_win(scan_win2294), .scan_win_std_dev(scan_win_std_dev[2294]), .feature_accum(feature_accums[2294]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2295]), .RECT1_Y(rectangle1_ys[2295]), .RECT1_WIDTH(rectangle1_widths[2295]), .RECT1_HEIGHT(rectangle1_heights[2295]), .RECT1_WEIGHT(rectangle1_weights[2295]), .RECT2_X(rectangle2_xs[2295]), .RECT2_Y(rectangle2_ys[2295]), .RECT2_WIDTH(rectangle2_widths[2295]), .RECT2_HEIGHT(rectangle2_heights[2295]), .RECT2_WEIGHT(rectangle2_weights[2295]), .RECT3_X(rectangle3_xs[2295]), .RECT3_Y(rectangle3_ys[2295]), .RECT3_WIDTH(rectangle3_widths[2295]), .RECT3_HEIGHT(rectangle3_heights[2295]), .RECT3_WEIGHT(rectangle3_weights[2295]), .FEAT_THRES(feature_thresholds[2295]), .FEAT_ABOVE(feature_aboves[2295]), .FEAT_BELOW(feature_belows[2295])) ac2295(.scan_win(scan_win2295), .scan_win_std_dev(scan_win_std_dev[2295]), .feature_accum(feature_accums[2295]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2296]), .RECT1_Y(rectangle1_ys[2296]), .RECT1_WIDTH(rectangle1_widths[2296]), .RECT1_HEIGHT(rectangle1_heights[2296]), .RECT1_WEIGHT(rectangle1_weights[2296]), .RECT2_X(rectangle2_xs[2296]), .RECT2_Y(rectangle2_ys[2296]), .RECT2_WIDTH(rectangle2_widths[2296]), .RECT2_HEIGHT(rectangle2_heights[2296]), .RECT2_WEIGHT(rectangle2_weights[2296]), .RECT3_X(rectangle3_xs[2296]), .RECT3_Y(rectangle3_ys[2296]), .RECT3_WIDTH(rectangle3_widths[2296]), .RECT3_HEIGHT(rectangle3_heights[2296]), .RECT3_WEIGHT(rectangle3_weights[2296]), .FEAT_THRES(feature_thresholds[2296]), .FEAT_ABOVE(feature_aboves[2296]), .FEAT_BELOW(feature_belows[2296])) ac2296(.scan_win(scan_win2296), .scan_win_std_dev(scan_win_std_dev[2296]), .feature_accum(feature_accums[2296]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2297]), .RECT1_Y(rectangle1_ys[2297]), .RECT1_WIDTH(rectangle1_widths[2297]), .RECT1_HEIGHT(rectangle1_heights[2297]), .RECT1_WEIGHT(rectangle1_weights[2297]), .RECT2_X(rectangle2_xs[2297]), .RECT2_Y(rectangle2_ys[2297]), .RECT2_WIDTH(rectangle2_widths[2297]), .RECT2_HEIGHT(rectangle2_heights[2297]), .RECT2_WEIGHT(rectangle2_weights[2297]), .RECT3_X(rectangle3_xs[2297]), .RECT3_Y(rectangle3_ys[2297]), .RECT3_WIDTH(rectangle3_widths[2297]), .RECT3_HEIGHT(rectangle3_heights[2297]), .RECT3_WEIGHT(rectangle3_weights[2297]), .FEAT_THRES(feature_thresholds[2297]), .FEAT_ABOVE(feature_aboves[2297]), .FEAT_BELOW(feature_belows[2297])) ac2297(.scan_win(scan_win2297), .scan_win_std_dev(scan_win_std_dev[2297]), .feature_accum(feature_accums[2297]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2298]), .RECT1_Y(rectangle1_ys[2298]), .RECT1_WIDTH(rectangle1_widths[2298]), .RECT1_HEIGHT(rectangle1_heights[2298]), .RECT1_WEIGHT(rectangle1_weights[2298]), .RECT2_X(rectangle2_xs[2298]), .RECT2_Y(rectangle2_ys[2298]), .RECT2_WIDTH(rectangle2_widths[2298]), .RECT2_HEIGHT(rectangle2_heights[2298]), .RECT2_WEIGHT(rectangle2_weights[2298]), .RECT3_X(rectangle3_xs[2298]), .RECT3_Y(rectangle3_ys[2298]), .RECT3_WIDTH(rectangle3_widths[2298]), .RECT3_HEIGHT(rectangle3_heights[2298]), .RECT3_WEIGHT(rectangle3_weights[2298]), .FEAT_THRES(feature_thresholds[2298]), .FEAT_ABOVE(feature_aboves[2298]), .FEAT_BELOW(feature_belows[2298])) ac2298(.scan_win(scan_win2298), .scan_win_std_dev(scan_win_std_dev[2298]), .feature_accum(feature_accums[2298]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2299]), .RECT1_Y(rectangle1_ys[2299]), .RECT1_WIDTH(rectangle1_widths[2299]), .RECT1_HEIGHT(rectangle1_heights[2299]), .RECT1_WEIGHT(rectangle1_weights[2299]), .RECT2_X(rectangle2_xs[2299]), .RECT2_Y(rectangle2_ys[2299]), .RECT2_WIDTH(rectangle2_widths[2299]), .RECT2_HEIGHT(rectangle2_heights[2299]), .RECT2_WEIGHT(rectangle2_weights[2299]), .RECT3_X(rectangle3_xs[2299]), .RECT3_Y(rectangle3_ys[2299]), .RECT3_WIDTH(rectangle3_widths[2299]), .RECT3_HEIGHT(rectangle3_heights[2299]), .RECT3_WEIGHT(rectangle3_weights[2299]), .FEAT_THRES(feature_thresholds[2299]), .FEAT_ABOVE(feature_aboves[2299]), .FEAT_BELOW(feature_belows[2299])) ac2299(.scan_win(scan_win2299), .scan_win_std_dev(scan_win_std_dev[2299]), .feature_accum(feature_accums[2299]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2300]), .RECT1_Y(rectangle1_ys[2300]), .RECT1_WIDTH(rectangle1_widths[2300]), .RECT1_HEIGHT(rectangle1_heights[2300]), .RECT1_WEIGHT(rectangle1_weights[2300]), .RECT2_X(rectangle2_xs[2300]), .RECT2_Y(rectangle2_ys[2300]), .RECT2_WIDTH(rectangle2_widths[2300]), .RECT2_HEIGHT(rectangle2_heights[2300]), .RECT2_WEIGHT(rectangle2_weights[2300]), .RECT3_X(rectangle3_xs[2300]), .RECT3_Y(rectangle3_ys[2300]), .RECT3_WIDTH(rectangle3_widths[2300]), .RECT3_HEIGHT(rectangle3_heights[2300]), .RECT3_WEIGHT(rectangle3_weights[2300]), .FEAT_THRES(feature_thresholds[2300]), .FEAT_ABOVE(feature_aboves[2300]), .FEAT_BELOW(feature_belows[2300])) ac2300(.scan_win(scan_win2300), .scan_win_std_dev(scan_win_std_dev[2300]), .feature_accum(feature_accums[2300]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2301]), .RECT1_Y(rectangle1_ys[2301]), .RECT1_WIDTH(rectangle1_widths[2301]), .RECT1_HEIGHT(rectangle1_heights[2301]), .RECT1_WEIGHT(rectangle1_weights[2301]), .RECT2_X(rectangle2_xs[2301]), .RECT2_Y(rectangle2_ys[2301]), .RECT2_WIDTH(rectangle2_widths[2301]), .RECT2_HEIGHT(rectangle2_heights[2301]), .RECT2_WEIGHT(rectangle2_weights[2301]), .RECT3_X(rectangle3_xs[2301]), .RECT3_Y(rectangle3_ys[2301]), .RECT3_WIDTH(rectangle3_widths[2301]), .RECT3_HEIGHT(rectangle3_heights[2301]), .RECT3_WEIGHT(rectangle3_weights[2301]), .FEAT_THRES(feature_thresholds[2301]), .FEAT_ABOVE(feature_aboves[2301]), .FEAT_BELOW(feature_belows[2301])) ac2301(.scan_win(scan_win2301), .scan_win_std_dev(scan_win_std_dev[2301]), .feature_accum(feature_accums[2301]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2302]), .RECT1_Y(rectangle1_ys[2302]), .RECT1_WIDTH(rectangle1_widths[2302]), .RECT1_HEIGHT(rectangle1_heights[2302]), .RECT1_WEIGHT(rectangle1_weights[2302]), .RECT2_X(rectangle2_xs[2302]), .RECT2_Y(rectangle2_ys[2302]), .RECT2_WIDTH(rectangle2_widths[2302]), .RECT2_HEIGHT(rectangle2_heights[2302]), .RECT2_WEIGHT(rectangle2_weights[2302]), .RECT3_X(rectangle3_xs[2302]), .RECT3_Y(rectangle3_ys[2302]), .RECT3_WIDTH(rectangle3_widths[2302]), .RECT3_HEIGHT(rectangle3_heights[2302]), .RECT3_WEIGHT(rectangle3_weights[2302]), .FEAT_THRES(feature_thresholds[2302]), .FEAT_ABOVE(feature_aboves[2302]), .FEAT_BELOW(feature_belows[2302])) ac2302(.scan_win(scan_win2302), .scan_win_std_dev(scan_win_std_dev[2302]), .feature_accum(feature_accums[2302]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2303]), .RECT1_Y(rectangle1_ys[2303]), .RECT1_WIDTH(rectangle1_widths[2303]), .RECT1_HEIGHT(rectangle1_heights[2303]), .RECT1_WEIGHT(rectangle1_weights[2303]), .RECT2_X(rectangle2_xs[2303]), .RECT2_Y(rectangle2_ys[2303]), .RECT2_WIDTH(rectangle2_widths[2303]), .RECT2_HEIGHT(rectangle2_heights[2303]), .RECT2_WEIGHT(rectangle2_weights[2303]), .RECT3_X(rectangle3_xs[2303]), .RECT3_Y(rectangle3_ys[2303]), .RECT3_WIDTH(rectangle3_widths[2303]), .RECT3_HEIGHT(rectangle3_heights[2303]), .RECT3_WEIGHT(rectangle3_weights[2303]), .FEAT_THRES(feature_thresholds[2303]), .FEAT_ABOVE(feature_aboves[2303]), .FEAT_BELOW(feature_belows[2303])) ac2303(.scan_win(scan_win2303), .scan_win_std_dev(scan_win_std_dev[2303]), .feature_accum(feature_accums[2303]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2304]), .RECT1_Y(rectangle1_ys[2304]), .RECT1_WIDTH(rectangle1_widths[2304]), .RECT1_HEIGHT(rectangle1_heights[2304]), .RECT1_WEIGHT(rectangle1_weights[2304]), .RECT2_X(rectangle2_xs[2304]), .RECT2_Y(rectangle2_ys[2304]), .RECT2_WIDTH(rectangle2_widths[2304]), .RECT2_HEIGHT(rectangle2_heights[2304]), .RECT2_WEIGHT(rectangle2_weights[2304]), .RECT3_X(rectangle3_xs[2304]), .RECT3_Y(rectangle3_ys[2304]), .RECT3_WIDTH(rectangle3_widths[2304]), .RECT3_HEIGHT(rectangle3_heights[2304]), .RECT3_WEIGHT(rectangle3_weights[2304]), .FEAT_THRES(feature_thresholds[2304]), .FEAT_ABOVE(feature_aboves[2304]), .FEAT_BELOW(feature_belows[2304])) ac2304(.scan_win(scan_win2304), .scan_win_std_dev(scan_win_std_dev[2304]), .feature_accum(feature_accums[2304]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2305]), .RECT1_Y(rectangle1_ys[2305]), .RECT1_WIDTH(rectangle1_widths[2305]), .RECT1_HEIGHT(rectangle1_heights[2305]), .RECT1_WEIGHT(rectangle1_weights[2305]), .RECT2_X(rectangle2_xs[2305]), .RECT2_Y(rectangle2_ys[2305]), .RECT2_WIDTH(rectangle2_widths[2305]), .RECT2_HEIGHT(rectangle2_heights[2305]), .RECT2_WEIGHT(rectangle2_weights[2305]), .RECT3_X(rectangle3_xs[2305]), .RECT3_Y(rectangle3_ys[2305]), .RECT3_WIDTH(rectangle3_widths[2305]), .RECT3_HEIGHT(rectangle3_heights[2305]), .RECT3_WEIGHT(rectangle3_weights[2305]), .FEAT_THRES(feature_thresholds[2305]), .FEAT_ABOVE(feature_aboves[2305]), .FEAT_BELOW(feature_belows[2305])) ac2305(.scan_win(scan_win2305), .scan_win_std_dev(scan_win_std_dev[2305]), .feature_accum(feature_accums[2305]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2306]), .RECT1_Y(rectangle1_ys[2306]), .RECT1_WIDTH(rectangle1_widths[2306]), .RECT1_HEIGHT(rectangle1_heights[2306]), .RECT1_WEIGHT(rectangle1_weights[2306]), .RECT2_X(rectangle2_xs[2306]), .RECT2_Y(rectangle2_ys[2306]), .RECT2_WIDTH(rectangle2_widths[2306]), .RECT2_HEIGHT(rectangle2_heights[2306]), .RECT2_WEIGHT(rectangle2_weights[2306]), .RECT3_X(rectangle3_xs[2306]), .RECT3_Y(rectangle3_ys[2306]), .RECT3_WIDTH(rectangle3_widths[2306]), .RECT3_HEIGHT(rectangle3_heights[2306]), .RECT3_WEIGHT(rectangle3_weights[2306]), .FEAT_THRES(feature_thresholds[2306]), .FEAT_ABOVE(feature_aboves[2306]), .FEAT_BELOW(feature_belows[2306])) ac2306(.scan_win(scan_win2306), .scan_win_std_dev(scan_win_std_dev[2306]), .feature_accum(feature_accums[2306]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2307]), .RECT1_Y(rectangle1_ys[2307]), .RECT1_WIDTH(rectangle1_widths[2307]), .RECT1_HEIGHT(rectangle1_heights[2307]), .RECT1_WEIGHT(rectangle1_weights[2307]), .RECT2_X(rectangle2_xs[2307]), .RECT2_Y(rectangle2_ys[2307]), .RECT2_WIDTH(rectangle2_widths[2307]), .RECT2_HEIGHT(rectangle2_heights[2307]), .RECT2_WEIGHT(rectangle2_weights[2307]), .RECT3_X(rectangle3_xs[2307]), .RECT3_Y(rectangle3_ys[2307]), .RECT3_WIDTH(rectangle3_widths[2307]), .RECT3_HEIGHT(rectangle3_heights[2307]), .RECT3_WEIGHT(rectangle3_weights[2307]), .FEAT_THRES(feature_thresholds[2307]), .FEAT_ABOVE(feature_aboves[2307]), .FEAT_BELOW(feature_belows[2307])) ac2307(.scan_win(scan_win2307), .scan_win_std_dev(scan_win_std_dev[2307]), .feature_accum(feature_accums[2307]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2308]), .RECT1_Y(rectangle1_ys[2308]), .RECT1_WIDTH(rectangle1_widths[2308]), .RECT1_HEIGHT(rectangle1_heights[2308]), .RECT1_WEIGHT(rectangle1_weights[2308]), .RECT2_X(rectangle2_xs[2308]), .RECT2_Y(rectangle2_ys[2308]), .RECT2_WIDTH(rectangle2_widths[2308]), .RECT2_HEIGHT(rectangle2_heights[2308]), .RECT2_WEIGHT(rectangle2_weights[2308]), .RECT3_X(rectangle3_xs[2308]), .RECT3_Y(rectangle3_ys[2308]), .RECT3_WIDTH(rectangle3_widths[2308]), .RECT3_HEIGHT(rectangle3_heights[2308]), .RECT3_WEIGHT(rectangle3_weights[2308]), .FEAT_THRES(feature_thresholds[2308]), .FEAT_ABOVE(feature_aboves[2308]), .FEAT_BELOW(feature_belows[2308])) ac2308(.scan_win(scan_win2308), .scan_win_std_dev(scan_win_std_dev[2308]), .feature_accum(feature_accums[2308]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2309]), .RECT1_Y(rectangle1_ys[2309]), .RECT1_WIDTH(rectangle1_widths[2309]), .RECT1_HEIGHT(rectangle1_heights[2309]), .RECT1_WEIGHT(rectangle1_weights[2309]), .RECT2_X(rectangle2_xs[2309]), .RECT2_Y(rectangle2_ys[2309]), .RECT2_WIDTH(rectangle2_widths[2309]), .RECT2_HEIGHT(rectangle2_heights[2309]), .RECT2_WEIGHT(rectangle2_weights[2309]), .RECT3_X(rectangle3_xs[2309]), .RECT3_Y(rectangle3_ys[2309]), .RECT3_WIDTH(rectangle3_widths[2309]), .RECT3_HEIGHT(rectangle3_heights[2309]), .RECT3_WEIGHT(rectangle3_weights[2309]), .FEAT_THRES(feature_thresholds[2309]), .FEAT_ABOVE(feature_aboves[2309]), .FEAT_BELOW(feature_belows[2309])) ac2309(.scan_win(scan_win2309), .scan_win_std_dev(scan_win_std_dev[2309]), .feature_accum(feature_accums[2309]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2310]), .RECT1_Y(rectangle1_ys[2310]), .RECT1_WIDTH(rectangle1_widths[2310]), .RECT1_HEIGHT(rectangle1_heights[2310]), .RECT1_WEIGHT(rectangle1_weights[2310]), .RECT2_X(rectangle2_xs[2310]), .RECT2_Y(rectangle2_ys[2310]), .RECT2_WIDTH(rectangle2_widths[2310]), .RECT2_HEIGHT(rectangle2_heights[2310]), .RECT2_WEIGHT(rectangle2_weights[2310]), .RECT3_X(rectangle3_xs[2310]), .RECT3_Y(rectangle3_ys[2310]), .RECT3_WIDTH(rectangle3_widths[2310]), .RECT3_HEIGHT(rectangle3_heights[2310]), .RECT3_WEIGHT(rectangle3_weights[2310]), .FEAT_THRES(feature_thresholds[2310]), .FEAT_ABOVE(feature_aboves[2310]), .FEAT_BELOW(feature_belows[2310])) ac2310(.scan_win(scan_win2310), .scan_win_std_dev(scan_win_std_dev[2310]), .feature_accum(feature_accums[2310]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2311]), .RECT1_Y(rectangle1_ys[2311]), .RECT1_WIDTH(rectangle1_widths[2311]), .RECT1_HEIGHT(rectangle1_heights[2311]), .RECT1_WEIGHT(rectangle1_weights[2311]), .RECT2_X(rectangle2_xs[2311]), .RECT2_Y(rectangle2_ys[2311]), .RECT2_WIDTH(rectangle2_widths[2311]), .RECT2_HEIGHT(rectangle2_heights[2311]), .RECT2_WEIGHT(rectangle2_weights[2311]), .RECT3_X(rectangle3_xs[2311]), .RECT3_Y(rectangle3_ys[2311]), .RECT3_WIDTH(rectangle3_widths[2311]), .RECT3_HEIGHT(rectangle3_heights[2311]), .RECT3_WEIGHT(rectangle3_weights[2311]), .FEAT_THRES(feature_thresholds[2311]), .FEAT_ABOVE(feature_aboves[2311]), .FEAT_BELOW(feature_belows[2311])) ac2311(.scan_win(scan_win2311), .scan_win_std_dev(scan_win_std_dev[2311]), .feature_accum(feature_accums[2311]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2312]), .RECT1_Y(rectangle1_ys[2312]), .RECT1_WIDTH(rectangle1_widths[2312]), .RECT1_HEIGHT(rectangle1_heights[2312]), .RECT1_WEIGHT(rectangle1_weights[2312]), .RECT2_X(rectangle2_xs[2312]), .RECT2_Y(rectangle2_ys[2312]), .RECT2_WIDTH(rectangle2_widths[2312]), .RECT2_HEIGHT(rectangle2_heights[2312]), .RECT2_WEIGHT(rectangle2_weights[2312]), .RECT3_X(rectangle3_xs[2312]), .RECT3_Y(rectangle3_ys[2312]), .RECT3_WIDTH(rectangle3_widths[2312]), .RECT3_HEIGHT(rectangle3_heights[2312]), .RECT3_WEIGHT(rectangle3_weights[2312]), .FEAT_THRES(feature_thresholds[2312]), .FEAT_ABOVE(feature_aboves[2312]), .FEAT_BELOW(feature_belows[2312])) ac2312(.scan_win(scan_win2312), .scan_win_std_dev(scan_win_std_dev[2312]), .feature_accum(feature_accums[2312]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2313]), .RECT1_Y(rectangle1_ys[2313]), .RECT1_WIDTH(rectangle1_widths[2313]), .RECT1_HEIGHT(rectangle1_heights[2313]), .RECT1_WEIGHT(rectangle1_weights[2313]), .RECT2_X(rectangle2_xs[2313]), .RECT2_Y(rectangle2_ys[2313]), .RECT2_WIDTH(rectangle2_widths[2313]), .RECT2_HEIGHT(rectangle2_heights[2313]), .RECT2_WEIGHT(rectangle2_weights[2313]), .RECT3_X(rectangle3_xs[2313]), .RECT3_Y(rectangle3_ys[2313]), .RECT3_WIDTH(rectangle3_widths[2313]), .RECT3_HEIGHT(rectangle3_heights[2313]), .RECT3_WEIGHT(rectangle3_weights[2313]), .FEAT_THRES(feature_thresholds[2313]), .FEAT_ABOVE(feature_aboves[2313]), .FEAT_BELOW(feature_belows[2313])) ac2313(.scan_win(scan_win2313), .scan_win_std_dev(scan_win_std_dev[2313]), .feature_accum(feature_accums[2313]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2314]), .RECT1_Y(rectangle1_ys[2314]), .RECT1_WIDTH(rectangle1_widths[2314]), .RECT1_HEIGHT(rectangle1_heights[2314]), .RECT1_WEIGHT(rectangle1_weights[2314]), .RECT2_X(rectangle2_xs[2314]), .RECT2_Y(rectangle2_ys[2314]), .RECT2_WIDTH(rectangle2_widths[2314]), .RECT2_HEIGHT(rectangle2_heights[2314]), .RECT2_WEIGHT(rectangle2_weights[2314]), .RECT3_X(rectangle3_xs[2314]), .RECT3_Y(rectangle3_ys[2314]), .RECT3_WIDTH(rectangle3_widths[2314]), .RECT3_HEIGHT(rectangle3_heights[2314]), .RECT3_WEIGHT(rectangle3_weights[2314]), .FEAT_THRES(feature_thresholds[2314]), .FEAT_ABOVE(feature_aboves[2314]), .FEAT_BELOW(feature_belows[2314])) ac2314(.scan_win(scan_win2314), .scan_win_std_dev(scan_win_std_dev[2314]), .feature_accum(feature_accums[2314]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2315]), .RECT1_Y(rectangle1_ys[2315]), .RECT1_WIDTH(rectangle1_widths[2315]), .RECT1_HEIGHT(rectangle1_heights[2315]), .RECT1_WEIGHT(rectangle1_weights[2315]), .RECT2_X(rectangle2_xs[2315]), .RECT2_Y(rectangle2_ys[2315]), .RECT2_WIDTH(rectangle2_widths[2315]), .RECT2_HEIGHT(rectangle2_heights[2315]), .RECT2_WEIGHT(rectangle2_weights[2315]), .RECT3_X(rectangle3_xs[2315]), .RECT3_Y(rectangle3_ys[2315]), .RECT3_WIDTH(rectangle3_widths[2315]), .RECT3_HEIGHT(rectangle3_heights[2315]), .RECT3_WEIGHT(rectangle3_weights[2315]), .FEAT_THRES(feature_thresholds[2315]), .FEAT_ABOVE(feature_aboves[2315]), .FEAT_BELOW(feature_belows[2315])) ac2315(.scan_win(scan_win2315), .scan_win_std_dev(scan_win_std_dev[2315]), .feature_accum(feature_accums[2315]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2316]), .RECT1_Y(rectangle1_ys[2316]), .RECT1_WIDTH(rectangle1_widths[2316]), .RECT1_HEIGHT(rectangle1_heights[2316]), .RECT1_WEIGHT(rectangle1_weights[2316]), .RECT2_X(rectangle2_xs[2316]), .RECT2_Y(rectangle2_ys[2316]), .RECT2_WIDTH(rectangle2_widths[2316]), .RECT2_HEIGHT(rectangle2_heights[2316]), .RECT2_WEIGHT(rectangle2_weights[2316]), .RECT3_X(rectangle3_xs[2316]), .RECT3_Y(rectangle3_ys[2316]), .RECT3_WIDTH(rectangle3_widths[2316]), .RECT3_HEIGHT(rectangle3_heights[2316]), .RECT3_WEIGHT(rectangle3_weights[2316]), .FEAT_THRES(feature_thresholds[2316]), .FEAT_ABOVE(feature_aboves[2316]), .FEAT_BELOW(feature_belows[2316])) ac2316(.scan_win(scan_win2316), .scan_win_std_dev(scan_win_std_dev[2316]), .feature_accum(feature_accums[2316]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2317]), .RECT1_Y(rectangle1_ys[2317]), .RECT1_WIDTH(rectangle1_widths[2317]), .RECT1_HEIGHT(rectangle1_heights[2317]), .RECT1_WEIGHT(rectangle1_weights[2317]), .RECT2_X(rectangle2_xs[2317]), .RECT2_Y(rectangle2_ys[2317]), .RECT2_WIDTH(rectangle2_widths[2317]), .RECT2_HEIGHT(rectangle2_heights[2317]), .RECT2_WEIGHT(rectangle2_weights[2317]), .RECT3_X(rectangle3_xs[2317]), .RECT3_Y(rectangle3_ys[2317]), .RECT3_WIDTH(rectangle3_widths[2317]), .RECT3_HEIGHT(rectangle3_heights[2317]), .RECT3_WEIGHT(rectangle3_weights[2317]), .FEAT_THRES(feature_thresholds[2317]), .FEAT_ABOVE(feature_aboves[2317]), .FEAT_BELOW(feature_belows[2317])) ac2317(.scan_win(scan_win2317), .scan_win_std_dev(scan_win_std_dev[2317]), .feature_accum(feature_accums[2317]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2318]), .RECT1_Y(rectangle1_ys[2318]), .RECT1_WIDTH(rectangle1_widths[2318]), .RECT1_HEIGHT(rectangle1_heights[2318]), .RECT1_WEIGHT(rectangle1_weights[2318]), .RECT2_X(rectangle2_xs[2318]), .RECT2_Y(rectangle2_ys[2318]), .RECT2_WIDTH(rectangle2_widths[2318]), .RECT2_HEIGHT(rectangle2_heights[2318]), .RECT2_WEIGHT(rectangle2_weights[2318]), .RECT3_X(rectangle3_xs[2318]), .RECT3_Y(rectangle3_ys[2318]), .RECT3_WIDTH(rectangle3_widths[2318]), .RECT3_HEIGHT(rectangle3_heights[2318]), .RECT3_WEIGHT(rectangle3_weights[2318]), .FEAT_THRES(feature_thresholds[2318]), .FEAT_ABOVE(feature_aboves[2318]), .FEAT_BELOW(feature_belows[2318])) ac2318(.scan_win(scan_win2318), .scan_win_std_dev(scan_win_std_dev[2318]), .feature_accum(feature_accums[2318]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2319]), .RECT1_Y(rectangle1_ys[2319]), .RECT1_WIDTH(rectangle1_widths[2319]), .RECT1_HEIGHT(rectangle1_heights[2319]), .RECT1_WEIGHT(rectangle1_weights[2319]), .RECT2_X(rectangle2_xs[2319]), .RECT2_Y(rectangle2_ys[2319]), .RECT2_WIDTH(rectangle2_widths[2319]), .RECT2_HEIGHT(rectangle2_heights[2319]), .RECT2_WEIGHT(rectangle2_weights[2319]), .RECT3_X(rectangle3_xs[2319]), .RECT3_Y(rectangle3_ys[2319]), .RECT3_WIDTH(rectangle3_widths[2319]), .RECT3_HEIGHT(rectangle3_heights[2319]), .RECT3_WEIGHT(rectangle3_weights[2319]), .FEAT_THRES(feature_thresholds[2319]), .FEAT_ABOVE(feature_aboves[2319]), .FEAT_BELOW(feature_belows[2319])) ac2319(.scan_win(scan_win2319), .scan_win_std_dev(scan_win_std_dev[2319]), .feature_accum(feature_accums[2319]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2320]), .RECT1_Y(rectangle1_ys[2320]), .RECT1_WIDTH(rectangle1_widths[2320]), .RECT1_HEIGHT(rectangle1_heights[2320]), .RECT1_WEIGHT(rectangle1_weights[2320]), .RECT2_X(rectangle2_xs[2320]), .RECT2_Y(rectangle2_ys[2320]), .RECT2_WIDTH(rectangle2_widths[2320]), .RECT2_HEIGHT(rectangle2_heights[2320]), .RECT2_WEIGHT(rectangle2_weights[2320]), .RECT3_X(rectangle3_xs[2320]), .RECT3_Y(rectangle3_ys[2320]), .RECT3_WIDTH(rectangle3_widths[2320]), .RECT3_HEIGHT(rectangle3_heights[2320]), .RECT3_WEIGHT(rectangle3_weights[2320]), .FEAT_THRES(feature_thresholds[2320]), .FEAT_ABOVE(feature_aboves[2320]), .FEAT_BELOW(feature_belows[2320])) ac2320(.scan_win(scan_win2320), .scan_win_std_dev(scan_win_std_dev[2320]), .feature_accum(feature_accums[2320]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2321]), .RECT1_Y(rectangle1_ys[2321]), .RECT1_WIDTH(rectangle1_widths[2321]), .RECT1_HEIGHT(rectangle1_heights[2321]), .RECT1_WEIGHT(rectangle1_weights[2321]), .RECT2_X(rectangle2_xs[2321]), .RECT2_Y(rectangle2_ys[2321]), .RECT2_WIDTH(rectangle2_widths[2321]), .RECT2_HEIGHT(rectangle2_heights[2321]), .RECT2_WEIGHT(rectangle2_weights[2321]), .RECT3_X(rectangle3_xs[2321]), .RECT3_Y(rectangle3_ys[2321]), .RECT3_WIDTH(rectangle3_widths[2321]), .RECT3_HEIGHT(rectangle3_heights[2321]), .RECT3_WEIGHT(rectangle3_weights[2321]), .FEAT_THRES(feature_thresholds[2321]), .FEAT_ABOVE(feature_aboves[2321]), .FEAT_BELOW(feature_belows[2321])) ac2321(.scan_win(scan_win2321), .scan_win_std_dev(scan_win_std_dev[2321]), .feature_accum(feature_accums[2321]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2322]), .RECT1_Y(rectangle1_ys[2322]), .RECT1_WIDTH(rectangle1_widths[2322]), .RECT1_HEIGHT(rectangle1_heights[2322]), .RECT1_WEIGHT(rectangle1_weights[2322]), .RECT2_X(rectangle2_xs[2322]), .RECT2_Y(rectangle2_ys[2322]), .RECT2_WIDTH(rectangle2_widths[2322]), .RECT2_HEIGHT(rectangle2_heights[2322]), .RECT2_WEIGHT(rectangle2_weights[2322]), .RECT3_X(rectangle3_xs[2322]), .RECT3_Y(rectangle3_ys[2322]), .RECT3_WIDTH(rectangle3_widths[2322]), .RECT3_HEIGHT(rectangle3_heights[2322]), .RECT3_WEIGHT(rectangle3_weights[2322]), .FEAT_THRES(feature_thresholds[2322]), .FEAT_ABOVE(feature_aboves[2322]), .FEAT_BELOW(feature_belows[2322])) ac2322(.scan_win(scan_win2322), .scan_win_std_dev(scan_win_std_dev[2322]), .feature_accum(feature_accums[2322]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2323]), .RECT1_Y(rectangle1_ys[2323]), .RECT1_WIDTH(rectangle1_widths[2323]), .RECT1_HEIGHT(rectangle1_heights[2323]), .RECT1_WEIGHT(rectangle1_weights[2323]), .RECT2_X(rectangle2_xs[2323]), .RECT2_Y(rectangle2_ys[2323]), .RECT2_WIDTH(rectangle2_widths[2323]), .RECT2_HEIGHT(rectangle2_heights[2323]), .RECT2_WEIGHT(rectangle2_weights[2323]), .RECT3_X(rectangle3_xs[2323]), .RECT3_Y(rectangle3_ys[2323]), .RECT3_WIDTH(rectangle3_widths[2323]), .RECT3_HEIGHT(rectangle3_heights[2323]), .RECT3_WEIGHT(rectangle3_weights[2323]), .FEAT_THRES(feature_thresholds[2323]), .FEAT_ABOVE(feature_aboves[2323]), .FEAT_BELOW(feature_belows[2323])) ac2323(.scan_win(scan_win2323), .scan_win_std_dev(scan_win_std_dev[2323]), .feature_accum(feature_accums[2323]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2324]), .RECT1_Y(rectangle1_ys[2324]), .RECT1_WIDTH(rectangle1_widths[2324]), .RECT1_HEIGHT(rectangle1_heights[2324]), .RECT1_WEIGHT(rectangle1_weights[2324]), .RECT2_X(rectangle2_xs[2324]), .RECT2_Y(rectangle2_ys[2324]), .RECT2_WIDTH(rectangle2_widths[2324]), .RECT2_HEIGHT(rectangle2_heights[2324]), .RECT2_WEIGHT(rectangle2_weights[2324]), .RECT3_X(rectangle3_xs[2324]), .RECT3_Y(rectangle3_ys[2324]), .RECT3_WIDTH(rectangle3_widths[2324]), .RECT3_HEIGHT(rectangle3_heights[2324]), .RECT3_WEIGHT(rectangle3_weights[2324]), .FEAT_THRES(feature_thresholds[2324]), .FEAT_ABOVE(feature_aboves[2324]), .FEAT_BELOW(feature_belows[2324])) ac2324(.scan_win(scan_win2324), .scan_win_std_dev(scan_win_std_dev[2324]), .feature_accum(feature_accums[2324]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2325]), .RECT1_Y(rectangle1_ys[2325]), .RECT1_WIDTH(rectangle1_widths[2325]), .RECT1_HEIGHT(rectangle1_heights[2325]), .RECT1_WEIGHT(rectangle1_weights[2325]), .RECT2_X(rectangle2_xs[2325]), .RECT2_Y(rectangle2_ys[2325]), .RECT2_WIDTH(rectangle2_widths[2325]), .RECT2_HEIGHT(rectangle2_heights[2325]), .RECT2_WEIGHT(rectangle2_weights[2325]), .RECT3_X(rectangle3_xs[2325]), .RECT3_Y(rectangle3_ys[2325]), .RECT3_WIDTH(rectangle3_widths[2325]), .RECT3_HEIGHT(rectangle3_heights[2325]), .RECT3_WEIGHT(rectangle3_weights[2325]), .FEAT_THRES(feature_thresholds[2325]), .FEAT_ABOVE(feature_aboves[2325]), .FEAT_BELOW(feature_belows[2325])) ac2325(.scan_win(scan_win2325), .scan_win_std_dev(scan_win_std_dev[2325]), .feature_accum(feature_accums[2325]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2326]), .RECT1_Y(rectangle1_ys[2326]), .RECT1_WIDTH(rectangle1_widths[2326]), .RECT1_HEIGHT(rectangle1_heights[2326]), .RECT1_WEIGHT(rectangle1_weights[2326]), .RECT2_X(rectangle2_xs[2326]), .RECT2_Y(rectangle2_ys[2326]), .RECT2_WIDTH(rectangle2_widths[2326]), .RECT2_HEIGHT(rectangle2_heights[2326]), .RECT2_WEIGHT(rectangle2_weights[2326]), .RECT3_X(rectangle3_xs[2326]), .RECT3_Y(rectangle3_ys[2326]), .RECT3_WIDTH(rectangle3_widths[2326]), .RECT3_HEIGHT(rectangle3_heights[2326]), .RECT3_WEIGHT(rectangle3_weights[2326]), .FEAT_THRES(feature_thresholds[2326]), .FEAT_ABOVE(feature_aboves[2326]), .FEAT_BELOW(feature_belows[2326])) ac2326(.scan_win(scan_win2326), .scan_win_std_dev(scan_win_std_dev[2326]), .feature_accum(feature_accums[2326]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2327]), .RECT1_Y(rectangle1_ys[2327]), .RECT1_WIDTH(rectangle1_widths[2327]), .RECT1_HEIGHT(rectangle1_heights[2327]), .RECT1_WEIGHT(rectangle1_weights[2327]), .RECT2_X(rectangle2_xs[2327]), .RECT2_Y(rectangle2_ys[2327]), .RECT2_WIDTH(rectangle2_widths[2327]), .RECT2_HEIGHT(rectangle2_heights[2327]), .RECT2_WEIGHT(rectangle2_weights[2327]), .RECT3_X(rectangle3_xs[2327]), .RECT3_Y(rectangle3_ys[2327]), .RECT3_WIDTH(rectangle3_widths[2327]), .RECT3_HEIGHT(rectangle3_heights[2327]), .RECT3_WEIGHT(rectangle3_weights[2327]), .FEAT_THRES(feature_thresholds[2327]), .FEAT_ABOVE(feature_aboves[2327]), .FEAT_BELOW(feature_belows[2327])) ac2327(.scan_win(scan_win2327), .scan_win_std_dev(scan_win_std_dev[2327]), .feature_accum(feature_accums[2327]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2328]), .RECT1_Y(rectangle1_ys[2328]), .RECT1_WIDTH(rectangle1_widths[2328]), .RECT1_HEIGHT(rectangle1_heights[2328]), .RECT1_WEIGHT(rectangle1_weights[2328]), .RECT2_X(rectangle2_xs[2328]), .RECT2_Y(rectangle2_ys[2328]), .RECT2_WIDTH(rectangle2_widths[2328]), .RECT2_HEIGHT(rectangle2_heights[2328]), .RECT2_WEIGHT(rectangle2_weights[2328]), .RECT3_X(rectangle3_xs[2328]), .RECT3_Y(rectangle3_ys[2328]), .RECT3_WIDTH(rectangle3_widths[2328]), .RECT3_HEIGHT(rectangle3_heights[2328]), .RECT3_WEIGHT(rectangle3_weights[2328]), .FEAT_THRES(feature_thresholds[2328]), .FEAT_ABOVE(feature_aboves[2328]), .FEAT_BELOW(feature_belows[2328])) ac2328(.scan_win(scan_win2328), .scan_win_std_dev(scan_win_std_dev[2328]), .feature_accum(feature_accums[2328]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2329]), .RECT1_Y(rectangle1_ys[2329]), .RECT1_WIDTH(rectangle1_widths[2329]), .RECT1_HEIGHT(rectangle1_heights[2329]), .RECT1_WEIGHT(rectangle1_weights[2329]), .RECT2_X(rectangle2_xs[2329]), .RECT2_Y(rectangle2_ys[2329]), .RECT2_WIDTH(rectangle2_widths[2329]), .RECT2_HEIGHT(rectangle2_heights[2329]), .RECT2_WEIGHT(rectangle2_weights[2329]), .RECT3_X(rectangle3_xs[2329]), .RECT3_Y(rectangle3_ys[2329]), .RECT3_WIDTH(rectangle3_widths[2329]), .RECT3_HEIGHT(rectangle3_heights[2329]), .RECT3_WEIGHT(rectangle3_weights[2329]), .FEAT_THRES(feature_thresholds[2329]), .FEAT_ABOVE(feature_aboves[2329]), .FEAT_BELOW(feature_belows[2329])) ac2329(.scan_win(scan_win2329), .scan_win_std_dev(scan_win_std_dev[2329]), .feature_accum(feature_accums[2329]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2330]), .RECT1_Y(rectangle1_ys[2330]), .RECT1_WIDTH(rectangle1_widths[2330]), .RECT1_HEIGHT(rectangle1_heights[2330]), .RECT1_WEIGHT(rectangle1_weights[2330]), .RECT2_X(rectangle2_xs[2330]), .RECT2_Y(rectangle2_ys[2330]), .RECT2_WIDTH(rectangle2_widths[2330]), .RECT2_HEIGHT(rectangle2_heights[2330]), .RECT2_WEIGHT(rectangle2_weights[2330]), .RECT3_X(rectangle3_xs[2330]), .RECT3_Y(rectangle3_ys[2330]), .RECT3_WIDTH(rectangle3_widths[2330]), .RECT3_HEIGHT(rectangle3_heights[2330]), .RECT3_WEIGHT(rectangle3_weights[2330]), .FEAT_THRES(feature_thresholds[2330]), .FEAT_ABOVE(feature_aboves[2330]), .FEAT_BELOW(feature_belows[2330])) ac2330(.scan_win(scan_win2330), .scan_win_std_dev(scan_win_std_dev[2330]), .feature_accum(feature_accums[2330]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2331]), .RECT1_Y(rectangle1_ys[2331]), .RECT1_WIDTH(rectangle1_widths[2331]), .RECT1_HEIGHT(rectangle1_heights[2331]), .RECT1_WEIGHT(rectangle1_weights[2331]), .RECT2_X(rectangle2_xs[2331]), .RECT2_Y(rectangle2_ys[2331]), .RECT2_WIDTH(rectangle2_widths[2331]), .RECT2_HEIGHT(rectangle2_heights[2331]), .RECT2_WEIGHT(rectangle2_weights[2331]), .RECT3_X(rectangle3_xs[2331]), .RECT3_Y(rectangle3_ys[2331]), .RECT3_WIDTH(rectangle3_widths[2331]), .RECT3_HEIGHT(rectangle3_heights[2331]), .RECT3_WEIGHT(rectangle3_weights[2331]), .FEAT_THRES(feature_thresholds[2331]), .FEAT_ABOVE(feature_aboves[2331]), .FEAT_BELOW(feature_belows[2331])) ac2331(.scan_win(scan_win2331), .scan_win_std_dev(scan_win_std_dev[2331]), .feature_accum(feature_accums[2331]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2332]), .RECT1_Y(rectangle1_ys[2332]), .RECT1_WIDTH(rectangle1_widths[2332]), .RECT1_HEIGHT(rectangle1_heights[2332]), .RECT1_WEIGHT(rectangle1_weights[2332]), .RECT2_X(rectangle2_xs[2332]), .RECT2_Y(rectangle2_ys[2332]), .RECT2_WIDTH(rectangle2_widths[2332]), .RECT2_HEIGHT(rectangle2_heights[2332]), .RECT2_WEIGHT(rectangle2_weights[2332]), .RECT3_X(rectangle3_xs[2332]), .RECT3_Y(rectangle3_ys[2332]), .RECT3_WIDTH(rectangle3_widths[2332]), .RECT3_HEIGHT(rectangle3_heights[2332]), .RECT3_WEIGHT(rectangle3_weights[2332]), .FEAT_THRES(feature_thresholds[2332]), .FEAT_ABOVE(feature_aboves[2332]), .FEAT_BELOW(feature_belows[2332])) ac2332(.scan_win(scan_win2332), .scan_win_std_dev(scan_win_std_dev[2332]), .feature_accum(feature_accums[2332]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2333]), .RECT1_Y(rectangle1_ys[2333]), .RECT1_WIDTH(rectangle1_widths[2333]), .RECT1_HEIGHT(rectangle1_heights[2333]), .RECT1_WEIGHT(rectangle1_weights[2333]), .RECT2_X(rectangle2_xs[2333]), .RECT2_Y(rectangle2_ys[2333]), .RECT2_WIDTH(rectangle2_widths[2333]), .RECT2_HEIGHT(rectangle2_heights[2333]), .RECT2_WEIGHT(rectangle2_weights[2333]), .RECT3_X(rectangle3_xs[2333]), .RECT3_Y(rectangle3_ys[2333]), .RECT3_WIDTH(rectangle3_widths[2333]), .RECT3_HEIGHT(rectangle3_heights[2333]), .RECT3_WEIGHT(rectangle3_weights[2333]), .FEAT_THRES(feature_thresholds[2333]), .FEAT_ABOVE(feature_aboves[2333]), .FEAT_BELOW(feature_belows[2333])) ac2333(.scan_win(scan_win2333), .scan_win_std_dev(scan_win_std_dev[2333]), .feature_accum(feature_accums[2333]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2334]), .RECT1_Y(rectangle1_ys[2334]), .RECT1_WIDTH(rectangle1_widths[2334]), .RECT1_HEIGHT(rectangle1_heights[2334]), .RECT1_WEIGHT(rectangle1_weights[2334]), .RECT2_X(rectangle2_xs[2334]), .RECT2_Y(rectangle2_ys[2334]), .RECT2_WIDTH(rectangle2_widths[2334]), .RECT2_HEIGHT(rectangle2_heights[2334]), .RECT2_WEIGHT(rectangle2_weights[2334]), .RECT3_X(rectangle3_xs[2334]), .RECT3_Y(rectangle3_ys[2334]), .RECT3_WIDTH(rectangle3_widths[2334]), .RECT3_HEIGHT(rectangle3_heights[2334]), .RECT3_WEIGHT(rectangle3_weights[2334]), .FEAT_THRES(feature_thresholds[2334]), .FEAT_ABOVE(feature_aboves[2334]), .FEAT_BELOW(feature_belows[2334])) ac2334(.scan_win(scan_win2334), .scan_win_std_dev(scan_win_std_dev[2334]), .feature_accum(feature_accums[2334]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2335]), .RECT1_Y(rectangle1_ys[2335]), .RECT1_WIDTH(rectangle1_widths[2335]), .RECT1_HEIGHT(rectangle1_heights[2335]), .RECT1_WEIGHT(rectangle1_weights[2335]), .RECT2_X(rectangle2_xs[2335]), .RECT2_Y(rectangle2_ys[2335]), .RECT2_WIDTH(rectangle2_widths[2335]), .RECT2_HEIGHT(rectangle2_heights[2335]), .RECT2_WEIGHT(rectangle2_weights[2335]), .RECT3_X(rectangle3_xs[2335]), .RECT3_Y(rectangle3_ys[2335]), .RECT3_WIDTH(rectangle3_widths[2335]), .RECT3_HEIGHT(rectangle3_heights[2335]), .RECT3_WEIGHT(rectangle3_weights[2335]), .FEAT_THRES(feature_thresholds[2335]), .FEAT_ABOVE(feature_aboves[2335]), .FEAT_BELOW(feature_belows[2335])) ac2335(.scan_win(scan_win2335), .scan_win_std_dev(scan_win_std_dev[2335]), .feature_accum(feature_accums[2335]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2336]), .RECT1_Y(rectangle1_ys[2336]), .RECT1_WIDTH(rectangle1_widths[2336]), .RECT1_HEIGHT(rectangle1_heights[2336]), .RECT1_WEIGHT(rectangle1_weights[2336]), .RECT2_X(rectangle2_xs[2336]), .RECT2_Y(rectangle2_ys[2336]), .RECT2_WIDTH(rectangle2_widths[2336]), .RECT2_HEIGHT(rectangle2_heights[2336]), .RECT2_WEIGHT(rectangle2_weights[2336]), .RECT3_X(rectangle3_xs[2336]), .RECT3_Y(rectangle3_ys[2336]), .RECT3_WIDTH(rectangle3_widths[2336]), .RECT3_HEIGHT(rectangle3_heights[2336]), .RECT3_WEIGHT(rectangle3_weights[2336]), .FEAT_THRES(feature_thresholds[2336]), .FEAT_ABOVE(feature_aboves[2336]), .FEAT_BELOW(feature_belows[2336])) ac2336(.scan_win(scan_win2336), .scan_win_std_dev(scan_win_std_dev[2336]), .feature_accum(feature_accums[2336]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2337]), .RECT1_Y(rectangle1_ys[2337]), .RECT1_WIDTH(rectangle1_widths[2337]), .RECT1_HEIGHT(rectangle1_heights[2337]), .RECT1_WEIGHT(rectangle1_weights[2337]), .RECT2_X(rectangle2_xs[2337]), .RECT2_Y(rectangle2_ys[2337]), .RECT2_WIDTH(rectangle2_widths[2337]), .RECT2_HEIGHT(rectangle2_heights[2337]), .RECT2_WEIGHT(rectangle2_weights[2337]), .RECT3_X(rectangle3_xs[2337]), .RECT3_Y(rectangle3_ys[2337]), .RECT3_WIDTH(rectangle3_widths[2337]), .RECT3_HEIGHT(rectangle3_heights[2337]), .RECT3_WEIGHT(rectangle3_weights[2337]), .FEAT_THRES(feature_thresholds[2337]), .FEAT_ABOVE(feature_aboves[2337]), .FEAT_BELOW(feature_belows[2337])) ac2337(.scan_win(scan_win2337), .scan_win_std_dev(scan_win_std_dev[2337]), .feature_accum(feature_accums[2337]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2338]), .RECT1_Y(rectangle1_ys[2338]), .RECT1_WIDTH(rectangle1_widths[2338]), .RECT1_HEIGHT(rectangle1_heights[2338]), .RECT1_WEIGHT(rectangle1_weights[2338]), .RECT2_X(rectangle2_xs[2338]), .RECT2_Y(rectangle2_ys[2338]), .RECT2_WIDTH(rectangle2_widths[2338]), .RECT2_HEIGHT(rectangle2_heights[2338]), .RECT2_WEIGHT(rectangle2_weights[2338]), .RECT3_X(rectangle3_xs[2338]), .RECT3_Y(rectangle3_ys[2338]), .RECT3_WIDTH(rectangle3_widths[2338]), .RECT3_HEIGHT(rectangle3_heights[2338]), .RECT3_WEIGHT(rectangle3_weights[2338]), .FEAT_THRES(feature_thresholds[2338]), .FEAT_ABOVE(feature_aboves[2338]), .FEAT_BELOW(feature_belows[2338])) ac2338(.scan_win(scan_win2338), .scan_win_std_dev(scan_win_std_dev[2338]), .feature_accum(feature_accums[2338]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2339]), .RECT1_Y(rectangle1_ys[2339]), .RECT1_WIDTH(rectangle1_widths[2339]), .RECT1_HEIGHT(rectangle1_heights[2339]), .RECT1_WEIGHT(rectangle1_weights[2339]), .RECT2_X(rectangle2_xs[2339]), .RECT2_Y(rectangle2_ys[2339]), .RECT2_WIDTH(rectangle2_widths[2339]), .RECT2_HEIGHT(rectangle2_heights[2339]), .RECT2_WEIGHT(rectangle2_weights[2339]), .RECT3_X(rectangle3_xs[2339]), .RECT3_Y(rectangle3_ys[2339]), .RECT3_WIDTH(rectangle3_widths[2339]), .RECT3_HEIGHT(rectangle3_heights[2339]), .RECT3_WEIGHT(rectangle3_weights[2339]), .FEAT_THRES(feature_thresholds[2339]), .FEAT_ABOVE(feature_aboves[2339]), .FEAT_BELOW(feature_belows[2339])) ac2339(.scan_win(scan_win2339), .scan_win_std_dev(scan_win_std_dev[2339]), .feature_accum(feature_accums[2339]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2340]), .RECT1_Y(rectangle1_ys[2340]), .RECT1_WIDTH(rectangle1_widths[2340]), .RECT1_HEIGHT(rectangle1_heights[2340]), .RECT1_WEIGHT(rectangle1_weights[2340]), .RECT2_X(rectangle2_xs[2340]), .RECT2_Y(rectangle2_ys[2340]), .RECT2_WIDTH(rectangle2_widths[2340]), .RECT2_HEIGHT(rectangle2_heights[2340]), .RECT2_WEIGHT(rectangle2_weights[2340]), .RECT3_X(rectangle3_xs[2340]), .RECT3_Y(rectangle3_ys[2340]), .RECT3_WIDTH(rectangle3_widths[2340]), .RECT3_HEIGHT(rectangle3_heights[2340]), .RECT3_WEIGHT(rectangle3_weights[2340]), .FEAT_THRES(feature_thresholds[2340]), .FEAT_ABOVE(feature_aboves[2340]), .FEAT_BELOW(feature_belows[2340])) ac2340(.scan_win(scan_win2340), .scan_win_std_dev(scan_win_std_dev[2340]), .feature_accum(feature_accums[2340]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2341]), .RECT1_Y(rectangle1_ys[2341]), .RECT1_WIDTH(rectangle1_widths[2341]), .RECT1_HEIGHT(rectangle1_heights[2341]), .RECT1_WEIGHT(rectangle1_weights[2341]), .RECT2_X(rectangle2_xs[2341]), .RECT2_Y(rectangle2_ys[2341]), .RECT2_WIDTH(rectangle2_widths[2341]), .RECT2_HEIGHT(rectangle2_heights[2341]), .RECT2_WEIGHT(rectangle2_weights[2341]), .RECT3_X(rectangle3_xs[2341]), .RECT3_Y(rectangle3_ys[2341]), .RECT3_WIDTH(rectangle3_widths[2341]), .RECT3_HEIGHT(rectangle3_heights[2341]), .RECT3_WEIGHT(rectangle3_weights[2341]), .FEAT_THRES(feature_thresholds[2341]), .FEAT_ABOVE(feature_aboves[2341]), .FEAT_BELOW(feature_belows[2341])) ac2341(.scan_win(scan_win2341), .scan_win_std_dev(scan_win_std_dev[2341]), .feature_accum(feature_accums[2341]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2342]), .RECT1_Y(rectangle1_ys[2342]), .RECT1_WIDTH(rectangle1_widths[2342]), .RECT1_HEIGHT(rectangle1_heights[2342]), .RECT1_WEIGHT(rectangle1_weights[2342]), .RECT2_X(rectangle2_xs[2342]), .RECT2_Y(rectangle2_ys[2342]), .RECT2_WIDTH(rectangle2_widths[2342]), .RECT2_HEIGHT(rectangle2_heights[2342]), .RECT2_WEIGHT(rectangle2_weights[2342]), .RECT3_X(rectangle3_xs[2342]), .RECT3_Y(rectangle3_ys[2342]), .RECT3_WIDTH(rectangle3_widths[2342]), .RECT3_HEIGHT(rectangle3_heights[2342]), .RECT3_WEIGHT(rectangle3_weights[2342]), .FEAT_THRES(feature_thresholds[2342]), .FEAT_ABOVE(feature_aboves[2342]), .FEAT_BELOW(feature_belows[2342])) ac2342(.scan_win(scan_win2342), .scan_win_std_dev(scan_win_std_dev[2342]), .feature_accum(feature_accums[2342]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2343]), .RECT1_Y(rectangle1_ys[2343]), .RECT1_WIDTH(rectangle1_widths[2343]), .RECT1_HEIGHT(rectangle1_heights[2343]), .RECT1_WEIGHT(rectangle1_weights[2343]), .RECT2_X(rectangle2_xs[2343]), .RECT2_Y(rectangle2_ys[2343]), .RECT2_WIDTH(rectangle2_widths[2343]), .RECT2_HEIGHT(rectangle2_heights[2343]), .RECT2_WEIGHT(rectangle2_weights[2343]), .RECT3_X(rectangle3_xs[2343]), .RECT3_Y(rectangle3_ys[2343]), .RECT3_WIDTH(rectangle3_widths[2343]), .RECT3_HEIGHT(rectangle3_heights[2343]), .RECT3_WEIGHT(rectangle3_weights[2343]), .FEAT_THRES(feature_thresholds[2343]), .FEAT_ABOVE(feature_aboves[2343]), .FEAT_BELOW(feature_belows[2343])) ac2343(.scan_win(scan_win2343), .scan_win_std_dev(scan_win_std_dev[2343]), .feature_accum(feature_accums[2343]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2344]), .RECT1_Y(rectangle1_ys[2344]), .RECT1_WIDTH(rectangle1_widths[2344]), .RECT1_HEIGHT(rectangle1_heights[2344]), .RECT1_WEIGHT(rectangle1_weights[2344]), .RECT2_X(rectangle2_xs[2344]), .RECT2_Y(rectangle2_ys[2344]), .RECT2_WIDTH(rectangle2_widths[2344]), .RECT2_HEIGHT(rectangle2_heights[2344]), .RECT2_WEIGHT(rectangle2_weights[2344]), .RECT3_X(rectangle3_xs[2344]), .RECT3_Y(rectangle3_ys[2344]), .RECT3_WIDTH(rectangle3_widths[2344]), .RECT3_HEIGHT(rectangle3_heights[2344]), .RECT3_WEIGHT(rectangle3_weights[2344]), .FEAT_THRES(feature_thresholds[2344]), .FEAT_ABOVE(feature_aboves[2344]), .FEAT_BELOW(feature_belows[2344])) ac2344(.scan_win(scan_win2344), .scan_win_std_dev(scan_win_std_dev[2344]), .feature_accum(feature_accums[2344]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2345]), .RECT1_Y(rectangle1_ys[2345]), .RECT1_WIDTH(rectangle1_widths[2345]), .RECT1_HEIGHT(rectangle1_heights[2345]), .RECT1_WEIGHT(rectangle1_weights[2345]), .RECT2_X(rectangle2_xs[2345]), .RECT2_Y(rectangle2_ys[2345]), .RECT2_WIDTH(rectangle2_widths[2345]), .RECT2_HEIGHT(rectangle2_heights[2345]), .RECT2_WEIGHT(rectangle2_weights[2345]), .RECT3_X(rectangle3_xs[2345]), .RECT3_Y(rectangle3_ys[2345]), .RECT3_WIDTH(rectangle3_widths[2345]), .RECT3_HEIGHT(rectangle3_heights[2345]), .RECT3_WEIGHT(rectangle3_weights[2345]), .FEAT_THRES(feature_thresholds[2345]), .FEAT_ABOVE(feature_aboves[2345]), .FEAT_BELOW(feature_belows[2345])) ac2345(.scan_win(scan_win2345), .scan_win_std_dev(scan_win_std_dev[2345]), .feature_accum(feature_accums[2345]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2346]), .RECT1_Y(rectangle1_ys[2346]), .RECT1_WIDTH(rectangle1_widths[2346]), .RECT1_HEIGHT(rectangle1_heights[2346]), .RECT1_WEIGHT(rectangle1_weights[2346]), .RECT2_X(rectangle2_xs[2346]), .RECT2_Y(rectangle2_ys[2346]), .RECT2_WIDTH(rectangle2_widths[2346]), .RECT2_HEIGHT(rectangle2_heights[2346]), .RECT2_WEIGHT(rectangle2_weights[2346]), .RECT3_X(rectangle3_xs[2346]), .RECT3_Y(rectangle3_ys[2346]), .RECT3_WIDTH(rectangle3_widths[2346]), .RECT3_HEIGHT(rectangle3_heights[2346]), .RECT3_WEIGHT(rectangle3_weights[2346]), .FEAT_THRES(feature_thresholds[2346]), .FEAT_ABOVE(feature_aboves[2346]), .FEAT_BELOW(feature_belows[2346])) ac2346(.scan_win(scan_win2346), .scan_win_std_dev(scan_win_std_dev[2346]), .feature_accum(feature_accums[2346]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2347]), .RECT1_Y(rectangle1_ys[2347]), .RECT1_WIDTH(rectangle1_widths[2347]), .RECT1_HEIGHT(rectangle1_heights[2347]), .RECT1_WEIGHT(rectangle1_weights[2347]), .RECT2_X(rectangle2_xs[2347]), .RECT2_Y(rectangle2_ys[2347]), .RECT2_WIDTH(rectangle2_widths[2347]), .RECT2_HEIGHT(rectangle2_heights[2347]), .RECT2_WEIGHT(rectangle2_weights[2347]), .RECT3_X(rectangle3_xs[2347]), .RECT3_Y(rectangle3_ys[2347]), .RECT3_WIDTH(rectangle3_widths[2347]), .RECT3_HEIGHT(rectangle3_heights[2347]), .RECT3_WEIGHT(rectangle3_weights[2347]), .FEAT_THRES(feature_thresholds[2347]), .FEAT_ABOVE(feature_aboves[2347]), .FEAT_BELOW(feature_belows[2347])) ac2347(.scan_win(scan_win2347), .scan_win_std_dev(scan_win_std_dev[2347]), .feature_accum(feature_accums[2347]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2348]), .RECT1_Y(rectangle1_ys[2348]), .RECT1_WIDTH(rectangle1_widths[2348]), .RECT1_HEIGHT(rectangle1_heights[2348]), .RECT1_WEIGHT(rectangle1_weights[2348]), .RECT2_X(rectangle2_xs[2348]), .RECT2_Y(rectangle2_ys[2348]), .RECT2_WIDTH(rectangle2_widths[2348]), .RECT2_HEIGHT(rectangle2_heights[2348]), .RECT2_WEIGHT(rectangle2_weights[2348]), .RECT3_X(rectangle3_xs[2348]), .RECT3_Y(rectangle3_ys[2348]), .RECT3_WIDTH(rectangle3_widths[2348]), .RECT3_HEIGHT(rectangle3_heights[2348]), .RECT3_WEIGHT(rectangle3_weights[2348]), .FEAT_THRES(feature_thresholds[2348]), .FEAT_ABOVE(feature_aboves[2348]), .FEAT_BELOW(feature_belows[2348])) ac2348(.scan_win(scan_win2348), .scan_win_std_dev(scan_win_std_dev[2348]), .feature_accum(feature_accums[2348]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2349]), .RECT1_Y(rectangle1_ys[2349]), .RECT1_WIDTH(rectangle1_widths[2349]), .RECT1_HEIGHT(rectangle1_heights[2349]), .RECT1_WEIGHT(rectangle1_weights[2349]), .RECT2_X(rectangle2_xs[2349]), .RECT2_Y(rectangle2_ys[2349]), .RECT2_WIDTH(rectangle2_widths[2349]), .RECT2_HEIGHT(rectangle2_heights[2349]), .RECT2_WEIGHT(rectangle2_weights[2349]), .RECT3_X(rectangle3_xs[2349]), .RECT3_Y(rectangle3_ys[2349]), .RECT3_WIDTH(rectangle3_widths[2349]), .RECT3_HEIGHT(rectangle3_heights[2349]), .RECT3_WEIGHT(rectangle3_weights[2349]), .FEAT_THRES(feature_thresholds[2349]), .FEAT_ABOVE(feature_aboves[2349]), .FEAT_BELOW(feature_belows[2349])) ac2349(.scan_win(scan_win2349), .scan_win_std_dev(scan_win_std_dev[2349]), .feature_accum(feature_accums[2349]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2350]), .RECT1_Y(rectangle1_ys[2350]), .RECT1_WIDTH(rectangle1_widths[2350]), .RECT1_HEIGHT(rectangle1_heights[2350]), .RECT1_WEIGHT(rectangle1_weights[2350]), .RECT2_X(rectangle2_xs[2350]), .RECT2_Y(rectangle2_ys[2350]), .RECT2_WIDTH(rectangle2_widths[2350]), .RECT2_HEIGHT(rectangle2_heights[2350]), .RECT2_WEIGHT(rectangle2_weights[2350]), .RECT3_X(rectangle3_xs[2350]), .RECT3_Y(rectangle3_ys[2350]), .RECT3_WIDTH(rectangle3_widths[2350]), .RECT3_HEIGHT(rectangle3_heights[2350]), .RECT3_WEIGHT(rectangle3_weights[2350]), .FEAT_THRES(feature_thresholds[2350]), .FEAT_ABOVE(feature_aboves[2350]), .FEAT_BELOW(feature_belows[2350])) ac2350(.scan_win(scan_win2350), .scan_win_std_dev(scan_win_std_dev[2350]), .feature_accum(feature_accums[2350]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2351]), .RECT1_Y(rectangle1_ys[2351]), .RECT1_WIDTH(rectangle1_widths[2351]), .RECT1_HEIGHT(rectangle1_heights[2351]), .RECT1_WEIGHT(rectangle1_weights[2351]), .RECT2_X(rectangle2_xs[2351]), .RECT2_Y(rectangle2_ys[2351]), .RECT2_WIDTH(rectangle2_widths[2351]), .RECT2_HEIGHT(rectangle2_heights[2351]), .RECT2_WEIGHT(rectangle2_weights[2351]), .RECT3_X(rectangle3_xs[2351]), .RECT3_Y(rectangle3_ys[2351]), .RECT3_WIDTH(rectangle3_widths[2351]), .RECT3_HEIGHT(rectangle3_heights[2351]), .RECT3_WEIGHT(rectangle3_weights[2351]), .FEAT_THRES(feature_thresholds[2351]), .FEAT_ABOVE(feature_aboves[2351]), .FEAT_BELOW(feature_belows[2351])) ac2351(.scan_win(scan_win2351), .scan_win_std_dev(scan_win_std_dev[2351]), .feature_accum(feature_accums[2351]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2352]), .RECT1_Y(rectangle1_ys[2352]), .RECT1_WIDTH(rectangle1_widths[2352]), .RECT1_HEIGHT(rectangle1_heights[2352]), .RECT1_WEIGHT(rectangle1_weights[2352]), .RECT2_X(rectangle2_xs[2352]), .RECT2_Y(rectangle2_ys[2352]), .RECT2_WIDTH(rectangle2_widths[2352]), .RECT2_HEIGHT(rectangle2_heights[2352]), .RECT2_WEIGHT(rectangle2_weights[2352]), .RECT3_X(rectangle3_xs[2352]), .RECT3_Y(rectangle3_ys[2352]), .RECT3_WIDTH(rectangle3_widths[2352]), .RECT3_HEIGHT(rectangle3_heights[2352]), .RECT3_WEIGHT(rectangle3_weights[2352]), .FEAT_THRES(feature_thresholds[2352]), .FEAT_ABOVE(feature_aboves[2352]), .FEAT_BELOW(feature_belows[2352])) ac2352(.scan_win(scan_win2352), .scan_win_std_dev(scan_win_std_dev[2352]), .feature_accum(feature_accums[2352]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2353]), .RECT1_Y(rectangle1_ys[2353]), .RECT1_WIDTH(rectangle1_widths[2353]), .RECT1_HEIGHT(rectangle1_heights[2353]), .RECT1_WEIGHT(rectangle1_weights[2353]), .RECT2_X(rectangle2_xs[2353]), .RECT2_Y(rectangle2_ys[2353]), .RECT2_WIDTH(rectangle2_widths[2353]), .RECT2_HEIGHT(rectangle2_heights[2353]), .RECT2_WEIGHT(rectangle2_weights[2353]), .RECT3_X(rectangle3_xs[2353]), .RECT3_Y(rectangle3_ys[2353]), .RECT3_WIDTH(rectangle3_widths[2353]), .RECT3_HEIGHT(rectangle3_heights[2353]), .RECT3_WEIGHT(rectangle3_weights[2353]), .FEAT_THRES(feature_thresholds[2353]), .FEAT_ABOVE(feature_aboves[2353]), .FEAT_BELOW(feature_belows[2353])) ac2353(.scan_win(scan_win2353), .scan_win_std_dev(scan_win_std_dev[2353]), .feature_accum(feature_accums[2353]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2354]), .RECT1_Y(rectangle1_ys[2354]), .RECT1_WIDTH(rectangle1_widths[2354]), .RECT1_HEIGHT(rectangle1_heights[2354]), .RECT1_WEIGHT(rectangle1_weights[2354]), .RECT2_X(rectangle2_xs[2354]), .RECT2_Y(rectangle2_ys[2354]), .RECT2_WIDTH(rectangle2_widths[2354]), .RECT2_HEIGHT(rectangle2_heights[2354]), .RECT2_WEIGHT(rectangle2_weights[2354]), .RECT3_X(rectangle3_xs[2354]), .RECT3_Y(rectangle3_ys[2354]), .RECT3_WIDTH(rectangle3_widths[2354]), .RECT3_HEIGHT(rectangle3_heights[2354]), .RECT3_WEIGHT(rectangle3_weights[2354]), .FEAT_THRES(feature_thresholds[2354]), .FEAT_ABOVE(feature_aboves[2354]), .FEAT_BELOW(feature_belows[2354])) ac2354(.scan_win(scan_win2354), .scan_win_std_dev(scan_win_std_dev[2354]), .feature_accum(feature_accums[2354]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2355]), .RECT1_Y(rectangle1_ys[2355]), .RECT1_WIDTH(rectangle1_widths[2355]), .RECT1_HEIGHT(rectangle1_heights[2355]), .RECT1_WEIGHT(rectangle1_weights[2355]), .RECT2_X(rectangle2_xs[2355]), .RECT2_Y(rectangle2_ys[2355]), .RECT2_WIDTH(rectangle2_widths[2355]), .RECT2_HEIGHT(rectangle2_heights[2355]), .RECT2_WEIGHT(rectangle2_weights[2355]), .RECT3_X(rectangle3_xs[2355]), .RECT3_Y(rectangle3_ys[2355]), .RECT3_WIDTH(rectangle3_widths[2355]), .RECT3_HEIGHT(rectangle3_heights[2355]), .RECT3_WEIGHT(rectangle3_weights[2355]), .FEAT_THRES(feature_thresholds[2355]), .FEAT_ABOVE(feature_aboves[2355]), .FEAT_BELOW(feature_belows[2355])) ac2355(.scan_win(scan_win2355), .scan_win_std_dev(scan_win_std_dev[2355]), .feature_accum(feature_accums[2355]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2356]), .RECT1_Y(rectangle1_ys[2356]), .RECT1_WIDTH(rectangle1_widths[2356]), .RECT1_HEIGHT(rectangle1_heights[2356]), .RECT1_WEIGHT(rectangle1_weights[2356]), .RECT2_X(rectangle2_xs[2356]), .RECT2_Y(rectangle2_ys[2356]), .RECT2_WIDTH(rectangle2_widths[2356]), .RECT2_HEIGHT(rectangle2_heights[2356]), .RECT2_WEIGHT(rectangle2_weights[2356]), .RECT3_X(rectangle3_xs[2356]), .RECT3_Y(rectangle3_ys[2356]), .RECT3_WIDTH(rectangle3_widths[2356]), .RECT3_HEIGHT(rectangle3_heights[2356]), .RECT3_WEIGHT(rectangle3_weights[2356]), .FEAT_THRES(feature_thresholds[2356]), .FEAT_ABOVE(feature_aboves[2356]), .FEAT_BELOW(feature_belows[2356])) ac2356(.scan_win(scan_win2356), .scan_win_std_dev(scan_win_std_dev[2356]), .feature_accum(feature_accums[2356]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2357]), .RECT1_Y(rectangle1_ys[2357]), .RECT1_WIDTH(rectangle1_widths[2357]), .RECT1_HEIGHT(rectangle1_heights[2357]), .RECT1_WEIGHT(rectangle1_weights[2357]), .RECT2_X(rectangle2_xs[2357]), .RECT2_Y(rectangle2_ys[2357]), .RECT2_WIDTH(rectangle2_widths[2357]), .RECT2_HEIGHT(rectangle2_heights[2357]), .RECT2_WEIGHT(rectangle2_weights[2357]), .RECT3_X(rectangle3_xs[2357]), .RECT3_Y(rectangle3_ys[2357]), .RECT3_WIDTH(rectangle3_widths[2357]), .RECT3_HEIGHT(rectangle3_heights[2357]), .RECT3_WEIGHT(rectangle3_weights[2357]), .FEAT_THRES(feature_thresholds[2357]), .FEAT_ABOVE(feature_aboves[2357]), .FEAT_BELOW(feature_belows[2357])) ac2357(.scan_win(scan_win2357), .scan_win_std_dev(scan_win_std_dev[2357]), .feature_accum(feature_accums[2357]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2358]), .RECT1_Y(rectangle1_ys[2358]), .RECT1_WIDTH(rectangle1_widths[2358]), .RECT1_HEIGHT(rectangle1_heights[2358]), .RECT1_WEIGHT(rectangle1_weights[2358]), .RECT2_X(rectangle2_xs[2358]), .RECT2_Y(rectangle2_ys[2358]), .RECT2_WIDTH(rectangle2_widths[2358]), .RECT2_HEIGHT(rectangle2_heights[2358]), .RECT2_WEIGHT(rectangle2_weights[2358]), .RECT3_X(rectangle3_xs[2358]), .RECT3_Y(rectangle3_ys[2358]), .RECT3_WIDTH(rectangle3_widths[2358]), .RECT3_HEIGHT(rectangle3_heights[2358]), .RECT3_WEIGHT(rectangle3_weights[2358]), .FEAT_THRES(feature_thresholds[2358]), .FEAT_ABOVE(feature_aboves[2358]), .FEAT_BELOW(feature_belows[2358])) ac2358(.scan_win(scan_win2358), .scan_win_std_dev(scan_win_std_dev[2358]), .feature_accum(feature_accums[2358]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2359]), .RECT1_Y(rectangle1_ys[2359]), .RECT1_WIDTH(rectangle1_widths[2359]), .RECT1_HEIGHT(rectangle1_heights[2359]), .RECT1_WEIGHT(rectangle1_weights[2359]), .RECT2_X(rectangle2_xs[2359]), .RECT2_Y(rectangle2_ys[2359]), .RECT2_WIDTH(rectangle2_widths[2359]), .RECT2_HEIGHT(rectangle2_heights[2359]), .RECT2_WEIGHT(rectangle2_weights[2359]), .RECT3_X(rectangle3_xs[2359]), .RECT3_Y(rectangle3_ys[2359]), .RECT3_WIDTH(rectangle3_widths[2359]), .RECT3_HEIGHT(rectangle3_heights[2359]), .RECT3_WEIGHT(rectangle3_weights[2359]), .FEAT_THRES(feature_thresholds[2359]), .FEAT_ABOVE(feature_aboves[2359]), .FEAT_BELOW(feature_belows[2359])) ac2359(.scan_win(scan_win2359), .scan_win_std_dev(scan_win_std_dev[2359]), .feature_accum(feature_accums[2359]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2360]), .RECT1_Y(rectangle1_ys[2360]), .RECT1_WIDTH(rectangle1_widths[2360]), .RECT1_HEIGHT(rectangle1_heights[2360]), .RECT1_WEIGHT(rectangle1_weights[2360]), .RECT2_X(rectangle2_xs[2360]), .RECT2_Y(rectangle2_ys[2360]), .RECT2_WIDTH(rectangle2_widths[2360]), .RECT2_HEIGHT(rectangle2_heights[2360]), .RECT2_WEIGHT(rectangle2_weights[2360]), .RECT3_X(rectangle3_xs[2360]), .RECT3_Y(rectangle3_ys[2360]), .RECT3_WIDTH(rectangle3_widths[2360]), .RECT3_HEIGHT(rectangle3_heights[2360]), .RECT3_WEIGHT(rectangle3_weights[2360]), .FEAT_THRES(feature_thresholds[2360]), .FEAT_ABOVE(feature_aboves[2360]), .FEAT_BELOW(feature_belows[2360])) ac2360(.scan_win(scan_win2360), .scan_win_std_dev(scan_win_std_dev[2360]), .feature_accum(feature_accums[2360]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2361]), .RECT1_Y(rectangle1_ys[2361]), .RECT1_WIDTH(rectangle1_widths[2361]), .RECT1_HEIGHT(rectangle1_heights[2361]), .RECT1_WEIGHT(rectangle1_weights[2361]), .RECT2_X(rectangle2_xs[2361]), .RECT2_Y(rectangle2_ys[2361]), .RECT2_WIDTH(rectangle2_widths[2361]), .RECT2_HEIGHT(rectangle2_heights[2361]), .RECT2_WEIGHT(rectangle2_weights[2361]), .RECT3_X(rectangle3_xs[2361]), .RECT3_Y(rectangle3_ys[2361]), .RECT3_WIDTH(rectangle3_widths[2361]), .RECT3_HEIGHT(rectangle3_heights[2361]), .RECT3_WEIGHT(rectangle3_weights[2361]), .FEAT_THRES(feature_thresholds[2361]), .FEAT_ABOVE(feature_aboves[2361]), .FEAT_BELOW(feature_belows[2361])) ac2361(.scan_win(scan_win2361), .scan_win_std_dev(scan_win_std_dev[2361]), .feature_accum(feature_accums[2361]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2362]), .RECT1_Y(rectangle1_ys[2362]), .RECT1_WIDTH(rectangle1_widths[2362]), .RECT1_HEIGHT(rectangle1_heights[2362]), .RECT1_WEIGHT(rectangle1_weights[2362]), .RECT2_X(rectangle2_xs[2362]), .RECT2_Y(rectangle2_ys[2362]), .RECT2_WIDTH(rectangle2_widths[2362]), .RECT2_HEIGHT(rectangle2_heights[2362]), .RECT2_WEIGHT(rectangle2_weights[2362]), .RECT3_X(rectangle3_xs[2362]), .RECT3_Y(rectangle3_ys[2362]), .RECT3_WIDTH(rectangle3_widths[2362]), .RECT3_HEIGHT(rectangle3_heights[2362]), .RECT3_WEIGHT(rectangle3_weights[2362]), .FEAT_THRES(feature_thresholds[2362]), .FEAT_ABOVE(feature_aboves[2362]), .FEAT_BELOW(feature_belows[2362])) ac2362(.scan_win(scan_win2362), .scan_win_std_dev(scan_win_std_dev[2362]), .feature_accum(feature_accums[2362]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2363]), .RECT1_Y(rectangle1_ys[2363]), .RECT1_WIDTH(rectangle1_widths[2363]), .RECT1_HEIGHT(rectangle1_heights[2363]), .RECT1_WEIGHT(rectangle1_weights[2363]), .RECT2_X(rectangle2_xs[2363]), .RECT2_Y(rectangle2_ys[2363]), .RECT2_WIDTH(rectangle2_widths[2363]), .RECT2_HEIGHT(rectangle2_heights[2363]), .RECT2_WEIGHT(rectangle2_weights[2363]), .RECT3_X(rectangle3_xs[2363]), .RECT3_Y(rectangle3_ys[2363]), .RECT3_WIDTH(rectangle3_widths[2363]), .RECT3_HEIGHT(rectangle3_heights[2363]), .RECT3_WEIGHT(rectangle3_weights[2363]), .FEAT_THRES(feature_thresholds[2363]), .FEAT_ABOVE(feature_aboves[2363]), .FEAT_BELOW(feature_belows[2363])) ac2363(.scan_win(scan_win2363), .scan_win_std_dev(scan_win_std_dev[2363]), .feature_accum(feature_accums[2363]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2364]), .RECT1_Y(rectangle1_ys[2364]), .RECT1_WIDTH(rectangle1_widths[2364]), .RECT1_HEIGHT(rectangle1_heights[2364]), .RECT1_WEIGHT(rectangle1_weights[2364]), .RECT2_X(rectangle2_xs[2364]), .RECT2_Y(rectangle2_ys[2364]), .RECT2_WIDTH(rectangle2_widths[2364]), .RECT2_HEIGHT(rectangle2_heights[2364]), .RECT2_WEIGHT(rectangle2_weights[2364]), .RECT3_X(rectangle3_xs[2364]), .RECT3_Y(rectangle3_ys[2364]), .RECT3_WIDTH(rectangle3_widths[2364]), .RECT3_HEIGHT(rectangle3_heights[2364]), .RECT3_WEIGHT(rectangle3_weights[2364]), .FEAT_THRES(feature_thresholds[2364]), .FEAT_ABOVE(feature_aboves[2364]), .FEAT_BELOW(feature_belows[2364])) ac2364(.scan_win(scan_win2364), .scan_win_std_dev(scan_win_std_dev[2364]), .feature_accum(feature_accums[2364]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2365]), .RECT1_Y(rectangle1_ys[2365]), .RECT1_WIDTH(rectangle1_widths[2365]), .RECT1_HEIGHT(rectangle1_heights[2365]), .RECT1_WEIGHT(rectangle1_weights[2365]), .RECT2_X(rectangle2_xs[2365]), .RECT2_Y(rectangle2_ys[2365]), .RECT2_WIDTH(rectangle2_widths[2365]), .RECT2_HEIGHT(rectangle2_heights[2365]), .RECT2_WEIGHT(rectangle2_weights[2365]), .RECT3_X(rectangle3_xs[2365]), .RECT3_Y(rectangle3_ys[2365]), .RECT3_WIDTH(rectangle3_widths[2365]), .RECT3_HEIGHT(rectangle3_heights[2365]), .RECT3_WEIGHT(rectangle3_weights[2365]), .FEAT_THRES(feature_thresholds[2365]), .FEAT_ABOVE(feature_aboves[2365]), .FEAT_BELOW(feature_belows[2365])) ac2365(.scan_win(scan_win2365), .scan_win_std_dev(scan_win_std_dev[2365]), .feature_accum(feature_accums[2365]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2366]), .RECT1_Y(rectangle1_ys[2366]), .RECT1_WIDTH(rectangle1_widths[2366]), .RECT1_HEIGHT(rectangle1_heights[2366]), .RECT1_WEIGHT(rectangle1_weights[2366]), .RECT2_X(rectangle2_xs[2366]), .RECT2_Y(rectangle2_ys[2366]), .RECT2_WIDTH(rectangle2_widths[2366]), .RECT2_HEIGHT(rectangle2_heights[2366]), .RECT2_WEIGHT(rectangle2_weights[2366]), .RECT3_X(rectangle3_xs[2366]), .RECT3_Y(rectangle3_ys[2366]), .RECT3_WIDTH(rectangle3_widths[2366]), .RECT3_HEIGHT(rectangle3_heights[2366]), .RECT3_WEIGHT(rectangle3_weights[2366]), .FEAT_THRES(feature_thresholds[2366]), .FEAT_ABOVE(feature_aboves[2366]), .FEAT_BELOW(feature_belows[2366])) ac2366(.scan_win(scan_win2366), .scan_win_std_dev(scan_win_std_dev[2366]), .feature_accum(feature_accums[2366]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2367]), .RECT1_Y(rectangle1_ys[2367]), .RECT1_WIDTH(rectangle1_widths[2367]), .RECT1_HEIGHT(rectangle1_heights[2367]), .RECT1_WEIGHT(rectangle1_weights[2367]), .RECT2_X(rectangle2_xs[2367]), .RECT2_Y(rectangle2_ys[2367]), .RECT2_WIDTH(rectangle2_widths[2367]), .RECT2_HEIGHT(rectangle2_heights[2367]), .RECT2_WEIGHT(rectangle2_weights[2367]), .RECT3_X(rectangle3_xs[2367]), .RECT3_Y(rectangle3_ys[2367]), .RECT3_WIDTH(rectangle3_widths[2367]), .RECT3_HEIGHT(rectangle3_heights[2367]), .RECT3_WEIGHT(rectangle3_weights[2367]), .FEAT_THRES(feature_thresholds[2367]), .FEAT_ABOVE(feature_aboves[2367]), .FEAT_BELOW(feature_belows[2367])) ac2367(.scan_win(scan_win2367), .scan_win_std_dev(scan_win_std_dev[2367]), .feature_accum(feature_accums[2367]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2368]), .RECT1_Y(rectangle1_ys[2368]), .RECT1_WIDTH(rectangle1_widths[2368]), .RECT1_HEIGHT(rectangle1_heights[2368]), .RECT1_WEIGHT(rectangle1_weights[2368]), .RECT2_X(rectangle2_xs[2368]), .RECT2_Y(rectangle2_ys[2368]), .RECT2_WIDTH(rectangle2_widths[2368]), .RECT2_HEIGHT(rectangle2_heights[2368]), .RECT2_WEIGHT(rectangle2_weights[2368]), .RECT3_X(rectangle3_xs[2368]), .RECT3_Y(rectangle3_ys[2368]), .RECT3_WIDTH(rectangle3_widths[2368]), .RECT3_HEIGHT(rectangle3_heights[2368]), .RECT3_WEIGHT(rectangle3_weights[2368]), .FEAT_THRES(feature_thresholds[2368]), .FEAT_ABOVE(feature_aboves[2368]), .FEAT_BELOW(feature_belows[2368])) ac2368(.scan_win(scan_win2368), .scan_win_std_dev(scan_win_std_dev[2368]), .feature_accum(feature_accums[2368]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2369]), .RECT1_Y(rectangle1_ys[2369]), .RECT1_WIDTH(rectangle1_widths[2369]), .RECT1_HEIGHT(rectangle1_heights[2369]), .RECT1_WEIGHT(rectangle1_weights[2369]), .RECT2_X(rectangle2_xs[2369]), .RECT2_Y(rectangle2_ys[2369]), .RECT2_WIDTH(rectangle2_widths[2369]), .RECT2_HEIGHT(rectangle2_heights[2369]), .RECT2_WEIGHT(rectangle2_weights[2369]), .RECT3_X(rectangle3_xs[2369]), .RECT3_Y(rectangle3_ys[2369]), .RECT3_WIDTH(rectangle3_widths[2369]), .RECT3_HEIGHT(rectangle3_heights[2369]), .RECT3_WEIGHT(rectangle3_weights[2369]), .FEAT_THRES(feature_thresholds[2369]), .FEAT_ABOVE(feature_aboves[2369]), .FEAT_BELOW(feature_belows[2369])) ac2369(.scan_win(scan_win2369), .scan_win_std_dev(scan_win_std_dev[2369]), .feature_accum(feature_accums[2369]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2370]), .RECT1_Y(rectangle1_ys[2370]), .RECT1_WIDTH(rectangle1_widths[2370]), .RECT1_HEIGHT(rectangle1_heights[2370]), .RECT1_WEIGHT(rectangle1_weights[2370]), .RECT2_X(rectangle2_xs[2370]), .RECT2_Y(rectangle2_ys[2370]), .RECT2_WIDTH(rectangle2_widths[2370]), .RECT2_HEIGHT(rectangle2_heights[2370]), .RECT2_WEIGHT(rectangle2_weights[2370]), .RECT3_X(rectangle3_xs[2370]), .RECT3_Y(rectangle3_ys[2370]), .RECT3_WIDTH(rectangle3_widths[2370]), .RECT3_HEIGHT(rectangle3_heights[2370]), .RECT3_WEIGHT(rectangle3_weights[2370]), .FEAT_THRES(feature_thresholds[2370]), .FEAT_ABOVE(feature_aboves[2370]), .FEAT_BELOW(feature_belows[2370])) ac2370(.scan_win(scan_win2370), .scan_win_std_dev(scan_win_std_dev[2370]), .feature_accum(feature_accums[2370]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2371]), .RECT1_Y(rectangle1_ys[2371]), .RECT1_WIDTH(rectangle1_widths[2371]), .RECT1_HEIGHT(rectangle1_heights[2371]), .RECT1_WEIGHT(rectangle1_weights[2371]), .RECT2_X(rectangle2_xs[2371]), .RECT2_Y(rectangle2_ys[2371]), .RECT2_WIDTH(rectangle2_widths[2371]), .RECT2_HEIGHT(rectangle2_heights[2371]), .RECT2_WEIGHT(rectangle2_weights[2371]), .RECT3_X(rectangle3_xs[2371]), .RECT3_Y(rectangle3_ys[2371]), .RECT3_WIDTH(rectangle3_widths[2371]), .RECT3_HEIGHT(rectangle3_heights[2371]), .RECT3_WEIGHT(rectangle3_weights[2371]), .FEAT_THRES(feature_thresholds[2371]), .FEAT_ABOVE(feature_aboves[2371]), .FEAT_BELOW(feature_belows[2371])) ac2371(.scan_win(scan_win2371), .scan_win_std_dev(scan_win_std_dev[2371]), .feature_accum(feature_accums[2371]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2372]), .RECT1_Y(rectangle1_ys[2372]), .RECT1_WIDTH(rectangle1_widths[2372]), .RECT1_HEIGHT(rectangle1_heights[2372]), .RECT1_WEIGHT(rectangle1_weights[2372]), .RECT2_X(rectangle2_xs[2372]), .RECT2_Y(rectangle2_ys[2372]), .RECT2_WIDTH(rectangle2_widths[2372]), .RECT2_HEIGHT(rectangle2_heights[2372]), .RECT2_WEIGHT(rectangle2_weights[2372]), .RECT3_X(rectangle3_xs[2372]), .RECT3_Y(rectangle3_ys[2372]), .RECT3_WIDTH(rectangle3_widths[2372]), .RECT3_HEIGHT(rectangle3_heights[2372]), .RECT3_WEIGHT(rectangle3_weights[2372]), .FEAT_THRES(feature_thresholds[2372]), .FEAT_ABOVE(feature_aboves[2372]), .FEAT_BELOW(feature_belows[2372])) ac2372(.scan_win(scan_win2372), .scan_win_std_dev(scan_win_std_dev[2372]), .feature_accum(feature_accums[2372]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2373]), .RECT1_Y(rectangle1_ys[2373]), .RECT1_WIDTH(rectangle1_widths[2373]), .RECT1_HEIGHT(rectangle1_heights[2373]), .RECT1_WEIGHT(rectangle1_weights[2373]), .RECT2_X(rectangle2_xs[2373]), .RECT2_Y(rectangle2_ys[2373]), .RECT2_WIDTH(rectangle2_widths[2373]), .RECT2_HEIGHT(rectangle2_heights[2373]), .RECT2_WEIGHT(rectangle2_weights[2373]), .RECT3_X(rectangle3_xs[2373]), .RECT3_Y(rectangle3_ys[2373]), .RECT3_WIDTH(rectangle3_widths[2373]), .RECT3_HEIGHT(rectangle3_heights[2373]), .RECT3_WEIGHT(rectangle3_weights[2373]), .FEAT_THRES(feature_thresholds[2373]), .FEAT_ABOVE(feature_aboves[2373]), .FEAT_BELOW(feature_belows[2373])) ac2373(.scan_win(scan_win2373), .scan_win_std_dev(scan_win_std_dev[2373]), .feature_accum(feature_accums[2373]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2374]), .RECT1_Y(rectangle1_ys[2374]), .RECT1_WIDTH(rectangle1_widths[2374]), .RECT1_HEIGHT(rectangle1_heights[2374]), .RECT1_WEIGHT(rectangle1_weights[2374]), .RECT2_X(rectangle2_xs[2374]), .RECT2_Y(rectangle2_ys[2374]), .RECT2_WIDTH(rectangle2_widths[2374]), .RECT2_HEIGHT(rectangle2_heights[2374]), .RECT2_WEIGHT(rectangle2_weights[2374]), .RECT3_X(rectangle3_xs[2374]), .RECT3_Y(rectangle3_ys[2374]), .RECT3_WIDTH(rectangle3_widths[2374]), .RECT3_HEIGHT(rectangle3_heights[2374]), .RECT3_WEIGHT(rectangle3_weights[2374]), .FEAT_THRES(feature_thresholds[2374]), .FEAT_ABOVE(feature_aboves[2374]), .FEAT_BELOW(feature_belows[2374])) ac2374(.scan_win(scan_win2374), .scan_win_std_dev(scan_win_std_dev[2374]), .feature_accum(feature_accums[2374]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2375]), .RECT1_Y(rectangle1_ys[2375]), .RECT1_WIDTH(rectangle1_widths[2375]), .RECT1_HEIGHT(rectangle1_heights[2375]), .RECT1_WEIGHT(rectangle1_weights[2375]), .RECT2_X(rectangle2_xs[2375]), .RECT2_Y(rectangle2_ys[2375]), .RECT2_WIDTH(rectangle2_widths[2375]), .RECT2_HEIGHT(rectangle2_heights[2375]), .RECT2_WEIGHT(rectangle2_weights[2375]), .RECT3_X(rectangle3_xs[2375]), .RECT3_Y(rectangle3_ys[2375]), .RECT3_WIDTH(rectangle3_widths[2375]), .RECT3_HEIGHT(rectangle3_heights[2375]), .RECT3_WEIGHT(rectangle3_weights[2375]), .FEAT_THRES(feature_thresholds[2375]), .FEAT_ABOVE(feature_aboves[2375]), .FEAT_BELOW(feature_belows[2375])) ac2375(.scan_win(scan_win2375), .scan_win_std_dev(scan_win_std_dev[2375]), .feature_accum(feature_accums[2375]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2376]), .RECT1_Y(rectangle1_ys[2376]), .RECT1_WIDTH(rectangle1_widths[2376]), .RECT1_HEIGHT(rectangle1_heights[2376]), .RECT1_WEIGHT(rectangle1_weights[2376]), .RECT2_X(rectangle2_xs[2376]), .RECT2_Y(rectangle2_ys[2376]), .RECT2_WIDTH(rectangle2_widths[2376]), .RECT2_HEIGHT(rectangle2_heights[2376]), .RECT2_WEIGHT(rectangle2_weights[2376]), .RECT3_X(rectangle3_xs[2376]), .RECT3_Y(rectangle3_ys[2376]), .RECT3_WIDTH(rectangle3_widths[2376]), .RECT3_HEIGHT(rectangle3_heights[2376]), .RECT3_WEIGHT(rectangle3_weights[2376]), .FEAT_THRES(feature_thresholds[2376]), .FEAT_ABOVE(feature_aboves[2376]), .FEAT_BELOW(feature_belows[2376])) ac2376(.scan_win(scan_win2376), .scan_win_std_dev(scan_win_std_dev[2376]), .feature_accum(feature_accums[2376]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2377]), .RECT1_Y(rectangle1_ys[2377]), .RECT1_WIDTH(rectangle1_widths[2377]), .RECT1_HEIGHT(rectangle1_heights[2377]), .RECT1_WEIGHT(rectangle1_weights[2377]), .RECT2_X(rectangle2_xs[2377]), .RECT2_Y(rectangle2_ys[2377]), .RECT2_WIDTH(rectangle2_widths[2377]), .RECT2_HEIGHT(rectangle2_heights[2377]), .RECT2_WEIGHT(rectangle2_weights[2377]), .RECT3_X(rectangle3_xs[2377]), .RECT3_Y(rectangle3_ys[2377]), .RECT3_WIDTH(rectangle3_widths[2377]), .RECT3_HEIGHT(rectangle3_heights[2377]), .RECT3_WEIGHT(rectangle3_weights[2377]), .FEAT_THRES(feature_thresholds[2377]), .FEAT_ABOVE(feature_aboves[2377]), .FEAT_BELOW(feature_belows[2377])) ac2377(.scan_win(scan_win2377), .scan_win_std_dev(scan_win_std_dev[2377]), .feature_accum(feature_accums[2377]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2378]), .RECT1_Y(rectangle1_ys[2378]), .RECT1_WIDTH(rectangle1_widths[2378]), .RECT1_HEIGHT(rectangle1_heights[2378]), .RECT1_WEIGHT(rectangle1_weights[2378]), .RECT2_X(rectangle2_xs[2378]), .RECT2_Y(rectangle2_ys[2378]), .RECT2_WIDTH(rectangle2_widths[2378]), .RECT2_HEIGHT(rectangle2_heights[2378]), .RECT2_WEIGHT(rectangle2_weights[2378]), .RECT3_X(rectangle3_xs[2378]), .RECT3_Y(rectangle3_ys[2378]), .RECT3_WIDTH(rectangle3_widths[2378]), .RECT3_HEIGHT(rectangle3_heights[2378]), .RECT3_WEIGHT(rectangle3_weights[2378]), .FEAT_THRES(feature_thresholds[2378]), .FEAT_ABOVE(feature_aboves[2378]), .FEAT_BELOW(feature_belows[2378])) ac2378(.scan_win(scan_win2378), .scan_win_std_dev(scan_win_std_dev[2378]), .feature_accum(feature_accums[2378]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2379]), .RECT1_Y(rectangle1_ys[2379]), .RECT1_WIDTH(rectangle1_widths[2379]), .RECT1_HEIGHT(rectangle1_heights[2379]), .RECT1_WEIGHT(rectangle1_weights[2379]), .RECT2_X(rectangle2_xs[2379]), .RECT2_Y(rectangle2_ys[2379]), .RECT2_WIDTH(rectangle2_widths[2379]), .RECT2_HEIGHT(rectangle2_heights[2379]), .RECT2_WEIGHT(rectangle2_weights[2379]), .RECT3_X(rectangle3_xs[2379]), .RECT3_Y(rectangle3_ys[2379]), .RECT3_WIDTH(rectangle3_widths[2379]), .RECT3_HEIGHT(rectangle3_heights[2379]), .RECT3_WEIGHT(rectangle3_weights[2379]), .FEAT_THRES(feature_thresholds[2379]), .FEAT_ABOVE(feature_aboves[2379]), .FEAT_BELOW(feature_belows[2379])) ac2379(.scan_win(scan_win2379), .scan_win_std_dev(scan_win_std_dev[2379]), .feature_accum(feature_accums[2379]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2380]), .RECT1_Y(rectangle1_ys[2380]), .RECT1_WIDTH(rectangle1_widths[2380]), .RECT1_HEIGHT(rectangle1_heights[2380]), .RECT1_WEIGHT(rectangle1_weights[2380]), .RECT2_X(rectangle2_xs[2380]), .RECT2_Y(rectangle2_ys[2380]), .RECT2_WIDTH(rectangle2_widths[2380]), .RECT2_HEIGHT(rectangle2_heights[2380]), .RECT2_WEIGHT(rectangle2_weights[2380]), .RECT3_X(rectangle3_xs[2380]), .RECT3_Y(rectangle3_ys[2380]), .RECT3_WIDTH(rectangle3_widths[2380]), .RECT3_HEIGHT(rectangle3_heights[2380]), .RECT3_WEIGHT(rectangle3_weights[2380]), .FEAT_THRES(feature_thresholds[2380]), .FEAT_ABOVE(feature_aboves[2380]), .FEAT_BELOW(feature_belows[2380])) ac2380(.scan_win(scan_win2380), .scan_win_std_dev(scan_win_std_dev[2380]), .feature_accum(feature_accums[2380]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2381]), .RECT1_Y(rectangle1_ys[2381]), .RECT1_WIDTH(rectangle1_widths[2381]), .RECT1_HEIGHT(rectangle1_heights[2381]), .RECT1_WEIGHT(rectangle1_weights[2381]), .RECT2_X(rectangle2_xs[2381]), .RECT2_Y(rectangle2_ys[2381]), .RECT2_WIDTH(rectangle2_widths[2381]), .RECT2_HEIGHT(rectangle2_heights[2381]), .RECT2_WEIGHT(rectangle2_weights[2381]), .RECT3_X(rectangle3_xs[2381]), .RECT3_Y(rectangle3_ys[2381]), .RECT3_WIDTH(rectangle3_widths[2381]), .RECT3_HEIGHT(rectangle3_heights[2381]), .RECT3_WEIGHT(rectangle3_weights[2381]), .FEAT_THRES(feature_thresholds[2381]), .FEAT_ABOVE(feature_aboves[2381]), .FEAT_BELOW(feature_belows[2381])) ac2381(.scan_win(scan_win2381), .scan_win_std_dev(scan_win_std_dev[2381]), .feature_accum(feature_accums[2381]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2382]), .RECT1_Y(rectangle1_ys[2382]), .RECT1_WIDTH(rectangle1_widths[2382]), .RECT1_HEIGHT(rectangle1_heights[2382]), .RECT1_WEIGHT(rectangle1_weights[2382]), .RECT2_X(rectangle2_xs[2382]), .RECT2_Y(rectangle2_ys[2382]), .RECT2_WIDTH(rectangle2_widths[2382]), .RECT2_HEIGHT(rectangle2_heights[2382]), .RECT2_WEIGHT(rectangle2_weights[2382]), .RECT3_X(rectangle3_xs[2382]), .RECT3_Y(rectangle3_ys[2382]), .RECT3_WIDTH(rectangle3_widths[2382]), .RECT3_HEIGHT(rectangle3_heights[2382]), .RECT3_WEIGHT(rectangle3_weights[2382]), .FEAT_THRES(feature_thresholds[2382]), .FEAT_ABOVE(feature_aboves[2382]), .FEAT_BELOW(feature_belows[2382])) ac2382(.scan_win(scan_win2382), .scan_win_std_dev(scan_win_std_dev[2382]), .feature_accum(feature_accums[2382]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2383]), .RECT1_Y(rectangle1_ys[2383]), .RECT1_WIDTH(rectangle1_widths[2383]), .RECT1_HEIGHT(rectangle1_heights[2383]), .RECT1_WEIGHT(rectangle1_weights[2383]), .RECT2_X(rectangle2_xs[2383]), .RECT2_Y(rectangle2_ys[2383]), .RECT2_WIDTH(rectangle2_widths[2383]), .RECT2_HEIGHT(rectangle2_heights[2383]), .RECT2_WEIGHT(rectangle2_weights[2383]), .RECT3_X(rectangle3_xs[2383]), .RECT3_Y(rectangle3_ys[2383]), .RECT3_WIDTH(rectangle3_widths[2383]), .RECT3_HEIGHT(rectangle3_heights[2383]), .RECT3_WEIGHT(rectangle3_weights[2383]), .FEAT_THRES(feature_thresholds[2383]), .FEAT_ABOVE(feature_aboves[2383]), .FEAT_BELOW(feature_belows[2383])) ac2383(.scan_win(scan_win2383), .scan_win_std_dev(scan_win_std_dev[2383]), .feature_accum(feature_accums[2383]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2384]), .RECT1_Y(rectangle1_ys[2384]), .RECT1_WIDTH(rectangle1_widths[2384]), .RECT1_HEIGHT(rectangle1_heights[2384]), .RECT1_WEIGHT(rectangle1_weights[2384]), .RECT2_X(rectangle2_xs[2384]), .RECT2_Y(rectangle2_ys[2384]), .RECT2_WIDTH(rectangle2_widths[2384]), .RECT2_HEIGHT(rectangle2_heights[2384]), .RECT2_WEIGHT(rectangle2_weights[2384]), .RECT3_X(rectangle3_xs[2384]), .RECT3_Y(rectangle3_ys[2384]), .RECT3_WIDTH(rectangle3_widths[2384]), .RECT3_HEIGHT(rectangle3_heights[2384]), .RECT3_WEIGHT(rectangle3_weights[2384]), .FEAT_THRES(feature_thresholds[2384]), .FEAT_ABOVE(feature_aboves[2384]), .FEAT_BELOW(feature_belows[2384])) ac2384(.scan_win(scan_win2384), .scan_win_std_dev(scan_win_std_dev[2384]), .feature_accum(feature_accums[2384]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2385]), .RECT1_Y(rectangle1_ys[2385]), .RECT1_WIDTH(rectangle1_widths[2385]), .RECT1_HEIGHT(rectangle1_heights[2385]), .RECT1_WEIGHT(rectangle1_weights[2385]), .RECT2_X(rectangle2_xs[2385]), .RECT2_Y(rectangle2_ys[2385]), .RECT2_WIDTH(rectangle2_widths[2385]), .RECT2_HEIGHT(rectangle2_heights[2385]), .RECT2_WEIGHT(rectangle2_weights[2385]), .RECT3_X(rectangle3_xs[2385]), .RECT3_Y(rectangle3_ys[2385]), .RECT3_WIDTH(rectangle3_widths[2385]), .RECT3_HEIGHT(rectangle3_heights[2385]), .RECT3_WEIGHT(rectangle3_weights[2385]), .FEAT_THRES(feature_thresholds[2385]), .FEAT_ABOVE(feature_aboves[2385]), .FEAT_BELOW(feature_belows[2385])) ac2385(.scan_win(scan_win2385), .scan_win_std_dev(scan_win_std_dev[2385]), .feature_accum(feature_accums[2385]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2386]), .RECT1_Y(rectangle1_ys[2386]), .RECT1_WIDTH(rectangle1_widths[2386]), .RECT1_HEIGHT(rectangle1_heights[2386]), .RECT1_WEIGHT(rectangle1_weights[2386]), .RECT2_X(rectangle2_xs[2386]), .RECT2_Y(rectangle2_ys[2386]), .RECT2_WIDTH(rectangle2_widths[2386]), .RECT2_HEIGHT(rectangle2_heights[2386]), .RECT2_WEIGHT(rectangle2_weights[2386]), .RECT3_X(rectangle3_xs[2386]), .RECT3_Y(rectangle3_ys[2386]), .RECT3_WIDTH(rectangle3_widths[2386]), .RECT3_HEIGHT(rectangle3_heights[2386]), .RECT3_WEIGHT(rectangle3_weights[2386]), .FEAT_THRES(feature_thresholds[2386]), .FEAT_ABOVE(feature_aboves[2386]), .FEAT_BELOW(feature_belows[2386])) ac2386(.scan_win(scan_win2386), .scan_win_std_dev(scan_win_std_dev[2386]), .feature_accum(feature_accums[2386]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2387]), .RECT1_Y(rectangle1_ys[2387]), .RECT1_WIDTH(rectangle1_widths[2387]), .RECT1_HEIGHT(rectangle1_heights[2387]), .RECT1_WEIGHT(rectangle1_weights[2387]), .RECT2_X(rectangle2_xs[2387]), .RECT2_Y(rectangle2_ys[2387]), .RECT2_WIDTH(rectangle2_widths[2387]), .RECT2_HEIGHT(rectangle2_heights[2387]), .RECT2_WEIGHT(rectangle2_weights[2387]), .RECT3_X(rectangle3_xs[2387]), .RECT3_Y(rectangle3_ys[2387]), .RECT3_WIDTH(rectangle3_widths[2387]), .RECT3_HEIGHT(rectangle3_heights[2387]), .RECT3_WEIGHT(rectangle3_weights[2387]), .FEAT_THRES(feature_thresholds[2387]), .FEAT_ABOVE(feature_aboves[2387]), .FEAT_BELOW(feature_belows[2387])) ac2387(.scan_win(scan_win2387), .scan_win_std_dev(scan_win_std_dev[2387]), .feature_accum(feature_accums[2387]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2388]), .RECT1_Y(rectangle1_ys[2388]), .RECT1_WIDTH(rectangle1_widths[2388]), .RECT1_HEIGHT(rectangle1_heights[2388]), .RECT1_WEIGHT(rectangle1_weights[2388]), .RECT2_X(rectangle2_xs[2388]), .RECT2_Y(rectangle2_ys[2388]), .RECT2_WIDTH(rectangle2_widths[2388]), .RECT2_HEIGHT(rectangle2_heights[2388]), .RECT2_WEIGHT(rectangle2_weights[2388]), .RECT3_X(rectangle3_xs[2388]), .RECT3_Y(rectangle3_ys[2388]), .RECT3_WIDTH(rectangle3_widths[2388]), .RECT3_HEIGHT(rectangle3_heights[2388]), .RECT3_WEIGHT(rectangle3_weights[2388]), .FEAT_THRES(feature_thresholds[2388]), .FEAT_ABOVE(feature_aboves[2388]), .FEAT_BELOW(feature_belows[2388])) ac2388(.scan_win(scan_win2388), .scan_win_std_dev(scan_win_std_dev[2388]), .feature_accum(feature_accums[2388]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2389]), .RECT1_Y(rectangle1_ys[2389]), .RECT1_WIDTH(rectangle1_widths[2389]), .RECT1_HEIGHT(rectangle1_heights[2389]), .RECT1_WEIGHT(rectangle1_weights[2389]), .RECT2_X(rectangle2_xs[2389]), .RECT2_Y(rectangle2_ys[2389]), .RECT2_WIDTH(rectangle2_widths[2389]), .RECT2_HEIGHT(rectangle2_heights[2389]), .RECT2_WEIGHT(rectangle2_weights[2389]), .RECT3_X(rectangle3_xs[2389]), .RECT3_Y(rectangle3_ys[2389]), .RECT3_WIDTH(rectangle3_widths[2389]), .RECT3_HEIGHT(rectangle3_heights[2389]), .RECT3_WEIGHT(rectangle3_weights[2389]), .FEAT_THRES(feature_thresholds[2389]), .FEAT_ABOVE(feature_aboves[2389]), .FEAT_BELOW(feature_belows[2389])) ac2389(.scan_win(scan_win2389), .scan_win_std_dev(scan_win_std_dev[2389]), .feature_accum(feature_accums[2389]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2390]), .RECT1_Y(rectangle1_ys[2390]), .RECT1_WIDTH(rectangle1_widths[2390]), .RECT1_HEIGHT(rectangle1_heights[2390]), .RECT1_WEIGHT(rectangle1_weights[2390]), .RECT2_X(rectangle2_xs[2390]), .RECT2_Y(rectangle2_ys[2390]), .RECT2_WIDTH(rectangle2_widths[2390]), .RECT2_HEIGHT(rectangle2_heights[2390]), .RECT2_WEIGHT(rectangle2_weights[2390]), .RECT3_X(rectangle3_xs[2390]), .RECT3_Y(rectangle3_ys[2390]), .RECT3_WIDTH(rectangle3_widths[2390]), .RECT3_HEIGHT(rectangle3_heights[2390]), .RECT3_WEIGHT(rectangle3_weights[2390]), .FEAT_THRES(feature_thresholds[2390]), .FEAT_ABOVE(feature_aboves[2390]), .FEAT_BELOW(feature_belows[2390])) ac2390(.scan_win(scan_win2390), .scan_win_std_dev(scan_win_std_dev[2390]), .feature_accum(feature_accums[2390]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2391]), .RECT1_Y(rectangle1_ys[2391]), .RECT1_WIDTH(rectangle1_widths[2391]), .RECT1_HEIGHT(rectangle1_heights[2391]), .RECT1_WEIGHT(rectangle1_weights[2391]), .RECT2_X(rectangle2_xs[2391]), .RECT2_Y(rectangle2_ys[2391]), .RECT2_WIDTH(rectangle2_widths[2391]), .RECT2_HEIGHT(rectangle2_heights[2391]), .RECT2_WEIGHT(rectangle2_weights[2391]), .RECT3_X(rectangle3_xs[2391]), .RECT3_Y(rectangle3_ys[2391]), .RECT3_WIDTH(rectangle3_widths[2391]), .RECT3_HEIGHT(rectangle3_heights[2391]), .RECT3_WEIGHT(rectangle3_weights[2391]), .FEAT_THRES(feature_thresholds[2391]), .FEAT_ABOVE(feature_aboves[2391]), .FEAT_BELOW(feature_belows[2391])) ac2391(.scan_win(scan_win2391), .scan_win_std_dev(scan_win_std_dev[2391]), .feature_accum(feature_accums[2391]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2392]), .RECT1_Y(rectangle1_ys[2392]), .RECT1_WIDTH(rectangle1_widths[2392]), .RECT1_HEIGHT(rectangle1_heights[2392]), .RECT1_WEIGHT(rectangle1_weights[2392]), .RECT2_X(rectangle2_xs[2392]), .RECT2_Y(rectangle2_ys[2392]), .RECT2_WIDTH(rectangle2_widths[2392]), .RECT2_HEIGHT(rectangle2_heights[2392]), .RECT2_WEIGHT(rectangle2_weights[2392]), .RECT3_X(rectangle3_xs[2392]), .RECT3_Y(rectangle3_ys[2392]), .RECT3_WIDTH(rectangle3_widths[2392]), .RECT3_HEIGHT(rectangle3_heights[2392]), .RECT3_WEIGHT(rectangle3_weights[2392]), .FEAT_THRES(feature_thresholds[2392]), .FEAT_ABOVE(feature_aboves[2392]), .FEAT_BELOW(feature_belows[2392])) ac2392(.scan_win(scan_win2392), .scan_win_std_dev(scan_win_std_dev[2392]), .feature_accum(feature_accums[2392]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2393]), .RECT1_Y(rectangle1_ys[2393]), .RECT1_WIDTH(rectangle1_widths[2393]), .RECT1_HEIGHT(rectangle1_heights[2393]), .RECT1_WEIGHT(rectangle1_weights[2393]), .RECT2_X(rectangle2_xs[2393]), .RECT2_Y(rectangle2_ys[2393]), .RECT2_WIDTH(rectangle2_widths[2393]), .RECT2_HEIGHT(rectangle2_heights[2393]), .RECT2_WEIGHT(rectangle2_weights[2393]), .RECT3_X(rectangle3_xs[2393]), .RECT3_Y(rectangle3_ys[2393]), .RECT3_WIDTH(rectangle3_widths[2393]), .RECT3_HEIGHT(rectangle3_heights[2393]), .RECT3_WEIGHT(rectangle3_weights[2393]), .FEAT_THRES(feature_thresholds[2393]), .FEAT_ABOVE(feature_aboves[2393]), .FEAT_BELOW(feature_belows[2393])) ac2393(.scan_win(scan_win2393), .scan_win_std_dev(scan_win_std_dev[2393]), .feature_accum(feature_accums[2393]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2394]), .RECT1_Y(rectangle1_ys[2394]), .RECT1_WIDTH(rectangle1_widths[2394]), .RECT1_HEIGHT(rectangle1_heights[2394]), .RECT1_WEIGHT(rectangle1_weights[2394]), .RECT2_X(rectangle2_xs[2394]), .RECT2_Y(rectangle2_ys[2394]), .RECT2_WIDTH(rectangle2_widths[2394]), .RECT2_HEIGHT(rectangle2_heights[2394]), .RECT2_WEIGHT(rectangle2_weights[2394]), .RECT3_X(rectangle3_xs[2394]), .RECT3_Y(rectangle3_ys[2394]), .RECT3_WIDTH(rectangle3_widths[2394]), .RECT3_HEIGHT(rectangle3_heights[2394]), .RECT3_WEIGHT(rectangle3_weights[2394]), .FEAT_THRES(feature_thresholds[2394]), .FEAT_ABOVE(feature_aboves[2394]), .FEAT_BELOW(feature_belows[2394])) ac2394(.scan_win(scan_win2394), .scan_win_std_dev(scan_win_std_dev[2394]), .feature_accum(feature_accums[2394]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2395]), .RECT1_Y(rectangle1_ys[2395]), .RECT1_WIDTH(rectangle1_widths[2395]), .RECT1_HEIGHT(rectangle1_heights[2395]), .RECT1_WEIGHT(rectangle1_weights[2395]), .RECT2_X(rectangle2_xs[2395]), .RECT2_Y(rectangle2_ys[2395]), .RECT2_WIDTH(rectangle2_widths[2395]), .RECT2_HEIGHT(rectangle2_heights[2395]), .RECT2_WEIGHT(rectangle2_weights[2395]), .RECT3_X(rectangle3_xs[2395]), .RECT3_Y(rectangle3_ys[2395]), .RECT3_WIDTH(rectangle3_widths[2395]), .RECT3_HEIGHT(rectangle3_heights[2395]), .RECT3_WEIGHT(rectangle3_weights[2395]), .FEAT_THRES(feature_thresholds[2395]), .FEAT_ABOVE(feature_aboves[2395]), .FEAT_BELOW(feature_belows[2395])) ac2395(.scan_win(scan_win2395), .scan_win_std_dev(scan_win_std_dev[2395]), .feature_accum(feature_accums[2395]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2396]), .RECT1_Y(rectangle1_ys[2396]), .RECT1_WIDTH(rectangle1_widths[2396]), .RECT1_HEIGHT(rectangle1_heights[2396]), .RECT1_WEIGHT(rectangle1_weights[2396]), .RECT2_X(rectangle2_xs[2396]), .RECT2_Y(rectangle2_ys[2396]), .RECT2_WIDTH(rectangle2_widths[2396]), .RECT2_HEIGHT(rectangle2_heights[2396]), .RECT2_WEIGHT(rectangle2_weights[2396]), .RECT3_X(rectangle3_xs[2396]), .RECT3_Y(rectangle3_ys[2396]), .RECT3_WIDTH(rectangle3_widths[2396]), .RECT3_HEIGHT(rectangle3_heights[2396]), .RECT3_WEIGHT(rectangle3_weights[2396]), .FEAT_THRES(feature_thresholds[2396]), .FEAT_ABOVE(feature_aboves[2396]), .FEAT_BELOW(feature_belows[2396])) ac2396(.scan_win(scan_win2396), .scan_win_std_dev(scan_win_std_dev[2396]), .feature_accum(feature_accums[2396]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2397]), .RECT1_Y(rectangle1_ys[2397]), .RECT1_WIDTH(rectangle1_widths[2397]), .RECT1_HEIGHT(rectangle1_heights[2397]), .RECT1_WEIGHT(rectangle1_weights[2397]), .RECT2_X(rectangle2_xs[2397]), .RECT2_Y(rectangle2_ys[2397]), .RECT2_WIDTH(rectangle2_widths[2397]), .RECT2_HEIGHT(rectangle2_heights[2397]), .RECT2_WEIGHT(rectangle2_weights[2397]), .RECT3_X(rectangle3_xs[2397]), .RECT3_Y(rectangle3_ys[2397]), .RECT3_WIDTH(rectangle3_widths[2397]), .RECT3_HEIGHT(rectangle3_heights[2397]), .RECT3_WEIGHT(rectangle3_weights[2397]), .FEAT_THRES(feature_thresholds[2397]), .FEAT_ABOVE(feature_aboves[2397]), .FEAT_BELOW(feature_belows[2397])) ac2397(.scan_win(scan_win2397), .scan_win_std_dev(scan_win_std_dev[2397]), .feature_accum(feature_accums[2397]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2398]), .RECT1_Y(rectangle1_ys[2398]), .RECT1_WIDTH(rectangle1_widths[2398]), .RECT1_HEIGHT(rectangle1_heights[2398]), .RECT1_WEIGHT(rectangle1_weights[2398]), .RECT2_X(rectangle2_xs[2398]), .RECT2_Y(rectangle2_ys[2398]), .RECT2_WIDTH(rectangle2_widths[2398]), .RECT2_HEIGHT(rectangle2_heights[2398]), .RECT2_WEIGHT(rectangle2_weights[2398]), .RECT3_X(rectangle3_xs[2398]), .RECT3_Y(rectangle3_ys[2398]), .RECT3_WIDTH(rectangle3_widths[2398]), .RECT3_HEIGHT(rectangle3_heights[2398]), .RECT3_WEIGHT(rectangle3_weights[2398]), .FEAT_THRES(feature_thresholds[2398]), .FEAT_ABOVE(feature_aboves[2398]), .FEAT_BELOW(feature_belows[2398])) ac2398(.scan_win(scan_win2398), .scan_win_std_dev(scan_win_std_dev[2398]), .feature_accum(feature_accums[2398]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2399]), .RECT1_Y(rectangle1_ys[2399]), .RECT1_WIDTH(rectangle1_widths[2399]), .RECT1_HEIGHT(rectangle1_heights[2399]), .RECT1_WEIGHT(rectangle1_weights[2399]), .RECT2_X(rectangle2_xs[2399]), .RECT2_Y(rectangle2_ys[2399]), .RECT2_WIDTH(rectangle2_widths[2399]), .RECT2_HEIGHT(rectangle2_heights[2399]), .RECT2_WEIGHT(rectangle2_weights[2399]), .RECT3_X(rectangle3_xs[2399]), .RECT3_Y(rectangle3_ys[2399]), .RECT3_WIDTH(rectangle3_widths[2399]), .RECT3_HEIGHT(rectangle3_heights[2399]), .RECT3_WEIGHT(rectangle3_weights[2399]), .FEAT_THRES(feature_thresholds[2399]), .FEAT_ABOVE(feature_aboves[2399]), .FEAT_BELOW(feature_belows[2399])) ac2399(.scan_win(scan_win2399), .scan_win_std_dev(scan_win_std_dev[2399]), .feature_accum(feature_accums[2399]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2400]), .RECT1_Y(rectangle1_ys[2400]), .RECT1_WIDTH(rectangle1_widths[2400]), .RECT1_HEIGHT(rectangle1_heights[2400]), .RECT1_WEIGHT(rectangle1_weights[2400]), .RECT2_X(rectangle2_xs[2400]), .RECT2_Y(rectangle2_ys[2400]), .RECT2_WIDTH(rectangle2_widths[2400]), .RECT2_HEIGHT(rectangle2_heights[2400]), .RECT2_WEIGHT(rectangle2_weights[2400]), .RECT3_X(rectangle3_xs[2400]), .RECT3_Y(rectangle3_ys[2400]), .RECT3_WIDTH(rectangle3_widths[2400]), .RECT3_HEIGHT(rectangle3_heights[2400]), .RECT3_WEIGHT(rectangle3_weights[2400]), .FEAT_THRES(feature_thresholds[2400]), .FEAT_ABOVE(feature_aboves[2400]), .FEAT_BELOW(feature_belows[2400])) ac2400(.scan_win(scan_win2400), .scan_win_std_dev(scan_win_std_dev[2400]), .feature_accum(feature_accums[2400]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2401]), .RECT1_Y(rectangle1_ys[2401]), .RECT1_WIDTH(rectangle1_widths[2401]), .RECT1_HEIGHT(rectangle1_heights[2401]), .RECT1_WEIGHT(rectangle1_weights[2401]), .RECT2_X(rectangle2_xs[2401]), .RECT2_Y(rectangle2_ys[2401]), .RECT2_WIDTH(rectangle2_widths[2401]), .RECT2_HEIGHT(rectangle2_heights[2401]), .RECT2_WEIGHT(rectangle2_weights[2401]), .RECT3_X(rectangle3_xs[2401]), .RECT3_Y(rectangle3_ys[2401]), .RECT3_WIDTH(rectangle3_widths[2401]), .RECT3_HEIGHT(rectangle3_heights[2401]), .RECT3_WEIGHT(rectangle3_weights[2401]), .FEAT_THRES(feature_thresholds[2401]), .FEAT_ABOVE(feature_aboves[2401]), .FEAT_BELOW(feature_belows[2401])) ac2401(.scan_win(scan_win2401), .scan_win_std_dev(scan_win_std_dev[2401]), .feature_accum(feature_accums[2401]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2402]), .RECT1_Y(rectangle1_ys[2402]), .RECT1_WIDTH(rectangle1_widths[2402]), .RECT1_HEIGHT(rectangle1_heights[2402]), .RECT1_WEIGHT(rectangle1_weights[2402]), .RECT2_X(rectangle2_xs[2402]), .RECT2_Y(rectangle2_ys[2402]), .RECT2_WIDTH(rectangle2_widths[2402]), .RECT2_HEIGHT(rectangle2_heights[2402]), .RECT2_WEIGHT(rectangle2_weights[2402]), .RECT3_X(rectangle3_xs[2402]), .RECT3_Y(rectangle3_ys[2402]), .RECT3_WIDTH(rectangle3_widths[2402]), .RECT3_HEIGHT(rectangle3_heights[2402]), .RECT3_WEIGHT(rectangle3_weights[2402]), .FEAT_THRES(feature_thresholds[2402]), .FEAT_ABOVE(feature_aboves[2402]), .FEAT_BELOW(feature_belows[2402])) ac2402(.scan_win(scan_win2402), .scan_win_std_dev(scan_win_std_dev[2402]), .feature_accum(feature_accums[2402]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2403]), .RECT1_Y(rectangle1_ys[2403]), .RECT1_WIDTH(rectangle1_widths[2403]), .RECT1_HEIGHT(rectangle1_heights[2403]), .RECT1_WEIGHT(rectangle1_weights[2403]), .RECT2_X(rectangle2_xs[2403]), .RECT2_Y(rectangle2_ys[2403]), .RECT2_WIDTH(rectangle2_widths[2403]), .RECT2_HEIGHT(rectangle2_heights[2403]), .RECT2_WEIGHT(rectangle2_weights[2403]), .RECT3_X(rectangle3_xs[2403]), .RECT3_Y(rectangle3_ys[2403]), .RECT3_WIDTH(rectangle3_widths[2403]), .RECT3_HEIGHT(rectangle3_heights[2403]), .RECT3_WEIGHT(rectangle3_weights[2403]), .FEAT_THRES(feature_thresholds[2403]), .FEAT_ABOVE(feature_aboves[2403]), .FEAT_BELOW(feature_belows[2403])) ac2403(.scan_win(scan_win2403), .scan_win_std_dev(scan_win_std_dev[2403]), .feature_accum(feature_accums[2403]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2404]), .RECT1_Y(rectangle1_ys[2404]), .RECT1_WIDTH(rectangle1_widths[2404]), .RECT1_HEIGHT(rectangle1_heights[2404]), .RECT1_WEIGHT(rectangle1_weights[2404]), .RECT2_X(rectangle2_xs[2404]), .RECT2_Y(rectangle2_ys[2404]), .RECT2_WIDTH(rectangle2_widths[2404]), .RECT2_HEIGHT(rectangle2_heights[2404]), .RECT2_WEIGHT(rectangle2_weights[2404]), .RECT3_X(rectangle3_xs[2404]), .RECT3_Y(rectangle3_ys[2404]), .RECT3_WIDTH(rectangle3_widths[2404]), .RECT3_HEIGHT(rectangle3_heights[2404]), .RECT3_WEIGHT(rectangle3_weights[2404]), .FEAT_THRES(feature_thresholds[2404]), .FEAT_ABOVE(feature_aboves[2404]), .FEAT_BELOW(feature_belows[2404])) ac2404(.scan_win(scan_win2404), .scan_win_std_dev(scan_win_std_dev[2404]), .feature_accum(feature_accums[2404]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2405]), .RECT1_Y(rectangle1_ys[2405]), .RECT1_WIDTH(rectangle1_widths[2405]), .RECT1_HEIGHT(rectangle1_heights[2405]), .RECT1_WEIGHT(rectangle1_weights[2405]), .RECT2_X(rectangle2_xs[2405]), .RECT2_Y(rectangle2_ys[2405]), .RECT2_WIDTH(rectangle2_widths[2405]), .RECT2_HEIGHT(rectangle2_heights[2405]), .RECT2_WEIGHT(rectangle2_weights[2405]), .RECT3_X(rectangle3_xs[2405]), .RECT3_Y(rectangle3_ys[2405]), .RECT3_WIDTH(rectangle3_widths[2405]), .RECT3_HEIGHT(rectangle3_heights[2405]), .RECT3_WEIGHT(rectangle3_weights[2405]), .FEAT_THRES(feature_thresholds[2405]), .FEAT_ABOVE(feature_aboves[2405]), .FEAT_BELOW(feature_belows[2405])) ac2405(.scan_win(scan_win2405), .scan_win_std_dev(scan_win_std_dev[2405]), .feature_accum(feature_accums[2405]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2406]), .RECT1_Y(rectangle1_ys[2406]), .RECT1_WIDTH(rectangle1_widths[2406]), .RECT1_HEIGHT(rectangle1_heights[2406]), .RECT1_WEIGHT(rectangle1_weights[2406]), .RECT2_X(rectangle2_xs[2406]), .RECT2_Y(rectangle2_ys[2406]), .RECT2_WIDTH(rectangle2_widths[2406]), .RECT2_HEIGHT(rectangle2_heights[2406]), .RECT2_WEIGHT(rectangle2_weights[2406]), .RECT3_X(rectangle3_xs[2406]), .RECT3_Y(rectangle3_ys[2406]), .RECT3_WIDTH(rectangle3_widths[2406]), .RECT3_HEIGHT(rectangle3_heights[2406]), .RECT3_WEIGHT(rectangle3_weights[2406]), .FEAT_THRES(feature_thresholds[2406]), .FEAT_ABOVE(feature_aboves[2406]), .FEAT_BELOW(feature_belows[2406])) ac2406(.scan_win(scan_win2406), .scan_win_std_dev(scan_win_std_dev[2406]), .feature_accum(feature_accums[2406]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2407]), .RECT1_Y(rectangle1_ys[2407]), .RECT1_WIDTH(rectangle1_widths[2407]), .RECT1_HEIGHT(rectangle1_heights[2407]), .RECT1_WEIGHT(rectangle1_weights[2407]), .RECT2_X(rectangle2_xs[2407]), .RECT2_Y(rectangle2_ys[2407]), .RECT2_WIDTH(rectangle2_widths[2407]), .RECT2_HEIGHT(rectangle2_heights[2407]), .RECT2_WEIGHT(rectangle2_weights[2407]), .RECT3_X(rectangle3_xs[2407]), .RECT3_Y(rectangle3_ys[2407]), .RECT3_WIDTH(rectangle3_widths[2407]), .RECT3_HEIGHT(rectangle3_heights[2407]), .RECT3_WEIGHT(rectangle3_weights[2407]), .FEAT_THRES(feature_thresholds[2407]), .FEAT_ABOVE(feature_aboves[2407]), .FEAT_BELOW(feature_belows[2407])) ac2407(.scan_win(scan_win2407), .scan_win_std_dev(scan_win_std_dev[2407]), .feature_accum(feature_accums[2407]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2408]), .RECT1_Y(rectangle1_ys[2408]), .RECT1_WIDTH(rectangle1_widths[2408]), .RECT1_HEIGHT(rectangle1_heights[2408]), .RECT1_WEIGHT(rectangle1_weights[2408]), .RECT2_X(rectangle2_xs[2408]), .RECT2_Y(rectangle2_ys[2408]), .RECT2_WIDTH(rectangle2_widths[2408]), .RECT2_HEIGHT(rectangle2_heights[2408]), .RECT2_WEIGHT(rectangle2_weights[2408]), .RECT3_X(rectangle3_xs[2408]), .RECT3_Y(rectangle3_ys[2408]), .RECT3_WIDTH(rectangle3_widths[2408]), .RECT3_HEIGHT(rectangle3_heights[2408]), .RECT3_WEIGHT(rectangle3_weights[2408]), .FEAT_THRES(feature_thresholds[2408]), .FEAT_ABOVE(feature_aboves[2408]), .FEAT_BELOW(feature_belows[2408])) ac2408(.scan_win(scan_win2408), .scan_win_std_dev(scan_win_std_dev[2408]), .feature_accum(feature_accums[2408]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2409]), .RECT1_Y(rectangle1_ys[2409]), .RECT1_WIDTH(rectangle1_widths[2409]), .RECT1_HEIGHT(rectangle1_heights[2409]), .RECT1_WEIGHT(rectangle1_weights[2409]), .RECT2_X(rectangle2_xs[2409]), .RECT2_Y(rectangle2_ys[2409]), .RECT2_WIDTH(rectangle2_widths[2409]), .RECT2_HEIGHT(rectangle2_heights[2409]), .RECT2_WEIGHT(rectangle2_weights[2409]), .RECT3_X(rectangle3_xs[2409]), .RECT3_Y(rectangle3_ys[2409]), .RECT3_WIDTH(rectangle3_widths[2409]), .RECT3_HEIGHT(rectangle3_heights[2409]), .RECT3_WEIGHT(rectangle3_weights[2409]), .FEAT_THRES(feature_thresholds[2409]), .FEAT_ABOVE(feature_aboves[2409]), .FEAT_BELOW(feature_belows[2409])) ac2409(.scan_win(scan_win2409), .scan_win_std_dev(scan_win_std_dev[2409]), .feature_accum(feature_accums[2409]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2410]), .RECT1_Y(rectangle1_ys[2410]), .RECT1_WIDTH(rectangle1_widths[2410]), .RECT1_HEIGHT(rectangle1_heights[2410]), .RECT1_WEIGHT(rectangle1_weights[2410]), .RECT2_X(rectangle2_xs[2410]), .RECT2_Y(rectangle2_ys[2410]), .RECT2_WIDTH(rectangle2_widths[2410]), .RECT2_HEIGHT(rectangle2_heights[2410]), .RECT2_WEIGHT(rectangle2_weights[2410]), .RECT3_X(rectangle3_xs[2410]), .RECT3_Y(rectangle3_ys[2410]), .RECT3_WIDTH(rectangle3_widths[2410]), .RECT3_HEIGHT(rectangle3_heights[2410]), .RECT3_WEIGHT(rectangle3_weights[2410]), .FEAT_THRES(feature_thresholds[2410]), .FEAT_ABOVE(feature_aboves[2410]), .FEAT_BELOW(feature_belows[2410])) ac2410(.scan_win(scan_win2410), .scan_win_std_dev(scan_win_std_dev[2410]), .feature_accum(feature_accums[2410]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2411]), .RECT1_Y(rectangle1_ys[2411]), .RECT1_WIDTH(rectangle1_widths[2411]), .RECT1_HEIGHT(rectangle1_heights[2411]), .RECT1_WEIGHT(rectangle1_weights[2411]), .RECT2_X(rectangle2_xs[2411]), .RECT2_Y(rectangle2_ys[2411]), .RECT2_WIDTH(rectangle2_widths[2411]), .RECT2_HEIGHT(rectangle2_heights[2411]), .RECT2_WEIGHT(rectangle2_weights[2411]), .RECT3_X(rectangle3_xs[2411]), .RECT3_Y(rectangle3_ys[2411]), .RECT3_WIDTH(rectangle3_widths[2411]), .RECT3_HEIGHT(rectangle3_heights[2411]), .RECT3_WEIGHT(rectangle3_weights[2411]), .FEAT_THRES(feature_thresholds[2411]), .FEAT_ABOVE(feature_aboves[2411]), .FEAT_BELOW(feature_belows[2411])) ac2411(.scan_win(scan_win2411), .scan_win_std_dev(scan_win_std_dev[2411]), .feature_accum(feature_accums[2411]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2412]), .RECT1_Y(rectangle1_ys[2412]), .RECT1_WIDTH(rectangle1_widths[2412]), .RECT1_HEIGHT(rectangle1_heights[2412]), .RECT1_WEIGHT(rectangle1_weights[2412]), .RECT2_X(rectangle2_xs[2412]), .RECT2_Y(rectangle2_ys[2412]), .RECT2_WIDTH(rectangle2_widths[2412]), .RECT2_HEIGHT(rectangle2_heights[2412]), .RECT2_WEIGHT(rectangle2_weights[2412]), .RECT3_X(rectangle3_xs[2412]), .RECT3_Y(rectangle3_ys[2412]), .RECT3_WIDTH(rectangle3_widths[2412]), .RECT3_HEIGHT(rectangle3_heights[2412]), .RECT3_WEIGHT(rectangle3_weights[2412]), .FEAT_THRES(feature_thresholds[2412]), .FEAT_ABOVE(feature_aboves[2412]), .FEAT_BELOW(feature_belows[2412])) ac2412(.scan_win(scan_win2412), .scan_win_std_dev(scan_win_std_dev[2412]), .feature_accum(feature_accums[2412]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2413]), .RECT1_Y(rectangle1_ys[2413]), .RECT1_WIDTH(rectangle1_widths[2413]), .RECT1_HEIGHT(rectangle1_heights[2413]), .RECT1_WEIGHT(rectangle1_weights[2413]), .RECT2_X(rectangle2_xs[2413]), .RECT2_Y(rectangle2_ys[2413]), .RECT2_WIDTH(rectangle2_widths[2413]), .RECT2_HEIGHT(rectangle2_heights[2413]), .RECT2_WEIGHT(rectangle2_weights[2413]), .RECT3_X(rectangle3_xs[2413]), .RECT3_Y(rectangle3_ys[2413]), .RECT3_WIDTH(rectangle3_widths[2413]), .RECT3_HEIGHT(rectangle3_heights[2413]), .RECT3_WEIGHT(rectangle3_weights[2413]), .FEAT_THRES(feature_thresholds[2413]), .FEAT_ABOVE(feature_aboves[2413]), .FEAT_BELOW(feature_belows[2413])) ac2413(.scan_win(scan_win2413), .scan_win_std_dev(scan_win_std_dev[2413]), .feature_accum(feature_accums[2413]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2414]), .RECT1_Y(rectangle1_ys[2414]), .RECT1_WIDTH(rectangle1_widths[2414]), .RECT1_HEIGHT(rectangle1_heights[2414]), .RECT1_WEIGHT(rectangle1_weights[2414]), .RECT2_X(rectangle2_xs[2414]), .RECT2_Y(rectangle2_ys[2414]), .RECT2_WIDTH(rectangle2_widths[2414]), .RECT2_HEIGHT(rectangle2_heights[2414]), .RECT2_WEIGHT(rectangle2_weights[2414]), .RECT3_X(rectangle3_xs[2414]), .RECT3_Y(rectangle3_ys[2414]), .RECT3_WIDTH(rectangle3_widths[2414]), .RECT3_HEIGHT(rectangle3_heights[2414]), .RECT3_WEIGHT(rectangle3_weights[2414]), .FEAT_THRES(feature_thresholds[2414]), .FEAT_ABOVE(feature_aboves[2414]), .FEAT_BELOW(feature_belows[2414])) ac2414(.scan_win(scan_win2414), .scan_win_std_dev(scan_win_std_dev[2414]), .feature_accum(feature_accums[2414]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2415]), .RECT1_Y(rectangle1_ys[2415]), .RECT1_WIDTH(rectangle1_widths[2415]), .RECT1_HEIGHT(rectangle1_heights[2415]), .RECT1_WEIGHT(rectangle1_weights[2415]), .RECT2_X(rectangle2_xs[2415]), .RECT2_Y(rectangle2_ys[2415]), .RECT2_WIDTH(rectangle2_widths[2415]), .RECT2_HEIGHT(rectangle2_heights[2415]), .RECT2_WEIGHT(rectangle2_weights[2415]), .RECT3_X(rectangle3_xs[2415]), .RECT3_Y(rectangle3_ys[2415]), .RECT3_WIDTH(rectangle3_widths[2415]), .RECT3_HEIGHT(rectangle3_heights[2415]), .RECT3_WEIGHT(rectangle3_weights[2415]), .FEAT_THRES(feature_thresholds[2415]), .FEAT_ABOVE(feature_aboves[2415]), .FEAT_BELOW(feature_belows[2415])) ac2415(.scan_win(scan_win2415), .scan_win_std_dev(scan_win_std_dev[2415]), .feature_accum(feature_accums[2415]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2416]), .RECT1_Y(rectangle1_ys[2416]), .RECT1_WIDTH(rectangle1_widths[2416]), .RECT1_HEIGHT(rectangle1_heights[2416]), .RECT1_WEIGHT(rectangle1_weights[2416]), .RECT2_X(rectangle2_xs[2416]), .RECT2_Y(rectangle2_ys[2416]), .RECT2_WIDTH(rectangle2_widths[2416]), .RECT2_HEIGHT(rectangle2_heights[2416]), .RECT2_WEIGHT(rectangle2_weights[2416]), .RECT3_X(rectangle3_xs[2416]), .RECT3_Y(rectangle3_ys[2416]), .RECT3_WIDTH(rectangle3_widths[2416]), .RECT3_HEIGHT(rectangle3_heights[2416]), .RECT3_WEIGHT(rectangle3_weights[2416]), .FEAT_THRES(feature_thresholds[2416]), .FEAT_ABOVE(feature_aboves[2416]), .FEAT_BELOW(feature_belows[2416])) ac2416(.scan_win(scan_win2416), .scan_win_std_dev(scan_win_std_dev[2416]), .feature_accum(feature_accums[2416]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2417]), .RECT1_Y(rectangle1_ys[2417]), .RECT1_WIDTH(rectangle1_widths[2417]), .RECT1_HEIGHT(rectangle1_heights[2417]), .RECT1_WEIGHT(rectangle1_weights[2417]), .RECT2_X(rectangle2_xs[2417]), .RECT2_Y(rectangle2_ys[2417]), .RECT2_WIDTH(rectangle2_widths[2417]), .RECT2_HEIGHT(rectangle2_heights[2417]), .RECT2_WEIGHT(rectangle2_weights[2417]), .RECT3_X(rectangle3_xs[2417]), .RECT3_Y(rectangle3_ys[2417]), .RECT3_WIDTH(rectangle3_widths[2417]), .RECT3_HEIGHT(rectangle3_heights[2417]), .RECT3_WEIGHT(rectangle3_weights[2417]), .FEAT_THRES(feature_thresholds[2417]), .FEAT_ABOVE(feature_aboves[2417]), .FEAT_BELOW(feature_belows[2417])) ac2417(.scan_win(scan_win2417), .scan_win_std_dev(scan_win_std_dev[2417]), .feature_accum(feature_accums[2417]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2418]), .RECT1_Y(rectangle1_ys[2418]), .RECT1_WIDTH(rectangle1_widths[2418]), .RECT1_HEIGHT(rectangle1_heights[2418]), .RECT1_WEIGHT(rectangle1_weights[2418]), .RECT2_X(rectangle2_xs[2418]), .RECT2_Y(rectangle2_ys[2418]), .RECT2_WIDTH(rectangle2_widths[2418]), .RECT2_HEIGHT(rectangle2_heights[2418]), .RECT2_WEIGHT(rectangle2_weights[2418]), .RECT3_X(rectangle3_xs[2418]), .RECT3_Y(rectangle3_ys[2418]), .RECT3_WIDTH(rectangle3_widths[2418]), .RECT3_HEIGHT(rectangle3_heights[2418]), .RECT3_WEIGHT(rectangle3_weights[2418]), .FEAT_THRES(feature_thresholds[2418]), .FEAT_ABOVE(feature_aboves[2418]), .FEAT_BELOW(feature_belows[2418])) ac2418(.scan_win(scan_win2418), .scan_win_std_dev(scan_win_std_dev[2418]), .feature_accum(feature_accums[2418]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2419]), .RECT1_Y(rectangle1_ys[2419]), .RECT1_WIDTH(rectangle1_widths[2419]), .RECT1_HEIGHT(rectangle1_heights[2419]), .RECT1_WEIGHT(rectangle1_weights[2419]), .RECT2_X(rectangle2_xs[2419]), .RECT2_Y(rectangle2_ys[2419]), .RECT2_WIDTH(rectangle2_widths[2419]), .RECT2_HEIGHT(rectangle2_heights[2419]), .RECT2_WEIGHT(rectangle2_weights[2419]), .RECT3_X(rectangle3_xs[2419]), .RECT3_Y(rectangle3_ys[2419]), .RECT3_WIDTH(rectangle3_widths[2419]), .RECT3_HEIGHT(rectangle3_heights[2419]), .RECT3_WEIGHT(rectangle3_weights[2419]), .FEAT_THRES(feature_thresholds[2419]), .FEAT_ABOVE(feature_aboves[2419]), .FEAT_BELOW(feature_belows[2419])) ac2419(.scan_win(scan_win2419), .scan_win_std_dev(scan_win_std_dev[2419]), .feature_accum(feature_accums[2419]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2420]), .RECT1_Y(rectangle1_ys[2420]), .RECT1_WIDTH(rectangle1_widths[2420]), .RECT1_HEIGHT(rectangle1_heights[2420]), .RECT1_WEIGHT(rectangle1_weights[2420]), .RECT2_X(rectangle2_xs[2420]), .RECT2_Y(rectangle2_ys[2420]), .RECT2_WIDTH(rectangle2_widths[2420]), .RECT2_HEIGHT(rectangle2_heights[2420]), .RECT2_WEIGHT(rectangle2_weights[2420]), .RECT3_X(rectangle3_xs[2420]), .RECT3_Y(rectangle3_ys[2420]), .RECT3_WIDTH(rectangle3_widths[2420]), .RECT3_HEIGHT(rectangle3_heights[2420]), .RECT3_WEIGHT(rectangle3_weights[2420]), .FEAT_THRES(feature_thresholds[2420]), .FEAT_ABOVE(feature_aboves[2420]), .FEAT_BELOW(feature_belows[2420])) ac2420(.scan_win(scan_win2420), .scan_win_std_dev(scan_win_std_dev[2420]), .feature_accum(feature_accums[2420]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2421]), .RECT1_Y(rectangle1_ys[2421]), .RECT1_WIDTH(rectangle1_widths[2421]), .RECT1_HEIGHT(rectangle1_heights[2421]), .RECT1_WEIGHT(rectangle1_weights[2421]), .RECT2_X(rectangle2_xs[2421]), .RECT2_Y(rectangle2_ys[2421]), .RECT2_WIDTH(rectangle2_widths[2421]), .RECT2_HEIGHT(rectangle2_heights[2421]), .RECT2_WEIGHT(rectangle2_weights[2421]), .RECT3_X(rectangle3_xs[2421]), .RECT3_Y(rectangle3_ys[2421]), .RECT3_WIDTH(rectangle3_widths[2421]), .RECT3_HEIGHT(rectangle3_heights[2421]), .RECT3_WEIGHT(rectangle3_weights[2421]), .FEAT_THRES(feature_thresholds[2421]), .FEAT_ABOVE(feature_aboves[2421]), .FEAT_BELOW(feature_belows[2421])) ac2421(.scan_win(scan_win2421), .scan_win_std_dev(scan_win_std_dev[2421]), .feature_accum(feature_accums[2421]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2422]), .RECT1_Y(rectangle1_ys[2422]), .RECT1_WIDTH(rectangle1_widths[2422]), .RECT1_HEIGHT(rectangle1_heights[2422]), .RECT1_WEIGHT(rectangle1_weights[2422]), .RECT2_X(rectangle2_xs[2422]), .RECT2_Y(rectangle2_ys[2422]), .RECT2_WIDTH(rectangle2_widths[2422]), .RECT2_HEIGHT(rectangle2_heights[2422]), .RECT2_WEIGHT(rectangle2_weights[2422]), .RECT3_X(rectangle3_xs[2422]), .RECT3_Y(rectangle3_ys[2422]), .RECT3_WIDTH(rectangle3_widths[2422]), .RECT3_HEIGHT(rectangle3_heights[2422]), .RECT3_WEIGHT(rectangle3_weights[2422]), .FEAT_THRES(feature_thresholds[2422]), .FEAT_ABOVE(feature_aboves[2422]), .FEAT_BELOW(feature_belows[2422])) ac2422(.scan_win(scan_win2422), .scan_win_std_dev(scan_win_std_dev[2422]), .feature_accum(feature_accums[2422]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2423]), .RECT1_Y(rectangle1_ys[2423]), .RECT1_WIDTH(rectangle1_widths[2423]), .RECT1_HEIGHT(rectangle1_heights[2423]), .RECT1_WEIGHT(rectangle1_weights[2423]), .RECT2_X(rectangle2_xs[2423]), .RECT2_Y(rectangle2_ys[2423]), .RECT2_WIDTH(rectangle2_widths[2423]), .RECT2_HEIGHT(rectangle2_heights[2423]), .RECT2_WEIGHT(rectangle2_weights[2423]), .RECT3_X(rectangle3_xs[2423]), .RECT3_Y(rectangle3_ys[2423]), .RECT3_WIDTH(rectangle3_widths[2423]), .RECT3_HEIGHT(rectangle3_heights[2423]), .RECT3_WEIGHT(rectangle3_weights[2423]), .FEAT_THRES(feature_thresholds[2423]), .FEAT_ABOVE(feature_aboves[2423]), .FEAT_BELOW(feature_belows[2423])) ac2423(.scan_win(scan_win2423), .scan_win_std_dev(scan_win_std_dev[2423]), .feature_accum(feature_accums[2423]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2424]), .RECT1_Y(rectangle1_ys[2424]), .RECT1_WIDTH(rectangle1_widths[2424]), .RECT1_HEIGHT(rectangle1_heights[2424]), .RECT1_WEIGHT(rectangle1_weights[2424]), .RECT2_X(rectangle2_xs[2424]), .RECT2_Y(rectangle2_ys[2424]), .RECT2_WIDTH(rectangle2_widths[2424]), .RECT2_HEIGHT(rectangle2_heights[2424]), .RECT2_WEIGHT(rectangle2_weights[2424]), .RECT3_X(rectangle3_xs[2424]), .RECT3_Y(rectangle3_ys[2424]), .RECT3_WIDTH(rectangle3_widths[2424]), .RECT3_HEIGHT(rectangle3_heights[2424]), .RECT3_WEIGHT(rectangle3_weights[2424]), .FEAT_THRES(feature_thresholds[2424]), .FEAT_ABOVE(feature_aboves[2424]), .FEAT_BELOW(feature_belows[2424])) ac2424(.scan_win(scan_win2424), .scan_win_std_dev(scan_win_std_dev[2424]), .feature_accum(feature_accums[2424]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2425]), .RECT1_Y(rectangle1_ys[2425]), .RECT1_WIDTH(rectangle1_widths[2425]), .RECT1_HEIGHT(rectangle1_heights[2425]), .RECT1_WEIGHT(rectangle1_weights[2425]), .RECT2_X(rectangle2_xs[2425]), .RECT2_Y(rectangle2_ys[2425]), .RECT2_WIDTH(rectangle2_widths[2425]), .RECT2_HEIGHT(rectangle2_heights[2425]), .RECT2_WEIGHT(rectangle2_weights[2425]), .RECT3_X(rectangle3_xs[2425]), .RECT3_Y(rectangle3_ys[2425]), .RECT3_WIDTH(rectangle3_widths[2425]), .RECT3_HEIGHT(rectangle3_heights[2425]), .RECT3_WEIGHT(rectangle3_weights[2425]), .FEAT_THRES(feature_thresholds[2425]), .FEAT_ABOVE(feature_aboves[2425]), .FEAT_BELOW(feature_belows[2425])) ac2425(.scan_win(scan_win2425), .scan_win_std_dev(scan_win_std_dev[2425]), .feature_accum(feature_accums[2425]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2426]), .RECT1_Y(rectangle1_ys[2426]), .RECT1_WIDTH(rectangle1_widths[2426]), .RECT1_HEIGHT(rectangle1_heights[2426]), .RECT1_WEIGHT(rectangle1_weights[2426]), .RECT2_X(rectangle2_xs[2426]), .RECT2_Y(rectangle2_ys[2426]), .RECT2_WIDTH(rectangle2_widths[2426]), .RECT2_HEIGHT(rectangle2_heights[2426]), .RECT2_WEIGHT(rectangle2_weights[2426]), .RECT3_X(rectangle3_xs[2426]), .RECT3_Y(rectangle3_ys[2426]), .RECT3_WIDTH(rectangle3_widths[2426]), .RECT3_HEIGHT(rectangle3_heights[2426]), .RECT3_WEIGHT(rectangle3_weights[2426]), .FEAT_THRES(feature_thresholds[2426]), .FEAT_ABOVE(feature_aboves[2426]), .FEAT_BELOW(feature_belows[2426])) ac2426(.scan_win(scan_win2426), .scan_win_std_dev(scan_win_std_dev[2426]), .feature_accum(feature_accums[2426]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2427]), .RECT1_Y(rectangle1_ys[2427]), .RECT1_WIDTH(rectangle1_widths[2427]), .RECT1_HEIGHT(rectangle1_heights[2427]), .RECT1_WEIGHT(rectangle1_weights[2427]), .RECT2_X(rectangle2_xs[2427]), .RECT2_Y(rectangle2_ys[2427]), .RECT2_WIDTH(rectangle2_widths[2427]), .RECT2_HEIGHT(rectangle2_heights[2427]), .RECT2_WEIGHT(rectangle2_weights[2427]), .RECT3_X(rectangle3_xs[2427]), .RECT3_Y(rectangle3_ys[2427]), .RECT3_WIDTH(rectangle3_widths[2427]), .RECT3_HEIGHT(rectangle3_heights[2427]), .RECT3_WEIGHT(rectangle3_weights[2427]), .FEAT_THRES(feature_thresholds[2427]), .FEAT_ABOVE(feature_aboves[2427]), .FEAT_BELOW(feature_belows[2427])) ac2427(.scan_win(scan_win2427), .scan_win_std_dev(scan_win_std_dev[2427]), .feature_accum(feature_accums[2427]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2428]), .RECT1_Y(rectangle1_ys[2428]), .RECT1_WIDTH(rectangle1_widths[2428]), .RECT1_HEIGHT(rectangle1_heights[2428]), .RECT1_WEIGHT(rectangle1_weights[2428]), .RECT2_X(rectangle2_xs[2428]), .RECT2_Y(rectangle2_ys[2428]), .RECT2_WIDTH(rectangle2_widths[2428]), .RECT2_HEIGHT(rectangle2_heights[2428]), .RECT2_WEIGHT(rectangle2_weights[2428]), .RECT3_X(rectangle3_xs[2428]), .RECT3_Y(rectangle3_ys[2428]), .RECT3_WIDTH(rectangle3_widths[2428]), .RECT3_HEIGHT(rectangle3_heights[2428]), .RECT3_WEIGHT(rectangle3_weights[2428]), .FEAT_THRES(feature_thresholds[2428]), .FEAT_ABOVE(feature_aboves[2428]), .FEAT_BELOW(feature_belows[2428])) ac2428(.scan_win(scan_win2428), .scan_win_std_dev(scan_win_std_dev[2428]), .feature_accum(feature_accums[2428]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2429]), .RECT1_Y(rectangle1_ys[2429]), .RECT1_WIDTH(rectangle1_widths[2429]), .RECT1_HEIGHT(rectangle1_heights[2429]), .RECT1_WEIGHT(rectangle1_weights[2429]), .RECT2_X(rectangle2_xs[2429]), .RECT2_Y(rectangle2_ys[2429]), .RECT2_WIDTH(rectangle2_widths[2429]), .RECT2_HEIGHT(rectangle2_heights[2429]), .RECT2_WEIGHT(rectangle2_weights[2429]), .RECT3_X(rectangle3_xs[2429]), .RECT3_Y(rectangle3_ys[2429]), .RECT3_WIDTH(rectangle3_widths[2429]), .RECT3_HEIGHT(rectangle3_heights[2429]), .RECT3_WEIGHT(rectangle3_weights[2429]), .FEAT_THRES(feature_thresholds[2429]), .FEAT_ABOVE(feature_aboves[2429]), .FEAT_BELOW(feature_belows[2429])) ac2429(.scan_win(scan_win2429), .scan_win_std_dev(scan_win_std_dev[2429]), .feature_accum(feature_accums[2429]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2430]), .RECT1_Y(rectangle1_ys[2430]), .RECT1_WIDTH(rectangle1_widths[2430]), .RECT1_HEIGHT(rectangle1_heights[2430]), .RECT1_WEIGHT(rectangle1_weights[2430]), .RECT2_X(rectangle2_xs[2430]), .RECT2_Y(rectangle2_ys[2430]), .RECT2_WIDTH(rectangle2_widths[2430]), .RECT2_HEIGHT(rectangle2_heights[2430]), .RECT2_WEIGHT(rectangle2_weights[2430]), .RECT3_X(rectangle3_xs[2430]), .RECT3_Y(rectangle3_ys[2430]), .RECT3_WIDTH(rectangle3_widths[2430]), .RECT3_HEIGHT(rectangle3_heights[2430]), .RECT3_WEIGHT(rectangle3_weights[2430]), .FEAT_THRES(feature_thresholds[2430]), .FEAT_ABOVE(feature_aboves[2430]), .FEAT_BELOW(feature_belows[2430])) ac2430(.scan_win(scan_win2430), .scan_win_std_dev(scan_win_std_dev[2430]), .feature_accum(feature_accums[2430]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2431]), .RECT1_Y(rectangle1_ys[2431]), .RECT1_WIDTH(rectangle1_widths[2431]), .RECT1_HEIGHT(rectangle1_heights[2431]), .RECT1_WEIGHT(rectangle1_weights[2431]), .RECT2_X(rectangle2_xs[2431]), .RECT2_Y(rectangle2_ys[2431]), .RECT2_WIDTH(rectangle2_widths[2431]), .RECT2_HEIGHT(rectangle2_heights[2431]), .RECT2_WEIGHT(rectangle2_weights[2431]), .RECT3_X(rectangle3_xs[2431]), .RECT3_Y(rectangle3_ys[2431]), .RECT3_WIDTH(rectangle3_widths[2431]), .RECT3_HEIGHT(rectangle3_heights[2431]), .RECT3_WEIGHT(rectangle3_weights[2431]), .FEAT_THRES(feature_thresholds[2431]), .FEAT_ABOVE(feature_aboves[2431]), .FEAT_BELOW(feature_belows[2431])) ac2431(.scan_win(scan_win2431), .scan_win_std_dev(scan_win_std_dev[2431]), .feature_accum(feature_accums[2431]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2432]), .RECT1_Y(rectangle1_ys[2432]), .RECT1_WIDTH(rectangle1_widths[2432]), .RECT1_HEIGHT(rectangle1_heights[2432]), .RECT1_WEIGHT(rectangle1_weights[2432]), .RECT2_X(rectangle2_xs[2432]), .RECT2_Y(rectangle2_ys[2432]), .RECT2_WIDTH(rectangle2_widths[2432]), .RECT2_HEIGHT(rectangle2_heights[2432]), .RECT2_WEIGHT(rectangle2_weights[2432]), .RECT3_X(rectangle3_xs[2432]), .RECT3_Y(rectangle3_ys[2432]), .RECT3_WIDTH(rectangle3_widths[2432]), .RECT3_HEIGHT(rectangle3_heights[2432]), .RECT3_WEIGHT(rectangle3_weights[2432]), .FEAT_THRES(feature_thresholds[2432]), .FEAT_ABOVE(feature_aboves[2432]), .FEAT_BELOW(feature_belows[2432])) ac2432(.scan_win(scan_win2432), .scan_win_std_dev(scan_win_std_dev[2432]), .feature_accum(feature_accums[2432]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2433]), .RECT1_Y(rectangle1_ys[2433]), .RECT1_WIDTH(rectangle1_widths[2433]), .RECT1_HEIGHT(rectangle1_heights[2433]), .RECT1_WEIGHT(rectangle1_weights[2433]), .RECT2_X(rectangle2_xs[2433]), .RECT2_Y(rectangle2_ys[2433]), .RECT2_WIDTH(rectangle2_widths[2433]), .RECT2_HEIGHT(rectangle2_heights[2433]), .RECT2_WEIGHT(rectangle2_weights[2433]), .RECT3_X(rectangle3_xs[2433]), .RECT3_Y(rectangle3_ys[2433]), .RECT3_WIDTH(rectangle3_widths[2433]), .RECT3_HEIGHT(rectangle3_heights[2433]), .RECT3_WEIGHT(rectangle3_weights[2433]), .FEAT_THRES(feature_thresholds[2433]), .FEAT_ABOVE(feature_aboves[2433]), .FEAT_BELOW(feature_belows[2433])) ac2433(.scan_win(scan_win2433), .scan_win_std_dev(scan_win_std_dev[2433]), .feature_accum(feature_accums[2433]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2434]), .RECT1_Y(rectangle1_ys[2434]), .RECT1_WIDTH(rectangle1_widths[2434]), .RECT1_HEIGHT(rectangle1_heights[2434]), .RECT1_WEIGHT(rectangle1_weights[2434]), .RECT2_X(rectangle2_xs[2434]), .RECT2_Y(rectangle2_ys[2434]), .RECT2_WIDTH(rectangle2_widths[2434]), .RECT2_HEIGHT(rectangle2_heights[2434]), .RECT2_WEIGHT(rectangle2_weights[2434]), .RECT3_X(rectangle3_xs[2434]), .RECT3_Y(rectangle3_ys[2434]), .RECT3_WIDTH(rectangle3_widths[2434]), .RECT3_HEIGHT(rectangle3_heights[2434]), .RECT3_WEIGHT(rectangle3_weights[2434]), .FEAT_THRES(feature_thresholds[2434]), .FEAT_ABOVE(feature_aboves[2434]), .FEAT_BELOW(feature_belows[2434])) ac2434(.scan_win(scan_win2434), .scan_win_std_dev(scan_win_std_dev[2434]), .feature_accum(feature_accums[2434]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2435]), .RECT1_Y(rectangle1_ys[2435]), .RECT1_WIDTH(rectangle1_widths[2435]), .RECT1_HEIGHT(rectangle1_heights[2435]), .RECT1_WEIGHT(rectangle1_weights[2435]), .RECT2_X(rectangle2_xs[2435]), .RECT2_Y(rectangle2_ys[2435]), .RECT2_WIDTH(rectangle2_widths[2435]), .RECT2_HEIGHT(rectangle2_heights[2435]), .RECT2_WEIGHT(rectangle2_weights[2435]), .RECT3_X(rectangle3_xs[2435]), .RECT3_Y(rectangle3_ys[2435]), .RECT3_WIDTH(rectangle3_widths[2435]), .RECT3_HEIGHT(rectangle3_heights[2435]), .RECT3_WEIGHT(rectangle3_weights[2435]), .FEAT_THRES(feature_thresholds[2435]), .FEAT_ABOVE(feature_aboves[2435]), .FEAT_BELOW(feature_belows[2435])) ac2435(.scan_win(scan_win2435), .scan_win_std_dev(scan_win_std_dev[2435]), .feature_accum(feature_accums[2435]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2436]), .RECT1_Y(rectangle1_ys[2436]), .RECT1_WIDTH(rectangle1_widths[2436]), .RECT1_HEIGHT(rectangle1_heights[2436]), .RECT1_WEIGHT(rectangle1_weights[2436]), .RECT2_X(rectangle2_xs[2436]), .RECT2_Y(rectangle2_ys[2436]), .RECT2_WIDTH(rectangle2_widths[2436]), .RECT2_HEIGHT(rectangle2_heights[2436]), .RECT2_WEIGHT(rectangle2_weights[2436]), .RECT3_X(rectangle3_xs[2436]), .RECT3_Y(rectangle3_ys[2436]), .RECT3_WIDTH(rectangle3_widths[2436]), .RECT3_HEIGHT(rectangle3_heights[2436]), .RECT3_WEIGHT(rectangle3_weights[2436]), .FEAT_THRES(feature_thresholds[2436]), .FEAT_ABOVE(feature_aboves[2436]), .FEAT_BELOW(feature_belows[2436])) ac2436(.scan_win(scan_win2436), .scan_win_std_dev(scan_win_std_dev[2436]), .feature_accum(feature_accums[2436]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2437]), .RECT1_Y(rectangle1_ys[2437]), .RECT1_WIDTH(rectangle1_widths[2437]), .RECT1_HEIGHT(rectangle1_heights[2437]), .RECT1_WEIGHT(rectangle1_weights[2437]), .RECT2_X(rectangle2_xs[2437]), .RECT2_Y(rectangle2_ys[2437]), .RECT2_WIDTH(rectangle2_widths[2437]), .RECT2_HEIGHT(rectangle2_heights[2437]), .RECT2_WEIGHT(rectangle2_weights[2437]), .RECT3_X(rectangle3_xs[2437]), .RECT3_Y(rectangle3_ys[2437]), .RECT3_WIDTH(rectangle3_widths[2437]), .RECT3_HEIGHT(rectangle3_heights[2437]), .RECT3_WEIGHT(rectangle3_weights[2437]), .FEAT_THRES(feature_thresholds[2437]), .FEAT_ABOVE(feature_aboves[2437]), .FEAT_BELOW(feature_belows[2437])) ac2437(.scan_win(scan_win2437), .scan_win_std_dev(scan_win_std_dev[2437]), .feature_accum(feature_accums[2437]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2438]), .RECT1_Y(rectangle1_ys[2438]), .RECT1_WIDTH(rectangle1_widths[2438]), .RECT1_HEIGHT(rectangle1_heights[2438]), .RECT1_WEIGHT(rectangle1_weights[2438]), .RECT2_X(rectangle2_xs[2438]), .RECT2_Y(rectangle2_ys[2438]), .RECT2_WIDTH(rectangle2_widths[2438]), .RECT2_HEIGHT(rectangle2_heights[2438]), .RECT2_WEIGHT(rectangle2_weights[2438]), .RECT3_X(rectangle3_xs[2438]), .RECT3_Y(rectangle3_ys[2438]), .RECT3_WIDTH(rectangle3_widths[2438]), .RECT3_HEIGHT(rectangle3_heights[2438]), .RECT3_WEIGHT(rectangle3_weights[2438]), .FEAT_THRES(feature_thresholds[2438]), .FEAT_ABOVE(feature_aboves[2438]), .FEAT_BELOW(feature_belows[2438])) ac2438(.scan_win(scan_win2438), .scan_win_std_dev(scan_win_std_dev[2438]), .feature_accum(feature_accums[2438]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2439]), .RECT1_Y(rectangle1_ys[2439]), .RECT1_WIDTH(rectangle1_widths[2439]), .RECT1_HEIGHT(rectangle1_heights[2439]), .RECT1_WEIGHT(rectangle1_weights[2439]), .RECT2_X(rectangle2_xs[2439]), .RECT2_Y(rectangle2_ys[2439]), .RECT2_WIDTH(rectangle2_widths[2439]), .RECT2_HEIGHT(rectangle2_heights[2439]), .RECT2_WEIGHT(rectangle2_weights[2439]), .RECT3_X(rectangle3_xs[2439]), .RECT3_Y(rectangle3_ys[2439]), .RECT3_WIDTH(rectangle3_widths[2439]), .RECT3_HEIGHT(rectangle3_heights[2439]), .RECT3_WEIGHT(rectangle3_weights[2439]), .FEAT_THRES(feature_thresholds[2439]), .FEAT_ABOVE(feature_aboves[2439]), .FEAT_BELOW(feature_belows[2439])) ac2439(.scan_win(scan_win2439), .scan_win_std_dev(scan_win_std_dev[2439]), .feature_accum(feature_accums[2439]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2440]), .RECT1_Y(rectangle1_ys[2440]), .RECT1_WIDTH(rectangle1_widths[2440]), .RECT1_HEIGHT(rectangle1_heights[2440]), .RECT1_WEIGHT(rectangle1_weights[2440]), .RECT2_X(rectangle2_xs[2440]), .RECT2_Y(rectangle2_ys[2440]), .RECT2_WIDTH(rectangle2_widths[2440]), .RECT2_HEIGHT(rectangle2_heights[2440]), .RECT2_WEIGHT(rectangle2_weights[2440]), .RECT3_X(rectangle3_xs[2440]), .RECT3_Y(rectangle3_ys[2440]), .RECT3_WIDTH(rectangle3_widths[2440]), .RECT3_HEIGHT(rectangle3_heights[2440]), .RECT3_WEIGHT(rectangle3_weights[2440]), .FEAT_THRES(feature_thresholds[2440]), .FEAT_ABOVE(feature_aboves[2440]), .FEAT_BELOW(feature_belows[2440])) ac2440(.scan_win(scan_win2440), .scan_win_std_dev(scan_win_std_dev[2440]), .feature_accum(feature_accums[2440]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2441]), .RECT1_Y(rectangle1_ys[2441]), .RECT1_WIDTH(rectangle1_widths[2441]), .RECT1_HEIGHT(rectangle1_heights[2441]), .RECT1_WEIGHT(rectangle1_weights[2441]), .RECT2_X(rectangle2_xs[2441]), .RECT2_Y(rectangle2_ys[2441]), .RECT2_WIDTH(rectangle2_widths[2441]), .RECT2_HEIGHT(rectangle2_heights[2441]), .RECT2_WEIGHT(rectangle2_weights[2441]), .RECT3_X(rectangle3_xs[2441]), .RECT3_Y(rectangle3_ys[2441]), .RECT3_WIDTH(rectangle3_widths[2441]), .RECT3_HEIGHT(rectangle3_heights[2441]), .RECT3_WEIGHT(rectangle3_weights[2441]), .FEAT_THRES(feature_thresholds[2441]), .FEAT_ABOVE(feature_aboves[2441]), .FEAT_BELOW(feature_belows[2441])) ac2441(.scan_win(scan_win2441), .scan_win_std_dev(scan_win_std_dev[2441]), .feature_accum(feature_accums[2441]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2442]), .RECT1_Y(rectangle1_ys[2442]), .RECT1_WIDTH(rectangle1_widths[2442]), .RECT1_HEIGHT(rectangle1_heights[2442]), .RECT1_WEIGHT(rectangle1_weights[2442]), .RECT2_X(rectangle2_xs[2442]), .RECT2_Y(rectangle2_ys[2442]), .RECT2_WIDTH(rectangle2_widths[2442]), .RECT2_HEIGHT(rectangle2_heights[2442]), .RECT2_WEIGHT(rectangle2_weights[2442]), .RECT3_X(rectangle3_xs[2442]), .RECT3_Y(rectangle3_ys[2442]), .RECT3_WIDTH(rectangle3_widths[2442]), .RECT3_HEIGHT(rectangle3_heights[2442]), .RECT3_WEIGHT(rectangle3_weights[2442]), .FEAT_THRES(feature_thresholds[2442]), .FEAT_ABOVE(feature_aboves[2442]), .FEAT_BELOW(feature_belows[2442])) ac2442(.scan_win(scan_win2442), .scan_win_std_dev(scan_win_std_dev[2442]), .feature_accum(feature_accums[2442]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2443]), .RECT1_Y(rectangle1_ys[2443]), .RECT1_WIDTH(rectangle1_widths[2443]), .RECT1_HEIGHT(rectangle1_heights[2443]), .RECT1_WEIGHT(rectangle1_weights[2443]), .RECT2_X(rectangle2_xs[2443]), .RECT2_Y(rectangle2_ys[2443]), .RECT2_WIDTH(rectangle2_widths[2443]), .RECT2_HEIGHT(rectangle2_heights[2443]), .RECT2_WEIGHT(rectangle2_weights[2443]), .RECT3_X(rectangle3_xs[2443]), .RECT3_Y(rectangle3_ys[2443]), .RECT3_WIDTH(rectangle3_widths[2443]), .RECT3_HEIGHT(rectangle3_heights[2443]), .RECT3_WEIGHT(rectangle3_weights[2443]), .FEAT_THRES(feature_thresholds[2443]), .FEAT_ABOVE(feature_aboves[2443]), .FEAT_BELOW(feature_belows[2443])) ac2443(.scan_win(scan_win2443), .scan_win_std_dev(scan_win_std_dev[2443]), .feature_accum(feature_accums[2443]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2444]), .RECT1_Y(rectangle1_ys[2444]), .RECT1_WIDTH(rectangle1_widths[2444]), .RECT1_HEIGHT(rectangle1_heights[2444]), .RECT1_WEIGHT(rectangle1_weights[2444]), .RECT2_X(rectangle2_xs[2444]), .RECT2_Y(rectangle2_ys[2444]), .RECT2_WIDTH(rectangle2_widths[2444]), .RECT2_HEIGHT(rectangle2_heights[2444]), .RECT2_WEIGHT(rectangle2_weights[2444]), .RECT3_X(rectangle3_xs[2444]), .RECT3_Y(rectangle3_ys[2444]), .RECT3_WIDTH(rectangle3_widths[2444]), .RECT3_HEIGHT(rectangle3_heights[2444]), .RECT3_WEIGHT(rectangle3_weights[2444]), .FEAT_THRES(feature_thresholds[2444]), .FEAT_ABOVE(feature_aboves[2444]), .FEAT_BELOW(feature_belows[2444])) ac2444(.scan_win(scan_win2444), .scan_win_std_dev(scan_win_std_dev[2444]), .feature_accum(feature_accums[2444]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2445]), .RECT1_Y(rectangle1_ys[2445]), .RECT1_WIDTH(rectangle1_widths[2445]), .RECT1_HEIGHT(rectangle1_heights[2445]), .RECT1_WEIGHT(rectangle1_weights[2445]), .RECT2_X(rectangle2_xs[2445]), .RECT2_Y(rectangle2_ys[2445]), .RECT2_WIDTH(rectangle2_widths[2445]), .RECT2_HEIGHT(rectangle2_heights[2445]), .RECT2_WEIGHT(rectangle2_weights[2445]), .RECT3_X(rectangle3_xs[2445]), .RECT3_Y(rectangle3_ys[2445]), .RECT3_WIDTH(rectangle3_widths[2445]), .RECT3_HEIGHT(rectangle3_heights[2445]), .RECT3_WEIGHT(rectangle3_weights[2445]), .FEAT_THRES(feature_thresholds[2445]), .FEAT_ABOVE(feature_aboves[2445]), .FEAT_BELOW(feature_belows[2445])) ac2445(.scan_win(scan_win2445), .scan_win_std_dev(scan_win_std_dev[2445]), .feature_accum(feature_accums[2445]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2446]), .RECT1_Y(rectangle1_ys[2446]), .RECT1_WIDTH(rectangle1_widths[2446]), .RECT1_HEIGHT(rectangle1_heights[2446]), .RECT1_WEIGHT(rectangle1_weights[2446]), .RECT2_X(rectangle2_xs[2446]), .RECT2_Y(rectangle2_ys[2446]), .RECT2_WIDTH(rectangle2_widths[2446]), .RECT2_HEIGHT(rectangle2_heights[2446]), .RECT2_WEIGHT(rectangle2_weights[2446]), .RECT3_X(rectangle3_xs[2446]), .RECT3_Y(rectangle3_ys[2446]), .RECT3_WIDTH(rectangle3_widths[2446]), .RECT3_HEIGHT(rectangle3_heights[2446]), .RECT3_WEIGHT(rectangle3_weights[2446]), .FEAT_THRES(feature_thresholds[2446]), .FEAT_ABOVE(feature_aboves[2446]), .FEAT_BELOW(feature_belows[2446])) ac2446(.scan_win(scan_win2446), .scan_win_std_dev(scan_win_std_dev[2446]), .feature_accum(feature_accums[2446]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2447]), .RECT1_Y(rectangle1_ys[2447]), .RECT1_WIDTH(rectangle1_widths[2447]), .RECT1_HEIGHT(rectangle1_heights[2447]), .RECT1_WEIGHT(rectangle1_weights[2447]), .RECT2_X(rectangle2_xs[2447]), .RECT2_Y(rectangle2_ys[2447]), .RECT2_WIDTH(rectangle2_widths[2447]), .RECT2_HEIGHT(rectangle2_heights[2447]), .RECT2_WEIGHT(rectangle2_weights[2447]), .RECT3_X(rectangle3_xs[2447]), .RECT3_Y(rectangle3_ys[2447]), .RECT3_WIDTH(rectangle3_widths[2447]), .RECT3_HEIGHT(rectangle3_heights[2447]), .RECT3_WEIGHT(rectangle3_weights[2447]), .FEAT_THRES(feature_thresholds[2447]), .FEAT_ABOVE(feature_aboves[2447]), .FEAT_BELOW(feature_belows[2447])) ac2447(.scan_win(scan_win2447), .scan_win_std_dev(scan_win_std_dev[2447]), .feature_accum(feature_accums[2447]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2448]), .RECT1_Y(rectangle1_ys[2448]), .RECT1_WIDTH(rectangle1_widths[2448]), .RECT1_HEIGHT(rectangle1_heights[2448]), .RECT1_WEIGHT(rectangle1_weights[2448]), .RECT2_X(rectangle2_xs[2448]), .RECT2_Y(rectangle2_ys[2448]), .RECT2_WIDTH(rectangle2_widths[2448]), .RECT2_HEIGHT(rectangle2_heights[2448]), .RECT2_WEIGHT(rectangle2_weights[2448]), .RECT3_X(rectangle3_xs[2448]), .RECT3_Y(rectangle3_ys[2448]), .RECT3_WIDTH(rectangle3_widths[2448]), .RECT3_HEIGHT(rectangle3_heights[2448]), .RECT3_WEIGHT(rectangle3_weights[2448]), .FEAT_THRES(feature_thresholds[2448]), .FEAT_ABOVE(feature_aboves[2448]), .FEAT_BELOW(feature_belows[2448])) ac2448(.scan_win(scan_win2448), .scan_win_std_dev(scan_win_std_dev[2448]), .feature_accum(feature_accums[2448]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2449]), .RECT1_Y(rectangle1_ys[2449]), .RECT1_WIDTH(rectangle1_widths[2449]), .RECT1_HEIGHT(rectangle1_heights[2449]), .RECT1_WEIGHT(rectangle1_weights[2449]), .RECT2_X(rectangle2_xs[2449]), .RECT2_Y(rectangle2_ys[2449]), .RECT2_WIDTH(rectangle2_widths[2449]), .RECT2_HEIGHT(rectangle2_heights[2449]), .RECT2_WEIGHT(rectangle2_weights[2449]), .RECT3_X(rectangle3_xs[2449]), .RECT3_Y(rectangle3_ys[2449]), .RECT3_WIDTH(rectangle3_widths[2449]), .RECT3_HEIGHT(rectangle3_heights[2449]), .RECT3_WEIGHT(rectangle3_weights[2449]), .FEAT_THRES(feature_thresholds[2449]), .FEAT_ABOVE(feature_aboves[2449]), .FEAT_BELOW(feature_belows[2449])) ac2449(.scan_win(scan_win2449), .scan_win_std_dev(scan_win_std_dev[2449]), .feature_accum(feature_accums[2449]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2450]), .RECT1_Y(rectangle1_ys[2450]), .RECT1_WIDTH(rectangle1_widths[2450]), .RECT1_HEIGHT(rectangle1_heights[2450]), .RECT1_WEIGHT(rectangle1_weights[2450]), .RECT2_X(rectangle2_xs[2450]), .RECT2_Y(rectangle2_ys[2450]), .RECT2_WIDTH(rectangle2_widths[2450]), .RECT2_HEIGHT(rectangle2_heights[2450]), .RECT2_WEIGHT(rectangle2_weights[2450]), .RECT3_X(rectangle3_xs[2450]), .RECT3_Y(rectangle3_ys[2450]), .RECT3_WIDTH(rectangle3_widths[2450]), .RECT3_HEIGHT(rectangle3_heights[2450]), .RECT3_WEIGHT(rectangle3_weights[2450]), .FEAT_THRES(feature_thresholds[2450]), .FEAT_ABOVE(feature_aboves[2450]), .FEAT_BELOW(feature_belows[2450])) ac2450(.scan_win(scan_win2450), .scan_win_std_dev(scan_win_std_dev[2450]), .feature_accum(feature_accums[2450]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2451]), .RECT1_Y(rectangle1_ys[2451]), .RECT1_WIDTH(rectangle1_widths[2451]), .RECT1_HEIGHT(rectangle1_heights[2451]), .RECT1_WEIGHT(rectangle1_weights[2451]), .RECT2_X(rectangle2_xs[2451]), .RECT2_Y(rectangle2_ys[2451]), .RECT2_WIDTH(rectangle2_widths[2451]), .RECT2_HEIGHT(rectangle2_heights[2451]), .RECT2_WEIGHT(rectangle2_weights[2451]), .RECT3_X(rectangle3_xs[2451]), .RECT3_Y(rectangle3_ys[2451]), .RECT3_WIDTH(rectangle3_widths[2451]), .RECT3_HEIGHT(rectangle3_heights[2451]), .RECT3_WEIGHT(rectangle3_weights[2451]), .FEAT_THRES(feature_thresholds[2451]), .FEAT_ABOVE(feature_aboves[2451]), .FEAT_BELOW(feature_belows[2451])) ac2451(.scan_win(scan_win2451), .scan_win_std_dev(scan_win_std_dev[2451]), .feature_accum(feature_accums[2451]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2452]), .RECT1_Y(rectangle1_ys[2452]), .RECT1_WIDTH(rectangle1_widths[2452]), .RECT1_HEIGHT(rectangle1_heights[2452]), .RECT1_WEIGHT(rectangle1_weights[2452]), .RECT2_X(rectangle2_xs[2452]), .RECT2_Y(rectangle2_ys[2452]), .RECT2_WIDTH(rectangle2_widths[2452]), .RECT2_HEIGHT(rectangle2_heights[2452]), .RECT2_WEIGHT(rectangle2_weights[2452]), .RECT3_X(rectangle3_xs[2452]), .RECT3_Y(rectangle3_ys[2452]), .RECT3_WIDTH(rectangle3_widths[2452]), .RECT3_HEIGHT(rectangle3_heights[2452]), .RECT3_WEIGHT(rectangle3_weights[2452]), .FEAT_THRES(feature_thresholds[2452]), .FEAT_ABOVE(feature_aboves[2452]), .FEAT_BELOW(feature_belows[2452])) ac2452(.scan_win(scan_win2452), .scan_win_std_dev(scan_win_std_dev[2452]), .feature_accum(feature_accums[2452]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2453]), .RECT1_Y(rectangle1_ys[2453]), .RECT1_WIDTH(rectangle1_widths[2453]), .RECT1_HEIGHT(rectangle1_heights[2453]), .RECT1_WEIGHT(rectangle1_weights[2453]), .RECT2_X(rectangle2_xs[2453]), .RECT2_Y(rectangle2_ys[2453]), .RECT2_WIDTH(rectangle2_widths[2453]), .RECT2_HEIGHT(rectangle2_heights[2453]), .RECT2_WEIGHT(rectangle2_weights[2453]), .RECT3_X(rectangle3_xs[2453]), .RECT3_Y(rectangle3_ys[2453]), .RECT3_WIDTH(rectangle3_widths[2453]), .RECT3_HEIGHT(rectangle3_heights[2453]), .RECT3_WEIGHT(rectangle3_weights[2453]), .FEAT_THRES(feature_thresholds[2453]), .FEAT_ABOVE(feature_aboves[2453]), .FEAT_BELOW(feature_belows[2453])) ac2453(.scan_win(scan_win2453), .scan_win_std_dev(scan_win_std_dev[2453]), .feature_accum(feature_accums[2453]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2454]), .RECT1_Y(rectangle1_ys[2454]), .RECT1_WIDTH(rectangle1_widths[2454]), .RECT1_HEIGHT(rectangle1_heights[2454]), .RECT1_WEIGHT(rectangle1_weights[2454]), .RECT2_X(rectangle2_xs[2454]), .RECT2_Y(rectangle2_ys[2454]), .RECT2_WIDTH(rectangle2_widths[2454]), .RECT2_HEIGHT(rectangle2_heights[2454]), .RECT2_WEIGHT(rectangle2_weights[2454]), .RECT3_X(rectangle3_xs[2454]), .RECT3_Y(rectangle3_ys[2454]), .RECT3_WIDTH(rectangle3_widths[2454]), .RECT3_HEIGHT(rectangle3_heights[2454]), .RECT3_WEIGHT(rectangle3_weights[2454]), .FEAT_THRES(feature_thresholds[2454]), .FEAT_ABOVE(feature_aboves[2454]), .FEAT_BELOW(feature_belows[2454])) ac2454(.scan_win(scan_win2454), .scan_win_std_dev(scan_win_std_dev[2454]), .feature_accum(feature_accums[2454]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2455]), .RECT1_Y(rectangle1_ys[2455]), .RECT1_WIDTH(rectangle1_widths[2455]), .RECT1_HEIGHT(rectangle1_heights[2455]), .RECT1_WEIGHT(rectangle1_weights[2455]), .RECT2_X(rectangle2_xs[2455]), .RECT2_Y(rectangle2_ys[2455]), .RECT2_WIDTH(rectangle2_widths[2455]), .RECT2_HEIGHT(rectangle2_heights[2455]), .RECT2_WEIGHT(rectangle2_weights[2455]), .RECT3_X(rectangle3_xs[2455]), .RECT3_Y(rectangle3_ys[2455]), .RECT3_WIDTH(rectangle3_widths[2455]), .RECT3_HEIGHT(rectangle3_heights[2455]), .RECT3_WEIGHT(rectangle3_weights[2455]), .FEAT_THRES(feature_thresholds[2455]), .FEAT_ABOVE(feature_aboves[2455]), .FEAT_BELOW(feature_belows[2455])) ac2455(.scan_win(scan_win2455), .scan_win_std_dev(scan_win_std_dev[2455]), .feature_accum(feature_accums[2455]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2456]), .RECT1_Y(rectangle1_ys[2456]), .RECT1_WIDTH(rectangle1_widths[2456]), .RECT1_HEIGHT(rectangle1_heights[2456]), .RECT1_WEIGHT(rectangle1_weights[2456]), .RECT2_X(rectangle2_xs[2456]), .RECT2_Y(rectangle2_ys[2456]), .RECT2_WIDTH(rectangle2_widths[2456]), .RECT2_HEIGHT(rectangle2_heights[2456]), .RECT2_WEIGHT(rectangle2_weights[2456]), .RECT3_X(rectangle3_xs[2456]), .RECT3_Y(rectangle3_ys[2456]), .RECT3_WIDTH(rectangle3_widths[2456]), .RECT3_HEIGHT(rectangle3_heights[2456]), .RECT3_WEIGHT(rectangle3_weights[2456]), .FEAT_THRES(feature_thresholds[2456]), .FEAT_ABOVE(feature_aboves[2456]), .FEAT_BELOW(feature_belows[2456])) ac2456(.scan_win(scan_win2456), .scan_win_std_dev(scan_win_std_dev[2456]), .feature_accum(feature_accums[2456]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2457]), .RECT1_Y(rectangle1_ys[2457]), .RECT1_WIDTH(rectangle1_widths[2457]), .RECT1_HEIGHT(rectangle1_heights[2457]), .RECT1_WEIGHT(rectangle1_weights[2457]), .RECT2_X(rectangle2_xs[2457]), .RECT2_Y(rectangle2_ys[2457]), .RECT2_WIDTH(rectangle2_widths[2457]), .RECT2_HEIGHT(rectangle2_heights[2457]), .RECT2_WEIGHT(rectangle2_weights[2457]), .RECT3_X(rectangle3_xs[2457]), .RECT3_Y(rectangle3_ys[2457]), .RECT3_WIDTH(rectangle3_widths[2457]), .RECT3_HEIGHT(rectangle3_heights[2457]), .RECT3_WEIGHT(rectangle3_weights[2457]), .FEAT_THRES(feature_thresholds[2457]), .FEAT_ABOVE(feature_aboves[2457]), .FEAT_BELOW(feature_belows[2457])) ac2457(.scan_win(scan_win2457), .scan_win_std_dev(scan_win_std_dev[2457]), .feature_accum(feature_accums[2457]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2458]), .RECT1_Y(rectangle1_ys[2458]), .RECT1_WIDTH(rectangle1_widths[2458]), .RECT1_HEIGHT(rectangle1_heights[2458]), .RECT1_WEIGHT(rectangle1_weights[2458]), .RECT2_X(rectangle2_xs[2458]), .RECT2_Y(rectangle2_ys[2458]), .RECT2_WIDTH(rectangle2_widths[2458]), .RECT2_HEIGHT(rectangle2_heights[2458]), .RECT2_WEIGHT(rectangle2_weights[2458]), .RECT3_X(rectangle3_xs[2458]), .RECT3_Y(rectangle3_ys[2458]), .RECT3_WIDTH(rectangle3_widths[2458]), .RECT3_HEIGHT(rectangle3_heights[2458]), .RECT3_WEIGHT(rectangle3_weights[2458]), .FEAT_THRES(feature_thresholds[2458]), .FEAT_ABOVE(feature_aboves[2458]), .FEAT_BELOW(feature_belows[2458])) ac2458(.scan_win(scan_win2458), .scan_win_std_dev(scan_win_std_dev[2458]), .feature_accum(feature_accums[2458]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2459]), .RECT1_Y(rectangle1_ys[2459]), .RECT1_WIDTH(rectangle1_widths[2459]), .RECT1_HEIGHT(rectangle1_heights[2459]), .RECT1_WEIGHT(rectangle1_weights[2459]), .RECT2_X(rectangle2_xs[2459]), .RECT2_Y(rectangle2_ys[2459]), .RECT2_WIDTH(rectangle2_widths[2459]), .RECT2_HEIGHT(rectangle2_heights[2459]), .RECT2_WEIGHT(rectangle2_weights[2459]), .RECT3_X(rectangle3_xs[2459]), .RECT3_Y(rectangle3_ys[2459]), .RECT3_WIDTH(rectangle3_widths[2459]), .RECT3_HEIGHT(rectangle3_heights[2459]), .RECT3_WEIGHT(rectangle3_weights[2459]), .FEAT_THRES(feature_thresholds[2459]), .FEAT_ABOVE(feature_aboves[2459]), .FEAT_BELOW(feature_belows[2459])) ac2459(.scan_win(scan_win2459), .scan_win_std_dev(scan_win_std_dev[2459]), .feature_accum(feature_accums[2459]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2460]), .RECT1_Y(rectangle1_ys[2460]), .RECT1_WIDTH(rectangle1_widths[2460]), .RECT1_HEIGHT(rectangle1_heights[2460]), .RECT1_WEIGHT(rectangle1_weights[2460]), .RECT2_X(rectangle2_xs[2460]), .RECT2_Y(rectangle2_ys[2460]), .RECT2_WIDTH(rectangle2_widths[2460]), .RECT2_HEIGHT(rectangle2_heights[2460]), .RECT2_WEIGHT(rectangle2_weights[2460]), .RECT3_X(rectangle3_xs[2460]), .RECT3_Y(rectangle3_ys[2460]), .RECT3_WIDTH(rectangle3_widths[2460]), .RECT3_HEIGHT(rectangle3_heights[2460]), .RECT3_WEIGHT(rectangle3_weights[2460]), .FEAT_THRES(feature_thresholds[2460]), .FEAT_ABOVE(feature_aboves[2460]), .FEAT_BELOW(feature_belows[2460])) ac2460(.scan_win(scan_win2460), .scan_win_std_dev(scan_win_std_dev[2460]), .feature_accum(feature_accums[2460]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2461]), .RECT1_Y(rectangle1_ys[2461]), .RECT1_WIDTH(rectangle1_widths[2461]), .RECT1_HEIGHT(rectangle1_heights[2461]), .RECT1_WEIGHT(rectangle1_weights[2461]), .RECT2_X(rectangle2_xs[2461]), .RECT2_Y(rectangle2_ys[2461]), .RECT2_WIDTH(rectangle2_widths[2461]), .RECT2_HEIGHT(rectangle2_heights[2461]), .RECT2_WEIGHT(rectangle2_weights[2461]), .RECT3_X(rectangle3_xs[2461]), .RECT3_Y(rectangle3_ys[2461]), .RECT3_WIDTH(rectangle3_widths[2461]), .RECT3_HEIGHT(rectangle3_heights[2461]), .RECT3_WEIGHT(rectangle3_weights[2461]), .FEAT_THRES(feature_thresholds[2461]), .FEAT_ABOVE(feature_aboves[2461]), .FEAT_BELOW(feature_belows[2461])) ac2461(.scan_win(scan_win2461), .scan_win_std_dev(scan_win_std_dev[2461]), .feature_accum(feature_accums[2461]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2462]), .RECT1_Y(rectangle1_ys[2462]), .RECT1_WIDTH(rectangle1_widths[2462]), .RECT1_HEIGHT(rectangle1_heights[2462]), .RECT1_WEIGHT(rectangle1_weights[2462]), .RECT2_X(rectangle2_xs[2462]), .RECT2_Y(rectangle2_ys[2462]), .RECT2_WIDTH(rectangle2_widths[2462]), .RECT2_HEIGHT(rectangle2_heights[2462]), .RECT2_WEIGHT(rectangle2_weights[2462]), .RECT3_X(rectangle3_xs[2462]), .RECT3_Y(rectangle3_ys[2462]), .RECT3_WIDTH(rectangle3_widths[2462]), .RECT3_HEIGHT(rectangle3_heights[2462]), .RECT3_WEIGHT(rectangle3_weights[2462]), .FEAT_THRES(feature_thresholds[2462]), .FEAT_ABOVE(feature_aboves[2462]), .FEAT_BELOW(feature_belows[2462])) ac2462(.scan_win(scan_win2462), .scan_win_std_dev(scan_win_std_dev[2462]), .feature_accum(feature_accums[2462]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2463]), .RECT1_Y(rectangle1_ys[2463]), .RECT1_WIDTH(rectangle1_widths[2463]), .RECT1_HEIGHT(rectangle1_heights[2463]), .RECT1_WEIGHT(rectangle1_weights[2463]), .RECT2_X(rectangle2_xs[2463]), .RECT2_Y(rectangle2_ys[2463]), .RECT2_WIDTH(rectangle2_widths[2463]), .RECT2_HEIGHT(rectangle2_heights[2463]), .RECT2_WEIGHT(rectangle2_weights[2463]), .RECT3_X(rectangle3_xs[2463]), .RECT3_Y(rectangle3_ys[2463]), .RECT3_WIDTH(rectangle3_widths[2463]), .RECT3_HEIGHT(rectangle3_heights[2463]), .RECT3_WEIGHT(rectangle3_weights[2463]), .FEAT_THRES(feature_thresholds[2463]), .FEAT_ABOVE(feature_aboves[2463]), .FEAT_BELOW(feature_belows[2463])) ac2463(.scan_win(scan_win2463), .scan_win_std_dev(scan_win_std_dev[2463]), .feature_accum(feature_accums[2463]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2464]), .RECT1_Y(rectangle1_ys[2464]), .RECT1_WIDTH(rectangle1_widths[2464]), .RECT1_HEIGHT(rectangle1_heights[2464]), .RECT1_WEIGHT(rectangle1_weights[2464]), .RECT2_X(rectangle2_xs[2464]), .RECT2_Y(rectangle2_ys[2464]), .RECT2_WIDTH(rectangle2_widths[2464]), .RECT2_HEIGHT(rectangle2_heights[2464]), .RECT2_WEIGHT(rectangle2_weights[2464]), .RECT3_X(rectangle3_xs[2464]), .RECT3_Y(rectangle3_ys[2464]), .RECT3_WIDTH(rectangle3_widths[2464]), .RECT3_HEIGHT(rectangle3_heights[2464]), .RECT3_WEIGHT(rectangle3_weights[2464]), .FEAT_THRES(feature_thresholds[2464]), .FEAT_ABOVE(feature_aboves[2464]), .FEAT_BELOW(feature_belows[2464])) ac2464(.scan_win(scan_win2464), .scan_win_std_dev(scan_win_std_dev[2464]), .feature_accum(feature_accums[2464]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2465]), .RECT1_Y(rectangle1_ys[2465]), .RECT1_WIDTH(rectangle1_widths[2465]), .RECT1_HEIGHT(rectangle1_heights[2465]), .RECT1_WEIGHT(rectangle1_weights[2465]), .RECT2_X(rectangle2_xs[2465]), .RECT2_Y(rectangle2_ys[2465]), .RECT2_WIDTH(rectangle2_widths[2465]), .RECT2_HEIGHT(rectangle2_heights[2465]), .RECT2_WEIGHT(rectangle2_weights[2465]), .RECT3_X(rectangle3_xs[2465]), .RECT3_Y(rectangle3_ys[2465]), .RECT3_WIDTH(rectangle3_widths[2465]), .RECT3_HEIGHT(rectangle3_heights[2465]), .RECT3_WEIGHT(rectangle3_weights[2465]), .FEAT_THRES(feature_thresholds[2465]), .FEAT_ABOVE(feature_aboves[2465]), .FEAT_BELOW(feature_belows[2465])) ac2465(.scan_win(scan_win2465), .scan_win_std_dev(scan_win_std_dev[2465]), .feature_accum(feature_accums[2465]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2466]), .RECT1_Y(rectangle1_ys[2466]), .RECT1_WIDTH(rectangle1_widths[2466]), .RECT1_HEIGHT(rectangle1_heights[2466]), .RECT1_WEIGHT(rectangle1_weights[2466]), .RECT2_X(rectangle2_xs[2466]), .RECT2_Y(rectangle2_ys[2466]), .RECT2_WIDTH(rectangle2_widths[2466]), .RECT2_HEIGHT(rectangle2_heights[2466]), .RECT2_WEIGHT(rectangle2_weights[2466]), .RECT3_X(rectangle3_xs[2466]), .RECT3_Y(rectangle3_ys[2466]), .RECT3_WIDTH(rectangle3_widths[2466]), .RECT3_HEIGHT(rectangle3_heights[2466]), .RECT3_WEIGHT(rectangle3_weights[2466]), .FEAT_THRES(feature_thresholds[2466]), .FEAT_ABOVE(feature_aboves[2466]), .FEAT_BELOW(feature_belows[2466])) ac2466(.scan_win(scan_win2466), .scan_win_std_dev(scan_win_std_dev[2466]), .feature_accum(feature_accums[2466]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2467]), .RECT1_Y(rectangle1_ys[2467]), .RECT1_WIDTH(rectangle1_widths[2467]), .RECT1_HEIGHT(rectangle1_heights[2467]), .RECT1_WEIGHT(rectangle1_weights[2467]), .RECT2_X(rectangle2_xs[2467]), .RECT2_Y(rectangle2_ys[2467]), .RECT2_WIDTH(rectangle2_widths[2467]), .RECT2_HEIGHT(rectangle2_heights[2467]), .RECT2_WEIGHT(rectangle2_weights[2467]), .RECT3_X(rectangle3_xs[2467]), .RECT3_Y(rectangle3_ys[2467]), .RECT3_WIDTH(rectangle3_widths[2467]), .RECT3_HEIGHT(rectangle3_heights[2467]), .RECT3_WEIGHT(rectangle3_weights[2467]), .FEAT_THRES(feature_thresholds[2467]), .FEAT_ABOVE(feature_aboves[2467]), .FEAT_BELOW(feature_belows[2467])) ac2467(.scan_win(scan_win2467), .scan_win_std_dev(scan_win_std_dev[2467]), .feature_accum(feature_accums[2467]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2468]), .RECT1_Y(rectangle1_ys[2468]), .RECT1_WIDTH(rectangle1_widths[2468]), .RECT1_HEIGHT(rectangle1_heights[2468]), .RECT1_WEIGHT(rectangle1_weights[2468]), .RECT2_X(rectangle2_xs[2468]), .RECT2_Y(rectangle2_ys[2468]), .RECT2_WIDTH(rectangle2_widths[2468]), .RECT2_HEIGHT(rectangle2_heights[2468]), .RECT2_WEIGHT(rectangle2_weights[2468]), .RECT3_X(rectangle3_xs[2468]), .RECT3_Y(rectangle3_ys[2468]), .RECT3_WIDTH(rectangle3_widths[2468]), .RECT3_HEIGHT(rectangle3_heights[2468]), .RECT3_WEIGHT(rectangle3_weights[2468]), .FEAT_THRES(feature_thresholds[2468]), .FEAT_ABOVE(feature_aboves[2468]), .FEAT_BELOW(feature_belows[2468])) ac2468(.scan_win(scan_win2468), .scan_win_std_dev(scan_win_std_dev[2468]), .feature_accum(feature_accums[2468]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2469]), .RECT1_Y(rectangle1_ys[2469]), .RECT1_WIDTH(rectangle1_widths[2469]), .RECT1_HEIGHT(rectangle1_heights[2469]), .RECT1_WEIGHT(rectangle1_weights[2469]), .RECT2_X(rectangle2_xs[2469]), .RECT2_Y(rectangle2_ys[2469]), .RECT2_WIDTH(rectangle2_widths[2469]), .RECT2_HEIGHT(rectangle2_heights[2469]), .RECT2_WEIGHT(rectangle2_weights[2469]), .RECT3_X(rectangle3_xs[2469]), .RECT3_Y(rectangle3_ys[2469]), .RECT3_WIDTH(rectangle3_widths[2469]), .RECT3_HEIGHT(rectangle3_heights[2469]), .RECT3_WEIGHT(rectangle3_weights[2469]), .FEAT_THRES(feature_thresholds[2469]), .FEAT_ABOVE(feature_aboves[2469]), .FEAT_BELOW(feature_belows[2469])) ac2469(.scan_win(scan_win2469), .scan_win_std_dev(scan_win_std_dev[2469]), .feature_accum(feature_accums[2469]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2470]), .RECT1_Y(rectangle1_ys[2470]), .RECT1_WIDTH(rectangle1_widths[2470]), .RECT1_HEIGHT(rectangle1_heights[2470]), .RECT1_WEIGHT(rectangle1_weights[2470]), .RECT2_X(rectangle2_xs[2470]), .RECT2_Y(rectangle2_ys[2470]), .RECT2_WIDTH(rectangle2_widths[2470]), .RECT2_HEIGHT(rectangle2_heights[2470]), .RECT2_WEIGHT(rectangle2_weights[2470]), .RECT3_X(rectangle3_xs[2470]), .RECT3_Y(rectangle3_ys[2470]), .RECT3_WIDTH(rectangle3_widths[2470]), .RECT3_HEIGHT(rectangle3_heights[2470]), .RECT3_WEIGHT(rectangle3_weights[2470]), .FEAT_THRES(feature_thresholds[2470]), .FEAT_ABOVE(feature_aboves[2470]), .FEAT_BELOW(feature_belows[2470])) ac2470(.scan_win(scan_win2470), .scan_win_std_dev(scan_win_std_dev[2470]), .feature_accum(feature_accums[2470]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2471]), .RECT1_Y(rectangle1_ys[2471]), .RECT1_WIDTH(rectangle1_widths[2471]), .RECT1_HEIGHT(rectangle1_heights[2471]), .RECT1_WEIGHT(rectangle1_weights[2471]), .RECT2_X(rectangle2_xs[2471]), .RECT2_Y(rectangle2_ys[2471]), .RECT2_WIDTH(rectangle2_widths[2471]), .RECT2_HEIGHT(rectangle2_heights[2471]), .RECT2_WEIGHT(rectangle2_weights[2471]), .RECT3_X(rectangle3_xs[2471]), .RECT3_Y(rectangle3_ys[2471]), .RECT3_WIDTH(rectangle3_widths[2471]), .RECT3_HEIGHT(rectangle3_heights[2471]), .RECT3_WEIGHT(rectangle3_weights[2471]), .FEAT_THRES(feature_thresholds[2471]), .FEAT_ABOVE(feature_aboves[2471]), .FEAT_BELOW(feature_belows[2471])) ac2471(.scan_win(scan_win2471), .scan_win_std_dev(scan_win_std_dev[2471]), .feature_accum(feature_accums[2471]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2472]), .RECT1_Y(rectangle1_ys[2472]), .RECT1_WIDTH(rectangle1_widths[2472]), .RECT1_HEIGHT(rectangle1_heights[2472]), .RECT1_WEIGHT(rectangle1_weights[2472]), .RECT2_X(rectangle2_xs[2472]), .RECT2_Y(rectangle2_ys[2472]), .RECT2_WIDTH(rectangle2_widths[2472]), .RECT2_HEIGHT(rectangle2_heights[2472]), .RECT2_WEIGHT(rectangle2_weights[2472]), .RECT3_X(rectangle3_xs[2472]), .RECT3_Y(rectangle3_ys[2472]), .RECT3_WIDTH(rectangle3_widths[2472]), .RECT3_HEIGHT(rectangle3_heights[2472]), .RECT3_WEIGHT(rectangle3_weights[2472]), .FEAT_THRES(feature_thresholds[2472]), .FEAT_ABOVE(feature_aboves[2472]), .FEAT_BELOW(feature_belows[2472])) ac2472(.scan_win(scan_win2472), .scan_win_std_dev(scan_win_std_dev[2472]), .feature_accum(feature_accums[2472]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2473]), .RECT1_Y(rectangle1_ys[2473]), .RECT1_WIDTH(rectangle1_widths[2473]), .RECT1_HEIGHT(rectangle1_heights[2473]), .RECT1_WEIGHT(rectangle1_weights[2473]), .RECT2_X(rectangle2_xs[2473]), .RECT2_Y(rectangle2_ys[2473]), .RECT2_WIDTH(rectangle2_widths[2473]), .RECT2_HEIGHT(rectangle2_heights[2473]), .RECT2_WEIGHT(rectangle2_weights[2473]), .RECT3_X(rectangle3_xs[2473]), .RECT3_Y(rectangle3_ys[2473]), .RECT3_WIDTH(rectangle3_widths[2473]), .RECT3_HEIGHT(rectangle3_heights[2473]), .RECT3_WEIGHT(rectangle3_weights[2473]), .FEAT_THRES(feature_thresholds[2473]), .FEAT_ABOVE(feature_aboves[2473]), .FEAT_BELOW(feature_belows[2473])) ac2473(.scan_win(scan_win2473), .scan_win_std_dev(scan_win_std_dev[2473]), .feature_accum(feature_accums[2473]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2474]), .RECT1_Y(rectangle1_ys[2474]), .RECT1_WIDTH(rectangle1_widths[2474]), .RECT1_HEIGHT(rectangle1_heights[2474]), .RECT1_WEIGHT(rectangle1_weights[2474]), .RECT2_X(rectangle2_xs[2474]), .RECT2_Y(rectangle2_ys[2474]), .RECT2_WIDTH(rectangle2_widths[2474]), .RECT2_HEIGHT(rectangle2_heights[2474]), .RECT2_WEIGHT(rectangle2_weights[2474]), .RECT3_X(rectangle3_xs[2474]), .RECT3_Y(rectangle3_ys[2474]), .RECT3_WIDTH(rectangle3_widths[2474]), .RECT3_HEIGHT(rectangle3_heights[2474]), .RECT3_WEIGHT(rectangle3_weights[2474]), .FEAT_THRES(feature_thresholds[2474]), .FEAT_ABOVE(feature_aboves[2474]), .FEAT_BELOW(feature_belows[2474])) ac2474(.scan_win(scan_win2474), .scan_win_std_dev(scan_win_std_dev[2474]), .feature_accum(feature_accums[2474]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2475]), .RECT1_Y(rectangle1_ys[2475]), .RECT1_WIDTH(rectangle1_widths[2475]), .RECT1_HEIGHT(rectangle1_heights[2475]), .RECT1_WEIGHT(rectangle1_weights[2475]), .RECT2_X(rectangle2_xs[2475]), .RECT2_Y(rectangle2_ys[2475]), .RECT2_WIDTH(rectangle2_widths[2475]), .RECT2_HEIGHT(rectangle2_heights[2475]), .RECT2_WEIGHT(rectangle2_weights[2475]), .RECT3_X(rectangle3_xs[2475]), .RECT3_Y(rectangle3_ys[2475]), .RECT3_WIDTH(rectangle3_widths[2475]), .RECT3_HEIGHT(rectangle3_heights[2475]), .RECT3_WEIGHT(rectangle3_weights[2475]), .FEAT_THRES(feature_thresholds[2475]), .FEAT_ABOVE(feature_aboves[2475]), .FEAT_BELOW(feature_belows[2475])) ac2475(.scan_win(scan_win2475), .scan_win_std_dev(scan_win_std_dev[2475]), .feature_accum(feature_accums[2475]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2476]), .RECT1_Y(rectangle1_ys[2476]), .RECT1_WIDTH(rectangle1_widths[2476]), .RECT1_HEIGHT(rectangle1_heights[2476]), .RECT1_WEIGHT(rectangle1_weights[2476]), .RECT2_X(rectangle2_xs[2476]), .RECT2_Y(rectangle2_ys[2476]), .RECT2_WIDTH(rectangle2_widths[2476]), .RECT2_HEIGHT(rectangle2_heights[2476]), .RECT2_WEIGHT(rectangle2_weights[2476]), .RECT3_X(rectangle3_xs[2476]), .RECT3_Y(rectangle3_ys[2476]), .RECT3_WIDTH(rectangle3_widths[2476]), .RECT3_HEIGHT(rectangle3_heights[2476]), .RECT3_WEIGHT(rectangle3_weights[2476]), .FEAT_THRES(feature_thresholds[2476]), .FEAT_ABOVE(feature_aboves[2476]), .FEAT_BELOW(feature_belows[2476])) ac2476(.scan_win(scan_win2476), .scan_win_std_dev(scan_win_std_dev[2476]), .feature_accum(feature_accums[2476]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2477]), .RECT1_Y(rectangle1_ys[2477]), .RECT1_WIDTH(rectangle1_widths[2477]), .RECT1_HEIGHT(rectangle1_heights[2477]), .RECT1_WEIGHT(rectangle1_weights[2477]), .RECT2_X(rectangle2_xs[2477]), .RECT2_Y(rectangle2_ys[2477]), .RECT2_WIDTH(rectangle2_widths[2477]), .RECT2_HEIGHT(rectangle2_heights[2477]), .RECT2_WEIGHT(rectangle2_weights[2477]), .RECT3_X(rectangle3_xs[2477]), .RECT3_Y(rectangle3_ys[2477]), .RECT3_WIDTH(rectangle3_widths[2477]), .RECT3_HEIGHT(rectangle3_heights[2477]), .RECT3_WEIGHT(rectangle3_weights[2477]), .FEAT_THRES(feature_thresholds[2477]), .FEAT_ABOVE(feature_aboves[2477]), .FEAT_BELOW(feature_belows[2477])) ac2477(.scan_win(scan_win2477), .scan_win_std_dev(scan_win_std_dev[2477]), .feature_accum(feature_accums[2477]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2478]), .RECT1_Y(rectangle1_ys[2478]), .RECT1_WIDTH(rectangle1_widths[2478]), .RECT1_HEIGHT(rectangle1_heights[2478]), .RECT1_WEIGHT(rectangle1_weights[2478]), .RECT2_X(rectangle2_xs[2478]), .RECT2_Y(rectangle2_ys[2478]), .RECT2_WIDTH(rectangle2_widths[2478]), .RECT2_HEIGHT(rectangle2_heights[2478]), .RECT2_WEIGHT(rectangle2_weights[2478]), .RECT3_X(rectangle3_xs[2478]), .RECT3_Y(rectangle3_ys[2478]), .RECT3_WIDTH(rectangle3_widths[2478]), .RECT3_HEIGHT(rectangle3_heights[2478]), .RECT3_WEIGHT(rectangle3_weights[2478]), .FEAT_THRES(feature_thresholds[2478]), .FEAT_ABOVE(feature_aboves[2478]), .FEAT_BELOW(feature_belows[2478])) ac2478(.scan_win(scan_win2478), .scan_win_std_dev(scan_win_std_dev[2478]), .feature_accum(feature_accums[2478]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2479]), .RECT1_Y(rectangle1_ys[2479]), .RECT1_WIDTH(rectangle1_widths[2479]), .RECT1_HEIGHT(rectangle1_heights[2479]), .RECT1_WEIGHT(rectangle1_weights[2479]), .RECT2_X(rectangle2_xs[2479]), .RECT2_Y(rectangle2_ys[2479]), .RECT2_WIDTH(rectangle2_widths[2479]), .RECT2_HEIGHT(rectangle2_heights[2479]), .RECT2_WEIGHT(rectangle2_weights[2479]), .RECT3_X(rectangle3_xs[2479]), .RECT3_Y(rectangle3_ys[2479]), .RECT3_WIDTH(rectangle3_widths[2479]), .RECT3_HEIGHT(rectangle3_heights[2479]), .RECT3_WEIGHT(rectangle3_weights[2479]), .FEAT_THRES(feature_thresholds[2479]), .FEAT_ABOVE(feature_aboves[2479]), .FEAT_BELOW(feature_belows[2479])) ac2479(.scan_win(scan_win2479), .scan_win_std_dev(scan_win_std_dev[2479]), .feature_accum(feature_accums[2479]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2480]), .RECT1_Y(rectangle1_ys[2480]), .RECT1_WIDTH(rectangle1_widths[2480]), .RECT1_HEIGHT(rectangle1_heights[2480]), .RECT1_WEIGHT(rectangle1_weights[2480]), .RECT2_X(rectangle2_xs[2480]), .RECT2_Y(rectangle2_ys[2480]), .RECT2_WIDTH(rectangle2_widths[2480]), .RECT2_HEIGHT(rectangle2_heights[2480]), .RECT2_WEIGHT(rectangle2_weights[2480]), .RECT3_X(rectangle3_xs[2480]), .RECT3_Y(rectangle3_ys[2480]), .RECT3_WIDTH(rectangle3_widths[2480]), .RECT3_HEIGHT(rectangle3_heights[2480]), .RECT3_WEIGHT(rectangle3_weights[2480]), .FEAT_THRES(feature_thresholds[2480]), .FEAT_ABOVE(feature_aboves[2480]), .FEAT_BELOW(feature_belows[2480])) ac2480(.scan_win(scan_win2480), .scan_win_std_dev(scan_win_std_dev[2480]), .feature_accum(feature_accums[2480]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2481]), .RECT1_Y(rectangle1_ys[2481]), .RECT1_WIDTH(rectangle1_widths[2481]), .RECT1_HEIGHT(rectangle1_heights[2481]), .RECT1_WEIGHT(rectangle1_weights[2481]), .RECT2_X(rectangle2_xs[2481]), .RECT2_Y(rectangle2_ys[2481]), .RECT2_WIDTH(rectangle2_widths[2481]), .RECT2_HEIGHT(rectangle2_heights[2481]), .RECT2_WEIGHT(rectangle2_weights[2481]), .RECT3_X(rectangle3_xs[2481]), .RECT3_Y(rectangle3_ys[2481]), .RECT3_WIDTH(rectangle3_widths[2481]), .RECT3_HEIGHT(rectangle3_heights[2481]), .RECT3_WEIGHT(rectangle3_weights[2481]), .FEAT_THRES(feature_thresholds[2481]), .FEAT_ABOVE(feature_aboves[2481]), .FEAT_BELOW(feature_belows[2481])) ac2481(.scan_win(scan_win2481), .scan_win_std_dev(scan_win_std_dev[2481]), .feature_accum(feature_accums[2481]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2482]), .RECT1_Y(rectangle1_ys[2482]), .RECT1_WIDTH(rectangle1_widths[2482]), .RECT1_HEIGHT(rectangle1_heights[2482]), .RECT1_WEIGHT(rectangle1_weights[2482]), .RECT2_X(rectangle2_xs[2482]), .RECT2_Y(rectangle2_ys[2482]), .RECT2_WIDTH(rectangle2_widths[2482]), .RECT2_HEIGHT(rectangle2_heights[2482]), .RECT2_WEIGHT(rectangle2_weights[2482]), .RECT3_X(rectangle3_xs[2482]), .RECT3_Y(rectangle3_ys[2482]), .RECT3_WIDTH(rectangle3_widths[2482]), .RECT3_HEIGHT(rectangle3_heights[2482]), .RECT3_WEIGHT(rectangle3_weights[2482]), .FEAT_THRES(feature_thresholds[2482]), .FEAT_ABOVE(feature_aboves[2482]), .FEAT_BELOW(feature_belows[2482])) ac2482(.scan_win(scan_win2482), .scan_win_std_dev(scan_win_std_dev[2482]), .feature_accum(feature_accums[2482]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2483]), .RECT1_Y(rectangle1_ys[2483]), .RECT1_WIDTH(rectangle1_widths[2483]), .RECT1_HEIGHT(rectangle1_heights[2483]), .RECT1_WEIGHT(rectangle1_weights[2483]), .RECT2_X(rectangle2_xs[2483]), .RECT2_Y(rectangle2_ys[2483]), .RECT2_WIDTH(rectangle2_widths[2483]), .RECT2_HEIGHT(rectangle2_heights[2483]), .RECT2_WEIGHT(rectangle2_weights[2483]), .RECT3_X(rectangle3_xs[2483]), .RECT3_Y(rectangle3_ys[2483]), .RECT3_WIDTH(rectangle3_widths[2483]), .RECT3_HEIGHT(rectangle3_heights[2483]), .RECT3_WEIGHT(rectangle3_weights[2483]), .FEAT_THRES(feature_thresholds[2483]), .FEAT_ABOVE(feature_aboves[2483]), .FEAT_BELOW(feature_belows[2483])) ac2483(.scan_win(scan_win2483), .scan_win_std_dev(scan_win_std_dev[2483]), .feature_accum(feature_accums[2483]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2484]), .RECT1_Y(rectangle1_ys[2484]), .RECT1_WIDTH(rectangle1_widths[2484]), .RECT1_HEIGHT(rectangle1_heights[2484]), .RECT1_WEIGHT(rectangle1_weights[2484]), .RECT2_X(rectangle2_xs[2484]), .RECT2_Y(rectangle2_ys[2484]), .RECT2_WIDTH(rectangle2_widths[2484]), .RECT2_HEIGHT(rectangle2_heights[2484]), .RECT2_WEIGHT(rectangle2_weights[2484]), .RECT3_X(rectangle3_xs[2484]), .RECT3_Y(rectangle3_ys[2484]), .RECT3_WIDTH(rectangle3_widths[2484]), .RECT3_HEIGHT(rectangle3_heights[2484]), .RECT3_WEIGHT(rectangle3_weights[2484]), .FEAT_THRES(feature_thresholds[2484]), .FEAT_ABOVE(feature_aboves[2484]), .FEAT_BELOW(feature_belows[2484])) ac2484(.scan_win(scan_win2484), .scan_win_std_dev(scan_win_std_dev[2484]), .feature_accum(feature_accums[2484]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2485]), .RECT1_Y(rectangle1_ys[2485]), .RECT1_WIDTH(rectangle1_widths[2485]), .RECT1_HEIGHT(rectangle1_heights[2485]), .RECT1_WEIGHT(rectangle1_weights[2485]), .RECT2_X(rectangle2_xs[2485]), .RECT2_Y(rectangle2_ys[2485]), .RECT2_WIDTH(rectangle2_widths[2485]), .RECT2_HEIGHT(rectangle2_heights[2485]), .RECT2_WEIGHT(rectangle2_weights[2485]), .RECT3_X(rectangle3_xs[2485]), .RECT3_Y(rectangle3_ys[2485]), .RECT3_WIDTH(rectangle3_widths[2485]), .RECT3_HEIGHT(rectangle3_heights[2485]), .RECT3_WEIGHT(rectangle3_weights[2485]), .FEAT_THRES(feature_thresholds[2485]), .FEAT_ABOVE(feature_aboves[2485]), .FEAT_BELOW(feature_belows[2485])) ac2485(.scan_win(scan_win2485), .scan_win_std_dev(scan_win_std_dev[2485]), .feature_accum(feature_accums[2485]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2486]), .RECT1_Y(rectangle1_ys[2486]), .RECT1_WIDTH(rectangle1_widths[2486]), .RECT1_HEIGHT(rectangle1_heights[2486]), .RECT1_WEIGHT(rectangle1_weights[2486]), .RECT2_X(rectangle2_xs[2486]), .RECT2_Y(rectangle2_ys[2486]), .RECT2_WIDTH(rectangle2_widths[2486]), .RECT2_HEIGHT(rectangle2_heights[2486]), .RECT2_WEIGHT(rectangle2_weights[2486]), .RECT3_X(rectangle3_xs[2486]), .RECT3_Y(rectangle3_ys[2486]), .RECT3_WIDTH(rectangle3_widths[2486]), .RECT3_HEIGHT(rectangle3_heights[2486]), .RECT3_WEIGHT(rectangle3_weights[2486]), .FEAT_THRES(feature_thresholds[2486]), .FEAT_ABOVE(feature_aboves[2486]), .FEAT_BELOW(feature_belows[2486])) ac2486(.scan_win(scan_win2486), .scan_win_std_dev(scan_win_std_dev[2486]), .feature_accum(feature_accums[2486]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2487]), .RECT1_Y(rectangle1_ys[2487]), .RECT1_WIDTH(rectangle1_widths[2487]), .RECT1_HEIGHT(rectangle1_heights[2487]), .RECT1_WEIGHT(rectangle1_weights[2487]), .RECT2_X(rectangle2_xs[2487]), .RECT2_Y(rectangle2_ys[2487]), .RECT2_WIDTH(rectangle2_widths[2487]), .RECT2_HEIGHT(rectangle2_heights[2487]), .RECT2_WEIGHT(rectangle2_weights[2487]), .RECT3_X(rectangle3_xs[2487]), .RECT3_Y(rectangle3_ys[2487]), .RECT3_WIDTH(rectangle3_widths[2487]), .RECT3_HEIGHT(rectangle3_heights[2487]), .RECT3_WEIGHT(rectangle3_weights[2487]), .FEAT_THRES(feature_thresholds[2487]), .FEAT_ABOVE(feature_aboves[2487]), .FEAT_BELOW(feature_belows[2487])) ac2487(.scan_win(scan_win2487), .scan_win_std_dev(scan_win_std_dev[2487]), .feature_accum(feature_accums[2487]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2488]), .RECT1_Y(rectangle1_ys[2488]), .RECT1_WIDTH(rectangle1_widths[2488]), .RECT1_HEIGHT(rectangle1_heights[2488]), .RECT1_WEIGHT(rectangle1_weights[2488]), .RECT2_X(rectangle2_xs[2488]), .RECT2_Y(rectangle2_ys[2488]), .RECT2_WIDTH(rectangle2_widths[2488]), .RECT2_HEIGHT(rectangle2_heights[2488]), .RECT2_WEIGHT(rectangle2_weights[2488]), .RECT3_X(rectangle3_xs[2488]), .RECT3_Y(rectangle3_ys[2488]), .RECT3_WIDTH(rectangle3_widths[2488]), .RECT3_HEIGHT(rectangle3_heights[2488]), .RECT3_WEIGHT(rectangle3_weights[2488]), .FEAT_THRES(feature_thresholds[2488]), .FEAT_ABOVE(feature_aboves[2488]), .FEAT_BELOW(feature_belows[2488])) ac2488(.scan_win(scan_win2488), .scan_win_std_dev(scan_win_std_dev[2488]), .feature_accum(feature_accums[2488]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2489]), .RECT1_Y(rectangle1_ys[2489]), .RECT1_WIDTH(rectangle1_widths[2489]), .RECT1_HEIGHT(rectangle1_heights[2489]), .RECT1_WEIGHT(rectangle1_weights[2489]), .RECT2_X(rectangle2_xs[2489]), .RECT2_Y(rectangle2_ys[2489]), .RECT2_WIDTH(rectangle2_widths[2489]), .RECT2_HEIGHT(rectangle2_heights[2489]), .RECT2_WEIGHT(rectangle2_weights[2489]), .RECT3_X(rectangle3_xs[2489]), .RECT3_Y(rectangle3_ys[2489]), .RECT3_WIDTH(rectangle3_widths[2489]), .RECT3_HEIGHT(rectangle3_heights[2489]), .RECT3_WEIGHT(rectangle3_weights[2489]), .FEAT_THRES(feature_thresholds[2489]), .FEAT_ABOVE(feature_aboves[2489]), .FEAT_BELOW(feature_belows[2489])) ac2489(.scan_win(scan_win2489), .scan_win_std_dev(scan_win_std_dev[2489]), .feature_accum(feature_accums[2489]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2490]), .RECT1_Y(rectangle1_ys[2490]), .RECT1_WIDTH(rectangle1_widths[2490]), .RECT1_HEIGHT(rectangle1_heights[2490]), .RECT1_WEIGHT(rectangle1_weights[2490]), .RECT2_X(rectangle2_xs[2490]), .RECT2_Y(rectangle2_ys[2490]), .RECT2_WIDTH(rectangle2_widths[2490]), .RECT2_HEIGHT(rectangle2_heights[2490]), .RECT2_WEIGHT(rectangle2_weights[2490]), .RECT3_X(rectangle3_xs[2490]), .RECT3_Y(rectangle3_ys[2490]), .RECT3_WIDTH(rectangle3_widths[2490]), .RECT3_HEIGHT(rectangle3_heights[2490]), .RECT3_WEIGHT(rectangle3_weights[2490]), .FEAT_THRES(feature_thresholds[2490]), .FEAT_ABOVE(feature_aboves[2490]), .FEAT_BELOW(feature_belows[2490])) ac2490(.scan_win(scan_win2490), .scan_win_std_dev(scan_win_std_dev[2490]), .feature_accum(feature_accums[2490]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2491]), .RECT1_Y(rectangle1_ys[2491]), .RECT1_WIDTH(rectangle1_widths[2491]), .RECT1_HEIGHT(rectangle1_heights[2491]), .RECT1_WEIGHT(rectangle1_weights[2491]), .RECT2_X(rectangle2_xs[2491]), .RECT2_Y(rectangle2_ys[2491]), .RECT2_WIDTH(rectangle2_widths[2491]), .RECT2_HEIGHT(rectangle2_heights[2491]), .RECT2_WEIGHT(rectangle2_weights[2491]), .RECT3_X(rectangle3_xs[2491]), .RECT3_Y(rectangle3_ys[2491]), .RECT3_WIDTH(rectangle3_widths[2491]), .RECT3_HEIGHT(rectangle3_heights[2491]), .RECT3_WEIGHT(rectangle3_weights[2491]), .FEAT_THRES(feature_thresholds[2491]), .FEAT_ABOVE(feature_aboves[2491]), .FEAT_BELOW(feature_belows[2491])) ac2491(.scan_win(scan_win2491), .scan_win_std_dev(scan_win_std_dev[2491]), .feature_accum(feature_accums[2491]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2492]), .RECT1_Y(rectangle1_ys[2492]), .RECT1_WIDTH(rectangle1_widths[2492]), .RECT1_HEIGHT(rectangle1_heights[2492]), .RECT1_WEIGHT(rectangle1_weights[2492]), .RECT2_X(rectangle2_xs[2492]), .RECT2_Y(rectangle2_ys[2492]), .RECT2_WIDTH(rectangle2_widths[2492]), .RECT2_HEIGHT(rectangle2_heights[2492]), .RECT2_WEIGHT(rectangle2_weights[2492]), .RECT3_X(rectangle3_xs[2492]), .RECT3_Y(rectangle3_ys[2492]), .RECT3_WIDTH(rectangle3_widths[2492]), .RECT3_HEIGHT(rectangle3_heights[2492]), .RECT3_WEIGHT(rectangle3_weights[2492]), .FEAT_THRES(feature_thresholds[2492]), .FEAT_ABOVE(feature_aboves[2492]), .FEAT_BELOW(feature_belows[2492])) ac2492(.scan_win(scan_win2492), .scan_win_std_dev(scan_win_std_dev[2492]), .feature_accum(feature_accums[2492]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2493]), .RECT1_Y(rectangle1_ys[2493]), .RECT1_WIDTH(rectangle1_widths[2493]), .RECT1_HEIGHT(rectangle1_heights[2493]), .RECT1_WEIGHT(rectangle1_weights[2493]), .RECT2_X(rectangle2_xs[2493]), .RECT2_Y(rectangle2_ys[2493]), .RECT2_WIDTH(rectangle2_widths[2493]), .RECT2_HEIGHT(rectangle2_heights[2493]), .RECT2_WEIGHT(rectangle2_weights[2493]), .RECT3_X(rectangle3_xs[2493]), .RECT3_Y(rectangle3_ys[2493]), .RECT3_WIDTH(rectangle3_widths[2493]), .RECT3_HEIGHT(rectangle3_heights[2493]), .RECT3_WEIGHT(rectangle3_weights[2493]), .FEAT_THRES(feature_thresholds[2493]), .FEAT_ABOVE(feature_aboves[2493]), .FEAT_BELOW(feature_belows[2493])) ac2493(.scan_win(scan_win2493), .scan_win_std_dev(scan_win_std_dev[2493]), .feature_accum(feature_accums[2493]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2494]), .RECT1_Y(rectangle1_ys[2494]), .RECT1_WIDTH(rectangle1_widths[2494]), .RECT1_HEIGHT(rectangle1_heights[2494]), .RECT1_WEIGHT(rectangle1_weights[2494]), .RECT2_X(rectangle2_xs[2494]), .RECT2_Y(rectangle2_ys[2494]), .RECT2_WIDTH(rectangle2_widths[2494]), .RECT2_HEIGHT(rectangle2_heights[2494]), .RECT2_WEIGHT(rectangle2_weights[2494]), .RECT3_X(rectangle3_xs[2494]), .RECT3_Y(rectangle3_ys[2494]), .RECT3_WIDTH(rectangle3_widths[2494]), .RECT3_HEIGHT(rectangle3_heights[2494]), .RECT3_WEIGHT(rectangle3_weights[2494]), .FEAT_THRES(feature_thresholds[2494]), .FEAT_ABOVE(feature_aboves[2494]), .FEAT_BELOW(feature_belows[2494])) ac2494(.scan_win(scan_win2494), .scan_win_std_dev(scan_win_std_dev[2494]), .feature_accum(feature_accums[2494]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2495]), .RECT1_Y(rectangle1_ys[2495]), .RECT1_WIDTH(rectangle1_widths[2495]), .RECT1_HEIGHT(rectangle1_heights[2495]), .RECT1_WEIGHT(rectangle1_weights[2495]), .RECT2_X(rectangle2_xs[2495]), .RECT2_Y(rectangle2_ys[2495]), .RECT2_WIDTH(rectangle2_widths[2495]), .RECT2_HEIGHT(rectangle2_heights[2495]), .RECT2_WEIGHT(rectangle2_weights[2495]), .RECT3_X(rectangle3_xs[2495]), .RECT3_Y(rectangle3_ys[2495]), .RECT3_WIDTH(rectangle3_widths[2495]), .RECT3_HEIGHT(rectangle3_heights[2495]), .RECT3_WEIGHT(rectangle3_weights[2495]), .FEAT_THRES(feature_thresholds[2495]), .FEAT_ABOVE(feature_aboves[2495]), .FEAT_BELOW(feature_belows[2495])) ac2495(.scan_win(scan_win2495), .scan_win_std_dev(scan_win_std_dev[2495]), .feature_accum(feature_accums[2495]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2496]), .RECT1_Y(rectangle1_ys[2496]), .RECT1_WIDTH(rectangle1_widths[2496]), .RECT1_HEIGHT(rectangle1_heights[2496]), .RECT1_WEIGHT(rectangle1_weights[2496]), .RECT2_X(rectangle2_xs[2496]), .RECT2_Y(rectangle2_ys[2496]), .RECT2_WIDTH(rectangle2_widths[2496]), .RECT2_HEIGHT(rectangle2_heights[2496]), .RECT2_WEIGHT(rectangle2_weights[2496]), .RECT3_X(rectangle3_xs[2496]), .RECT3_Y(rectangle3_ys[2496]), .RECT3_WIDTH(rectangle3_widths[2496]), .RECT3_HEIGHT(rectangle3_heights[2496]), .RECT3_WEIGHT(rectangle3_weights[2496]), .FEAT_THRES(feature_thresholds[2496]), .FEAT_ABOVE(feature_aboves[2496]), .FEAT_BELOW(feature_belows[2496])) ac2496(.scan_win(scan_win2496), .scan_win_std_dev(scan_win_std_dev[2496]), .feature_accum(feature_accums[2496]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2497]), .RECT1_Y(rectangle1_ys[2497]), .RECT1_WIDTH(rectangle1_widths[2497]), .RECT1_HEIGHT(rectangle1_heights[2497]), .RECT1_WEIGHT(rectangle1_weights[2497]), .RECT2_X(rectangle2_xs[2497]), .RECT2_Y(rectangle2_ys[2497]), .RECT2_WIDTH(rectangle2_widths[2497]), .RECT2_HEIGHT(rectangle2_heights[2497]), .RECT2_WEIGHT(rectangle2_weights[2497]), .RECT3_X(rectangle3_xs[2497]), .RECT3_Y(rectangle3_ys[2497]), .RECT3_WIDTH(rectangle3_widths[2497]), .RECT3_HEIGHT(rectangle3_heights[2497]), .RECT3_WEIGHT(rectangle3_weights[2497]), .FEAT_THRES(feature_thresholds[2497]), .FEAT_ABOVE(feature_aboves[2497]), .FEAT_BELOW(feature_belows[2497])) ac2497(.scan_win(scan_win2497), .scan_win_std_dev(scan_win_std_dev[2497]), .feature_accum(feature_accums[2497]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2498]), .RECT1_Y(rectangle1_ys[2498]), .RECT1_WIDTH(rectangle1_widths[2498]), .RECT1_HEIGHT(rectangle1_heights[2498]), .RECT1_WEIGHT(rectangle1_weights[2498]), .RECT2_X(rectangle2_xs[2498]), .RECT2_Y(rectangle2_ys[2498]), .RECT2_WIDTH(rectangle2_widths[2498]), .RECT2_HEIGHT(rectangle2_heights[2498]), .RECT2_WEIGHT(rectangle2_weights[2498]), .RECT3_X(rectangle3_xs[2498]), .RECT3_Y(rectangle3_ys[2498]), .RECT3_WIDTH(rectangle3_widths[2498]), .RECT3_HEIGHT(rectangle3_heights[2498]), .RECT3_WEIGHT(rectangle3_weights[2498]), .FEAT_THRES(feature_thresholds[2498]), .FEAT_ABOVE(feature_aboves[2498]), .FEAT_BELOW(feature_belows[2498])) ac2498(.scan_win(scan_win2498), .scan_win_std_dev(scan_win_std_dev[2498]), .feature_accum(feature_accums[2498]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2499]), .RECT1_Y(rectangle1_ys[2499]), .RECT1_WIDTH(rectangle1_widths[2499]), .RECT1_HEIGHT(rectangle1_heights[2499]), .RECT1_WEIGHT(rectangle1_weights[2499]), .RECT2_X(rectangle2_xs[2499]), .RECT2_Y(rectangle2_ys[2499]), .RECT2_WIDTH(rectangle2_widths[2499]), .RECT2_HEIGHT(rectangle2_heights[2499]), .RECT2_WEIGHT(rectangle2_weights[2499]), .RECT3_X(rectangle3_xs[2499]), .RECT3_Y(rectangle3_ys[2499]), .RECT3_WIDTH(rectangle3_widths[2499]), .RECT3_HEIGHT(rectangle3_heights[2499]), .RECT3_WEIGHT(rectangle3_weights[2499]), .FEAT_THRES(feature_thresholds[2499]), .FEAT_ABOVE(feature_aboves[2499]), .FEAT_BELOW(feature_belows[2499])) ac2499(.scan_win(scan_win2499), .scan_win_std_dev(scan_win_std_dev[2499]), .feature_accum(feature_accums[2499]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2500]), .RECT1_Y(rectangle1_ys[2500]), .RECT1_WIDTH(rectangle1_widths[2500]), .RECT1_HEIGHT(rectangle1_heights[2500]), .RECT1_WEIGHT(rectangle1_weights[2500]), .RECT2_X(rectangle2_xs[2500]), .RECT2_Y(rectangle2_ys[2500]), .RECT2_WIDTH(rectangle2_widths[2500]), .RECT2_HEIGHT(rectangle2_heights[2500]), .RECT2_WEIGHT(rectangle2_weights[2500]), .RECT3_X(rectangle3_xs[2500]), .RECT3_Y(rectangle3_ys[2500]), .RECT3_WIDTH(rectangle3_widths[2500]), .RECT3_HEIGHT(rectangle3_heights[2500]), .RECT3_WEIGHT(rectangle3_weights[2500]), .FEAT_THRES(feature_thresholds[2500]), .FEAT_ABOVE(feature_aboves[2500]), .FEAT_BELOW(feature_belows[2500])) ac2500(.scan_win(scan_win2500), .scan_win_std_dev(scan_win_std_dev[2500]), .feature_accum(feature_accums[2500]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2501]), .RECT1_Y(rectangle1_ys[2501]), .RECT1_WIDTH(rectangle1_widths[2501]), .RECT1_HEIGHT(rectangle1_heights[2501]), .RECT1_WEIGHT(rectangle1_weights[2501]), .RECT2_X(rectangle2_xs[2501]), .RECT2_Y(rectangle2_ys[2501]), .RECT2_WIDTH(rectangle2_widths[2501]), .RECT2_HEIGHT(rectangle2_heights[2501]), .RECT2_WEIGHT(rectangle2_weights[2501]), .RECT3_X(rectangle3_xs[2501]), .RECT3_Y(rectangle3_ys[2501]), .RECT3_WIDTH(rectangle3_widths[2501]), .RECT3_HEIGHT(rectangle3_heights[2501]), .RECT3_WEIGHT(rectangle3_weights[2501]), .FEAT_THRES(feature_thresholds[2501]), .FEAT_ABOVE(feature_aboves[2501]), .FEAT_BELOW(feature_belows[2501])) ac2501(.scan_win(scan_win2501), .scan_win_std_dev(scan_win_std_dev[2501]), .feature_accum(feature_accums[2501]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2502]), .RECT1_Y(rectangle1_ys[2502]), .RECT1_WIDTH(rectangle1_widths[2502]), .RECT1_HEIGHT(rectangle1_heights[2502]), .RECT1_WEIGHT(rectangle1_weights[2502]), .RECT2_X(rectangle2_xs[2502]), .RECT2_Y(rectangle2_ys[2502]), .RECT2_WIDTH(rectangle2_widths[2502]), .RECT2_HEIGHT(rectangle2_heights[2502]), .RECT2_WEIGHT(rectangle2_weights[2502]), .RECT3_X(rectangle3_xs[2502]), .RECT3_Y(rectangle3_ys[2502]), .RECT3_WIDTH(rectangle3_widths[2502]), .RECT3_HEIGHT(rectangle3_heights[2502]), .RECT3_WEIGHT(rectangle3_weights[2502]), .FEAT_THRES(feature_thresholds[2502]), .FEAT_ABOVE(feature_aboves[2502]), .FEAT_BELOW(feature_belows[2502])) ac2502(.scan_win(scan_win2502), .scan_win_std_dev(scan_win_std_dev[2502]), .feature_accum(feature_accums[2502]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2503]), .RECT1_Y(rectangle1_ys[2503]), .RECT1_WIDTH(rectangle1_widths[2503]), .RECT1_HEIGHT(rectangle1_heights[2503]), .RECT1_WEIGHT(rectangle1_weights[2503]), .RECT2_X(rectangle2_xs[2503]), .RECT2_Y(rectangle2_ys[2503]), .RECT2_WIDTH(rectangle2_widths[2503]), .RECT2_HEIGHT(rectangle2_heights[2503]), .RECT2_WEIGHT(rectangle2_weights[2503]), .RECT3_X(rectangle3_xs[2503]), .RECT3_Y(rectangle3_ys[2503]), .RECT3_WIDTH(rectangle3_widths[2503]), .RECT3_HEIGHT(rectangle3_heights[2503]), .RECT3_WEIGHT(rectangle3_weights[2503]), .FEAT_THRES(feature_thresholds[2503]), .FEAT_ABOVE(feature_aboves[2503]), .FEAT_BELOW(feature_belows[2503])) ac2503(.scan_win(scan_win2503), .scan_win_std_dev(scan_win_std_dev[2503]), .feature_accum(feature_accums[2503]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2504]), .RECT1_Y(rectangle1_ys[2504]), .RECT1_WIDTH(rectangle1_widths[2504]), .RECT1_HEIGHT(rectangle1_heights[2504]), .RECT1_WEIGHT(rectangle1_weights[2504]), .RECT2_X(rectangle2_xs[2504]), .RECT2_Y(rectangle2_ys[2504]), .RECT2_WIDTH(rectangle2_widths[2504]), .RECT2_HEIGHT(rectangle2_heights[2504]), .RECT2_WEIGHT(rectangle2_weights[2504]), .RECT3_X(rectangle3_xs[2504]), .RECT3_Y(rectangle3_ys[2504]), .RECT3_WIDTH(rectangle3_widths[2504]), .RECT3_HEIGHT(rectangle3_heights[2504]), .RECT3_WEIGHT(rectangle3_weights[2504]), .FEAT_THRES(feature_thresholds[2504]), .FEAT_ABOVE(feature_aboves[2504]), .FEAT_BELOW(feature_belows[2504])) ac2504(.scan_win(scan_win2504), .scan_win_std_dev(scan_win_std_dev[2504]), .feature_accum(feature_accums[2504]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2505]), .RECT1_Y(rectangle1_ys[2505]), .RECT1_WIDTH(rectangle1_widths[2505]), .RECT1_HEIGHT(rectangle1_heights[2505]), .RECT1_WEIGHT(rectangle1_weights[2505]), .RECT2_X(rectangle2_xs[2505]), .RECT2_Y(rectangle2_ys[2505]), .RECT2_WIDTH(rectangle2_widths[2505]), .RECT2_HEIGHT(rectangle2_heights[2505]), .RECT2_WEIGHT(rectangle2_weights[2505]), .RECT3_X(rectangle3_xs[2505]), .RECT3_Y(rectangle3_ys[2505]), .RECT3_WIDTH(rectangle3_widths[2505]), .RECT3_HEIGHT(rectangle3_heights[2505]), .RECT3_WEIGHT(rectangle3_weights[2505]), .FEAT_THRES(feature_thresholds[2505]), .FEAT_ABOVE(feature_aboves[2505]), .FEAT_BELOW(feature_belows[2505])) ac2505(.scan_win(scan_win2505), .scan_win_std_dev(scan_win_std_dev[2505]), .feature_accum(feature_accums[2505]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2506]), .RECT1_Y(rectangle1_ys[2506]), .RECT1_WIDTH(rectangle1_widths[2506]), .RECT1_HEIGHT(rectangle1_heights[2506]), .RECT1_WEIGHT(rectangle1_weights[2506]), .RECT2_X(rectangle2_xs[2506]), .RECT2_Y(rectangle2_ys[2506]), .RECT2_WIDTH(rectangle2_widths[2506]), .RECT2_HEIGHT(rectangle2_heights[2506]), .RECT2_WEIGHT(rectangle2_weights[2506]), .RECT3_X(rectangle3_xs[2506]), .RECT3_Y(rectangle3_ys[2506]), .RECT3_WIDTH(rectangle3_widths[2506]), .RECT3_HEIGHT(rectangle3_heights[2506]), .RECT3_WEIGHT(rectangle3_weights[2506]), .FEAT_THRES(feature_thresholds[2506]), .FEAT_ABOVE(feature_aboves[2506]), .FEAT_BELOW(feature_belows[2506])) ac2506(.scan_win(scan_win2506), .scan_win_std_dev(scan_win_std_dev[2506]), .feature_accum(feature_accums[2506]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2507]), .RECT1_Y(rectangle1_ys[2507]), .RECT1_WIDTH(rectangle1_widths[2507]), .RECT1_HEIGHT(rectangle1_heights[2507]), .RECT1_WEIGHT(rectangle1_weights[2507]), .RECT2_X(rectangle2_xs[2507]), .RECT2_Y(rectangle2_ys[2507]), .RECT2_WIDTH(rectangle2_widths[2507]), .RECT2_HEIGHT(rectangle2_heights[2507]), .RECT2_WEIGHT(rectangle2_weights[2507]), .RECT3_X(rectangle3_xs[2507]), .RECT3_Y(rectangle3_ys[2507]), .RECT3_WIDTH(rectangle3_widths[2507]), .RECT3_HEIGHT(rectangle3_heights[2507]), .RECT3_WEIGHT(rectangle3_weights[2507]), .FEAT_THRES(feature_thresholds[2507]), .FEAT_ABOVE(feature_aboves[2507]), .FEAT_BELOW(feature_belows[2507])) ac2507(.scan_win(scan_win2507), .scan_win_std_dev(scan_win_std_dev[2507]), .feature_accum(feature_accums[2507]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2508]), .RECT1_Y(rectangle1_ys[2508]), .RECT1_WIDTH(rectangle1_widths[2508]), .RECT1_HEIGHT(rectangle1_heights[2508]), .RECT1_WEIGHT(rectangle1_weights[2508]), .RECT2_X(rectangle2_xs[2508]), .RECT2_Y(rectangle2_ys[2508]), .RECT2_WIDTH(rectangle2_widths[2508]), .RECT2_HEIGHT(rectangle2_heights[2508]), .RECT2_WEIGHT(rectangle2_weights[2508]), .RECT3_X(rectangle3_xs[2508]), .RECT3_Y(rectangle3_ys[2508]), .RECT3_WIDTH(rectangle3_widths[2508]), .RECT3_HEIGHT(rectangle3_heights[2508]), .RECT3_WEIGHT(rectangle3_weights[2508]), .FEAT_THRES(feature_thresholds[2508]), .FEAT_ABOVE(feature_aboves[2508]), .FEAT_BELOW(feature_belows[2508])) ac2508(.scan_win(scan_win2508), .scan_win_std_dev(scan_win_std_dev[2508]), .feature_accum(feature_accums[2508]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2509]), .RECT1_Y(rectangle1_ys[2509]), .RECT1_WIDTH(rectangle1_widths[2509]), .RECT1_HEIGHT(rectangle1_heights[2509]), .RECT1_WEIGHT(rectangle1_weights[2509]), .RECT2_X(rectangle2_xs[2509]), .RECT2_Y(rectangle2_ys[2509]), .RECT2_WIDTH(rectangle2_widths[2509]), .RECT2_HEIGHT(rectangle2_heights[2509]), .RECT2_WEIGHT(rectangle2_weights[2509]), .RECT3_X(rectangle3_xs[2509]), .RECT3_Y(rectangle3_ys[2509]), .RECT3_WIDTH(rectangle3_widths[2509]), .RECT3_HEIGHT(rectangle3_heights[2509]), .RECT3_WEIGHT(rectangle3_weights[2509]), .FEAT_THRES(feature_thresholds[2509]), .FEAT_ABOVE(feature_aboves[2509]), .FEAT_BELOW(feature_belows[2509])) ac2509(.scan_win(scan_win2509), .scan_win_std_dev(scan_win_std_dev[2509]), .feature_accum(feature_accums[2509]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2510]), .RECT1_Y(rectangle1_ys[2510]), .RECT1_WIDTH(rectangle1_widths[2510]), .RECT1_HEIGHT(rectangle1_heights[2510]), .RECT1_WEIGHT(rectangle1_weights[2510]), .RECT2_X(rectangle2_xs[2510]), .RECT2_Y(rectangle2_ys[2510]), .RECT2_WIDTH(rectangle2_widths[2510]), .RECT2_HEIGHT(rectangle2_heights[2510]), .RECT2_WEIGHT(rectangle2_weights[2510]), .RECT3_X(rectangle3_xs[2510]), .RECT3_Y(rectangle3_ys[2510]), .RECT3_WIDTH(rectangle3_widths[2510]), .RECT3_HEIGHT(rectangle3_heights[2510]), .RECT3_WEIGHT(rectangle3_weights[2510]), .FEAT_THRES(feature_thresholds[2510]), .FEAT_ABOVE(feature_aboves[2510]), .FEAT_BELOW(feature_belows[2510])) ac2510(.scan_win(scan_win2510), .scan_win_std_dev(scan_win_std_dev[2510]), .feature_accum(feature_accums[2510]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2511]), .RECT1_Y(rectangle1_ys[2511]), .RECT1_WIDTH(rectangle1_widths[2511]), .RECT1_HEIGHT(rectangle1_heights[2511]), .RECT1_WEIGHT(rectangle1_weights[2511]), .RECT2_X(rectangle2_xs[2511]), .RECT2_Y(rectangle2_ys[2511]), .RECT2_WIDTH(rectangle2_widths[2511]), .RECT2_HEIGHT(rectangle2_heights[2511]), .RECT2_WEIGHT(rectangle2_weights[2511]), .RECT3_X(rectangle3_xs[2511]), .RECT3_Y(rectangle3_ys[2511]), .RECT3_WIDTH(rectangle3_widths[2511]), .RECT3_HEIGHT(rectangle3_heights[2511]), .RECT3_WEIGHT(rectangle3_weights[2511]), .FEAT_THRES(feature_thresholds[2511]), .FEAT_ABOVE(feature_aboves[2511]), .FEAT_BELOW(feature_belows[2511])) ac2511(.scan_win(scan_win2511), .scan_win_std_dev(scan_win_std_dev[2511]), .feature_accum(feature_accums[2511]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2512]), .RECT1_Y(rectangle1_ys[2512]), .RECT1_WIDTH(rectangle1_widths[2512]), .RECT1_HEIGHT(rectangle1_heights[2512]), .RECT1_WEIGHT(rectangle1_weights[2512]), .RECT2_X(rectangle2_xs[2512]), .RECT2_Y(rectangle2_ys[2512]), .RECT2_WIDTH(rectangle2_widths[2512]), .RECT2_HEIGHT(rectangle2_heights[2512]), .RECT2_WEIGHT(rectangle2_weights[2512]), .RECT3_X(rectangle3_xs[2512]), .RECT3_Y(rectangle3_ys[2512]), .RECT3_WIDTH(rectangle3_widths[2512]), .RECT3_HEIGHT(rectangle3_heights[2512]), .RECT3_WEIGHT(rectangle3_weights[2512]), .FEAT_THRES(feature_thresholds[2512]), .FEAT_ABOVE(feature_aboves[2512]), .FEAT_BELOW(feature_belows[2512])) ac2512(.scan_win(scan_win2512), .scan_win_std_dev(scan_win_std_dev[2512]), .feature_accum(feature_accums[2512]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2513]), .RECT1_Y(rectangle1_ys[2513]), .RECT1_WIDTH(rectangle1_widths[2513]), .RECT1_HEIGHT(rectangle1_heights[2513]), .RECT1_WEIGHT(rectangle1_weights[2513]), .RECT2_X(rectangle2_xs[2513]), .RECT2_Y(rectangle2_ys[2513]), .RECT2_WIDTH(rectangle2_widths[2513]), .RECT2_HEIGHT(rectangle2_heights[2513]), .RECT2_WEIGHT(rectangle2_weights[2513]), .RECT3_X(rectangle3_xs[2513]), .RECT3_Y(rectangle3_ys[2513]), .RECT3_WIDTH(rectangle3_widths[2513]), .RECT3_HEIGHT(rectangle3_heights[2513]), .RECT3_WEIGHT(rectangle3_weights[2513]), .FEAT_THRES(feature_thresholds[2513]), .FEAT_ABOVE(feature_aboves[2513]), .FEAT_BELOW(feature_belows[2513])) ac2513(.scan_win(scan_win2513), .scan_win_std_dev(scan_win_std_dev[2513]), .feature_accum(feature_accums[2513]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2514]), .RECT1_Y(rectangle1_ys[2514]), .RECT1_WIDTH(rectangle1_widths[2514]), .RECT1_HEIGHT(rectangle1_heights[2514]), .RECT1_WEIGHT(rectangle1_weights[2514]), .RECT2_X(rectangle2_xs[2514]), .RECT2_Y(rectangle2_ys[2514]), .RECT2_WIDTH(rectangle2_widths[2514]), .RECT2_HEIGHT(rectangle2_heights[2514]), .RECT2_WEIGHT(rectangle2_weights[2514]), .RECT3_X(rectangle3_xs[2514]), .RECT3_Y(rectangle3_ys[2514]), .RECT3_WIDTH(rectangle3_widths[2514]), .RECT3_HEIGHT(rectangle3_heights[2514]), .RECT3_WEIGHT(rectangle3_weights[2514]), .FEAT_THRES(feature_thresholds[2514]), .FEAT_ABOVE(feature_aboves[2514]), .FEAT_BELOW(feature_belows[2514])) ac2514(.scan_win(scan_win2514), .scan_win_std_dev(scan_win_std_dev[2514]), .feature_accum(feature_accums[2514]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2515]), .RECT1_Y(rectangle1_ys[2515]), .RECT1_WIDTH(rectangle1_widths[2515]), .RECT1_HEIGHT(rectangle1_heights[2515]), .RECT1_WEIGHT(rectangle1_weights[2515]), .RECT2_X(rectangle2_xs[2515]), .RECT2_Y(rectangle2_ys[2515]), .RECT2_WIDTH(rectangle2_widths[2515]), .RECT2_HEIGHT(rectangle2_heights[2515]), .RECT2_WEIGHT(rectangle2_weights[2515]), .RECT3_X(rectangle3_xs[2515]), .RECT3_Y(rectangle3_ys[2515]), .RECT3_WIDTH(rectangle3_widths[2515]), .RECT3_HEIGHT(rectangle3_heights[2515]), .RECT3_WEIGHT(rectangle3_weights[2515]), .FEAT_THRES(feature_thresholds[2515]), .FEAT_ABOVE(feature_aboves[2515]), .FEAT_BELOW(feature_belows[2515])) ac2515(.scan_win(scan_win2515), .scan_win_std_dev(scan_win_std_dev[2515]), .feature_accum(feature_accums[2515]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2516]), .RECT1_Y(rectangle1_ys[2516]), .RECT1_WIDTH(rectangle1_widths[2516]), .RECT1_HEIGHT(rectangle1_heights[2516]), .RECT1_WEIGHT(rectangle1_weights[2516]), .RECT2_X(rectangle2_xs[2516]), .RECT2_Y(rectangle2_ys[2516]), .RECT2_WIDTH(rectangle2_widths[2516]), .RECT2_HEIGHT(rectangle2_heights[2516]), .RECT2_WEIGHT(rectangle2_weights[2516]), .RECT3_X(rectangle3_xs[2516]), .RECT3_Y(rectangle3_ys[2516]), .RECT3_WIDTH(rectangle3_widths[2516]), .RECT3_HEIGHT(rectangle3_heights[2516]), .RECT3_WEIGHT(rectangle3_weights[2516]), .FEAT_THRES(feature_thresholds[2516]), .FEAT_ABOVE(feature_aboves[2516]), .FEAT_BELOW(feature_belows[2516])) ac2516(.scan_win(scan_win2516), .scan_win_std_dev(scan_win_std_dev[2516]), .feature_accum(feature_accums[2516]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2517]), .RECT1_Y(rectangle1_ys[2517]), .RECT1_WIDTH(rectangle1_widths[2517]), .RECT1_HEIGHT(rectangle1_heights[2517]), .RECT1_WEIGHT(rectangle1_weights[2517]), .RECT2_X(rectangle2_xs[2517]), .RECT2_Y(rectangle2_ys[2517]), .RECT2_WIDTH(rectangle2_widths[2517]), .RECT2_HEIGHT(rectangle2_heights[2517]), .RECT2_WEIGHT(rectangle2_weights[2517]), .RECT3_X(rectangle3_xs[2517]), .RECT3_Y(rectangle3_ys[2517]), .RECT3_WIDTH(rectangle3_widths[2517]), .RECT3_HEIGHT(rectangle3_heights[2517]), .RECT3_WEIGHT(rectangle3_weights[2517]), .FEAT_THRES(feature_thresholds[2517]), .FEAT_ABOVE(feature_aboves[2517]), .FEAT_BELOW(feature_belows[2517])) ac2517(.scan_win(scan_win2517), .scan_win_std_dev(scan_win_std_dev[2517]), .feature_accum(feature_accums[2517]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2518]), .RECT1_Y(rectangle1_ys[2518]), .RECT1_WIDTH(rectangle1_widths[2518]), .RECT1_HEIGHT(rectangle1_heights[2518]), .RECT1_WEIGHT(rectangle1_weights[2518]), .RECT2_X(rectangle2_xs[2518]), .RECT2_Y(rectangle2_ys[2518]), .RECT2_WIDTH(rectangle2_widths[2518]), .RECT2_HEIGHT(rectangle2_heights[2518]), .RECT2_WEIGHT(rectangle2_weights[2518]), .RECT3_X(rectangle3_xs[2518]), .RECT3_Y(rectangle3_ys[2518]), .RECT3_WIDTH(rectangle3_widths[2518]), .RECT3_HEIGHT(rectangle3_heights[2518]), .RECT3_WEIGHT(rectangle3_weights[2518]), .FEAT_THRES(feature_thresholds[2518]), .FEAT_ABOVE(feature_aboves[2518]), .FEAT_BELOW(feature_belows[2518])) ac2518(.scan_win(scan_win2518), .scan_win_std_dev(scan_win_std_dev[2518]), .feature_accum(feature_accums[2518]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2519]), .RECT1_Y(rectangle1_ys[2519]), .RECT1_WIDTH(rectangle1_widths[2519]), .RECT1_HEIGHT(rectangle1_heights[2519]), .RECT1_WEIGHT(rectangle1_weights[2519]), .RECT2_X(rectangle2_xs[2519]), .RECT2_Y(rectangle2_ys[2519]), .RECT2_WIDTH(rectangle2_widths[2519]), .RECT2_HEIGHT(rectangle2_heights[2519]), .RECT2_WEIGHT(rectangle2_weights[2519]), .RECT3_X(rectangle3_xs[2519]), .RECT3_Y(rectangle3_ys[2519]), .RECT3_WIDTH(rectangle3_widths[2519]), .RECT3_HEIGHT(rectangle3_heights[2519]), .RECT3_WEIGHT(rectangle3_weights[2519]), .FEAT_THRES(feature_thresholds[2519]), .FEAT_ABOVE(feature_aboves[2519]), .FEAT_BELOW(feature_belows[2519])) ac2519(.scan_win(scan_win2519), .scan_win_std_dev(scan_win_std_dev[2519]), .feature_accum(feature_accums[2519]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2520]), .RECT1_Y(rectangle1_ys[2520]), .RECT1_WIDTH(rectangle1_widths[2520]), .RECT1_HEIGHT(rectangle1_heights[2520]), .RECT1_WEIGHT(rectangle1_weights[2520]), .RECT2_X(rectangle2_xs[2520]), .RECT2_Y(rectangle2_ys[2520]), .RECT2_WIDTH(rectangle2_widths[2520]), .RECT2_HEIGHT(rectangle2_heights[2520]), .RECT2_WEIGHT(rectangle2_weights[2520]), .RECT3_X(rectangle3_xs[2520]), .RECT3_Y(rectangle3_ys[2520]), .RECT3_WIDTH(rectangle3_widths[2520]), .RECT3_HEIGHT(rectangle3_heights[2520]), .RECT3_WEIGHT(rectangle3_weights[2520]), .FEAT_THRES(feature_thresholds[2520]), .FEAT_ABOVE(feature_aboves[2520]), .FEAT_BELOW(feature_belows[2520])) ac2520(.scan_win(scan_win2520), .scan_win_std_dev(scan_win_std_dev[2520]), .feature_accum(feature_accums[2520]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2521]), .RECT1_Y(rectangle1_ys[2521]), .RECT1_WIDTH(rectangle1_widths[2521]), .RECT1_HEIGHT(rectangle1_heights[2521]), .RECT1_WEIGHT(rectangle1_weights[2521]), .RECT2_X(rectangle2_xs[2521]), .RECT2_Y(rectangle2_ys[2521]), .RECT2_WIDTH(rectangle2_widths[2521]), .RECT2_HEIGHT(rectangle2_heights[2521]), .RECT2_WEIGHT(rectangle2_weights[2521]), .RECT3_X(rectangle3_xs[2521]), .RECT3_Y(rectangle3_ys[2521]), .RECT3_WIDTH(rectangle3_widths[2521]), .RECT3_HEIGHT(rectangle3_heights[2521]), .RECT3_WEIGHT(rectangle3_weights[2521]), .FEAT_THRES(feature_thresholds[2521]), .FEAT_ABOVE(feature_aboves[2521]), .FEAT_BELOW(feature_belows[2521])) ac2521(.scan_win(scan_win2521), .scan_win_std_dev(scan_win_std_dev[2521]), .feature_accum(feature_accums[2521]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2522]), .RECT1_Y(rectangle1_ys[2522]), .RECT1_WIDTH(rectangle1_widths[2522]), .RECT1_HEIGHT(rectangle1_heights[2522]), .RECT1_WEIGHT(rectangle1_weights[2522]), .RECT2_X(rectangle2_xs[2522]), .RECT2_Y(rectangle2_ys[2522]), .RECT2_WIDTH(rectangle2_widths[2522]), .RECT2_HEIGHT(rectangle2_heights[2522]), .RECT2_WEIGHT(rectangle2_weights[2522]), .RECT3_X(rectangle3_xs[2522]), .RECT3_Y(rectangle3_ys[2522]), .RECT3_WIDTH(rectangle3_widths[2522]), .RECT3_HEIGHT(rectangle3_heights[2522]), .RECT3_WEIGHT(rectangle3_weights[2522]), .FEAT_THRES(feature_thresholds[2522]), .FEAT_ABOVE(feature_aboves[2522]), .FEAT_BELOW(feature_belows[2522])) ac2522(.scan_win(scan_win2522), .scan_win_std_dev(scan_win_std_dev[2522]), .feature_accum(feature_accums[2522]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2523]), .RECT1_Y(rectangle1_ys[2523]), .RECT1_WIDTH(rectangle1_widths[2523]), .RECT1_HEIGHT(rectangle1_heights[2523]), .RECT1_WEIGHT(rectangle1_weights[2523]), .RECT2_X(rectangle2_xs[2523]), .RECT2_Y(rectangle2_ys[2523]), .RECT2_WIDTH(rectangle2_widths[2523]), .RECT2_HEIGHT(rectangle2_heights[2523]), .RECT2_WEIGHT(rectangle2_weights[2523]), .RECT3_X(rectangle3_xs[2523]), .RECT3_Y(rectangle3_ys[2523]), .RECT3_WIDTH(rectangle3_widths[2523]), .RECT3_HEIGHT(rectangle3_heights[2523]), .RECT3_WEIGHT(rectangle3_weights[2523]), .FEAT_THRES(feature_thresholds[2523]), .FEAT_ABOVE(feature_aboves[2523]), .FEAT_BELOW(feature_belows[2523])) ac2523(.scan_win(scan_win2523), .scan_win_std_dev(scan_win_std_dev[2523]), .feature_accum(feature_accums[2523]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2524]), .RECT1_Y(rectangle1_ys[2524]), .RECT1_WIDTH(rectangle1_widths[2524]), .RECT1_HEIGHT(rectangle1_heights[2524]), .RECT1_WEIGHT(rectangle1_weights[2524]), .RECT2_X(rectangle2_xs[2524]), .RECT2_Y(rectangle2_ys[2524]), .RECT2_WIDTH(rectangle2_widths[2524]), .RECT2_HEIGHT(rectangle2_heights[2524]), .RECT2_WEIGHT(rectangle2_weights[2524]), .RECT3_X(rectangle3_xs[2524]), .RECT3_Y(rectangle3_ys[2524]), .RECT3_WIDTH(rectangle3_widths[2524]), .RECT3_HEIGHT(rectangle3_heights[2524]), .RECT3_WEIGHT(rectangle3_weights[2524]), .FEAT_THRES(feature_thresholds[2524]), .FEAT_ABOVE(feature_aboves[2524]), .FEAT_BELOW(feature_belows[2524])) ac2524(.scan_win(scan_win2524), .scan_win_std_dev(scan_win_std_dev[2524]), .feature_accum(feature_accums[2524]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2525]), .RECT1_Y(rectangle1_ys[2525]), .RECT1_WIDTH(rectangle1_widths[2525]), .RECT1_HEIGHT(rectangle1_heights[2525]), .RECT1_WEIGHT(rectangle1_weights[2525]), .RECT2_X(rectangle2_xs[2525]), .RECT2_Y(rectangle2_ys[2525]), .RECT2_WIDTH(rectangle2_widths[2525]), .RECT2_HEIGHT(rectangle2_heights[2525]), .RECT2_WEIGHT(rectangle2_weights[2525]), .RECT3_X(rectangle3_xs[2525]), .RECT3_Y(rectangle3_ys[2525]), .RECT3_WIDTH(rectangle3_widths[2525]), .RECT3_HEIGHT(rectangle3_heights[2525]), .RECT3_WEIGHT(rectangle3_weights[2525]), .FEAT_THRES(feature_thresholds[2525]), .FEAT_ABOVE(feature_aboves[2525]), .FEAT_BELOW(feature_belows[2525])) ac2525(.scan_win(scan_win2525), .scan_win_std_dev(scan_win_std_dev[2525]), .feature_accum(feature_accums[2525]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2526]), .RECT1_Y(rectangle1_ys[2526]), .RECT1_WIDTH(rectangle1_widths[2526]), .RECT1_HEIGHT(rectangle1_heights[2526]), .RECT1_WEIGHT(rectangle1_weights[2526]), .RECT2_X(rectangle2_xs[2526]), .RECT2_Y(rectangle2_ys[2526]), .RECT2_WIDTH(rectangle2_widths[2526]), .RECT2_HEIGHT(rectangle2_heights[2526]), .RECT2_WEIGHT(rectangle2_weights[2526]), .RECT3_X(rectangle3_xs[2526]), .RECT3_Y(rectangle3_ys[2526]), .RECT3_WIDTH(rectangle3_widths[2526]), .RECT3_HEIGHT(rectangle3_heights[2526]), .RECT3_WEIGHT(rectangle3_weights[2526]), .FEAT_THRES(feature_thresholds[2526]), .FEAT_ABOVE(feature_aboves[2526]), .FEAT_BELOW(feature_belows[2526])) ac2526(.scan_win(scan_win2526), .scan_win_std_dev(scan_win_std_dev[2526]), .feature_accum(feature_accums[2526]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2527]), .RECT1_Y(rectangle1_ys[2527]), .RECT1_WIDTH(rectangle1_widths[2527]), .RECT1_HEIGHT(rectangle1_heights[2527]), .RECT1_WEIGHT(rectangle1_weights[2527]), .RECT2_X(rectangle2_xs[2527]), .RECT2_Y(rectangle2_ys[2527]), .RECT2_WIDTH(rectangle2_widths[2527]), .RECT2_HEIGHT(rectangle2_heights[2527]), .RECT2_WEIGHT(rectangle2_weights[2527]), .RECT3_X(rectangle3_xs[2527]), .RECT3_Y(rectangle3_ys[2527]), .RECT3_WIDTH(rectangle3_widths[2527]), .RECT3_HEIGHT(rectangle3_heights[2527]), .RECT3_WEIGHT(rectangle3_weights[2527]), .FEAT_THRES(feature_thresholds[2527]), .FEAT_ABOVE(feature_aboves[2527]), .FEAT_BELOW(feature_belows[2527])) ac2527(.scan_win(scan_win2527), .scan_win_std_dev(scan_win_std_dev[2527]), .feature_accum(feature_accums[2527]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2528]), .RECT1_Y(rectangle1_ys[2528]), .RECT1_WIDTH(rectangle1_widths[2528]), .RECT1_HEIGHT(rectangle1_heights[2528]), .RECT1_WEIGHT(rectangle1_weights[2528]), .RECT2_X(rectangle2_xs[2528]), .RECT2_Y(rectangle2_ys[2528]), .RECT2_WIDTH(rectangle2_widths[2528]), .RECT2_HEIGHT(rectangle2_heights[2528]), .RECT2_WEIGHT(rectangle2_weights[2528]), .RECT3_X(rectangle3_xs[2528]), .RECT3_Y(rectangle3_ys[2528]), .RECT3_WIDTH(rectangle3_widths[2528]), .RECT3_HEIGHT(rectangle3_heights[2528]), .RECT3_WEIGHT(rectangle3_weights[2528]), .FEAT_THRES(feature_thresholds[2528]), .FEAT_ABOVE(feature_aboves[2528]), .FEAT_BELOW(feature_belows[2528])) ac2528(.scan_win(scan_win2528), .scan_win_std_dev(scan_win_std_dev[2528]), .feature_accum(feature_accums[2528]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2529]), .RECT1_Y(rectangle1_ys[2529]), .RECT1_WIDTH(rectangle1_widths[2529]), .RECT1_HEIGHT(rectangle1_heights[2529]), .RECT1_WEIGHT(rectangle1_weights[2529]), .RECT2_X(rectangle2_xs[2529]), .RECT2_Y(rectangle2_ys[2529]), .RECT2_WIDTH(rectangle2_widths[2529]), .RECT2_HEIGHT(rectangle2_heights[2529]), .RECT2_WEIGHT(rectangle2_weights[2529]), .RECT3_X(rectangle3_xs[2529]), .RECT3_Y(rectangle3_ys[2529]), .RECT3_WIDTH(rectangle3_widths[2529]), .RECT3_HEIGHT(rectangle3_heights[2529]), .RECT3_WEIGHT(rectangle3_weights[2529]), .FEAT_THRES(feature_thresholds[2529]), .FEAT_ABOVE(feature_aboves[2529]), .FEAT_BELOW(feature_belows[2529])) ac2529(.scan_win(scan_win2529), .scan_win_std_dev(scan_win_std_dev[2529]), .feature_accum(feature_accums[2529]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2530]), .RECT1_Y(rectangle1_ys[2530]), .RECT1_WIDTH(rectangle1_widths[2530]), .RECT1_HEIGHT(rectangle1_heights[2530]), .RECT1_WEIGHT(rectangle1_weights[2530]), .RECT2_X(rectangle2_xs[2530]), .RECT2_Y(rectangle2_ys[2530]), .RECT2_WIDTH(rectangle2_widths[2530]), .RECT2_HEIGHT(rectangle2_heights[2530]), .RECT2_WEIGHT(rectangle2_weights[2530]), .RECT3_X(rectangle3_xs[2530]), .RECT3_Y(rectangle3_ys[2530]), .RECT3_WIDTH(rectangle3_widths[2530]), .RECT3_HEIGHT(rectangle3_heights[2530]), .RECT3_WEIGHT(rectangle3_weights[2530]), .FEAT_THRES(feature_thresholds[2530]), .FEAT_ABOVE(feature_aboves[2530]), .FEAT_BELOW(feature_belows[2530])) ac2530(.scan_win(scan_win2530), .scan_win_std_dev(scan_win_std_dev[2530]), .feature_accum(feature_accums[2530]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2531]), .RECT1_Y(rectangle1_ys[2531]), .RECT1_WIDTH(rectangle1_widths[2531]), .RECT1_HEIGHT(rectangle1_heights[2531]), .RECT1_WEIGHT(rectangle1_weights[2531]), .RECT2_X(rectangle2_xs[2531]), .RECT2_Y(rectangle2_ys[2531]), .RECT2_WIDTH(rectangle2_widths[2531]), .RECT2_HEIGHT(rectangle2_heights[2531]), .RECT2_WEIGHT(rectangle2_weights[2531]), .RECT3_X(rectangle3_xs[2531]), .RECT3_Y(rectangle3_ys[2531]), .RECT3_WIDTH(rectangle3_widths[2531]), .RECT3_HEIGHT(rectangle3_heights[2531]), .RECT3_WEIGHT(rectangle3_weights[2531]), .FEAT_THRES(feature_thresholds[2531]), .FEAT_ABOVE(feature_aboves[2531]), .FEAT_BELOW(feature_belows[2531])) ac2531(.scan_win(scan_win2531), .scan_win_std_dev(scan_win_std_dev[2531]), .feature_accum(feature_accums[2531]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2532]), .RECT1_Y(rectangle1_ys[2532]), .RECT1_WIDTH(rectangle1_widths[2532]), .RECT1_HEIGHT(rectangle1_heights[2532]), .RECT1_WEIGHT(rectangle1_weights[2532]), .RECT2_X(rectangle2_xs[2532]), .RECT2_Y(rectangle2_ys[2532]), .RECT2_WIDTH(rectangle2_widths[2532]), .RECT2_HEIGHT(rectangle2_heights[2532]), .RECT2_WEIGHT(rectangle2_weights[2532]), .RECT3_X(rectangle3_xs[2532]), .RECT3_Y(rectangle3_ys[2532]), .RECT3_WIDTH(rectangle3_widths[2532]), .RECT3_HEIGHT(rectangle3_heights[2532]), .RECT3_WEIGHT(rectangle3_weights[2532]), .FEAT_THRES(feature_thresholds[2532]), .FEAT_ABOVE(feature_aboves[2532]), .FEAT_BELOW(feature_belows[2532])) ac2532(.scan_win(scan_win2532), .scan_win_std_dev(scan_win_std_dev[2532]), .feature_accum(feature_accums[2532]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2533]), .RECT1_Y(rectangle1_ys[2533]), .RECT1_WIDTH(rectangle1_widths[2533]), .RECT1_HEIGHT(rectangle1_heights[2533]), .RECT1_WEIGHT(rectangle1_weights[2533]), .RECT2_X(rectangle2_xs[2533]), .RECT2_Y(rectangle2_ys[2533]), .RECT2_WIDTH(rectangle2_widths[2533]), .RECT2_HEIGHT(rectangle2_heights[2533]), .RECT2_WEIGHT(rectangle2_weights[2533]), .RECT3_X(rectangle3_xs[2533]), .RECT3_Y(rectangle3_ys[2533]), .RECT3_WIDTH(rectangle3_widths[2533]), .RECT3_HEIGHT(rectangle3_heights[2533]), .RECT3_WEIGHT(rectangle3_weights[2533]), .FEAT_THRES(feature_thresholds[2533]), .FEAT_ABOVE(feature_aboves[2533]), .FEAT_BELOW(feature_belows[2533])) ac2533(.scan_win(scan_win2533), .scan_win_std_dev(scan_win_std_dev[2533]), .feature_accum(feature_accums[2533]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2534]), .RECT1_Y(rectangle1_ys[2534]), .RECT1_WIDTH(rectangle1_widths[2534]), .RECT1_HEIGHT(rectangle1_heights[2534]), .RECT1_WEIGHT(rectangle1_weights[2534]), .RECT2_X(rectangle2_xs[2534]), .RECT2_Y(rectangle2_ys[2534]), .RECT2_WIDTH(rectangle2_widths[2534]), .RECT2_HEIGHT(rectangle2_heights[2534]), .RECT2_WEIGHT(rectangle2_weights[2534]), .RECT3_X(rectangle3_xs[2534]), .RECT3_Y(rectangle3_ys[2534]), .RECT3_WIDTH(rectangle3_widths[2534]), .RECT3_HEIGHT(rectangle3_heights[2534]), .RECT3_WEIGHT(rectangle3_weights[2534]), .FEAT_THRES(feature_thresholds[2534]), .FEAT_ABOVE(feature_aboves[2534]), .FEAT_BELOW(feature_belows[2534])) ac2534(.scan_win(scan_win2534), .scan_win_std_dev(scan_win_std_dev[2534]), .feature_accum(feature_accums[2534]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2535]), .RECT1_Y(rectangle1_ys[2535]), .RECT1_WIDTH(rectangle1_widths[2535]), .RECT1_HEIGHT(rectangle1_heights[2535]), .RECT1_WEIGHT(rectangle1_weights[2535]), .RECT2_X(rectangle2_xs[2535]), .RECT2_Y(rectangle2_ys[2535]), .RECT2_WIDTH(rectangle2_widths[2535]), .RECT2_HEIGHT(rectangle2_heights[2535]), .RECT2_WEIGHT(rectangle2_weights[2535]), .RECT3_X(rectangle3_xs[2535]), .RECT3_Y(rectangle3_ys[2535]), .RECT3_WIDTH(rectangle3_widths[2535]), .RECT3_HEIGHT(rectangle3_heights[2535]), .RECT3_WEIGHT(rectangle3_weights[2535]), .FEAT_THRES(feature_thresholds[2535]), .FEAT_ABOVE(feature_aboves[2535]), .FEAT_BELOW(feature_belows[2535])) ac2535(.scan_win(scan_win2535), .scan_win_std_dev(scan_win_std_dev[2535]), .feature_accum(feature_accums[2535]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2536]), .RECT1_Y(rectangle1_ys[2536]), .RECT1_WIDTH(rectangle1_widths[2536]), .RECT1_HEIGHT(rectangle1_heights[2536]), .RECT1_WEIGHT(rectangle1_weights[2536]), .RECT2_X(rectangle2_xs[2536]), .RECT2_Y(rectangle2_ys[2536]), .RECT2_WIDTH(rectangle2_widths[2536]), .RECT2_HEIGHT(rectangle2_heights[2536]), .RECT2_WEIGHT(rectangle2_weights[2536]), .RECT3_X(rectangle3_xs[2536]), .RECT3_Y(rectangle3_ys[2536]), .RECT3_WIDTH(rectangle3_widths[2536]), .RECT3_HEIGHT(rectangle3_heights[2536]), .RECT3_WEIGHT(rectangle3_weights[2536]), .FEAT_THRES(feature_thresholds[2536]), .FEAT_ABOVE(feature_aboves[2536]), .FEAT_BELOW(feature_belows[2536])) ac2536(.scan_win(scan_win2536), .scan_win_std_dev(scan_win_std_dev[2536]), .feature_accum(feature_accums[2536]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2537]), .RECT1_Y(rectangle1_ys[2537]), .RECT1_WIDTH(rectangle1_widths[2537]), .RECT1_HEIGHT(rectangle1_heights[2537]), .RECT1_WEIGHT(rectangle1_weights[2537]), .RECT2_X(rectangle2_xs[2537]), .RECT2_Y(rectangle2_ys[2537]), .RECT2_WIDTH(rectangle2_widths[2537]), .RECT2_HEIGHT(rectangle2_heights[2537]), .RECT2_WEIGHT(rectangle2_weights[2537]), .RECT3_X(rectangle3_xs[2537]), .RECT3_Y(rectangle3_ys[2537]), .RECT3_WIDTH(rectangle3_widths[2537]), .RECT3_HEIGHT(rectangle3_heights[2537]), .RECT3_WEIGHT(rectangle3_weights[2537]), .FEAT_THRES(feature_thresholds[2537]), .FEAT_ABOVE(feature_aboves[2537]), .FEAT_BELOW(feature_belows[2537])) ac2537(.scan_win(scan_win2537), .scan_win_std_dev(scan_win_std_dev[2537]), .feature_accum(feature_accums[2537]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2538]), .RECT1_Y(rectangle1_ys[2538]), .RECT1_WIDTH(rectangle1_widths[2538]), .RECT1_HEIGHT(rectangle1_heights[2538]), .RECT1_WEIGHT(rectangle1_weights[2538]), .RECT2_X(rectangle2_xs[2538]), .RECT2_Y(rectangle2_ys[2538]), .RECT2_WIDTH(rectangle2_widths[2538]), .RECT2_HEIGHT(rectangle2_heights[2538]), .RECT2_WEIGHT(rectangle2_weights[2538]), .RECT3_X(rectangle3_xs[2538]), .RECT3_Y(rectangle3_ys[2538]), .RECT3_WIDTH(rectangle3_widths[2538]), .RECT3_HEIGHT(rectangle3_heights[2538]), .RECT3_WEIGHT(rectangle3_weights[2538]), .FEAT_THRES(feature_thresholds[2538]), .FEAT_ABOVE(feature_aboves[2538]), .FEAT_BELOW(feature_belows[2538])) ac2538(.scan_win(scan_win2538), .scan_win_std_dev(scan_win_std_dev[2538]), .feature_accum(feature_accums[2538]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2539]), .RECT1_Y(rectangle1_ys[2539]), .RECT1_WIDTH(rectangle1_widths[2539]), .RECT1_HEIGHT(rectangle1_heights[2539]), .RECT1_WEIGHT(rectangle1_weights[2539]), .RECT2_X(rectangle2_xs[2539]), .RECT2_Y(rectangle2_ys[2539]), .RECT2_WIDTH(rectangle2_widths[2539]), .RECT2_HEIGHT(rectangle2_heights[2539]), .RECT2_WEIGHT(rectangle2_weights[2539]), .RECT3_X(rectangle3_xs[2539]), .RECT3_Y(rectangle3_ys[2539]), .RECT3_WIDTH(rectangle3_widths[2539]), .RECT3_HEIGHT(rectangle3_heights[2539]), .RECT3_WEIGHT(rectangle3_weights[2539]), .FEAT_THRES(feature_thresholds[2539]), .FEAT_ABOVE(feature_aboves[2539]), .FEAT_BELOW(feature_belows[2539])) ac2539(.scan_win(scan_win2539), .scan_win_std_dev(scan_win_std_dev[2539]), .feature_accum(feature_accums[2539]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2540]), .RECT1_Y(rectangle1_ys[2540]), .RECT1_WIDTH(rectangle1_widths[2540]), .RECT1_HEIGHT(rectangle1_heights[2540]), .RECT1_WEIGHT(rectangle1_weights[2540]), .RECT2_X(rectangle2_xs[2540]), .RECT2_Y(rectangle2_ys[2540]), .RECT2_WIDTH(rectangle2_widths[2540]), .RECT2_HEIGHT(rectangle2_heights[2540]), .RECT2_WEIGHT(rectangle2_weights[2540]), .RECT3_X(rectangle3_xs[2540]), .RECT3_Y(rectangle3_ys[2540]), .RECT3_WIDTH(rectangle3_widths[2540]), .RECT3_HEIGHT(rectangle3_heights[2540]), .RECT3_WEIGHT(rectangle3_weights[2540]), .FEAT_THRES(feature_thresholds[2540]), .FEAT_ABOVE(feature_aboves[2540]), .FEAT_BELOW(feature_belows[2540])) ac2540(.scan_win(scan_win2540), .scan_win_std_dev(scan_win_std_dev[2540]), .feature_accum(feature_accums[2540]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2541]), .RECT1_Y(rectangle1_ys[2541]), .RECT1_WIDTH(rectangle1_widths[2541]), .RECT1_HEIGHT(rectangle1_heights[2541]), .RECT1_WEIGHT(rectangle1_weights[2541]), .RECT2_X(rectangle2_xs[2541]), .RECT2_Y(rectangle2_ys[2541]), .RECT2_WIDTH(rectangle2_widths[2541]), .RECT2_HEIGHT(rectangle2_heights[2541]), .RECT2_WEIGHT(rectangle2_weights[2541]), .RECT3_X(rectangle3_xs[2541]), .RECT3_Y(rectangle3_ys[2541]), .RECT3_WIDTH(rectangle3_widths[2541]), .RECT3_HEIGHT(rectangle3_heights[2541]), .RECT3_WEIGHT(rectangle3_weights[2541]), .FEAT_THRES(feature_thresholds[2541]), .FEAT_ABOVE(feature_aboves[2541]), .FEAT_BELOW(feature_belows[2541])) ac2541(.scan_win(scan_win2541), .scan_win_std_dev(scan_win_std_dev[2541]), .feature_accum(feature_accums[2541]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2542]), .RECT1_Y(rectangle1_ys[2542]), .RECT1_WIDTH(rectangle1_widths[2542]), .RECT1_HEIGHT(rectangle1_heights[2542]), .RECT1_WEIGHT(rectangle1_weights[2542]), .RECT2_X(rectangle2_xs[2542]), .RECT2_Y(rectangle2_ys[2542]), .RECT2_WIDTH(rectangle2_widths[2542]), .RECT2_HEIGHT(rectangle2_heights[2542]), .RECT2_WEIGHT(rectangle2_weights[2542]), .RECT3_X(rectangle3_xs[2542]), .RECT3_Y(rectangle3_ys[2542]), .RECT3_WIDTH(rectangle3_widths[2542]), .RECT3_HEIGHT(rectangle3_heights[2542]), .RECT3_WEIGHT(rectangle3_weights[2542]), .FEAT_THRES(feature_thresholds[2542]), .FEAT_ABOVE(feature_aboves[2542]), .FEAT_BELOW(feature_belows[2542])) ac2542(.scan_win(scan_win2542), .scan_win_std_dev(scan_win_std_dev[2542]), .feature_accum(feature_accums[2542]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2543]), .RECT1_Y(rectangle1_ys[2543]), .RECT1_WIDTH(rectangle1_widths[2543]), .RECT1_HEIGHT(rectangle1_heights[2543]), .RECT1_WEIGHT(rectangle1_weights[2543]), .RECT2_X(rectangle2_xs[2543]), .RECT2_Y(rectangle2_ys[2543]), .RECT2_WIDTH(rectangle2_widths[2543]), .RECT2_HEIGHT(rectangle2_heights[2543]), .RECT2_WEIGHT(rectangle2_weights[2543]), .RECT3_X(rectangle3_xs[2543]), .RECT3_Y(rectangle3_ys[2543]), .RECT3_WIDTH(rectangle3_widths[2543]), .RECT3_HEIGHT(rectangle3_heights[2543]), .RECT3_WEIGHT(rectangle3_weights[2543]), .FEAT_THRES(feature_thresholds[2543]), .FEAT_ABOVE(feature_aboves[2543]), .FEAT_BELOW(feature_belows[2543])) ac2543(.scan_win(scan_win2543), .scan_win_std_dev(scan_win_std_dev[2543]), .feature_accum(feature_accums[2543]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2544]), .RECT1_Y(rectangle1_ys[2544]), .RECT1_WIDTH(rectangle1_widths[2544]), .RECT1_HEIGHT(rectangle1_heights[2544]), .RECT1_WEIGHT(rectangle1_weights[2544]), .RECT2_X(rectangle2_xs[2544]), .RECT2_Y(rectangle2_ys[2544]), .RECT2_WIDTH(rectangle2_widths[2544]), .RECT2_HEIGHT(rectangle2_heights[2544]), .RECT2_WEIGHT(rectangle2_weights[2544]), .RECT3_X(rectangle3_xs[2544]), .RECT3_Y(rectangle3_ys[2544]), .RECT3_WIDTH(rectangle3_widths[2544]), .RECT3_HEIGHT(rectangle3_heights[2544]), .RECT3_WEIGHT(rectangle3_weights[2544]), .FEAT_THRES(feature_thresholds[2544]), .FEAT_ABOVE(feature_aboves[2544]), .FEAT_BELOW(feature_belows[2544])) ac2544(.scan_win(scan_win2544), .scan_win_std_dev(scan_win_std_dev[2544]), .feature_accum(feature_accums[2544]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2545]), .RECT1_Y(rectangle1_ys[2545]), .RECT1_WIDTH(rectangle1_widths[2545]), .RECT1_HEIGHT(rectangle1_heights[2545]), .RECT1_WEIGHT(rectangle1_weights[2545]), .RECT2_X(rectangle2_xs[2545]), .RECT2_Y(rectangle2_ys[2545]), .RECT2_WIDTH(rectangle2_widths[2545]), .RECT2_HEIGHT(rectangle2_heights[2545]), .RECT2_WEIGHT(rectangle2_weights[2545]), .RECT3_X(rectangle3_xs[2545]), .RECT3_Y(rectangle3_ys[2545]), .RECT3_WIDTH(rectangle3_widths[2545]), .RECT3_HEIGHT(rectangle3_heights[2545]), .RECT3_WEIGHT(rectangle3_weights[2545]), .FEAT_THRES(feature_thresholds[2545]), .FEAT_ABOVE(feature_aboves[2545]), .FEAT_BELOW(feature_belows[2545])) ac2545(.scan_win(scan_win2545), .scan_win_std_dev(scan_win_std_dev[2545]), .feature_accum(feature_accums[2545]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2546]), .RECT1_Y(rectangle1_ys[2546]), .RECT1_WIDTH(rectangle1_widths[2546]), .RECT1_HEIGHT(rectangle1_heights[2546]), .RECT1_WEIGHT(rectangle1_weights[2546]), .RECT2_X(rectangle2_xs[2546]), .RECT2_Y(rectangle2_ys[2546]), .RECT2_WIDTH(rectangle2_widths[2546]), .RECT2_HEIGHT(rectangle2_heights[2546]), .RECT2_WEIGHT(rectangle2_weights[2546]), .RECT3_X(rectangle3_xs[2546]), .RECT3_Y(rectangle3_ys[2546]), .RECT3_WIDTH(rectangle3_widths[2546]), .RECT3_HEIGHT(rectangle3_heights[2546]), .RECT3_WEIGHT(rectangle3_weights[2546]), .FEAT_THRES(feature_thresholds[2546]), .FEAT_ABOVE(feature_aboves[2546]), .FEAT_BELOW(feature_belows[2546])) ac2546(.scan_win(scan_win2546), .scan_win_std_dev(scan_win_std_dev[2546]), .feature_accum(feature_accums[2546]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2547]), .RECT1_Y(rectangle1_ys[2547]), .RECT1_WIDTH(rectangle1_widths[2547]), .RECT1_HEIGHT(rectangle1_heights[2547]), .RECT1_WEIGHT(rectangle1_weights[2547]), .RECT2_X(rectangle2_xs[2547]), .RECT2_Y(rectangle2_ys[2547]), .RECT2_WIDTH(rectangle2_widths[2547]), .RECT2_HEIGHT(rectangle2_heights[2547]), .RECT2_WEIGHT(rectangle2_weights[2547]), .RECT3_X(rectangle3_xs[2547]), .RECT3_Y(rectangle3_ys[2547]), .RECT3_WIDTH(rectangle3_widths[2547]), .RECT3_HEIGHT(rectangle3_heights[2547]), .RECT3_WEIGHT(rectangle3_weights[2547]), .FEAT_THRES(feature_thresholds[2547]), .FEAT_ABOVE(feature_aboves[2547]), .FEAT_BELOW(feature_belows[2547])) ac2547(.scan_win(scan_win2547), .scan_win_std_dev(scan_win_std_dev[2547]), .feature_accum(feature_accums[2547]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2548]), .RECT1_Y(rectangle1_ys[2548]), .RECT1_WIDTH(rectangle1_widths[2548]), .RECT1_HEIGHT(rectangle1_heights[2548]), .RECT1_WEIGHT(rectangle1_weights[2548]), .RECT2_X(rectangle2_xs[2548]), .RECT2_Y(rectangle2_ys[2548]), .RECT2_WIDTH(rectangle2_widths[2548]), .RECT2_HEIGHT(rectangle2_heights[2548]), .RECT2_WEIGHT(rectangle2_weights[2548]), .RECT3_X(rectangle3_xs[2548]), .RECT3_Y(rectangle3_ys[2548]), .RECT3_WIDTH(rectangle3_widths[2548]), .RECT3_HEIGHT(rectangle3_heights[2548]), .RECT3_WEIGHT(rectangle3_weights[2548]), .FEAT_THRES(feature_thresholds[2548]), .FEAT_ABOVE(feature_aboves[2548]), .FEAT_BELOW(feature_belows[2548])) ac2548(.scan_win(scan_win2548), .scan_win_std_dev(scan_win_std_dev[2548]), .feature_accum(feature_accums[2548]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2549]), .RECT1_Y(rectangle1_ys[2549]), .RECT1_WIDTH(rectangle1_widths[2549]), .RECT1_HEIGHT(rectangle1_heights[2549]), .RECT1_WEIGHT(rectangle1_weights[2549]), .RECT2_X(rectangle2_xs[2549]), .RECT2_Y(rectangle2_ys[2549]), .RECT2_WIDTH(rectangle2_widths[2549]), .RECT2_HEIGHT(rectangle2_heights[2549]), .RECT2_WEIGHT(rectangle2_weights[2549]), .RECT3_X(rectangle3_xs[2549]), .RECT3_Y(rectangle3_ys[2549]), .RECT3_WIDTH(rectangle3_widths[2549]), .RECT3_HEIGHT(rectangle3_heights[2549]), .RECT3_WEIGHT(rectangle3_weights[2549]), .FEAT_THRES(feature_thresholds[2549]), .FEAT_ABOVE(feature_aboves[2549]), .FEAT_BELOW(feature_belows[2549])) ac2549(.scan_win(scan_win2549), .scan_win_std_dev(scan_win_std_dev[2549]), .feature_accum(feature_accums[2549]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2550]), .RECT1_Y(rectangle1_ys[2550]), .RECT1_WIDTH(rectangle1_widths[2550]), .RECT1_HEIGHT(rectangle1_heights[2550]), .RECT1_WEIGHT(rectangle1_weights[2550]), .RECT2_X(rectangle2_xs[2550]), .RECT2_Y(rectangle2_ys[2550]), .RECT2_WIDTH(rectangle2_widths[2550]), .RECT2_HEIGHT(rectangle2_heights[2550]), .RECT2_WEIGHT(rectangle2_weights[2550]), .RECT3_X(rectangle3_xs[2550]), .RECT3_Y(rectangle3_ys[2550]), .RECT3_WIDTH(rectangle3_widths[2550]), .RECT3_HEIGHT(rectangle3_heights[2550]), .RECT3_WEIGHT(rectangle3_weights[2550]), .FEAT_THRES(feature_thresholds[2550]), .FEAT_ABOVE(feature_aboves[2550]), .FEAT_BELOW(feature_belows[2550])) ac2550(.scan_win(scan_win2550), .scan_win_std_dev(scan_win_std_dev[2550]), .feature_accum(feature_accums[2550]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2551]), .RECT1_Y(rectangle1_ys[2551]), .RECT1_WIDTH(rectangle1_widths[2551]), .RECT1_HEIGHT(rectangle1_heights[2551]), .RECT1_WEIGHT(rectangle1_weights[2551]), .RECT2_X(rectangle2_xs[2551]), .RECT2_Y(rectangle2_ys[2551]), .RECT2_WIDTH(rectangle2_widths[2551]), .RECT2_HEIGHT(rectangle2_heights[2551]), .RECT2_WEIGHT(rectangle2_weights[2551]), .RECT3_X(rectangle3_xs[2551]), .RECT3_Y(rectangle3_ys[2551]), .RECT3_WIDTH(rectangle3_widths[2551]), .RECT3_HEIGHT(rectangle3_heights[2551]), .RECT3_WEIGHT(rectangle3_weights[2551]), .FEAT_THRES(feature_thresholds[2551]), .FEAT_ABOVE(feature_aboves[2551]), .FEAT_BELOW(feature_belows[2551])) ac2551(.scan_win(scan_win2551), .scan_win_std_dev(scan_win_std_dev[2551]), .feature_accum(feature_accums[2551]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2552]), .RECT1_Y(rectangle1_ys[2552]), .RECT1_WIDTH(rectangle1_widths[2552]), .RECT1_HEIGHT(rectangle1_heights[2552]), .RECT1_WEIGHT(rectangle1_weights[2552]), .RECT2_X(rectangle2_xs[2552]), .RECT2_Y(rectangle2_ys[2552]), .RECT2_WIDTH(rectangle2_widths[2552]), .RECT2_HEIGHT(rectangle2_heights[2552]), .RECT2_WEIGHT(rectangle2_weights[2552]), .RECT3_X(rectangle3_xs[2552]), .RECT3_Y(rectangle3_ys[2552]), .RECT3_WIDTH(rectangle3_widths[2552]), .RECT3_HEIGHT(rectangle3_heights[2552]), .RECT3_WEIGHT(rectangle3_weights[2552]), .FEAT_THRES(feature_thresholds[2552]), .FEAT_ABOVE(feature_aboves[2552]), .FEAT_BELOW(feature_belows[2552])) ac2552(.scan_win(scan_win2552), .scan_win_std_dev(scan_win_std_dev[2552]), .feature_accum(feature_accums[2552]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2553]), .RECT1_Y(rectangle1_ys[2553]), .RECT1_WIDTH(rectangle1_widths[2553]), .RECT1_HEIGHT(rectangle1_heights[2553]), .RECT1_WEIGHT(rectangle1_weights[2553]), .RECT2_X(rectangle2_xs[2553]), .RECT2_Y(rectangle2_ys[2553]), .RECT2_WIDTH(rectangle2_widths[2553]), .RECT2_HEIGHT(rectangle2_heights[2553]), .RECT2_WEIGHT(rectangle2_weights[2553]), .RECT3_X(rectangle3_xs[2553]), .RECT3_Y(rectangle3_ys[2553]), .RECT3_WIDTH(rectangle3_widths[2553]), .RECT3_HEIGHT(rectangle3_heights[2553]), .RECT3_WEIGHT(rectangle3_weights[2553]), .FEAT_THRES(feature_thresholds[2553]), .FEAT_ABOVE(feature_aboves[2553]), .FEAT_BELOW(feature_belows[2553])) ac2553(.scan_win(scan_win2553), .scan_win_std_dev(scan_win_std_dev[2553]), .feature_accum(feature_accums[2553]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2554]), .RECT1_Y(rectangle1_ys[2554]), .RECT1_WIDTH(rectangle1_widths[2554]), .RECT1_HEIGHT(rectangle1_heights[2554]), .RECT1_WEIGHT(rectangle1_weights[2554]), .RECT2_X(rectangle2_xs[2554]), .RECT2_Y(rectangle2_ys[2554]), .RECT2_WIDTH(rectangle2_widths[2554]), .RECT2_HEIGHT(rectangle2_heights[2554]), .RECT2_WEIGHT(rectangle2_weights[2554]), .RECT3_X(rectangle3_xs[2554]), .RECT3_Y(rectangle3_ys[2554]), .RECT3_WIDTH(rectangle3_widths[2554]), .RECT3_HEIGHT(rectangle3_heights[2554]), .RECT3_WEIGHT(rectangle3_weights[2554]), .FEAT_THRES(feature_thresholds[2554]), .FEAT_ABOVE(feature_aboves[2554]), .FEAT_BELOW(feature_belows[2554])) ac2554(.scan_win(scan_win2554), .scan_win_std_dev(scan_win_std_dev[2554]), .feature_accum(feature_accums[2554]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2555]), .RECT1_Y(rectangle1_ys[2555]), .RECT1_WIDTH(rectangle1_widths[2555]), .RECT1_HEIGHT(rectangle1_heights[2555]), .RECT1_WEIGHT(rectangle1_weights[2555]), .RECT2_X(rectangle2_xs[2555]), .RECT2_Y(rectangle2_ys[2555]), .RECT2_WIDTH(rectangle2_widths[2555]), .RECT2_HEIGHT(rectangle2_heights[2555]), .RECT2_WEIGHT(rectangle2_weights[2555]), .RECT3_X(rectangle3_xs[2555]), .RECT3_Y(rectangle3_ys[2555]), .RECT3_WIDTH(rectangle3_widths[2555]), .RECT3_HEIGHT(rectangle3_heights[2555]), .RECT3_WEIGHT(rectangle3_weights[2555]), .FEAT_THRES(feature_thresholds[2555]), .FEAT_ABOVE(feature_aboves[2555]), .FEAT_BELOW(feature_belows[2555])) ac2555(.scan_win(scan_win2555), .scan_win_std_dev(scan_win_std_dev[2555]), .feature_accum(feature_accums[2555]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2556]), .RECT1_Y(rectangle1_ys[2556]), .RECT1_WIDTH(rectangle1_widths[2556]), .RECT1_HEIGHT(rectangle1_heights[2556]), .RECT1_WEIGHT(rectangle1_weights[2556]), .RECT2_X(rectangle2_xs[2556]), .RECT2_Y(rectangle2_ys[2556]), .RECT2_WIDTH(rectangle2_widths[2556]), .RECT2_HEIGHT(rectangle2_heights[2556]), .RECT2_WEIGHT(rectangle2_weights[2556]), .RECT3_X(rectangle3_xs[2556]), .RECT3_Y(rectangle3_ys[2556]), .RECT3_WIDTH(rectangle3_widths[2556]), .RECT3_HEIGHT(rectangle3_heights[2556]), .RECT3_WEIGHT(rectangle3_weights[2556]), .FEAT_THRES(feature_thresholds[2556]), .FEAT_ABOVE(feature_aboves[2556]), .FEAT_BELOW(feature_belows[2556])) ac2556(.scan_win(scan_win2556), .scan_win_std_dev(scan_win_std_dev[2556]), .feature_accum(feature_accums[2556]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2557]), .RECT1_Y(rectangle1_ys[2557]), .RECT1_WIDTH(rectangle1_widths[2557]), .RECT1_HEIGHT(rectangle1_heights[2557]), .RECT1_WEIGHT(rectangle1_weights[2557]), .RECT2_X(rectangle2_xs[2557]), .RECT2_Y(rectangle2_ys[2557]), .RECT2_WIDTH(rectangle2_widths[2557]), .RECT2_HEIGHT(rectangle2_heights[2557]), .RECT2_WEIGHT(rectangle2_weights[2557]), .RECT3_X(rectangle3_xs[2557]), .RECT3_Y(rectangle3_ys[2557]), .RECT3_WIDTH(rectangle3_widths[2557]), .RECT3_HEIGHT(rectangle3_heights[2557]), .RECT3_WEIGHT(rectangle3_weights[2557]), .FEAT_THRES(feature_thresholds[2557]), .FEAT_ABOVE(feature_aboves[2557]), .FEAT_BELOW(feature_belows[2557])) ac2557(.scan_win(scan_win2557), .scan_win_std_dev(scan_win_std_dev[2557]), .feature_accum(feature_accums[2557]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2558]), .RECT1_Y(rectangle1_ys[2558]), .RECT1_WIDTH(rectangle1_widths[2558]), .RECT1_HEIGHT(rectangle1_heights[2558]), .RECT1_WEIGHT(rectangle1_weights[2558]), .RECT2_X(rectangle2_xs[2558]), .RECT2_Y(rectangle2_ys[2558]), .RECT2_WIDTH(rectangle2_widths[2558]), .RECT2_HEIGHT(rectangle2_heights[2558]), .RECT2_WEIGHT(rectangle2_weights[2558]), .RECT3_X(rectangle3_xs[2558]), .RECT3_Y(rectangle3_ys[2558]), .RECT3_WIDTH(rectangle3_widths[2558]), .RECT3_HEIGHT(rectangle3_heights[2558]), .RECT3_WEIGHT(rectangle3_weights[2558]), .FEAT_THRES(feature_thresholds[2558]), .FEAT_ABOVE(feature_aboves[2558]), .FEAT_BELOW(feature_belows[2558])) ac2558(.scan_win(scan_win2558), .scan_win_std_dev(scan_win_std_dev[2558]), .feature_accum(feature_accums[2558]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2559]), .RECT1_Y(rectangle1_ys[2559]), .RECT1_WIDTH(rectangle1_widths[2559]), .RECT1_HEIGHT(rectangle1_heights[2559]), .RECT1_WEIGHT(rectangle1_weights[2559]), .RECT2_X(rectangle2_xs[2559]), .RECT2_Y(rectangle2_ys[2559]), .RECT2_WIDTH(rectangle2_widths[2559]), .RECT2_HEIGHT(rectangle2_heights[2559]), .RECT2_WEIGHT(rectangle2_weights[2559]), .RECT3_X(rectangle3_xs[2559]), .RECT3_Y(rectangle3_ys[2559]), .RECT3_WIDTH(rectangle3_widths[2559]), .RECT3_HEIGHT(rectangle3_heights[2559]), .RECT3_WEIGHT(rectangle3_weights[2559]), .FEAT_THRES(feature_thresholds[2559]), .FEAT_ABOVE(feature_aboves[2559]), .FEAT_BELOW(feature_belows[2559])) ac2559(.scan_win(scan_win2559), .scan_win_std_dev(scan_win_std_dev[2559]), .feature_accum(feature_accums[2559]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2560]), .RECT1_Y(rectangle1_ys[2560]), .RECT1_WIDTH(rectangle1_widths[2560]), .RECT1_HEIGHT(rectangle1_heights[2560]), .RECT1_WEIGHT(rectangle1_weights[2560]), .RECT2_X(rectangle2_xs[2560]), .RECT2_Y(rectangle2_ys[2560]), .RECT2_WIDTH(rectangle2_widths[2560]), .RECT2_HEIGHT(rectangle2_heights[2560]), .RECT2_WEIGHT(rectangle2_weights[2560]), .RECT3_X(rectangle3_xs[2560]), .RECT3_Y(rectangle3_ys[2560]), .RECT3_WIDTH(rectangle3_widths[2560]), .RECT3_HEIGHT(rectangle3_heights[2560]), .RECT3_WEIGHT(rectangle3_weights[2560]), .FEAT_THRES(feature_thresholds[2560]), .FEAT_ABOVE(feature_aboves[2560]), .FEAT_BELOW(feature_belows[2560])) ac2560(.scan_win(scan_win2560), .scan_win_std_dev(scan_win_std_dev[2560]), .feature_accum(feature_accums[2560]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2561]), .RECT1_Y(rectangle1_ys[2561]), .RECT1_WIDTH(rectangle1_widths[2561]), .RECT1_HEIGHT(rectangle1_heights[2561]), .RECT1_WEIGHT(rectangle1_weights[2561]), .RECT2_X(rectangle2_xs[2561]), .RECT2_Y(rectangle2_ys[2561]), .RECT2_WIDTH(rectangle2_widths[2561]), .RECT2_HEIGHT(rectangle2_heights[2561]), .RECT2_WEIGHT(rectangle2_weights[2561]), .RECT3_X(rectangle3_xs[2561]), .RECT3_Y(rectangle3_ys[2561]), .RECT3_WIDTH(rectangle3_widths[2561]), .RECT3_HEIGHT(rectangle3_heights[2561]), .RECT3_WEIGHT(rectangle3_weights[2561]), .FEAT_THRES(feature_thresholds[2561]), .FEAT_ABOVE(feature_aboves[2561]), .FEAT_BELOW(feature_belows[2561])) ac2561(.scan_win(scan_win2561), .scan_win_std_dev(scan_win_std_dev[2561]), .feature_accum(feature_accums[2561]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2562]), .RECT1_Y(rectangle1_ys[2562]), .RECT1_WIDTH(rectangle1_widths[2562]), .RECT1_HEIGHT(rectangle1_heights[2562]), .RECT1_WEIGHT(rectangle1_weights[2562]), .RECT2_X(rectangle2_xs[2562]), .RECT2_Y(rectangle2_ys[2562]), .RECT2_WIDTH(rectangle2_widths[2562]), .RECT2_HEIGHT(rectangle2_heights[2562]), .RECT2_WEIGHT(rectangle2_weights[2562]), .RECT3_X(rectangle3_xs[2562]), .RECT3_Y(rectangle3_ys[2562]), .RECT3_WIDTH(rectangle3_widths[2562]), .RECT3_HEIGHT(rectangle3_heights[2562]), .RECT3_WEIGHT(rectangle3_weights[2562]), .FEAT_THRES(feature_thresholds[2562]), .FEAT_ABOVE(feature_aboves[2562]), .FEAT_BELOW(feature_belows[2562])) ac2562(.scan_win(scan_win2562), .scan_win_std_dev(scan_win_std_dev[2562]), .feature_accum(feature_accums[2562]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2563]), .RECT1_Y(rectangle1_ys[2563]), .RECT1_WIDTH(rectangle1_widths[2563]), .RECT1_HEIGHT(rectangle1_heights[2563]), .RECT1_WEIGHT(rectangle1_weights[2563]), .RECT2_X(rectangle2_xs[2563]), .RECT2_Y(rectangle2_ys[2563]), .RECT2_WIDTH(rectangle2_widths[2563]), .RECT2_HEIGHT(rectangle2_heights[2563]), .RECT2_WEIGHT(rectangle2_weights[2563]), .RECT3_X(rectangle3_xs[2563]), .RECT3_Y(rectangle3_ys[2563]), .RECT3_WIDTH(rectangle3_widths[2563]), .RECT3_HEIGHT(rectangle3_heights[2563]), .RECT3_WEIGHT(rectangle3_weights[2563]), .FEAT_THRES(feature_thresholds[2563]), .FEAT_ABOVE(feature_aboves[2563]), .FEAT_BELOW(feature_belows[2563])) ac2563(.scan_win(scan_win2563), .scan_win_std_dev(scan_win_std_dev[2563]), .feature_accum(feature_accums[2563]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2564]), .RECT1_Y(rectangle1_ys[2564]), .RECT1_WIDTH(rectangle1_widths[2564]), .RECT1_HEIGHT(rectangle1_heights[2564]), .RECT1_WEIGHT(rectangle1_weights[2564]), .RECT2_X(rectangle2_xs[2564]), .RECT2_Y(rectangle2_ys[2564]), .RECT2_WIDTH(rectangle2_widths[2564]), .RECT2_HEIGHT(rectangle2_heights[2564]), .RECT2_WEIGHT(rectangle2_weights[2564]), .RECT3_X(rectangle3_xs[2564]), .RECT3_Y(rectangle3_ys[2564]), .RECT3_WIDTH(rectangle3_widths[2564]), .RECT3_HEIGHT(rectangle3_heights[2564]), .RECT3_WEIGHT(rectangle3_weights[2564]), .FEAT_THRES(feature_thresholds[2564]), .FEAT_ABOVE(feature_aboves[2564]), .FEAT_BELOW(feature_belows[2564])) ac2564(.scan_win(scan_win2564), .scan_win_std_dev(scan_win_std_dev[2564]), .feature_accum(feature_accums[2564]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2565]), .RECT1_Y(rectangle1_ys[2565]), .RECT1_WIDTH(rectangle1_widths[2565]), .RECT1_HEIGHT(rectangle1_heights[2565]), .RECT1_WEIGHT(rectangle1_weights[2565]), .RECT2_X(rectangle2_xs[2565]), .RECT2_Y(rectangle2_ys[2565]), .RECT2_WIDTH(rectangle2_widths[2565]), .RECT2_HEIGHT(rectangle2_heights[2565]), .RECT2_WEIGHT(rectangle2_weights[2565]), .RECT3_X(rectangle3_xs[2565]), .RECT3_Y(rectangle3_ys[2565]), .RECT3_WIDTH(rectangle3_widths[2565]), .RECT3_HEIGHT(rectangle3_heights[2565]), .RECT3_WEIGHT(rectangle3_weights[2565]), .FEAT_THRES(feature_thresholds[2565]), .FEAT_ABOVE(feature_aboves[2565]), .FEAT_BELOW(feature_belows[2565])) ac2565(.scan_win(scan_win2565), .scan_win_std_dev(scan_win_std_dev[2565]), .feature_accum(feature_accums[2565]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2566]), .RECT1_Y(rectangle1_ys[2566]), .RECT1_WIDTH(rectangle1_widths[2566]), .RECT1_HEIGHT(rectangle1_heights[2566]), .RECT1_WEIGHT(rectangle1_weights[2566]), .RECT2_X(rectangle2_xs[2566]), .RECT2_Y(rectangle2_ys[2566]), .RECT2_WIDTH(rectangle2_widths[2566]), .RECT2_HEIGHT(rectangle2_heights[2566]), .RECT2_WEIGHT(rectangle2_weights[2566]), .RECT3_X(rectangle3_xs[2566]), .RECT3_Y(rectangle3_ys[2566]), .RECT3_WIDTH(rectangle3_widths[2566]), .RECT3_HEIGHT(rectangle3_heights[2566]), .RECT3_WEIGHT(rectangle3_weights[2566]), .FEAT_THRES(feature_thresholds[2566]), .FEAT_ABOVE(feature_aboves[2566]), .FEAT_BELOW(feature_belows[2566])) ac2566(.scan_win(scan_win2566), .scan_win_std_dev(scan_win_std_dev[2566]), .feature_accum(feature_accums[2566]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2567]), .RECT1_Y(rectangle1_ys[2567]), .RECT1_WIDTH(rectangle1_widths[2567]), .RECT1_HEIGHT(rectangle1_heights[2567]), .RECT1_WEIGHT(rectangle1_weights[2567]), .RECT2_X(rectangle2_xs[2567]), .RECT2_Y(rectangle2_ys[2567]), .RECT2_WIDTH(rectangle2_widths[2567]), .RECT2_HEIGHT(rectangle2_heights[2567]), .RECT2_WEIGHT(rectangle2_weights[2567]), .RECT3_X(rectangle3_xs[2567]), .RECT3_Y(rectangle3_ys[2567]), .RECT3_WIDTH(rectangle3_widths[2567]), .RECT3_HEIGHT(rectangle3_heights[2567]), .RECT3_WEIGHT(rectangle3_weights[2567]), .FEAT_THRES(feature_thresholds[2567]), .FEAT_ABOVE(feature_aboves[2567]), .FEAT_BELOW(feature_belows[2567])) ac2567(.scan_win(scan_win2567), .scan_win_std_dev(scan_win_std_dev[2567]), .feature_accum(feature_accums[2567]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2568]), .RECT1_Y(rectangle1_ys[2568]), .RECT1_WIDTH(rectangle1_widths[2568]), .RECT1_HEIGHT(rectangle1_heights[2568]), .RECT1_WEIGHT(rectangle1_weights[2568]), .RECT2_X(rectangle2_xs[2568]), .RECT2_Y(rectangle2_ys[2568]), .RECT2_WIDTH(rectangle2_widths[2568]), .RECT2_HEIGHT(rectangle2_heights[2568]), .RECT2_WEIGHT(rectangle2_weights[2568]), .RECT3_X(rectangle3_xs[2568]), .RECT3_Y(rectangle3_ys[2568]), .RECT3_WIDTH(rectangle3_widths[2568]), .RECT3_HEIGHT(rectangle3_heights[2568]), .RECT3_WEIGHT(rectangle3_weights[2568]), .FEAT_THRES(feature_thresholds[2568]), .FEAT_ABOVE(feature_aboves[2568]), .FEAT_BELOW(feature_belows[2568])) ac2568(.scan_win(scan_win2568), .scan_win_std_dev(scan_win_std_dev[2568]), .feature_accum(feature_accums[2568]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2569]), .RECT1_Y(rectangle1_ys[2569]), .RECT1_WIDTH(rectangle1_widths[2569]), .RECT1_HEIGHT(rectangle1_heights[2569]), .RECT1_WEIGHT(rectangle1_weights[2569]), .RECT2_X(rectangle2_xs[2569]), .RECT2_Y(rectangle2_ys[2569]), .RECT2_WIDTH(rectangle2_widths[2569]), .RECT2_HEIGHT(rectangle2_heights[2569]), .RECT2_WEIGHT(rectangle2_weights[2569]), .RECT3_X(rectangle3_xs[2569]), .RECT3_Y(rectangle3_ys[2569]), .RECT3_WIDTH(rectangle3_widths[2569]), .RECT3_HEIGHT(rectangle3_heights[2569]), .RECT3_WEIGHT(rectangle3_weights[2569]), .FEAT_THRES(feature_thresholds[2569]), .FEAT_ABOVE(feature_aboves[2569]), .FEAT_BELOW(feature_belows[2569])) ac2569(.scan_win(scan_win2569), .scan_win_std_dev(scan_win_std_dev[2569]), .feature_accum(feature_accums[2569]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2570]), .RECT1_Y(rectangle1_ys[2570]), .RECT1_WIDTH(rectangle1_widths[2570]), .RECT1_HEIGHT(rectangle1_heights[2570]), .RECT1_WEIGHT(rectangle1_weights[2570]), .RECT2_X(rectangle2_xs[2570]), .RECT2_Y(rectangle2_ys[2570]), .RECT2_WIDTH(rectangle2_widths[2570]), .RECT2_HEIGHT(rectangle2_heights[2570]), .RECT2_WEIGHT(rectangle2_weights[2570]), .RECT3_X(rectangle3_xs[2570]), .RECT3_Y(rectangle3_ys[2570]), .RECT3_WIDTH(rectangle3_widths[2570]), .RECT3_HEIGHT(rectangle3_heights[2570]), .RECT3_WEIGHT(rectangle3_weights[2570]), .FEAT_THRES(feature_thresholds[2570]), .FEAT_ABOVE(feature_aboves[2570]), .FEAT_BELOW(feature_belows[2570])) ac2570(.scan_win(scan_win2570), .scan_win_std_dev(scan_win_std_dev[2570]), .feature_accum(feature_accums[2570]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2571]), .RECT1_Y(rectangle1_ys[2571]), .RECT1_WIDTH(rectangle1_widths[2571]), .RECT1_HEIGHT(rectangle1_heights[2571]), .RECT1_WEIGHT(rectangle1_weights[2571]), .RECT2_X(rectangle2_xs[2571]), .RECT2_Y(rectangle2_ys[2571]), .RECT2_WIDTH(rectangle2_widths[2571]), .RECT2_HEIGHT(rectangle2_heights[2571]), .RECT2_WEIGHT(rectangle2_weights[2571]), .RECT3_X(rectangle3_xs[2571]), .RECT3_Y(rectangle3_ys[2571]), .RECT3_WIDTH(rectangle3_widths[2571]), .RECT3_HEIGHT(rectangle3_heights[2571]), .RECT3_WEIGHT(rectangle3_weights[2571]), .FEAT_THRES(feature_thresholds[2571]), .FEAT_ABOVE(feature_aboves[2571]), .FEAT_BELOW(feature_belows[2571])) ac2571(.scan_win(scan_win2571), .scan_win_std_dev(scan_win_std_dev[2571]), .feature_accum(feature_accums[2571]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2572]), .RECT1_Y(rectangle1_ys[2572]), .RECT1_WIDTH(rectangle1_widths[2572]), .RECT1_HEIGHT(rectangle1_heights[2572]), .RECT1_WEIGHT(rectangle1_weights[2572]), .RECT2_X(rectangle2_xs[2572]), .RECT2_Y(rectangle2_ys[2572]), .RECT2_WIDTH(rectangle2_widths[2572]), .RECT2_HEIGHT(rectangle2_heights[2572]), .RECT2_WEIGHT(rectangle2_weights[2572]), .RECT3_X(rectangle3_xs[2572]), .RECT3_Y(rectangle3_ys[2572]), .RECT3_WIDTH(rectangle3_widths[2572]), .RECT3_HEIGHT(rectangle3_heights[2572]), .RECT3_WEIGHT(rectangle3_weights[2572]), .FEAT_THRES(feature_thresholds[2572]), .FEAT_ABOVE(feature_aboves[2572]), .FEAT_BELOW(feature_belows[2572])) ac2572(.scan_win(scan_win2572), .scan_win_std_dev(scan_win_std_dev[2572]), .feature_accum(feature_accums[2572]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2573]), .RECT1_Y(rectangle1_ys[2573]), .RECT1_WIDTH(rectangle1_widths[2573]), .RECT1_HEIGHT(rectangle1_heights[2573]), .RECT1_WEIGHT(rectangle1_weights[2573]), .RECT2_X(rectangle2_xs[2573]), .RECT2_Y(rectangle2_ys[2573]), .RECT2_WIDTH(rectangle2_widths[2573]), .RECT2_HEIGHT(rectangle2_heights[2573]), .RECT2_WEIGHT(rectangle2_weights[2573]), .RECT3_X(rectangle3_xs[2573]), .RECT3_Y(rectangle3_ys[2573]), .RECT3_WIDTH(rectangle3_widths[2573]), .RECT3_HEIGHT(rectangle3_heights[2573]), .RECT3_WEIGHT(rectangle3_weights[2573]), .FEAT_THRES(feature_thresholds[2573]), .FEAT_ABOVE(feature_aboves[2573]), .FEAT_BELOW(feature_belows[2573])) ac2573(.scan_win(scan_win2573), .scan_win_std_dev(scan_win_std_dev[2573]), .feature_accum(feature_accums[2573]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2574]), .RECT1_Y(rectangle1_ys[2574]), .RECT1_WIDTH(rectangle1_widths[2574]), .RECT1_HEIGHT(rectangle1_heights[2574]), .RECT1_WEIGHT(rectangle1_weights[2574]), .RECT2_X(rectangle2_xs[2574]), .RECT2_Y(rectangle2_ys[2574]), .RECT2_WIDTH(rectangle2_widths[2574]), .RECT2_HEIGHT(rectangle2_heights[2574]), .RECT2_WEIGHT(rectangle2_weights[2574]), .RECT3_X(rectangle3_xs[2574]), .RECT3_Y(rectangle3_ys[2574]), .RECT3_WIDTH(rectangle3_widths[2574]), .RECT3_HEIGHT(rectangle3_heights[2574]), .RECT3_WEIGHT(rectangle3_weights[2574]), .FEAT_THRES(feature_thresholds[2574]), .FEAT_ABOVE(feature_aboves[2574]), .FEAT_BELOW(feature_belows[2574])) ac2574(.scan_win(scan_win2574), .scan_win_std_dev(scan_win_std_dev[2574]), .feature_accum(feature_accums[2574]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2575]), .RECT1_Y(rectangle1_ys[2575]), .RECT1_WIDTH(rectangle1_widths[2575]), .RECT1_HEIGHT(rectangle1_heights[2575]), .RECT1_WEIGHT(rectangle1_weights[2575]), .RECT2_X(rectangle2_xs[2575]), .RECT2_Y(rectangle2_ys[2575]), .RECT2_WIDTH(rectangle2_widths[2575]), .RECT2_HEIGHT(rectangle2_heights[2575]), .RECT2_WEIGHT(rectangle2_weights[2575]), .RECT3_X(rectangle3_xs[2575]), .RECT3_Y(rectangle3_ys[2575]), .RECT3_WIDTH(rectangle3_widths[2575]), .RECT3_HEIGHT(rectangle3_heights[2575]), .RECT3_WEIGHT(rectangle3_weights[2575]), .FEAT_THRES(feature_thresholds[2575]), .FEAT_ABOVE(feature_aboves[2575]), .FEAT_BELOW(feature_belows[2575])) ac2575(.scan_win(scan_win2575), .scan_win_std_dev(scan_win_std_dev[2575]), .feature_accum(feature_accums[2575]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2576]), .RECT1_Y(rectangle1_ys[2576]), .RECT1_WIDTH(rectangle1_widths[2576]), .RECT1_HEIGHT(rectangle1_heights[2576]), .RECT1_WEIGHT(rectangle1_weights[2576]), .RECT2_X(rectangle2_xs[2576]), .RECT2_Y(rectangle2_ys[2576]), .RECT2_WIDTH(rectangle2_widths[2576]), .RECT2_HEIGHT(rectangle2_heights[2576]), .RECT2_WEIGHT(rectangle2_weights[2576]), .RECT3_X(rectangle3_xs[2576]), .RECT3_Y(rectangle3_ys[2576]), .RECT3_WIDTH(rectangle3_widths[2576]), .RECT3_HEIGHT(rectangle3_heights[2576]), .RECT3_WEIGHT(rectangle3_weights[2576]), .FEAT_THRES(feature_thresholds[2576]), .FEAT_ABOVE(feature_aboves[2576]), .FEAT_BELOW(feature_belows[2576])) ac2576(.scan_win(scan_win2576), .scan_win_std_dev(scan_win_std_dev[2576]), .feature_accum(feature_accums[2576]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2577]), .RECT1_Y(rectangle1_ys[2577]), .RECT1_WIDTH(rectangle1_widths[2577]), .RECT1_HEIGHT(rectangle1_heights[2577]), .RECT1_WEIGHT(rectangle1_weights[2577]), .RECT2_X(rectangle2_xs[2577]), .RECT2_Y(rectangle2_ys[2577]), .RECT2_WIDTH(rectangle2_widths[2577]), .RECT2_HEIGHT(rectangle2_heights[2577]), .RECT2_WEIGHT(rectangle2_weights[2577]), .RECT3_X(rectangle3_xs[2577]), .RECT3_Y(rectangle3_ys[2577]), .RECT3_WIDTH(rectangle3_widths[2577]), .RECT3_HEIGHT(rectangle3_heights[2577]), .RECT3_WEIGHT(rectangle3_weights[2577]), .FEAT_THRES(feature_thresholds[2577]), .FEAT_ABOVE(feature_aboves[2577]), .FEAT_BELOW(feature_belows[2577])) ac2577(.scan_win(scan_win2577), .scan_win_std_dev(scan_win_std_dev[2577]), .feature_accum(feature_accums[2577]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2578]), .RECT1_Y(rectangle1_ys[2578]), .RECT1_WIDTH(rectangle1_widths[2578]), .RECT1_HEIGHT(rectangle1_heights[2578]), .RECT1_WEIGHT(rectangle1_weights[2578]), .RECT2_X(rectangle2_xs[2578]), .RECT2_Y(rectangle2_ys[2578]), .RECT2_WIDTH(rectangle2_widths[2578]), .RECT2_HEIGHT(rectangle2_heights[2578]), .RECT2_WEIGHT(rectangle2_weights[2578]), .RECT3_X(rectangle3_xs[2578]), .RECT3_Y(rectangle3_ys[2578]), .RECT3_WIDTH(rectangle3_widths[2578]), .RECT3_HEIGHT(rectangle3_heights[2578]), .RECT3_WEIGHT(rectangle3_weights[2578]), .FEAT_THRES(feature_thresholds[2578]), .FEAT_ABOVE(feature_aboves[2578]), .FEAT_BELOW(feature_belows[2578])) ac2578(.scan_win(scan_win2578), .scan_win_std_dev(scan_win_std_dev[2578]), .feature_accum(feature_accums[2578]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2579]), .RECT1_Y(rectangle1_ys[2579]), .RECT1_WIDTH(rectangle1_widths[2579]), .RECT1_HEIGHT(rectangle1_heights[2579]), .RECT1_WEIGHT(rectangle1_weights[2579]), .RECT2_X(rectangle2_xs[2579]), .RECT2_Y(rectangle2_ys[2579]), .RECT2_WIDTH(rectangle2_widths[2579]), .RECT2_HEIGHT(rectangle2_heights[2579]), .RECT2_WEIGHT(rectangle2_weights[2579]), .RECT3_X(rectangle3_xs[2579]), .RECT3_Y(rectangle3_ys[2579]), .RECT3_WIDTH(rectangle3_widths[2579]), .RECT3_HEIGHT(rectangle3_heights[2579]), .RECT3_WEIGHT(rectangle3_weights[2579]), .FEAT_THRES(feature_thresholds[2579]), .FEAT_ABOVE(feature_aboves[2579]), .FEAT_BELOW(feature_belows[2579])) ac2579(.scan_win(scan_win2579), .scan_win_std_dev(scan_win_std_dev[2579]), .feature_accum(feature_accums[2579]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2580]), .RECT1_Y(rectangle1_ys[2580]), .RECT1_WIDTH(rectangle1_widths[2580]), .RECT1_HEIGHT(rectangle1_heights[2580]), .RECT1_WEIGHT(rectangle1_weights[2580]), .RECT2_X(rectangle2_xs[2580]), .RECT2_Y(rectangle2_ys[2580]), .RECT2_WIDTH(rectangle2_widths[2580]), .RECT2_HEIGHT(rectangle2_heights[2580]), .RECT2_WEIGHT(rectangle2_weights[2580]), .RECT3_X(rectangle3_xs[2580]), .RECT3_Y(rectangle3_ys[2580]), .RECT3_WIDTH(rectangle3_widths[2580]), .RECT3_HEIGHT(rectangle3_heights[2580]), .RECT3_WEIGHT(rectangle3_weights[2580]), .FEAT_THRES(feature_thresholds[2580]), .FEAT_ABOVE(feature_aboves[2580]), .FEAT_BELOW(feature_belows[2580])) ac2580(.scan_win(scan_win2580), .scan_win_std_dev(scan_win_std_dev[2580]), .feature_accum(feature_accums[2580]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2581]), .RECT1_Y(rectangle1_ys[2581]), .RECT1_WIDTH(rectangle1_widths[2581]), .RECT1_HEIGHT(rectangle1_heights[2581]), .RECT1_WEIGHT(rectangle1_weights[2581]), .RECT2_X(rectangle2_xs[2581]), .RECT2_Y(rectangle2_ys[2581]), .RECT2_WIDTH(rectangle2_widths[2581]), .RECT2_HEIGHT(rectangle2_heights[2581]), .RECT2_WEIGHT(rectangle2_weights[2581]), .RECT3_X(rectangle3_xs[2581]), .RECT3_Y(rectangle3_ys[2581]), .RECT3_WIDTH(rectangle3_widths[2581]), .RECT3_HEIGHT(rectangle3_heights[2581]), .RECT3_WEIGHT(rectangle3_weights[2581]), .FEAT_THRES(feature_thresholds[2581]), .FEAT_ABOVE(feature_aboves[2581]), .FEAT_BELOW(feature_belows[2581])) ac2581(.scan_win(scan_win2581), .scan_win_std_dev(scan_win_std_dev[2581]), .feature_accum(feature_accums[2581]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2582]), .RECT1_Y(rectangle1_ys[2582]), .RECT1_WIDTH(rectangle1_widths[2582]), .RECT1_HEIGHT(rectangle1_heights[2582]), .RECT1_WEIGHT(rectangle1_weights[2582]), .RECT2_X(rectangle2_xs[2582]), .RECT2_Y(rectangle2_ys[2582]), .RECT2_WIDTH(rectangle2_widths[2582]), .RECT2_HEIGHT(rectangle2_heights[2582]), .RECT2_WEIGHT(rectangle2_weights[2582]), .RECT3_X(rectangle3_xs[2582]), .RECT3_Y(rectangle3_ys[2582]), .RECT3_WIDTH(rectangle3_widths[2582]), .RECT3_HEIGHT(rectangle3_heights[2582]), .RECT3_WEIGHT(rectangle3_weights[2582]), .FEAT_THRES(feature_thresholds[2582]), .FEAT_ABOVE(feature_aboves[2582]), .FEAT_BELOW(feature_belows[2582])) ac2582(.scan_win(scan_win2582), .scan_win_std_dev(scan_win_std_dev[2582]), .feature_accum(feature_accums[2582]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2583]), .RECT1_Y(rectangle1_ys[2583]), .RECT1_WIDTH(rectangle1_widths[2583]), .RECT1_HEIGHT(rectangle1_heights[2583]), .RECT1_WEIGHT(rectangle1_weights[2583]), .RECT2_X(rectangle2_xs[2583]), .RECT2_Y(rectangle2_ys[2583]), .RECT2_WIDTH(rectangle2_widths[2583]), .RECT2_HEIGHT(rectangle2_heights[2583]), .RECT2_WEIGHT(rectangle2_weights[2583]), .RECT3_X(rectangle3_xs[2583]), .RECT3_Y(rectangle3_ys[2583]), .RECT3_WIDTH(rectangle3_widths[2583]), .RECT3_HEIGHT(rectangle3_heights[2583]), .RECT3_WEIGHT(rectangle3_weights[2583]), .FEAT_THRES(feature_thresholds[2583]), .FEAT_ABOVE(feature_aboves[2583]), .FEAT_BELOW(feature_belows[2583])) ac2583(.scan_win(scan_win2583), .scan_win_std_dev(scan_win_std_dev[2583]), .feature_accum(feature_accums[2583]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2584]), .RECT1_Y(rectangle1_ys[2584]), .RECT1_WIDTH(rectangle1_widths[2584]), .RECT1_HEIGHT(rectangle1_heights[2584]), .RECT1_WEIGHT(rectangle1_weights[2584]), .RECT2_X(rectangle2_xs[2584]), .RECT2_Y(rectangle2_ys[2584]), .RECT2_WIDTH(rectangle2_widths[2584]), .RECT2_HEIGHT(rectangle2_heights[2584]), .RECT2_WEIGHT(rectangle2_weights[2584]), .RECT3_X(rectangle3_xs[2584]), .RECT3_Y(rectangle3_ys[2584]), .RECT3_WIDTH(rectangle3_widths[2584]), .RECT3_HEIGHT(rectangle3_heights[2584]), .RECT3_WEIGHT(rectangle3_weights[2584]), .FEAT_THRES(feature_thresholds[2584]), .FEAT_ABOVE(feature_aboves[2584]), .FEAT_BELOW(feature_belows[2584])) ac2584(.scan_win(scan_win2584), .scan_win_std_dev(scan_win_std_dev[2584]), .feature_accum(feature_accums[2584]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2585]), .RECT1_Y(rectangle1_ys[2585]), .RECT1_WIDTH(rectangle1_widths[2585]), .RECT1_HEIGHT(rectangle1_heights[2585]), .RECT1_WEIGHT(rectangle1_weights[2585]), .RECT2_X(rectangle2_xs[2585]), .RECT2_Y(rectangle2_ys[2585]), .RECT2_WIDTH(rectangle2_widths[2585]), .RECT2_HEIGHT(rectangle2_heights[2585]), .RECT2_WEIGHT(rectangle2_weights[2585]), .RECT3_X(rectangle3_xs[2585]), .RECT3_Y(rectangle3_ys[2585]), .RECT3_WIDTH(rectangle3_widths[2585]), .RECT3_HEIGHT(rectangle3_heights[2585]), .RECT3_WEIGHT(rectangle3_weights[2585]), .FEAT_THRES(feature_thresholds[2585]), .FEAT_ABOVE(feature_aboves[2585]), .FEAT_BELOW(feature_belows[2585])) ac2585(.scan_win(scan_win2585), .scan_win_std_dev(scan_win_std_dev[2585]), .feature_accum(feature_accums[2585]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2586]), .RECT1_Y(rectangle1_ys[2586]), .RECT1_WIDTH(rectangle1_widths[2586]), .RECT1_HEIGHT(rectangle1_heights[2586]), .RECT1_WEIGHT(rectangle1_weights[2586]), .RECT2_X(rectangle2_xs[2586]), .RECT2_Y(rectangle2_ys[2586]), .RECT2_WIDTH(rectangle2_widths[2586]), .RECT2_HEIGHT(rectangle2_heights[2586]), .RECT2_WEIGHT(rectangle2_weights[2586]), .RECT3_X(rectangle3_xs[2586]), .RECT3_Y(rectangle3_ys[2586]), .RECT3_WIDTH(rectangle3_widths[2586]), .RECT3_HEIGHT(rectangle3_heights[2586]), .RECT3_WEIGHT(rectangle3_weights[2586]), .FEAT_THRES(feature_thresholds[2586]), .FEAT_ABOVE(feature_aboves[2586]), .FEAT_BELOW(feature_belows[2586])) ac2586(.scan_win(scan_win2586), .scan_win_std_dev(scan_win_std_dev[2586]), .feature_accum(feature_accums[2586]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2587]), .RECT1_Y(rectangle1_ys[2587]), .RECT1_WIDTH(rectangle1_widths[2587]), .RECT1_HEIGHT(rectangle1_heights[2587]), .RECT1_WEIGHT(rectangle1_weights[2587]), .RECT2_X(rectangle2_xs[2587]), .RECT2_Y(rectangle2_ys[2587]), .RECT2_WIDTH(rectangle2_widths[2587]), .RECT2_HEIGHT(rectangle2_heights[2587]), .RECT2_WEIGHT(rectangle2_weights[2587]), .RECT3_X(rectangle3_xs[2587]), .RECT3_Y(rectangle3_ys[2587]), .RECT3_WIDTH(rectangle3_widths[2587]), .RECT3_HEIGHT(rectangle3_heights[2587]), .RECT3_WEIGHT(rectangle3_weights[2587]), .FEAT_THRES(feature_thresholds[2587]), .FEAT_ABOVE(feature_aboves[2587]), .FEAT_BELOW(feature_belows[2587])) ac2587(.scan_win(scan_win2587), .scan_win_std_dev(scan_win_std_dev[2587]), .feature_accum(feature_accums[2587]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2588]), .RECT1_Y(rectangle1_ys[2588]), .RECT1_WIDTH(rectangle1_widths[2588]), .RECT1_HEIGHT(rectangle1_heights[2588]), .RECT1_WEIGHT(rectangle1_weights[2588]), .RECT2_X(rectangle2_xs[2588]), .RECT2_Y(rectangle2_ys[2588]), .RECT2_WIDTH(rectangle2_widths[2588]), .RECT2_HEIGHT(rectangle2_heights[2588]), .RECT2_WEIGHT(rectangle2_weights[2588]), .RECT3_X(rectangle3_xs[2588]), .RECT3_Y(rectangle3_ys[2588]), .RECT3_WIDTH(rectangle3_widths[2588]), .RECT3_HEIGHT(rectangle3_heights[2588]), .RECT3_WEIGHT(rectangle3_weights[2588]), .FEAT_THRES(feature_thresholds[2588]), .FEAT_ABOVE(feature_aboves[2588]), .FEAT_BELOW(feature_belows[2588])) ac2588(.scan_win(scan_win2588), .scan_win_std_dev(scan_win_std_dev[2588]), .feature_accum(feature_accums[2588]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2589]), .RECT1_Y(rectangle1_ys[2589]), .RECT1_WIDTH(rectangle1_widths[2589]), .RECT1_HEIGHT(rectangle1_heights[2589]), .RECT1_WEIGHT(rectangle1_weights[2589]), .RECT2_X(rectangle2_xs[2589]), .RECT2_Y(rectangle2_ys[2589]), .RECT2_WIDTH(rectangle2_widths[2589]), .RECT2_HEIGHT(rectangle2_heights[2589]), .RECT2_WEIGHT(rectangle2_weights[2589]), .RECT3_X(rectangle3_xs[2589]), .RECT3_Y(rectangle3_ys[2589]), .RECT3_WIDTH(rectangle3_widths[2589]), .RECT3_HEIGHT(rectangle3_heights[2589]), .RECT3_WEIGHT(rectangle3_weights[2589]), .FEAT_THRES(feature_thresholds[2589]), .FEAT_ABOVE(feature_aboves[2589]), .FEAT_BELOW(feature_belows[2589])) ac2589(.scan_win(scan_win2589), .scan_win_std_dev(scan_win_std_dev[2589]), .feature_accum(feature_accums[2589]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2590]), .RECT1_Y(rectangle1_ys[2590]), .RECT1_WIDTH(rectangle1_widths[2590]), .RECT1_HEIGHT(rectangle1_heights[2590]), .RECT1_WEIGHT(rectangle1_weights[2590]), .RECT2_X(rectangle2_xs[2590]), .RECT2_Y(rectangle2_ys[2590]), .RECT2_WIDTH(rectangle2_widths[2590]), .RECT2_HEIGHT(rectangle2_heights[2590]), .RECT2_WEIGHT(rectangle2_weights[2590]), .RECT3_X(rectangle3_xs[2590]), .RECT3_Y(rectangle3_ys[2590]), .RECT3_WIDTH(rectangle3_widths[2590]), .RECT3_HEIGHT(rectangle3_heights[2590]), .RECT3_WEIGHT(rectangle3_weights[2590]), .FEAT_THRES(feature_thresholds[2590]), .FEAT_ABOVE(feature_aboves[2590]), .FEAT_BELOW(feature_belows[2590])) ac2590(.scan_win(scan_win2590), .scan_win_std_dev(scan_win_std_dev[2590]), .feature_accum(feature_accums[2590]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2591]), .RECT1_Y(rectangle1_ys[2591]), .RECT1_WIDTH(rectangle1_widths[2591]), .RECT1_HEIGHT(rectangle1_heights[2591]), .RECT1_WEIGHT(rectangle1_weights[2591]), .RECT2_X(rectangle2_xs[2591]), .RECT2_Y(rectangle2_ys[2591]), .RECT2_WIDTH(rectangle2_widths[2591]), .RECT2_HEIGHT(rectangle2_heights[2591]), .RECT2_WEIGHT(rectangle2_weights[2591]), .RECT3_X(rectangle3_xs[2591]), .RECT3_Y(rectangle3_ys[2591]), .RECT3_WIDTH(rectangle3_widths[2591]), .RECT3_HEIGHT(rectangle3_heights[2591]), .RECT3_WEIGHT(rectangle3_weights[2591]), .FEAT_THRES(feature_thresholds[2591]), .FEAT_ABOVE(feature_aboves[2591]), .FEAT_BELOW(feature_belows[2591])) ac2591(.scan_win(scan_win2591), .scan_win_std_dev(scan_win_std_dev[2591]), .feature_accum(feature_accums[2591]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2592]), .RECT1_Y(rectangle1_ys[2592]), .RECT1_WIDTH(rectangle1_widths[2592]), .RECT1_HEIGHT(rectangle1_heights[2592]), .RECT1_WEIGHT(rectangle1_weights[2592]), .RECT2_X(rectangle2_xs[2592]), .RECT2_Y(rectangle2_ys[2592]), .RECT2_WIDTH(rectangle2_widths[2592]), .RECT2_HEIGHT(rectangle2_heights[2592]), .RECT2_WEIGHT(rectangle2_weights[2592]), .RECT3_X(rectangle3_xs[2592]), .RECT3_Y(rectangle3_ys[2592]), .RECT3_WIDTH(rectangle3_widths[2592]), .RECT3_HEIGHT(rectangle3_heights[2592]), .RECT3_WEIGHT(rectangle3_weights[2592]), .FEAT_THRES(feature_thresholds[2592]), .FEAT_ABOVE(feature_aboves[2592]), .FEAT_BELOW(feature_belows[2592])) ac2592(.scan_win(scan_win2592), .scan_win_std_dev(scan_win_std_dev[2592]), .feature_accum(feature_accums[2592]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2593]), .RECT1_Y(rectangle1_ys[2593]), .RECT1_WIDTH(rectangle1_widths[2593]), .RECT1_HEIGHT(rectangle1_heights[2593]), .RECT1_WEIGHT(rectangle1_weights[2593]), .RECT2_X(rectangle2_xs[2593]), .RECT2_Y(rectangle2_ys[2593]), .RECT2_WIDTH(rectangle2_widths[2593]), .RECT2_HEIGHT(rectangle2_heights[2593]), .RECT2_WEIGHT(rectangle2_weights[2593]), .RECT3_X(rectangle3_xs[2593]), .RECT3_Y(rectangle3_ys[2593]), .RECT3_WIDTH(rectangle3_widths[2593]), .RECT3_HEIGHT(rectangle3_heights[2593]), .RECT3_WEIGHT(rectangle3_weights[2593]), .FEAT_THRES(feature_thresholds[2593]), .FEAT_ABOVE(feature_aboves[2593]), .FEAT_BELOW(feature_belows[2593])) ac2593(.scan_win(scan_win2593), .scan_win_std_dev(scan_win_std_dev[2593]), .feature_accum(feature_accums[2593]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2594]), .RECT1_Y(rectangle1_ys[2594]), .RECT1_WIDTH(rectangle1_widths[2594]), .RECT1_HEIGHT(rectangle1_heights[2594]), .RECT1_WEIGHT(rectangle1_weights[2594]), .RECT2_X(rectangle2_xs[2594]), .RECT2_Y(rectangle2_ys[2594]), .RECT2_WIDTH(rectangle2_widths[2594]), .RECT2_HEIGHT(rectangle2_heights[2594]), .RECT2_WEIGHT(rectangle2_weights[2594]), .RECT3_X(rectangle3_xs[2594]), .RECT3_Y(rectangle3_ys[2594]), .RECT3_WIDTH(rectangle3_widths[2594]), .RECT3_HEIGHT(rectangle3_heights[2594]), .RECT3_WEIGHT(rectangle3_weights[2594]), .FEAT_THRES(feature_thresholds[2594]), .FEAT_ABOVE(feature_aboves[2594]), .FEAT_BELOW(feature_belows[2594])) ac2594(.scan_win(scan_win2594), .scan_win_std_dev(scan_win_std_dev[2594]), .feature_accum(feature_accums[2594]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2595]), .RECT1_Y(rectangle1_ys[2595]), .RECT1_WIDTH(rectangle1_widths[2595]), .RECT1_HEIGHT(rectangle1_heights[2595]), .RECT1_WEIGHT(rectangle1_weights[2595]), .RECT2_X(rectangle2_xs[2595]), .RECT2_Y(rectangle2_ys[2595]), .RECT2_WIDTH(rectangle2_widths[2595]), .RECT2_HEIGHT(rectangle2_heights[2595]), .RECT2_WEIGHT(rectangle2_weights[2595]), .RECT3_X(rectangle3_xs[2595]), .RECT3_Y(rectangle3_ys[2595]), .RECT3_WIDTH(rectangle3_widths[2595]), .RECT3_HEIGHT(rectangle3_heights[2595]), .RECT3_WEIGHT(rectangle3_weights[2595]), .FEAT_THRES(feature_thresholds[2595]), .FEAT_ABOVE(feature_aboves[2595]), .FEAT_BELOW(feature_belows[2595])) ac2595(.scan_win(scan_win2595), .scan_win_std_dev(scan_win_std_dev[2595]), .feature_accum(feature_accums[2595]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2596]), .RECT1_Y(rectangle1_ys[2596]), .RECT1_WIDTH(rectangle1_widths[2596]), .RECT1_HEIGHT(rectangle1_heights[2596]), .RECT1_WEIGHT(rectangle1_weights[2596]), .RECT2_X(rectangle2_xs[2596]), .RECT2_Y(rectangle2_ys[2596]), .RECT2_WIDTH(rectangle2_widths[2596]), .RECT2_HEIGHT(rectangle2_heights[2596]), .RECT2_WEIGHT(rectangle2_weights[2596]), .RECT3_X(rectangle3_xs[2596]), .RECT3_Y(rectangle3_ys[2596]), .RECT3_WIDTH(rectangle3_widths[2596]), .RECT3_HEIGHT(rectangle3_heights[2596]), .RECT3_WEIGHT(rectangle3_weights[2596]), .FEAT_THRES(feature_thresholds[2596]), .FEAT_ABOVE(feature_aboves[2596]), .FEAT_BELOW(feature_belows[2596])) ac2596(.scan_win(scan_win2596), .scan_win_std_dev(scan_win_std_dev[2596]), .feature_accum(feature_accums[2596]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2597]), .RECT1_Y(rectangle1_ys[2597]), .RECT1_WIDTH(rectangle1_widths[2597]), .RECT1_HEIGHT(rectangle1_heights[2597]), .RECT1_WEIGHT(rectangle1_weights[2597]), .RECT2_X(rectangle2_xs[2597]), .RECT2_Y(rectangle2_ys[2597]), .RECT2_WIDTH(rectangle2_widths[2597]), .RECT2_HEIGHT(rectangle2_heights[2597]), .RECT2_WEIGHT(rectangle2_weights[2597]), .RECT3_X(rectangle3_xs[2597]), .RECT3_Y(rectangle3_ys[2597]), .RECT3_WIDTH(rectangle3_widths[2597]), .RECT3_HEIGHT(rectangle3_heights[2597]), .RECT3_WEIGHT(rectangle3_weights[2597]), .FEAT_THRES(feature_thresholds[2597]), .FEAT_ABOVE(feature_aboves[2597]), .FEAT_BELOW(feature_belows[2597])) ac2597(.scan_win(scan_win2597), .scan_win_std_dev(scan_win_std_dev[2597]), .feature_accum(feature_accums[2597]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2598]), .RECT1_Y(rectangle1_ys[2598]), .RECT1_WIDTH(rectangle1_widths[2598]), .RECT1_HEIGHT(rectangle1_heights[2598]), .RECT1_WEIGHT(rectangle1_weights[2598]), .RECT2_X(rectangle2_xs[2598]), .RECT2_Y(rectangle2_ys[2598]), .RECT2_WIDTH(rectangle2_widths[2598]), .RECT2_HEIGHT(rectangle2_heights[2598]), .RECT2_WEIGHT(rectangle2_weights[2598]), .RECT3_X(rectangle3_xs[2598]), .RECT3_Y(rectangle3_ys[2598]), .RECT3_WIDTH(rectangle3_widths[2598]), .RECT3_HEIGHT(rectangle3_heights[2598]), .RECT3_WEIGHT(rectangle3_weights[2598]), .FEAT_THRES(feature_thresholds[2598]), .FEAT_ABOVE(feature_aboves[2598]), .FEAT_BELOW(feature_belows[2598])) ac2598(.scan_win(scan_win2598), .scan_win_std_dev(scan_win_std_dev[2598]), .feature_accum(feature_accums[2598]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2599]), .RECT1_Y(rectangle1_ys[2599]), .RECT1_WIDTH(rectangle1_widths[2599]), .RECT1_HEIGHT(rectangle1_heights[2599]), .RECT1_WEIGHT(rectangle1_weights[2599]), .RECT2_X(rectangle2_xs[2599]), .RECT2_Y(rectangle2_ys[2599]), .RECT2_WIDTH(rectangle2_widths[2599]), .RECT2_HEIGHT(rectangle2_heights[2599]), .RECT2_WEIGHT(rectangle2_weights[2599]), .RECT3_X(rectangle3_xs[2599]), .RECT3_Y(rectangle3_ys[2599]), .RECT3_WIDTH(rectangle3_widths[2599]), .RECT3_HEIGHT(rectangle3_heights[2599]), .RECT3_WEIGHT(rectangle3_weights[2599]), .FEAT_THRES(feature_thresholds[2599]), .FEAT_ABOVE(feature_aboves[2599]), .FEAT_BELOW(feature_belows[2599])) ac2599(.scan_win(scan_win2599), .scan_win_std_dev(scan_win_std_dev[2599]), .feature_accum(feature_accums[2599]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2600]), .RECT1_Y(rectangle1_ys[2600]), .RECT1_WIDTH(rectangle1_widths[2600]), .RECT1_HEIGHT(rectangle1_heights[2600]), .RECT1_WEIGHT(rectangle1_weights[2600]), .RECT2_X(rectangle2_xs[2600]), .RECT2_Y(rectangle2_ys[2600]), .RECT2_WIDTH(rectangle2_widths[2600]), .RECT2_HEIGHT(rectangle2_heights[2600]), .RECT2_WEIGHT(rectangle2_weights[2600]), .RECT3_X(rectangle3_xs[2600]), .RECT3_Y(rectangle3_ys[2600]), .RECT3_WIDTH(rectangle3_widths[2600]), .RECT3_HEIGHT(rectangle3_heights[2600]), .RECT3_WEIGHT(rectangle3_weights[2600]), .FEAT_THRES(feature_thresholds[2600]), .FEAT_ABOVE(feature_aboves[2600]), .FEAT_BELOW(feature_belows[2600])) ac2600(.scan_win(scan_win2600), .scan_win_std_dev(scan_win_std_dev[2600]), .feature_accum(feature_accums[2600]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2601]), .RECT1_Y(rectangle1_ys[2601]), .RECT1_WIDTH(rectangle1_widths[2601]), .RECT1_HEIGHT(rectangle1_heights[2601]), .RECT1_WEIGHT(rectangle1_weights[2601]), .RECT2_X(rectangle2_xs[2601]), .RECT2_Y(rectangle2_ys[2601]), .RECT2_WIDTH(rectangle2_widths[2601]), .RECT2_HEIGHT(rectangle2_heights[2601]), .RECT2_WEIGHT(rectangle2_weights[2601]), .RECT3_X(rectangle3_xs[2601]), .RECT3_Y(rectangle3_ys[2601]), .RECT3_WIDTH(rectangle3_widths[2601]), .RECT3_HEIGHT(rectangle3_heights[2601]), .RECT3_WEIGHT(rectangle3_weights[2601]), .FEAT_THRES(feature_thresholds[2601]), .FEAT_ABOVE(feature_aboves[2601]), .FEAT_BELOW(feature_belows[2601])) ac2601(.scan_win(scan_win2601), .scan_win_std_dev(scan_win_std_dev[2601]), .feature_accum(feature_accums[2601]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2602]), .RECT1_Y(rectangle1_ys[2602]), .RECT1_WIDTH(rectangle1_widths[2602]), .RECT1_HEIGHT(rectangle1_heights[2602]), .RECT1_WEIGHT(rectangle1_weights[2602]), .RECT2_X(rectangle2_xs[2602]), .RECT2_Y(rectangle2_ys[2602]), .RECT2_WIDTH(rectangle2_widths[2602]), .RECT2_HEIGHT(rectangle2_heights[2602]), .RECT2_WEIGHT(rectangle2_weights[2602]), .RECT3_X(rectangle3_xs[2602]), .RECT3_Y(rectangle3_ys[2602]), .RECT3_WIDTH(rectangle3_widths[2602]), .RECT3_HEIGHT(rectangle3_heights[2602]), .RECT3_WEIGHT(rectangle3_weights[2602]), .FEAT_THRES(feature_thresholds[2602]), .FEAT_ABOVE(feature_aboves[2602]), .FEAT_BELOW(feature_belows[2602])) ac2602(.scan_win(scan_win2602), .scan_win_std_dev(scan_win_std_dev[2602]), .feature_accum(feature_accums[2602]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2603]), .RECT1_Y(rectangle1_ys[2603]), .RECT1_WIDTH(rectangle1_widths[2603]), .RECT1_HEIGHT(rectangle1_heights[2603]), .RECT1_WEIGHT(rectangle1_weights[2603]), .RECT2_X(rectangle2_xs[2603]), .RECT2_Y(rectangle2_ys[2603]), .RECT2_WIDTH(rectangle2_widths[2603]), .RECT2_HEIGHT(rectangle2_heights[2603]), .RECT2_WEIGHT(rectangle2_weights[2603]), .RECT3_X(rectangle3_xs[2603]), .RECT3_Y(rectangle3_ys[2603]), .RECT3_WIDTH(rectangle3_widths[2603]), .RECT3_HEIGHT(rectangle3_heights[2603]), .RECT3_WEIGHT(rectangle3_weights[2603]), .FEAT_THRES(feature_thresholds[2603]), .FEAT_ABOVE(feature_aboves[2603]), .FEAT_BELOW(feature_belows[2603])) ac2603(.scan_win(scan_win2603), .scan_win_std_dev(scan_win_std_dev[2603]), .feature_accum(feature_accums[2603]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2604]), .RECT1_Y(rectangle1_ys[2604]), .RECT1_WIDTH(rectangle1_widths[2604]), .RECT1_HEIGHT(rectangle1_heights[2604]), .RECT1_WEIGHT(rectangle1_weights[2604]), .RECT2_X(rectangle2_xs[2604]), .RECT2_Y(rectangle2_ys[2604]), .RECT2_WIDTH(rectangle2_widths[2604]), .RECT2_HEIGHT(rectangle2_heights[2604]), .RECT2_WEIGHT(rectangle2_weights[2604]), .RECT3_X(rectangle3_xs[2604]), .RECT3_Y(rectangle3_ys[2604]), .RECT3_WIDTH(rectangle3_widths[2604]), .RECT3_HEIGHT(rectangle3_heights[2604]), .RECT3_WEIGHT(rectangle3_weights[2604]), .FEAT_THRES(feature_thresholds[2604]), .FEAT_ABOVE(feature_aboves[2604]), .FEAT_BELOW(feature_belows[2604])) ac2604(.scan_win(scan_win2604), .scan_win_std_dev(scan_win_std_dev[2604]), .feature_accum(feature_accums[2604]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2605]), .RECT1_Y(rectangle1_ys[2605]), .RECT1_WIDTH(rectangle1_widths[2605]), .RECT1_HEIGHT(rectangle1_heights[2605]), .RECT1_WEIGHT(rectangle1_weights[2605]), .RECT2_X(rectangle2_xs[2605]), .RECT2_Y(rectangle2_ys[2605]), .RECT2_WIDTH(rectangle2_widths[2605]), .RECT2_HEIGHT(rectangle2_heights[2605]), .RECT2_WEIGHT(rectangle2_weights[2605]), .RECT3_X(rectangle3_xs[2605]), .RECT3_Y(rectangle3_ys[2605]), .RECT3_WIDTH(rectangle3_widths[2605]), .RECT3_HEIGHT(rectangle3_heights[2605]), .RECT3_WEIGHT(rectangle3_weights[2605]), .FEAT_THRES(feature_thresholds[2605]), .FEAT_ABOVE(feature_aboves[2605]), .FEAT_BELOW(feature_belows[2605])) ac2605(.scan_win(scan_win2605), .scan_win_std_dev(scan_win_std_dev[2605]), .feature_accum(feature_accums[2605]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2606]), .RECT1_Y(rectangle1_ys[2606]), .RECT1_WIDTH(rectangle1_widths[2606]), .RECT1_HEIGHT(rectangle1_heights[2606]), .RECT1_WEIGHT(rectangle1_weights[2606]), .RECT2_X(rectangle2_xs[2606]), .RECT2_Y(rectangle2_ys[2606]), .RECT2_WIDTH(rectangle2_widths[2606]), .RECT2_HEIGHT(rectangle2_heights[2606]), .RECT2_WEIGHT(rectangle2_weights[2606]), .RECT3_X(rectangle3_xs[2606]), .RECT3_Y(rectangle3_ys[2606]), .RECT3_WIDTH(rectangle3_widths[2606]), .RECT3_HEIGHT(rectangle3_heights[2606]), .RECT3_WEIGHT(rectangle3_weights[2606]), .FEAT_THRES(feature_thresholds[2606]), .FEAT_ABOVE(feature_aboves[2606]), .FEAT_BELOW(feature_belows[2606])) ac2606(.scan_win(scan_win2606), .scan_win_std_dev(scan_win_std_dev[2606]), .feature_accum(feature_accums[2606]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2607]), .RECT1_Y(rectangle1_ys[2607]), .RECT1_WIDTH(rectangle1_widths[2607]), .RECT1_HEIGHT(rectangle1_heights[2607]), .RECT1_WEIGHT(rectangle1_weights[2607]), .RECT2_X(rectangle2_xs[2607]), .RECT2_Y(rectangle2_ys[2607]), .RECT2_WIDTH(rectangle2_widths[2607]), .RECT2_HEIGHT(rectangle2_heights[2607]), .RECT2_WEIGHT(rectangle2_weights[2607]), .RECT3_X(rectangle3_xs[2607]), .RECT3_Y(rectangle3_ys[2607]), .RECT3_WIDTH(rectangle3_widths[2607]), .RECT3_HEIGHT(rectangle3_heights[2607]), .RECT3_WEIGHT(rectangle3_weights[2607]), .FEAT_THRES(feature_thresholds[2607]), .FEAT_ABOVE(feature_aboves[2607]), .FEAT_BELOW(feature_belows[2607])) ac2607(.scan_win(scan_win2607), .scan_win_std_dev(scan_win_std_dev[2607]), .feature_accum(feature_accums[2607]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2608]), .RECT1_Y(rectangle1_ys[2608]), .RECT1_WIDTH(rectangle1_widths[2608]), .RECT1_HEIGHT(rectangle1_heights[2608]), .RECT1_WEIGHT(rectangle1_weights[2608]), .RECT2_X(rectangle2_xs[2608]), .RECT2_Y(rectangle2_ys[2608]), .RECT2_WIDTH(rectangle2_widths[2608]), .RECT2_HEIGHT(rectangle2_heights[2608]), .RECT2_WEIGHT(rectangle2_weights[2608]), .RECT3_X(rectangle3_xs[2608]), .RECT3_Y(rectangle3_ys[2608]), .RECT3_WIDTH(rectangle3_widths[2608]), .RECT3_HEIGHT(rectangle3_heights[2608]), .RECT3_WEIGHT(rectangle3_weights[2608]), .FEAT_THRES(feature_thresholds[2608]), .FEAT_ABOVE(feature_aboves[2608]), .FEAT_BELOW(feature_belows[2608])) ac2608(.scan_win(scan_win2608), .scan_win_std_dev(scan_win_std_dev[2608]), .feature_accum(feature_accums[2608]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2609]), .RECT1_Y(rectangle1_ys[2609]), .RECT1_WIDTH(rectangle1_widths[2609]), .RECT1_HEIGHT(rectangle1_heights[2609]), .RECT1_WEIGHT(rectangle1_weights[2609]), .RECT2_X(rectangle2_xs[2609]), .RECT2_Y(rectangle2_ys[2609]), .RECT2_WIDTH(rectangle2_widths[2609]), .RECT2_HEIGHT(rectangle2_heights[2609]), .RECT2_WEIGHT(rectangle2_weights[2609]), .RECT3_X(rectangle3_xs[2609]), .RECT3_Y(rectangle3_ys[2609]), .RECT3_WIDTH(rectangle3_widths[2609]), .RECT3_HEIGHT(rectangle3_heights[2609]), .RECT3_WEIGHT(rectangle3_weights[2609]), .FEAT_THRES(feature_thresholds[2609]), .FEAT_ABOVE(feature_aboves[2609]), .FEAT_BELOW(feature_belows[2609])) ac2609(.scan_win(scan_win2609), .scan_win_std_dev(scan_win_std_dev[2609]), .feature_accum(feature_accums[2609]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2610]), .RECT1_Y(rectangle1_ys[2610]), .RECT1_WIDTH(rectangle1_widths[2610]), .RECT1_HEIGHT(rectangle1_heights[2610]), .RECT1_WEIGHT(rectangle1_weights[2610]), .RECT2_X(rectangle2_xs[2610]), .RECT2_Y(rectangle2_ys[2610]), .RECT2_WIDTH(rectangle2_widths[2610]), .RECT2_HEIGHT(rectangle2_heights[2610]), .RECT2_WEIGHT(rectangle2_weights[2610]), .RECT3_X(rectangle3_xs[2610]), .RECT3_Y(rectangle3_ys[2610]), .RECT3_WIDTH(rectangle3_widths[2610]), .RECT3_HEIGHT(rectangle3_heights[2610]), .RECT3_WEIGHT(rectangle3_weights[2610]), .FEAT_THRES(feature_thresholds[2610]), .FEAT_ABOVE(feature_aboves[2610]), .FEAT_BELOW(feature_belows[2610])) ac2610(.scan_win(scan_win2610), .scan_win_std_dev(scan_win_std_dev[2610]), .feature_accum(feature_accums[2610]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2611]), .RECT1_Y(rectangle1_ys[2611]), .RECT1_WIDTH(rectangle1_widths[2611]), .RECT1_HEIGHT(rectangle1_heights[2611]), .RECT1_WEIGHT(rectangle1_weights[2611]), .RECT2_X(rectangle2_xs[2611]), .RECT2_Y(rectangle2_ys[2611]), .RECT2_WIDTH(rectangle2_widths[2611]), .RECT2_HEIGHT(rectangle2_heights[2611]), .RECT2_WEIGHT(rectangle2_weights[2611]), .RECT3_X(rectangle3_xs[2611]), .RECT3_Y(rectangle3_ys[2611]), .RECT3_WIDTH(rectangle3_widths[2611]), .RECT3_HEIGHT(rectangle3_heights[2611]), .RECT3_WEIGHT(rectangle3_weights[2611]), .FEAT_THRES(feature_thresholds[2611]), .FEAT_ABOVE(feature_aboves[2611]), .FEAT_BELOW(feature_belows[2611])) ac2611(.scan_win(scan_win2611), .scan_win_std_dev(scan_win_std_dev[2611]), .feature_accum(feature_accums[2611]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2612]), .RECT1_Y(rectangle1_ys[2612]), .RECT1_WIDTH(rectangle1_widths[2612]), .RECT1_HEIGHT(rectangle1_heights[2612]), .RECT1_WEIGHT(rectangle1_weights[2612]), .RECT2_X(rectangle2_xs[2612]), .RECT2_Y(rectangle2_ys[2612]), .RECT2_WIDTH(rectangle2_widths[2612]), .RECT2_HEIGHT(rectangle2_heights[2612]), .RECT2_WEIGHT(rectangle2_weights[2612]), .RECT3_X(rectangle3_xs[2612]), .RECT3_Y(rectangle3_ys[2612]), .RECT3_WIDTH(rectangle3_widths[2612]), .RECT3_HEIGHT(rectangle3_heights[2612]), .RECT3_WEIGHT(rectangle3_weights[2612]), .FEAT_THRES(feature_thresholds[2612]), .FEAT_ABOVE(feature_aboves[2612]), .FEAT_BELOW(feature_belows[2612])) ac2612(.scan_win(scan_win2612), .scan_win_std_dev(scan_win_std_dev[2612]), .feature_accum(feature_accums[2612]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2613]), .RECT1_Y(rectangle1_ys[2613]), .RECT1_WIDTH(rectangle1_widths[2613]), .RECT1_HEIGHT(rectangle1_heights[2613]), .RECT1_WEIGHT(rectangle1_weights[2613]), .RECT2_X(rectangle2_xs[2613]), .RECT2_Y(rectangle2_ys[2613]), .RECT2_WIDTH(rectangle2_widths[2613]), .RECT2_HEIGHT(rectangle2_heights[2613]), .RECT2_WEIGHT(rectangle2_weights[2613]), .RECT3_X(rectangle3_xs[2613]), .RECT3_Y(rectangle3_ys[2613]), .RECT3_WIDTH(rectangle3_widths[2613]), .RECT3_HEIGHT(rectangle3_heights[2613]), .RECT3_WEIGHT(rectangle3_weights[2613]), .FEAT_THRES(feature_thresholds[2613]), .FEAT_ABOVE(feature_aboves[2613]), .FEAT_BELOW(feature_belows[2613])) ac2613(.scan_win(scan_win2613), .scan_win_std_dev(scan_win_std_dev[2613]), .feature_accum(feature_accums[2613]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2614]), .RECT1_Y(rectangle1_ys[2614]), .RECT1_WIDTH(rectangle1_widths[2614]), .RECT1_HEIGHT(rectangle1_heights[2614]), .RECT1_WEIGHT(rectangle1_weights[2614]), .RECT2_X(rectangle2_xs[2614]), .RECT2_Y(rectangle2_ys[2614]), .RECT2_WIDTH(rectangle2_widths[2614]), .RECT2_HEIGHT(rectangle2_heights[2614]), .RECT2_WEIGHT(rectangle2_weights[2614]), .RECT3_X(rectangle3_xs[2614]), .RECT3_Y(rectangle3_ys[2614]), .RECT3_WIDTH(rectangle3_widths[2614]), .RECT3_HEIGHT(rectangle3_heights[2614]), .RECT3_WEIGHT(rectangle3_weights[2614]), .FEAT_THRES(feature_thresholds[2614]), .FEAT_ABOVE(feature_aboves[2614]), .FEAT_BELOW(feature_belows[2614])) ac2614(.scan_win(scan_win2614), .scan_win_std_dev(scan_win_std_dev[2614]), .feature_accum(feature_accums[2614]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2615]), .RECT1_Y(rectangle1_ys[2615]), .RECT1_WIDTH(rectangle1_widths[2615]), .RECT1_HEIGHT(rectangle1_heights[2615]), .RECT1_WEIGHT(rectangle1_weights[2615]), .RECT2_X(rectangle2_xs[2615]), .RECT2_Y(rectangle2_ys[2615]), .RECT2_WIDTH(rectangle2_widths[2615]), .RECT2_HEIGHT(rectangle2_heights[2615]), .RECT2_WEIGHT(rectangle2_weights[2615]), .RECT3_X(rectangle3_xs[2615]), .RECT3_Y(rectangle3_ys[2615]), .RECT3_WIDTH(rectangle3_widths[2615]), .RECT3_HEIGHT(rectangle3_heights[2615]), .RECT3_WEIGHT(rectangle3_weights[2615]), .FEAT_THRES(feature_thresholds[2615]), .FEAT_ABOVE(feature_aboves[2615]), .FEAT_BELOW(feature_belows[2615])) ac2615(.scan_win(scan_win2615), .scan_win_std_dev(scan_win_std_dev[2615]), .feature_accum(feature_accums[2615]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2616]), .RECT1_Y(rectangle1_ys[2616]), .RECT1_WIDTH(rectangle1_widths[2616]), .RECT1_HEIGHT(rectangle1_heights[2616]), .RECT1_WEIGHT(rectangle1_weights[2616]), .RECT2_X(rectangle2_xs[2616]), .RECT2_Y(rectangle2_ys[2616]), .RECT2_WIDTH(rectangle2_widths[2616]), .RECT2_HEIGHT(rectangle2_heights[2616]), .RECT2_WEIGHT(rectangle2_weights[2616]), .RECT3_X(rectangle3_xs[2616]), .RECT3_Y(rectangle3_ys[2616]), .RECT3_WIDTH(rectangle3_widths[2616]), .RECT3_HEIGHT(rectangle3_heights[2616]), .RECT3_WEIGHT(rectangle3_weights[2616]), .FEAT_THRES(feature_thresholds[2616]), .FEAT_ABOVE(feature_aboves[2616]), .FEAT_BELOW(feature_belows[2616])) ac2616(.scan_win(scan_win2616), .scan_win_std_dev(scan_win_std_dev[2616]), .feature_accum(feature_accums[2616]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2617]), .RECT1_Y(rectangle1_ys[2617]), .RECT1_WIDTH(rectangle1_widths[2617]), .RECT1_HEIGHT(rectangle1_heights[2617]), .RECT1_WEIGHT(rectangle1_weights[2617]), .RECT2_X(rectangle2_xs[2617]), .RECT2_Y(rectangle2_ys[2617]), .RECT2_WIDTH(rectangle2_widths[2617]), .RECT2_HEIGHT(rectangle2_heights[2617]), .RECT2_WEIGHT(rectangle2_weights[2617]), .RECT3_X(rectangle3_xs[2617]), .RECT3_Y(rectangle3_ys[2617]), .RECT3_WIDTH(rectangle3_widths[2617]), .RECT3_HEIGHT(rectangle3_heights[2617]), .RECT3_WEIGHT(rectangle3_weights[2617]), .FEAT_THRES(feature_thresholds[2617]), .FEAT_ABOVE(feature_aboves[2617]), .FEAT_BELOW(feature_belows[2617])) ac2617(.scan_win(scan_win2617), .scan_win_std_dev(scan_win_std_dev[2617]), .feature_accum(feature_accums[2617]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2618]), .RECT1_Y(rectangle1_ys[2618]), .RECT1_WIDTH(rectangle1_widths[2618]), .RECT1_HEIGHT(rectangle1_heights[2618]), .RECT1_WEIGHT(rectangle1_weights[2618]), .RECT2_X(rectangle2_xs[2618]), .RECT2_Y(rectangle2_ys[2618]), .RECT2_WIDTH(rectangle2_widths[2618]), .RECT2_HEIGHT(rectangle2_heights[2618]), .RECT2_WEIGHT(rectangle2_weights[2618]), .RECT3_X(rectangle3_xs[2618]), .RECT3_Y(rectangle3_ys[2618]), .RECT3_WIDTH(rectangle3_widths[2618]), .RECT3_HEIGHT(rectangle3_heights[2618]), .RECT3_WEIGHT(rectangle3_weights[2618]), .FEAT_THRES(feature_thresholds[2618]), .FEAT_ABOVE(feature_aboves[2618]), .FEAT_BELOW(feature_belows[2618])) ac2618(.scan_win(scan_win2618), .scan_win_std_dev(scan_win_std_dev[2618]), .feature_accum(feature_accums[2618]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2619]), .RECT1_Y(rectangle1_ys[2619]), .RECT1_WIDTH(rectangle1_widths[2619]), .RECT1_HEIGHT(rectangle1_heights[2619]), .RECT1_WEIGHT(rectangle1_weights[2619]), .RECT2_X(rectangle2_xs[2619]), .RECT2_Y(rectangle2_ys[2619]), .RECT2_WIDTH(rectangle2_widths[2619]), .RECT2_HEIGHT(rectangle2_heights[2619]), .RECT2_WEIGHT(rectangle2_weights[2619]), .RECT3_X(rectangle3_xs[2619]), .RECT3_Y(rectangle3_ys[2619]), .RECT3_WIDTH(rectangle3_widths[2619]), .RECT3_HEIGHT(rectangle3_heights[2619]), .RECT3_WEIGHT(rectangle3_weights[2619]), .FEAT_THRES(feature_thresholds[2619]), .FEAT_ABOVE(feature_aboves[2619]), .FEAT_BELOW(feature_belows[2619])) ac2619(.scan_win(scan_win2619), .scan_win_std_dev(scan_win_std_dev[2619]), .feature_accum(feature_accums[2619]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2620]), .RECT1_Y(rectangle1_ys[2620]), .RECT1_WIDTH(rectangle1_widths[2620]), .RECT1_HEIGHT(rectangle1_heights[2620]), .RECT1_WEIGHT(rectangle1_weights[2620]), .RECT2_X(rectangle2_xs[2620]), .RECT2_Y(rectangle2_ys[2620]), .RECT2_WIDTH(rectangle2_widths[2620]), .RECT2_HEIGHT(rectangle2_heights[2620]), .RECT2_WEIGHT(rectangle2_weights[2620]), .RECT3_X(rectangle3_xs[2620]), .RECT3_Y(rectangle3_ys[2620]), .RECT3_WIDTH(rectangle3_widths[2620]), .RECT3_HEIGHT(rectangle3_heights[2620]), .RECT3_WEIGHT(rectangle3_weights[2620]), .FEAT_THRES(feature_thresholds[2620]), .FEAT_ABOVE(feature_aboves[2620]), .FEAT_BELOW(feature_belows[2620])) ac2620(.scan_win(scan_win2620), .scan_win_std_dev(scan_win_std_dev[2620]), .feature_accum(feature_accums[2620]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2621]), .RECT1_Y(rectangle1_ys[2621]), .RECT1_WIDTH(rectangle1_widths[2621]), .RECT1_HEIGHT(rectangle1_heights[2621]), .RECT1_WEIGHT(rectangle1_weights[2621]), .RECT2_X(rectangle2_xs[2621]), .RECT2_Y(rectangle2_ys[2621]), .RECT2_WIDTH(rectangle2_widths[2621]), .RECT2_HEIGHT(rectangle2_heights[2621]), .RECT2_WEIGHT(rectangle2_weights[2621]), .RECT3_X(rectangle3_xs[2621]), .RECT3_Y(rectangle3_ys[2621]), .RECT3_WIDTH(rectangle3_widths[2621]), .RECT3_HEIGHT(rectangle3_heights[2621]), .RECT3_WEIGHT(rectangle3_weights[2621]), .FEAT_THRES(feature_thresholds[2621]), .FEAT_ABOVE(feature_aboves[2621]), .FEAT_BELOW(feature_belows[2621])) ac2621(.scan_win(scan_win2621), .scan_win_std_dev(scan_win_std_dev[2621]), .feature_accum(feature_accums[2621]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2622]), .RECT1_Y(rectangle1_ys[2622]), .RECT1_WIDTH(rectangle1_widths[2622]), .RECT1_HEIGHT(rectangle1_heights[2622]), .RECT1_WEIGHT(rectangle1_weights[2622]), .RECT2_X(rectangle2_xs[2622]), .RECT2_Y(rectangle2_ys[2622]), .RECT2_WIDTH(rectangle2_widths[2622]), .RECT2_HEIGHT(rectangle2_heights[2622]), .RECT2_WEIGHT(rectangle2_weights[2622]), .RECT3_X(rectangle3_xs[2622]), .RECT3_Y(rectangle3_ys[2622]), .RECT3_WIDTH(rectangle3_widths[2622]), .RECT3_HEIGHT(rectangle3_heights[2622]), .RECT3_WEIGHT(rectangle3_weights[2622]), .FEAT_THRES(feature_thresholds[2622]), .FEAT_ABOVE(feature_aboves[2622]), .FEAT_BELOW(feature_belows[2622])) ac2622(.scan_win(scan_win2622), .scan_win_std_dev(scan_win_std_dev[2622]), .feature_accum(feature_accums[2622]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2623]), .RECT1_Y(rectangle1_ys[2623]), .RECT1_WIDTH(rectangle1_widths[2623]), .RECT1_HEIGHT(rectangle1_heights[2623]), .RECT1_WEIGHT(rectangle1_weights[2623]), .RECT2_X(rectangle2_xs[2623]), .RECT2_Y(rectangle2_ys[2623]), .RECT2_WIDTH(rectangle2_widths[2623]), .RECT2_HEIGHT(rectangle2_heights[2623]), .RECT2_WEIGHT(rectangle2_weights[2623]), .RECT3_X(rectangle3_xs[2623]), .RECT3_Y(rectangle3_ys[2623]), .RECT3_WIDTH(rectangle3_widths[2623]), .RECT3_HEIGHT(rectangle3_heights[2623]), .RECT3_WEIGHT(rectangle3_weights[2623]), .FEAT_THRES(feature_thresholds[2623]), .FEAT_ABOVE(feature_aboves[2623]), .FEAT_BELOW(feature_belows[2623])) ac2623(.scan_win(scan_win2623), .scan_win_std_dev(scan_win_std_dev[2623]), .feature_accum(feature_accums[2623]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2624]), .RECT1_Y(rectangle1_ys[2624]), .RECT1_WIDTH(rectangle1_widths[2624]), .RECT1_HEIGHT(rectangle1_heights[2624]), .RECT1_WEIGHT(rectangle1_weights[2624]), .RECT2_X(rectangle2_xs[2624]), .RECT2_Y(rectangle2_ys[2624]), .RECT2_WIDTH(rectangle2_widths[2624]), .RECT2_HEIGHT(rectangle2_heights[2624]), .RECT2_WEIGHT(rectangle2_weights[2624]), .RECT3_X(rectangle3_xs[2624]), .RECT3_Y(rectangle3_ys[2624]), .RECT3_WIDTH(rectangle3_widths[2624]), .RECT3_HEIGHT(rectangle3_heights[2624]), .RECT3_WEIGHT(rectangle3_weights[2624]), .FEAT_THRES(feature_thresholds[2624]), .FEAT_ABOVE(feature_aboves[2624]), .FEAT_BELOW(feature_belows[2624])) ac2624(.scan_win(scan_win2624), .scan_win_std_dev(scan_win_std_dev[2624]), .feature_accum(feature_accums[2624]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2625]), .RECT1_Y(rectangle1_ys[2625]), .RECT1_WIDTH(rectangle1_widths[2625]), .RECT1_HEIGHT(rectangle1_heights[2625]), .RECT1_WEIGHT(rectangle1_weights[2625]), .RECT2_X(rectangle2_xs[2625]), .RECT2_Y(rectangle2_ys[2625]), .RECT2_WIDTH(rectangle2_widths[2625]), .RECT2_HEIGHT(rectangle2_heights[2625]), .RECT2_WEIGHT(rectangle2_weights[2625]), .RECT3_X(rectangle3_xs[2625]), .RECT3_Y(rectangle3_ys[2625]), .RECT3_WIDTH(rectangle3_widths[2625]), .RECT3_HEIGHT(rectangle3_heights[2625]), .RECT3_WEIGHT(rectangle3_weights[2625]), .FEAT_THRES(feature_thresholds[2625]), .FEAT_ABOVE(feature_aboves[2625]), .FEAT_BELOW(feature_belows[2625])) ac2625(.scan_win(scan_win2625), .scan_win_std_dev(scan_win_std_dev[2625]), .feature_accum(feature_accums[2625]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2626]), .RECT1_Y(rectangle1_ys[2626]), .RECT1_WIDTH(rectangle1_widths[2626]), .RECT1_HEIGHT(rectangle1_heights[2626]), .RECT1_WEIGHT(rectangle1_weights[2626]), .RECT2_X(rectangle2_xs[2626]), .RECT2_Y(rectangle2_ys[2626]), .RECT2_WIDTH(rectangle2_widths[2626]), .RECT2_HEIGHT(rectangle2_heights[2626]), .RECT2_WEIGHT(rectangle2_weights[2626]), .RECT3_X(rectangle3_xs[2626]), .RECT3_Y(rectangle3_ys[2626]), .RECT3_WIDTH(rectangle3_widths[2626]), .RECT3_HEIGHT(rectangle3_heights[2626]), .RECT3_WEIGHT(rectangle3_weights[2626]), .FEAT_THRES(feature_thresholds[2626]), .FEAT_ABOVE(feature_aboves[2626]), .FEAT_BELOW(feature_belows[2626])) ac2626(.scan_win(scan_win2626), .scan_win_std_dev(scan_win_std_dev[2626]), .feature_accum(feature_accums[2626]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2627]), .RECT1_Y(rectangle1_ys[2627]), .RECT1_WIDTH(rectangle1_widths[2627]), .RECT1_HEIGHT(rectangle1_heights[2627]), .RECT1_WEIGHT(rectangle1_weights[2627]), .RECT2_X(rectangle2_xs[2627]), .RECT2_Y(rectangle2_ys[2627]), .RECT2_WIDTH(rectangle2_widths[2627]), .RECT2_HEIGHT(rectangle2_heights[2627]), .RECT2_WEIGHT(rectangle2_weights[2627]), .RECT3_X(rectangle3_xs[2627]), .RECT3_Y(rectangle3_ys[2627]), .RECT3_WIDTH(rectangle3_widths[2627]), .RECT3_HEIGHT(rectangle3_heights[2627]), .RECT3_WEIGHT(rectangle3_weights[2627]), .FEAT_THRES(feature_thresholds[2627]), .FEAT_ABOVE(feature_aboves[2627]), .FEAT_BELOW(feature_belows[2627])) ac2627(.scan_win(scan_win2627), .scan_win_std_dev(scan_win_std_dev[2627]), .feature_accum(feature_accums[2627]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2628]), .RECT1_Y(rectangle1_ys[2628]), .RECT1_WIDTH(rectangle1_widths[2628]), .RECT1_HEIGHT(rectangle1_heights[2628]), .RECT1_WEIGHT(rectangle1_weights[2628]), .RECT2_X(rectangle2_xs[2628]), .RECT2_Y(rectangle2_ys[2628]), .RECT2_WIDTH(rectangle2_widths[2628]), .RECT2_HEIGHT(rectangle2_heights[2628]), .RECT2_WEIGHT(rectangle2_weights[2628]), .RECT3_X(rectangle3_xs[2628]), .RECT3_Y(rectangle3_ys[2628]), .RECT3_WIDTH(rectangle3_widths[2628]), .RECT3_HEIGHT(rectangle3_heights[2628]), .RECT3_WEIGHT(rectangle3_weights[2628]), .FEAT_THRES(feature_thresholds[2628]), .FEAT_ABOVE(feature_aboves[2628]), .FEAT_BELOW(feature_belows[2628])) ac2628(.scan_win(scan_win2628), .scan_win_std_dev(scan_win_std_dev[2628]), .feature_accum(feature_accums[2628]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2629]), .RECT1_Y(rectangle1_ys[2629]), .RECT1_WIDTH(rectangle1_widths[2629]), .RECT1_HEIGHT(rectangle1_heights[2629]), .RECT1_WEIGHT(rectangle1_weights[2629]), .RECT2_X(rectangle2_xs[2629]), .RECT2_Y(rectangle2_ys[2629]), .RECT2_WIDTH(rectangle2_widths[2629]), .RECT2_HEIGHT(rectangle2_heights[2629]), .RECT2_WEIGHT(rectangle2_weights[2629]), .RECT3_X(rectangle3_xs[2629]), .RECT3_Y(rectangle3_ys[2629]), .RECT3_WIDTH(rectangle3_widths[2629]), .RECT3_HEIGHT(rectangle3_heights[2629]), .RECT3_WEIGHT(rectangle3_weights[2629]), .FEAT_THRES(feature_thresholds[2629]), .FEAT_ABOVE(feature_aboves[2629]), .FEAT_BELOW(feature_belows[2629])) ac2629(.scan_win(scan_win2629), .scan_win_std_dev(scan_win_std_dev[2629]), .feature_accum(feature_accums[2629]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2630]), .RECT1_Y(rectangle1_ys[2630]), .RECT1_WIDTH(rectangle1_widths[2630]), .RECT1_HEIGHT(rectangle1_heights[2630]), .RECT1_WEIGHT(rectangle1_weights[2630]), .RECT2_X(rectangle2_xs[2630]), .RECT2_Y(rectangle2_ys[2630]), .RECT2_WIDTH(rectangle2_widths[2630]), .RECT2_HEIGHT(rectangle2_heights[2630]), .RECT2_WEIGHT(rectangle2_weights[2630]), .RECT3_X(rectangle3_xs[2630]), .RECT3_Y(rectangle3_ys[2630]), .RECT3_WIDTH(rectangle3_widths[2630]), .RECT3_HEIGHT(rectangle3_heights[2630]), .RECT3_WEIGHT(rectangle3_weights[2630]), .FEAT_THRES(feature_thresholds[2630]), .FEAT_ABOVE(feature_aboves[2630]), .FEAT_BELOW(feature_belows[2630])) ac2630(.scan_win(scan_win2630), .scan_win_std_dev(scan_win_std_dev[2630]), .feature_accum(feature_accums[2630]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2631]), .RECT1_Y(rectangle1_ys[2631]), .RECT1_WIDTH(rectangle1_widths[2631]), .RECT1_HEIGHT(rectangle1_heights[2631]), .RECT1_WEIGHT(rectangle1_weights[2631]), .RECT2_X(rectangle2_xs[2631]), .RECT2_Y(rectangle2_ys[2631]), .RECT2_WIDTH(rectangle2_widths[2631]), .RECT2_HEIGHT(rectangle2_heights[2631]), .RECT2_WEIGHT(rectangle2_weights[2631]), .RECT3_X(rectangle3_xs[2631]), .RECT3_Y(rectangle3_ys[2631]), .RECT3_WIDTH(rectangle3_widths[2631]), .RECT3_HEIGHT(rectangle3_heights[2631]), .RECT3_WEIGHT(rectangle3_weights[2631]), .FEAT_THRES(feature_thresholds[2631]), .FEAT_ABOVE(feature_aboves[2631]), .FEAT_BELOW(feature_belows[2631])) ac2631(.scan_win(scan_win2631), .scan_win_std_dev(scan_win_std_dev[2631]), .feature_accum(feature_accums[2631]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2632]), .RECT1_Y(rectangle1_ys[2632]), .RECT1_WIDTH(rectangle1_widths[2632]), .RECT1_HEIGHT(rectangle1_heights[2632]), .RECT1_WEIGHT(rectangle1_weights[2632]), .RECT2_X(rectangle2_xs[2632]), .RECT2_Y(rectangle2_ys[2632]), .RECT2_WIDTH(rectangle2_widths[2632]), .RECT2_HEIGHT(rectangle2_heights[2632]), .RECT2_WEIGHT(rectangle2_weights[2632]), .RECT3_X(rectangle3_xs[2632]), .RECT3_Y(rectangle3_ys[2632]), .RECT3_WIDTH(rectangle3_widths[2632]), .RECT3_HEIGHT(rectangle3_heights[2632]), .RECT3_WEIGHT(rectangle3_weights[2632]), .FEAT_THRES(feature_thresholds[2632]), .FEAT_ABOVE(feature_aboves[2632]), .FEAT_BELOW(feature_belows[2632])) ac2632(.scan_win(scan_win2632), .scan_win_std_dev(scan_win_std_dev[2632]), .feature_accum(feature_accums[2632]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2633]), .RECT1_Y(rectangle1_ys[2633]), .RECT1_WIDTH(rectangle1_widths[2633]), .RECT1_HEIGHT(rectangle1_heights[2633]), .RECT1_WEIGHT(rectangle1_weights[2633]), .RECT2_X(rectangle2_xs[2633]), .RECT2_Y(rectangle2_ys[2633]), .RECT2_WIDTH(rectangle2_widths[2633]), .RECT2_HEIGHT(rectangle2_heights[2633]), .RECT2_WEIGHT(rectangle2_weights[2633]), .RECT3_X(rectangle3_xs[2633]), .RECT3_Y(rectangle3_ys[2633]), .RECT3_WIDTH(rectangle3_widths[2633]), .RECT3_HEIGHT(rectangle3_heights[2633]), .RECT3_WEIGHT(rectangle3_weights[2633]), .FEAT_THRES(feature_thresholds[2633]), .FEAT_ABOVE(feature_aboves[2633]), .FEAT_BELOW(feature_belows[2633])) ac2633(.scan_win(scan_win2633), .scan_win_std_dev(scan_win_std_dev[2633]), .feature_accum(feature_accums[2633]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2634]), .RECT1_Y(rectangle1_ys[2634]), .RECT1_WIDTH(rectangle1_widths[2634]), .RECT1_HEIGHT(rectangle1_heights[2634]), .RECT1_WEIGHT(rectangle1_weights[2634]), .RECT2_X(rectangle2_xs[2634]), .RECT2_Y(rectangle2_ys[2634]), .RECT2_WIDTH(rectangle2_widths[2634]), .RECT2_HEIGHT(rectangle2_heights[2634]), .RECT2_WEIGHT(rectangle2_weights[2634]), .RECT3_X(rectangle3_xs[2634]), .RECT3_Y(rectangle3_ys[2634]), .RECT3_WIDTH(rectangle3_widths[2634]), .RECT3_HEIGHT(rectangle3_heights[2634]), .RECT3_WEIGHT(rectangle3_weights[2634]), .FEAT_THRES(feature_thresholds[2634]), .FEAT_ABOVE(feature_aboves[2634]), .FEAT_BELOW(feature_belows[2634])) ac2634(.scan_win(scan_win2634), .scan_win_std_dev(scan_win_std_dev[2634]), .feature_accum(feature_accums[2634]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2635]), .RECT1_Y(rectangle1_ys[2635]), .RECT1_WIDTH(rectangle1_widths[2635]), .RECT1_HEIGHT(rectangle1_heights[2635]), .RECT1_WEIGHT(rectangle1_weights[2635]), .RECT2_X(rectangle2_xs[2635]), .RECT2_Y(rectangle2_ys[2635]), .RECT2_WIDTH(rectangle2_widths[2635]), .RECT2_HEIGHT(rectangle2_heights[2635]), .RECT2_WEIGHT(rectangle2_weights[2635]), .RECT3_X(rectangle3_xs[2635]), .RECT3_Y(rectangle3_ys[2635]), .RECT3_WIDTH(rectangle3_widths[2635]), .RECT3_HEIGHT(rectangle3_heights[2635]), .RECT3_WEIGHT(rectangle3_weights[2635]), .FEAT_THRES(feature_thresholds[2635]), .FEAT_ABOVE(feature_aboves[2635]), .FEAT_BELOW(feature_belows[2635])) ac2635(.scan_win(scan_win2635), .scan_win_std_dev(scan_win_std_dev[2635]), .feature_accum(feature_accums[2635]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2636]), .RECT1_Y(rectangle1_ys[2636]), .RECT1_WIDTH(rectangle1_widths[2636]), .RECT1_HEIGHT(rectangle1_heights[2636]), .RECT1_WEIGHT(rectangle1_weights[2636]), .RECT2_X(rectangle2_xs[2636]), .RECT2_Y(rectangle2_ys[2636]), .RECT2_WIDTH(rectangle2_widths[2636]), .RECT2_HEIGHT(rectangle2_heights[2636]), .RECT2_WEIGHT(rectangle2_weights[2636]), .RECT3_X(rectangle3_xs[2636]), .RECT3_Y(rectangle3_ys[2636]), .RECT3_WIDTH(rectangle3_widths[2636]), .RECT3_HEIGHT(rectangle3_heights[2636]), .RECT3_WEIGHT(rectangle3_weights[2636]), .FEAT_THRES(feature_thresholds[2636]), .FEAT_ABOVE(feature_aboves[2636]), .FEAT_BELOW(feature_belows[2636])) ac2636(.scan_win(scan_win2636), .scan_win_std_dev(scan_win_std_dev[2636]), .feature_accum(feature_accums[2636]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2637]), .RECT1_Y(rectangle1_ys[2637]), .RECT1_WIDTH(rectangle1_widths[2637]), .RECT1_HEIGHT(rectangle1_heights[2637]), .RECT1_WEIGHT(rectangle1_weights[2637]), .RECT2_X(rectangle2_xs[2637]), .RECT2_Y(rectangle2_ys[2637]), .RECT2_WIDTH(rectangle2_widths[2637]), .RECT2_HEIGHT(rectangle2_heights[2637]), .RECT2_WEIGHT(rectangle2_weights[2637]), .RECT3_X(rectangle3_xs[2637]), .RECT3_Y(rectangle3_ys[2637]), .RECT3_WIDTH(rectangle3_widths[2637]), .RECT3_HEIGHT(rectangle3_heights[2637]), .RECT3_WEIGHT(rectangle3_weights[2637]), .FEAT_THRES(feature_thresholds[2637]), .FEAT_ABOVE(feature_aboves[2637]), .FEAT_BELOW(feature_belows[2637])) ac2637(.scan_win(scan_win2637), .scan_win_std_dev(scan_win_std_dev[2637]), .feature_accum(feature_accums[2637]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2638]), .RECT1_Y(rectangle1_ys[2638]), .RECT1_WIDTH(rectangle1_widths[2638]), .RECT1_HEIGHT(rectangle1_heights[2638]), .RECT1_WEIGHT(rectangle1_weights[2638]), .RECT2_X(rectangle2_xs[2638]), .RECT2_Y(rectangle2_ys[2638]), .RECT2_WIDTH(rectangle2_widths[2638]), .RECT2_HEIGHT(rectangle2_heights[2638]), .RECT2_WEIGHT(rectangle2_weights[2638]), .RECT3_X(rectangle3_xs[2638]), .RECT3_Y(rectangle3_ys[2638]), .RECT3_WIDTH(rectangle3_widths[2638]), .RECT3_HEIGHT(rectangle3_heights[2638]), .RECT3_WEIGHT(rectangle3_weights[2638]), .FEAT_THRES(feature_thresholds[2638]), .FEAT_ABOVE(feature_aboves[2638]), .FEAT_BELOW(feature_belows[2638])) ac2638(.scan_win(scan_win2638), .scan_win_std_dev(scan_win_std_dev[2638]), .feature_accum(feature_accums[2638]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2639]), .RECT1_Y(rectangle1_ys[2639]), .RECT1_WIDTH(rectangle1_widths[2639]), .RECT1_HEIGHT(rectangle1_heights[2639]), .RECT1_WEIGHT(rectangle1_weights[2639]), .RECT2_X(rectangle2_xs[2639]), .RECT2_Y(rectangle2_ys[2639]), .RECT2_WIDTH(rectangle2_widths[2639]), .RECT2_HEIGHT(rectangle2_heights[2639]), .RECT2_WEIGHT(rectangle2_weights[2639]), .RECT3_X(rectangle3_xs[2639]), .RECT3_Y(rectangle3_ys[2639]), .RECT3_WIDTH(rectangle3_widths[2639]), .RECT3_HEIGHT(rectangle3_heights[2639]), .RECT3_WEIGHT(rectangle3_weights[2639]), .FEAT_THRES(feature_thresholds[2639]), .FEAT_ABOVE(feature_aboves[2639]), .FEAT_BELOW(feature_belows[2639])) ac2639(.scan_win(scan_win2639), .scan_win_std_dev(scan_win_std_dev[2639]), .feature_accum(feature_accums[2639]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2640]), .RECT1_Y(rectangle1_ys[2640]), .RECT1_WIDTH(rectangle1_widths[2640]), .RECT1_HEIGHT(rectangle1_heights[2640]), .RECT1_WEIGHT(rectangle1_weights[2640]), .RECT2_X(rectangle2_xs[2640]), .RECT2_Y(rectangle2_ys[2640]), .RECT2_WIDTH(rectangle2_widths[2640]), .RECT2_HEIGHT(rectangle2_heights[2640]), .RECT2_WEIGHT(rectangle2_weights[2640]), .RECT3_X(rectangle3_xs[2640]), .RECT3_Y(rectangle3_ys[2640]), .RECT3_WIDTH(rectangle3_widths[2640]), .RECT3_HEIGHT(rectangle3_heights[2640]), .RECT3_WEIGHT(rectangle3_weights[2640]), .FEAT_THRES(feature_thresholds[2640]), .FEAT_ABOVE(feature_aboves[2640]), .FEAT_BELOW(feature_belows[2640])) ac2640(.scan_win(scan_win2640), .scan_win_std_dev(scan_win_std_dev[2640]), .feature_accum(feature_accums[2640]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2641]), .RECT1_Y(rectangle1_ys[2641]), .RECT1_WIDTH(rectangle1_widths[2641]), .RECT1_HEIGHT(rectangle1_heights[2641]), .RECT1_WEIGHT(rectangle1_weights[2641]), .RECT2_X(rectangle2_xs[2641]), .RECT2_Y(rectangle2_ys[2641]), .RECT2_WIDTH(rectangle2_widths[2641]), .RECT2_HEIGHT(rectangle2_heights[2641]), .RECT2_WEIGHT(rectangle2_weights[2641]), .RECT3_X(rectangle3_xs[2641]), .RECT3_Y(rectangle3_ys[2641]), .RECT3_WIDTH(rectangle3_widths[2641]), .RECT3_HEIGHT(rectangle3_heights[2641]), .RECT3_WEIGHT(rectangle3_weights[2641]), .FEAT_THRES(feature_thresholds[2641]), .FEAT_ABOVE(feature_aboves[2641]), .FEAT_BELOW(feature_belows[2641])) ac2641(.scan_win(scan_win2641), .scan_win_std_dev(scan_win_std_dev[2641]), .feature_accum(feature_accums[2641]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2642]), .RECT1_Y(rectangle1_ys[2642]), .RECT1_WIDTH(rectangle1_widths[2642]), .RECT1_HEIGHT(rectangle1_heights[2642]), .RECT1_WEIGHT(rectangle1_weights[2642]), .RECT2_X(rectangle2_xs[2642]), .RECT2_Y(rectangle2_ys[2642]), .RECT2_WIDTH(rectangle2_widths[2642]), .RECT2_HEIGHT(rectangle2_heights[2642]), .RECT2_WEIGHT(rectangle2_weights[2642]), .RECT3_X(rectangle3_xs[2642]), .RECT3_Y(rectangle3_ys[2642]), .RECT3_WIDTH(rectangle3_widths[2642]), .RECT3_HEIGHT(rectangle3_heights[2642]), .RECT3_WEIGHT(rectangle3_weights[2642]), .FEAT_THRES(feature_thresholds[2642]), .FEAT_ABOVE(feature_aboves[2642]), .FEAT_BELOW(feature_belows[2642])) ac2642(.scan_win(scan_win2642), .scan_win_std_dev(scan_win_std_dev[2642]), .feature_accum(feature_accums[2642]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2643]), .RECT1_Y(rectangle1_ys[2643]), .RECT1_WIDTH(rectangle1_widths[2643]), .RECT1_HEIGHT(rectangle1_heights[2643]), .RECT1_WEIGHT(rectangle1_weights[2643]), .RECT2_X(rectangle2_xs[2643]), .RECT2_Y(rectangle2_ys[2643]), .RECT2_WIDTH(rectangle2_widths[2643]), .RECT2_HEIGHT(rectangle2_heights[2643]), .RECT2_WEIGHT(rectangle2_weights[2643]), .RECT3_X(rectangle3_xs[2643]), .RECT3_Y(rectangle3_ys[2643]), .RECT3_WIDTH(rectangle3_widths[2643]), .RECT3_HEIGHT(rectangle3_heights[2643]), .RECT3_WEIGHT(rectangle3_weights[2643]), .FEAT_THRES(feature_thresholds[2643]), .FEAT_ABOVE(feature_aboves[2643]), .FEAT_BELOW(feature_belows[2643])) ac2643(.scan_win(scan_win2643), .scan_win_std_dev(scan_win_std_dev[2643]), .feature_accum(feature_accums[2643]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2644]), .RECT1_Y(rectangle1_ys[2644]), .RECT1_WIDTH(rectangle1_widths[2644]), .RECT1_HEIGHT(rectangle1_heights[2644]), .RECT1_WEIGHT(rectangle1_weights[2644]), .RECT2_X(rectangle2_xs[2644]), .RECT2_Y(rectangle2_ys[2644]), .RECT2_WIDTH(rectangle2_widths[2644]), .RECT2_HEIGHT(rectangle2_heights[2644]), .RECT2_WEIGHT(rectangle2_weights[2644]), .RECT3_X(rectangle3_xs[2644]), .RECT3_Y(rectangle3_ys[2644]), .RECT3_WIDTH(rectangle3_widths[2644]), .RECT3_HEIGHT(rectangle3_heights[2644]), .RECT3_WEIGHT(rectangle3_weights[2644]), .FEAT_THRES(feature_thresholds[2644]), .FEAT_ABOVE(feature_aboves[2644]), .FEAT_BELOW(feature_belows[2644])) ac2644(.scan_win(scan_win2644), .scan_win_std_dev(scan_win_std_dev[2644]), .feature_accum(feature_accums[2644]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2645]), .RECT1_Y(rectangle1_ys[2645]), .RECT1_WIDTH(rectangle1_widths[2645]), .RECT1_HEIGHT(rectangle1_heights[2645]), .RECT1_WEIGHT(rectangle1_weights[2645]), .RECT2_X(rectangle2_xs[2645]), .RECT2_Y(rectangle2_ys[2645]), .RECT2_WIDTH(rectangle2_widths[2645]), .RECT2_HEIGHT(rectangle2_heights[2645]), .RECT2_WEIGHT(rectangle2_weights[2645]), .RECT3_X(rectangle3_xs[2645]), .RECT3_Y(rectangle3_ys[2645]), .RECT3_WIDTH(rectangle3_widths[2645]), .RECT3_HEIGHT(rectangle3_heights[2645]), .RECT3_WEIGHT(rectangle3_weights[2645]), .FEAT_THRES(feature_thresholds[2645]), .FEAT_ABOVE(feature_aboves[2645]), .FEAT_BELOW(feature_belows[2645])) ac2645(.scan_win(scan_win2645), .scan_win_std_dev(scan_win_std_dev[2645]), .feature_accum(feature_accums[2645]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2646]), .RECT1_Y(rectangle1_ys[2646]), .RECT1_WIDTH(rectangle1_widths[2646]), .RECT1_HEIGHT(rectangle1_heights[2646]), .RECT1_WEIGHT(rectangle1_weights[2646]), .RECT2_X(rectangle2_xs[2646]), .RECT2_Y(rectangle2_ys[2646]), .RECT2_WIDTH(rectangle2_widths[2646]), .RECT2_HEIGHT(rectangle2_heights[2646]), .RECT2_WEIGHT(rectangle2_weights[2646]), .RECT3_X(rectangle3_xs[2646]), .RECT3_Y(rectangle3_ys[2646]), .RECT3_WIDTH(rectangle3_widths[2646]), .RECT3_HEIGHT(rectangle3_heights[2646]), .RECT3_WEIGHT(rectangle3_weights[2646]), .FEAT_THRES(feature_thresholds[2646]), .FEAT_ABOVE(feature_aboves[2646]), .FEAT_BELOW(feature_belows[2646])) ac2646(.scan_win(scan_win2646), .scan_win_std_dev(scan_win_std_dev[2646]), .feature_accum(feature_accums[2646]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2647]), .RECT1_Y(rectangle1_ys[2647]), .RECT1_WIDTH(rectangle1_widths[2647]), .RECT1_HEIGHT(rectangle1_heights[2647]), .RECT1_WEIGHT(rectangle1_weights[2647]), .RECT2_X(rectangle2_xs[2647]), .RECT2_Y(rectangle2_ys[2647]), .RECT2_WIDTH(rectangle2_widths[2647]), .RECT2_HEIGHT(rectangle2_heights[2647]), .RECT2_WEIGHT(rectangle2_weights[2647]), .RECT3_X(rectangle3_xs[2647]), .RECT3_Y(rectangle3_ys[2647]), .RECT3_WIDTH(rectangle3_widths[2647]), .RECT3_HEIGHT(rectangle3_heights[2647]), .RECT3_WEIGHT(rectangle3_weights[2647]), .FEAT_THRES(feature_thresholds[2647]), .FEAT_ABOVE(feature_aboves[2647]), .FEAT_BELOW(feature_belows[2647])) ac2647(.scan_win(scan_win2647), .scan_win_std_dev(scan_win_std_dev[2647]), .feature_accum(feature_accums[2647]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2648]), .RECT1_Y(rectangle1_ys[2648]), .RECT1_WIDTH(rectangle1_widths[2648]), .RECT1_HEIGHT(rectangle1_heights[2648]), .RECT1_WEIGHT(rectangle1_weights[2648]), .RECT2_X(rectangle2_xs[2648]), .RECT2_Y(rectangle2_ys[2648]), .RECT2_WIDTH(rectangle2_widths[2648]), .RECT2_HEIGHT(rectangle2_heights[2648]), .RECT2_WEIGHT(rectangle2_weights[2648]), .RECT3_X(rectangle3_xs[2648]), .RECT3_Y(rectangle3_ys[2648]), .RECT3_WIDTH(rectangle3_widths[2648]), .RECT3_HEIGHT(rectangle3_heights[2648]), .RECT3_WEIGHT(rectangle3_weights[2648]), .FEAT_THRES(feature_thresholds[2648]), .FEAT_ABOVE(feature_aboves[2648]), .FEAT_BELOW(feature_belows[2648])) ac2648(.scan_win(scan_win2648), .scan_win_std_dev(scan_win_std_dev[2648]), .feature_accum(feature_accums[2648]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2649]), .RECT1_Y(rectangle1_ys[2649]), .RECT1_WIDTH(rectangle1_widths[2649]), .RECT1_HEIGHT(rectangle1_heights[2649]), .RECT1_WEIGHT(rectangle1_weights[2649]), .RECT2_X(rectangle2_xs[2649]), .RECT2_Y(rectangle2_ys[2649]), .RECT2_WIDTH(rectangle2_widths[2649]), .RECT2_HEIGHT(rectangle2_heights[2649]), .RECT2_WEIGHT(rectangle2_weights[2649]), .RECT3_X(rectangle3_xs[2649]), .RECT3_Y(rectangle3_ys[2649]), .RECT3_WIDTH(rectangle3_widths[2649]), .RECT3_HEIGHT(rectangle3_heights[2649]), .RECT3_WEIGHT(rectangle3_weights[2649]), .FEAT_THRES(feature_thresholds[2649]), .FEAT_ABOVE(feature_aboves[2649]), .FEAT_BELOW(feature_belows[2649])) ac2649(.scan_win(scan_win2649), .scan_win_std_dev(scan_win_std_dev[2649]), .feature_accum(feature_accums[2649]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2650]), .RECT1_Y(rectangle1_ys[2650]), .RECT1_WIDTH(rectangle1_widths[2650]), .RECT1_HEIGHT(rectangle1_heights[2650]), .RECT1_WEIGHT(rectangle1_weights[2650]), .RECT2_X(rectangle2_xs[2650]), .RECT2_Y(rectangle2_ys[2650]), .RECT2_WIDTH(rectangle2_widths[2650]), .RECT2_HEIGHT(rectangle2_heights[2650]), .RECT2_WEIGHT(rectangle2_weights[2650]), .RECT3_X(rectangle3_xs[2650]), .RECT3_Y(rectangle3_ys[2650]), .RECT3_WIDTH(rectangle3_widths[2650]), .RECT3_HEIGHT(rectangle3_heights[2650]), .RECT3_WEIGHT(rectangle3_weights[2650]), .FEAT_THRES(feature_thresholds[2650]), .FEAT_ABOVE(feature_aboves[2650]), .FEAT_BELOW(feature_belows[2650])) ac2650(.scan_win(scan_win2650), .scan_win_std_dev(scan_win_std_dev[2650]), .feature_accum(feature_accums[2650]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2651]), .RECT1_Y(rectangle1_ys[2651]), .RECT1_WIDTH(rectangle1_widths[2651]), .RECT1_HEIGHT(rectangle1_heights[2651]), .RECT1_WEIGHT(rectangle1_weights[2651]), .RECT2_X(rectangle2_xs[2651]), .RECT2_Y(rectangle2_ys[2651]), .RECT2_WIDTH(rectangle2_widths[2651]), .RECT2_HEIGHT(rectangle2_heights[2651]), .RECT2_WEIGHT(rectangle2_weights[2651]), .RECT3_X(rectangle3_xs[2651]), .RECT3_Y(rectangle3_ys[2651]), .RECT3_WIDTH(rectangle3_widths[2651]), .RECT3_HEIGHT(rectangle3_heights[2651]), .RECT3_WEIGHT(rectangle3_weights[2651]), .FEAT_THRES(feature_thresholds[2651]), .FEAT_ABOVE(feature_aboves[2651]), .FEAT_BELOW(feature_belows[2651])) ac2651(.scan_win(scan_win2651), .scan_win_std_dev(scan_win_std_dev[2651]), .feature_accum(feature_accums[2651]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2652]), .RECT1_Y(rectangle1_ys[2652]), .RECT1_WIDTH(rectangle1_widths[2652]), .RECT1_HEIGHT(rectangle1_heights[2652]), .RECT1_WEIGHT(rectangle1_weights[2652]), .RECT2_X(rectangle2_xs[2652]), .RECT2_Y(rectangle2_ys[2652]), .RECT2_WIDTH(rectangle2_widths[2652]), .RECT2_HEIGHT(rectangle2_heights[2652]), .RECT2_WEIGHT(rectangle2_weights[2652]), .RECT3_X(rectangle3_xs[2652]), .RECT3_Y(rectangle3_ys[2652]), .RECT3_WIDTH(rectangle3_widths[2652]), .RECT3_HEIGHT(rectangle3_heights[2652]), .RECT3_WEIGHT(rectangle3_weights[2652]), .FEAT_THRES(feature_thresholds[2652]), .FEAT_ABOVE(feature_aboves[2652]), .FEAT_BELOW(feature_belows[2652])) ac2652(.scan_win(scan_win2652), .scan_win_std_dev(scan_win_std_dev[2652]), .feature_accum(feature_accums[2652]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2653]), .RECT1_Y(rectangle1_ys[2653]), .RECT1_WIDTH(rectangle1_widths[2653]), .RECT1_HEIGHT(rectangle1_heights[2653]), .RECT1_WEIGHT(rectangle1_weights[2653]), .RECT2_X(rectangle2_xs[2653]), .RECT2_Y(rectangle2_ys[2653]), .RECT2_WIDTH(rectangle2_widths[2653]), .RECT2_HEIGHT(rectangle2_heights[2653]), .RECT2_WEIGHT(rectangle2_weights[2653]), .RECT3_X(rectangle3_xs[2653]), .RECT3_Y(rectangle3_ys[2653]), .RECT3_WIDTH(rectangle3_widths[2653]), .RECT3_HEIGHT(rectangle3_heights[2653]), .RECT3_WEIGHT(rectangle3_weights[2653]), .FEAT_THRES(feature_thresholds[2653]), .FEAT_ABOVE(feature_aboves[2653]), .FEAT_BELOW(feature_belows[2653])) ac2653(.scan_win(scan_win2653), .scan_win_std_dev(scan_win_std_dev[2653]), .feature_accum(feature_accums[2653]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2654]), .RECT1_Y(rectangle1_ys[2654]), .RECT1_WIDTH(rectangle1_widths[2654]), .RECT1_HEIGHT(rectangle1_heights[2654]), .RECT1_WEIGHT(rectangle1_weights[2654]), .RECT2_X(rectangle2_xs[2654]), .RECT2_Y(rectangle2_ys[2654]), .RECT2_WIDTH(rectangle2_widths[2654]), .RECT2_HEIGHT(rectangle2_heights[2654]), .RECT2_WEIGHT(rectangle2_weights[2654]), .RECT3_X(rectangle3_xs[2654]), .RECT3_Y(rectangle3_ys[2654]), .RECT3_WIDTH(rectangle3_widths[2654]), .RECT3_HEIGHT(rectangle3_heights[2654]), .RECT3_WEIGHT(rectangle3_weights[2654]), .FEAT_THRES(feature_thresholds[2654]), .FEAT_ABOVE(feature_aboves[2654]), .FEAT_BELOW(feature_belows[2654])) ac2654(.scan_win(scan_win2654), .scan_win_std_dev(scan_win_std_dev[2654]), .feature_accum(feature_accums[2654]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2655]), .RECT1_Y(rectangle1_ys[2655]), .RECT1_WIDTH(rectangle1_widths[2655]), .RECT1_HEIGHT(rectangle1_heights[2655]), .RECT1_WEIGHT(rectangle1_weights[2655]), .RECT2_X(rectangle2_xs[2655]), .RECT2_Y(rectangle2_ys[2655]), .RECT2_WIDTH(rectangle2_widths[2655]), .RECT2_HEIGHT(rectangle2_heights[2655]), .RECT2_WEIGHT(rectangle2_weights[2655]), .RECT3_X(rectangle3_xs[2655]), .RECT3_Y(rectangle3_ys[2655]), .RECT3_WIDTH(rectangle3_widths[2655]), .RECT3_HEIGHT(rectangle3_heights[2655]), .RECT3_WEIGHT(rectangle3_weights[2655]), .FEAT_THRES(feature_thresholds[2655]), .FEAT_ABOVE(feature_aboves[2655]), .FEAT_BELOW(feature_belows[2655])) ac2655(.scan_win(scan_win2655), .scan_win_std_dev(scan_win_std_dev[2655]), .feature_accum(feature_accums[2655]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2656]), .RECT1_Y(rectangle1_ys[2656]), .RECT1_WIDTH(rectangle1_widths[2656]), .RECT1_HEIGHT(rectangle1_heights[2656]), .RECT1_WEIGHT(rectangle1_weights[2656]), .RECT2_X(rectangle2_xs[2656]), .RECT2_Y(rectangle2_ys[2656]), .RECT2_WIDTH(rectangle2_widths[2656]), .RECT2_HEIGHT(rectangle2_heights[2656]), .RECT2_WEIGHT(rectangle2_weights[2656]), .RECT3_X(rectangle3_xs[2656]), .RECT3_Y(rectangle3_ys[2656]), .RECT3_WIDTH(rectangle3_widths[2656]), .RECT3_HEIGHT(rectangle3_heights[2656]), .RECT3_WEIGHT(rectangle3_weights[2656]), .FEAT_THRES(feature_thresholds[2656]), .FEAT_ABOVE(feature_aboves[2656]), .FEAT_BELOW(feature_belows[2656])) ac2656(.scan_win(scan_win2656), .scan_win_std_dev(scan_win_std_dev[2656]), .feature_accum(feature_accums[2656]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2657]), .RECT1_Y(rectangle1_ys[2657]), .RECT1_WIDTH(rectangle1_widths[2657]), .RECT1_HEIGHT(rectangle1_heights[2657]), .RECT1_WEIGHT(rectangle1_weights[2657]), .RECT2_X(rectangle2_xs[2657]), .RECT2_Y(rectangle2_ys[2657]), .RECT2_WIDTH(rectangle2_widths[2657]), .RECT2_HEIGHT(rectangle2_heights[2657]), .RECT2_WEIGHT(rectangle2_weights[2657]), .RECT3_X(rectangle3_xs[2657]), .RECT3_Y(rectangle3_ys[2657]), .RECT3_WIDTH(rectangle3_widths[2657]), .RECT3_HEIGHT(rectangle3_heights[2657]), .RECT3_WEIGHT(rectangle3_weights[2657]), .FEAT_THRES(feature_thresholds[2657]), .FEAT_ABOVE(feature_aboves[2657]), .FEAT_BELOW(feature_belows[2657])) ac2657(.scan_win(scan_win2657), .scan_win_std_dev(scan_win_std_dev[2657]), .feature_accum(feature_accums[2657]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2658]), .RECT1_Y(rectangle1_ys[2658]), .RECT1_WIDTH(rectangle1_widths[2658]), .RECT1_HEIGHT(rectangle1_heights[2658]), .RECT1_WEIGHT(rectangle1_weights[2658]), .RECT2_X(rectangle2_xs[2658]), .RECT2_Y(rectangle2_ys[2658]), .RECT2_WIDTH(rectangle2_widths[2658]), .RECT2_HEIGHT(rectangle2_heights[2658]), .RECT2_WEIGHT(rectangle2_weights[2658]), .RECT3_X(rectangle3_xs[2658]), .RECT3_Y(rectangle3_ys[2658]), .RECT3_WIDTH(rectangle3_widths[2658]), .RECT3_HEIGHT(rectangle3_heights[2658]), .RECT3_WEIGHT(rectangle3_weights[2658]), .FEAT_THRES(feature_thresholds[2658]), .FEAT_ABOVE(feature_aboves[2658]), .FEAT_BELOW(feature_belows[2658])) ac2658(.scan_win(scan_win2658), .scan_win_std_dev(scan_win_std_dev[2658]), .feature_accum(feature_accums[2658]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2659]), .RECT1_Y(rectangle1_ys[2659]), .RECT1_WIDTH(rectangle1_widths[2659]), .RECT1_HEIGHT(rectangle1_heights[2659]), .RECT1_WEIGHT(rectangle1_weights[2659]), .RECT2_X(rectangle2_xs[2659]), .RECT2_Y(rectangle2_ys[2659]), .RECT2_WIDTH(rectangle2_widths[2659]), .RECT2_HEIGHT(rectangle2_heights[2659]), .RECT2_WEIGHT(rectangle2_weights[2659]), .RECT3_X(rectangle3_xs[2659]), .RECT3_Y(rectangle3_ys[2659]), .RECT3_WIDTH(rectangle3_widths[2659]), .RECT3_HEIGHT(rectangle3_heights[2659]), .RECT3_WEIGHT(rectangle3_weights[2659]), .FEAT_THRES(feature_thresholds[2659]), .FEAT_ABOVE(feature_aboves[2659]), .FEAT_BELOW(feature_belows[2659])) ac2659(.scan_win(scan_win2659), .scan_win_std_dev(scan_win_std_dev[2659]), .feature_accum(feature_accums[2659]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2660]), .RECT1_Y(rectangle1_ys[2660]), .RECT1_WIDTH(rectangle1_widths[2660]), .RECT1_HEIGHT(rectangle1_heights[2660]), .RECT1_WEIGHT(rectangle1_weights[2660]), .RECT2_X(rectangle2_xs[2660]), .RECT2_Y(rectangle2_ys[2660]), .RECT2_WIDTH(rectangle2_widths[2660]), .RECT2_HEIGHT(rectangle2_heights[2660]), .RECT2_WEIGHT(rectangle2_weights[2660]), .RECT3_X(rectangle3_xs[2660]), .RECT3_Y(rectangle3_ys[2660]), .RECT3_WIDTH(rectangle3_widths[2660]), .RECT3_HEIGHT(rectangle3_heights[2660]), .RECT3_WEIGHT(rectangle3_weights[2660]), .FEAT_THRES(feature_thresholds[2660]), .FEAT_ABOVE(feature_aboves[2660]), .FEAT_BELOW(feature_belows[2660])) ac2660(.scan_win(scan_win2660), .scan_win_std_dev(scan_win_std_dev[2660]), .feature_accum(feature_accums[2660]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2661]), .RECT1_Y(rectangle1_ys[2661]), .RECT1_WIDTH(rectangle1_widths[2661]), .RECT1_HEIGHT(rectangle1_heights[2661]), .RECT1_WEIGHT(rectangle1_weights[2661]), .RECT2_X(rectangle2_xs[2661]), .RECT2_Y(rectangle2_ys[2661]), .RECT2_WIDTH(rectangle2_widths[2661]), .RECT2_HEIGHT(rectangle2_heights[2661]), .RECT2_WEIGHT(rectangle2_weights[2661]), .RECT3_X(rectangle3_xs[2661]), .RECT3_Y(rectangle3_ys[2661]), .RECT3_WIDTH(rectangle3_widths[2661]), .RECT3_HEIGHT(rectangle3_heights[2661]), .RECT3_WEIGHT(rectangle3_weights[2661]), .FEAT_THRES(feature_thresholds[2661]), .FEAT_ABOVE(feature_aboves[2661]), .FEAT_BELOW(feature_belows[2661])) ac2661(.scan_win(scan_win2661), .scan_win_std_dev(scan_win_std_dev[2661]), .feature_accum(feature_accums[2661]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2662]), .RECT1_Y(rectangle1_ys[2662]), .RECT1_WIDTH(rectangle1_widths[2662]), .RECT1_HEIGHT(rectangle1_heights[2662]), .RECT1_WEIGHT(rectangle1_weights[2662]), .RECT2_X(rectangle2_xs[2662]), .RECT2_Y(rectangle2_ys[2662]), .RECT2_WIDTH(rectangle2_widths[2662]), .RECT2_HEIGHT(rectangle2_heights[2662]), .RECT2_WEIGHT(rectangle2_weights[2662]), .RECT3_X(rectangle3_xs[2662]), .RECT3_Y(rectangle3_ys[2662]), .RECT3_WIDTH(rectangle3_widths[2662]), .RECT3_HEIGHT(rectangle3_heights[2662]), .RECT3_WEIGHT(rectangle3_weights[2662]), .FEAT_THRES(feature_thresholds[2662]), .FEAT_ABOVE(feature_aboves[2662]), .FEAT_BELOW(feature_belows[2662])) ac2662(.scan_win(scan_win2662), .scan_win_std_dev(scan_win_std_dev[2662]), .feature_accum(feature_accums[2662]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2663]), .RECT1_Y(rectangle1_ys[2663]), .RECT1_WIDTH(rectangle1_widths[2663]), .RECT1_HEIGHT(rectangle1_heights[2663]), .RECT1_WEIGHT(rectangle1_weights[2663]), .RECT2_X(rectangle2_xs[2663]), .RECT2_Y(rectangle2_ys[2663]), .RECT2_WIDTH(rectangle2_widths[2663]), .RECT2_HEIGHT(rectangle2_heights[2663]), .RECT2_WEIGHT(rectangle2_weights[2663]), .RECT3_X(rectangle3_xs[2663]), .RECT3_Y(rectangle3_ys[2663]), .RECT3_WIDTH(rectangle3_widths[2663]), .RECT3_HEIGHT(rectangle3_heights[2663]), .RECT3_WEIGHT(rectangle3_weights[2663]), .FEAT_THRES(feature_thresholds[2663]), .FEAT_ABOVE(feature_aboves[2663]), .FEAT_BELOW(feature_belows[2663])) ac2663(.scan_win(scan_win2663), .scan_win_std_dev(scan_win_std_dev[2663]), .feature_accum(feature_accums[2663]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2664]), .RECT1_Y(rectangle1_ys[2664]), .RECT1_WIDTH(rectangle1_widths[2664]), .RECT1_HEIGHT(rectangle1_heights[2664]), .RECT1_WEIGHT(rectangle1_weights[2664]), .RECT2_X(rectangle2_xs[2664]), .RECT2_Y(rectangle2_ys[2664]), .RECT2_WIDTH(rectangle2_widths[2664]), .RECT2_HEIGHT(rectangle2_heights[2664]), .RECT2_WEIGHT(rectangle2_weights[2664]), .RECT3_X(rectangle3_xs[2664]), .RECT3_Y(rectangle3_ys[2664]), .RECT3_WIDTH(rectangle3_widths[2664]), .RECT3_HEIGHT(rectangle3_heights[2664]), .RECT3_WEIGHT(rectangle3_weights[2664]), .FEAT_THRES(feature_thresholds[2664]), .FEAT_ABOVE(feature_aboves[2664]), .FEAT_BELOW(feature_belows[2664])) ac2664(.scan_win(scan_win2664), .scan_win_std_dev(scan_win_std_dev[2664]), .feature_accum(feature_accums[2664]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2665]), .RECT1_Y(rectangle1_ys[2665]), .RECT1_WIDTH(rectangle1_widths[2665]), .RECT1_HEIGHT(rectangle1_heights[2665]), .RECT1_WEIGHT(rectangle1_weights[2665]), .RECT2_X(rectangle2_xs[2665]), .RECT2_Y(rectangle2_ys[2665]), .RECT2_WIDTH(rectangle2_widths[2665]), .RECT2_HEIGHT(rectangle2_heights[2665]), .RECT2_WEIGHT(rectangle2_weights[2665]), .RECT3_X(rectangle3_xs[2665]), .RECT3_Y(rectangle3_ys[2665]), .RECT3_WIDTH(rectangle3_widths[2665]), .RECT3_HEIGHT(rectangle3_heights[2665]), .RECT3_WEIGHT(rectangle3_weights[2665]), .FEAT_THRES(feature_thresholds[2665]), .FEAT_ABOVE(feature_aboves[2665]), .FEAT_BELOW(feature_belows[2665])) ac2665(.scan_win(scan_win2665), .scan_win_std_dev(scan_win_std_dev[2665]), .feature_accum(feature_accums[2665]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2666]), .RECT1_Y(rectangle1_ys[2666]), .RECT1_WIDTH(rectangle1_widths[2666]), .RECT1_HEIGHT(rectangle1_heights[2666]), .RECT1_WEIGHT(rectangle1_weights[2666]), .RECT2_X(rectangle2_xs[2666]), .RECT2_Y(rectangle2_ys[2666]), .RECT2_WIDTH(rectangle2_widths[2666]), .RECT2_HEIGHT(rectangle2_heights[2666]), .RECT2_WEIGHT(rectangle2_weights[2666]), .RECT3_X(rectangle3_xs[2666]), .RECT3_Y(rectangle3_ys[2666]), .RECT3_WIDTH(rectangle3_widths[2666]), .RECT3_HEIGHT(rectangle3_heights[2666]), .RECT3_WEIGHT(rectangle3_weights[2666]), .FEAT_THRES(feature_thresholds[2666]), .FEAT_ABOVE(feature_aboves[2666]), .FEAT_BELOW(feature_belows[2666])) ac2666(.scan_win(scan_win2666), .scan_win_std_dev(scan_win_std_dev[2666]), .feature_accum(feature_accums[2666]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2667]), .RECT1_Y(rectangle1_ys[2667]), .RECT1_WIDTH(rectangle1_widths[2667]), .RECT1_HEIGHT(rectangle1_heights[2667]), .RECT1_WEIGHT(rectangle1_weights[2667]), .RECT2_X(rectangle2_xs[2667]), .RECT2_Y(rectangle2_ys[2667]), .RECT2_WIDTH(rectangle2_widths[2667]), .RECT2_HEIGHT(rectangle2_heights[2667]), .RECT2_WEIGHT(rectangle2_weights[2667]), .RECT3_X(rectangle3_xs[2667]), .RECT3_Y(rectangle3_ys[2667]), .RECT3_WIDTH(rectangle3_widths[2667]), .RECT3_HEIGHT(rectangle3_heights[2667]), .RECT3_WEIGHT(rectangle3_weights[2667]), .FEAT_THRES(feature_thresholds[2667]), .FEAT_ABOVE(feature_aboves[2667]), .FEAT_BELOW(feature_belows[2667])) ac2667(.scan_win(scan_win2667), .scan_win_std_dev(scan_win_std_dev[2667]), .feature_accum(feature_accums[2667]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2668]), .RECT1_Y(rectangle1_ys[2668]), .RECT1_WIDTH(rectangle1_widths[2668]), .RECT1_HEIGHT(rectangle1_heights[2668]), .RECT1_WEIGHT(rectangle1_weights[2668]), .RECT2_X(rectangle2_xs[2668]), .RECT2_Y(rectangle2_ys[2668]), .RECT2_WIDTH(rectangle2_widths[2668]), .RECT2_HEIGHT(rectangle2_heights[2668]), .RECT2_WEIGHT(rectangle2_weights[2668]), .RECT3_X(rectangle3_xs[2668]), .RECT3_Y(rectangle3_ys[2668]), .RECT3_WIDTH(rectangle3_widths[2668]), .RECT3_HEIGHT(rectangle3_heights[2668]), .RECT3_WEIGHT(rectangle3_weights[2668]), .FEAT_THRES(feature_thresholds[2668]), .FEAT_ABOVE(feature_aboves[2668]), .FEAT_BELOW(feature_belows[2668])) ac2668(.scan_win(scan_win2668), .scan_win_std_dev(scan_win_std_dev[2668]), .feature_accum(feature_accums[2668]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2669]), .RECT1_Y(rectangle1_ys[2669]), .RECT1_WIDTH(rectangle1_widths[2669]), .RECT1_HEIGHT(rectangle1_heights[2669]), .RECT1_WEIGHT(rectangle1_weights[2669]), .RECT2_X(rectangle2_xs[2669]), .RECT2_Y(rectangle2_ys[2669]), .RECT2_WIDTH(rectangle2_widths[2669]), .RECT2_HEIGHT(rectangle2_heights[2669]), .RECT2_WEIGHT(rectangle2_weights[2669]), .RECT3_X(rectangle3_xs[2669]), .RECT3_Y(rectangle3_ys[2669]), .RECT3_WIDTH(rectangle3_widths[2669]), .RECT3_HEIGHT(rectangle3_heights[2669]), .RECT3_WEIGHT(rectangle3_weights[2669]), .FEAT_THRES(feature_thresholds[2669]), .FEAT_ABOVE(feature_aboves[2669]), .FEAT_BELOW(feature_belows[2669])) ac2669(.scan_win(scan_win2669), .scan_win_std_dev(scan_win_std_dev[2669]), .feature_accum(feature_accums[2669]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2670]), .RECT1_Y(rectangle1_ys[2670]), .RECT1_WIDTH(rectangle1_widths[2670]), .RECT1_HEIGHT(rectangle1_heights[2670]), .RECT1_WEIGHT(rectangle1_weights[2670]), .RECT2_X(rectangle2_xs[2670]), .RECT2_Y(rectangle2_ys[2670]), .RECT2_WIDTH(rectangle2_widths[2670]), .RECT2_HEIGHT(rectangle2_heights[2670]), .RECT2_WEIGHT(rectangle2_weights[2670]), .RECT3_X(rectangle3_xs[2670]), .RECT3_Y(rectangle3_ys[2670]), .RECT3_WIDTH(rectangle3_widths[2670]), .RECT3_HEIGHT(rectangle3_heights[2670]), .RECT3_WEIGHT(rectangle3_weights[2670]), .FEAT_THRES(feature_thresholds[2670]), .FEAT_ABOVE(feature_aboves[2670]), .FEAT_BELOW(feature_belows[2670])) ac2670(.scan_win(scan_win2670), .scan_win_std_dev(scan_win_std_dev[2670]), .feature_accum(feature_accums[2670]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2671]), .RECT1_Y(rectangle1_ys[2671]), .RECT1_WIDTH(rectangle1_widths[2671]), .RECT1_HEIGHT(rectangle1_heights[2671]), .RECT1_WEIGHT(rectangle1_weights[2671]), .RECT2_X(rectangle2_xs[2671]), .RECT2_Y(rectangle2_ys[2671]), .RECT2_WIDTH(rectangle2_widths[2671]), .RECT2_HEIGHT(rectangle2_heights[2671]), .RECT2_WEIGHT(rectangle2_weights[2671]), .RECT3_X(rectangle3_xs[2671]), .RECT3_Y(rectangle3_ys[2671]), .RECT3_WIDTH(rectangle3_widths[2671]), .RECT3_HEIGHT(rectangle3_heights[2671]), .RECT3_WEIGHT(rectangle3_weights[2671]), .FEAT_THRES(feature_thresholds[2671]), .FEAT_ABOVE(feature_aboves[2671]), .FEAT_BELOW(feature_belows[2671])) ac2671(.scan_win(scan_win2671), .scan_win_std_dev(scan_win_std_dev[2671]), .feature_accum(feature_accums[2671]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2672]), .RECT1_Y(rectangle1_ys[2672]), .RECT1_WIDTH(rectangle1_widths[2672]), .RECT1_HEIGHT(rectangle1_heights[2672]), .RECT1_WEIGHT(rectangle1_weights[2672]), .RECT2_X(rectangle2_xs[2672]), .RECT2_Y(rectangle2_ys[2672]), .RECT2_WIDTH(rectangle2_widths[2672]), .RECT2_HEIGHT(rectangle2_heights[2672]), .RECT2_WEIGHT(rectangle2_weights[2672]), .RECT3_X(rectangle3_xs[2672]), .RECT3_Y(rectangle3_ys[2672]), .RECT3_WIDTH(rectangle3_widths[2672]), .RECT3_HEIGHT(rectangle3_heights[2672]), .RECT3_WEIGHT(rectangle3_weights[2672]), .FEAT_THRES(feature_thresholds[2672]), .FEAT_ABOVE(feature_aboves[2672]), .FEAT_BELOW(feature_belows[2672])) ac2672(.scan_win(scan_win2672), .scan_win_std_dev(scan_win_std_dev[2672]), .feature_accum(feature_accums[2672]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2673]), .RECT1_Y(rectangle1_ys[2673]), .RECT1_WIDTH(rectangle1_widths[2673]), .RECT1_HEIGHT(rectangle1_heights[2673]), .RECT1_WEIGHT(rectangle1_weights[2673]), .RECT2_X(rectangle2_xs[2673]), .RECT2_Y(rectangle2_ys[2673]), .RECT2_WIDTH(rectangle2_widths[2673]), .RECT2_HEIGHT(rectangle2_heights[2673]), .RECT2_WEIGHT(rectangle2_weights[2673]), .RECT3_X(rectangle3_xs[2673]), .RECT3_Y(rectangle3_ys[2673]), .RECT3_WIDTH(rectangle3_widths[2673]), .RECT3_HEIGHT(rectangle3_heights[2673]), .RECT3_WEIGHT(rectangle3_weights[2673]), .FEAT_THRES(feature_thresholds[2673]), .FEAT_ABOVE(feature_aboves[2673]), .FEAT_BELOW(feature_belows[2673])) ac2673(.scan_win(scan_win2673), .scan_win_std_dev(scan_win_std_dev[2673]), .feature_accum(feature_accums[2673]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2674]), .RECT1_Y(rectangle1_ys[2674]), .RECT1_WIDTH(rectangle1_widths[2674]), .RECT1_HEIGHT(rectangle1_heights[2674]), .RECT1_WEIGHT(rectangle1_weights[2674]), .RECT2_X(rectangle2_xs[2674]), .RECT2_Y(rectangle2_ys[2674]), .RECT2_WIDTH(rectangle2_widths[2674]), .RECT2_HEIGHT(rectangle2_heights[2674]), .RECT2_WEIGHT(rectangle2_weights[2674]), .RECT3_X(rectangle3_xs[2674]), .RECT3_Y(rectangle3_ys[2674]), .RECT3_WIDTH(rectangle3_widths[2674]), .RECT3_HEIGHT(rectangle3_heights[2674]), .RECT3_WEIGHT(rectangle3_weights[2674]), .FEAT_THRES(feature_thresholds[2674]), .FEAT_ABOVE(feature_aboves[2674]), .FEAT_BELOW(feature_belows[2674])) ac2674(.scan_win(scan_win2674), .scan_win_std_dev(scan_win_std_dev[2674]), .feature_accum(feature_accums[2674]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2675]), .RECT1_Y(rectangle1_ys[2675]), .RECT1_WIDTH(rectangle1_widths[2675]), .RECT1_HEIGHT(rectangle1_heights[2675]), .RECT1_WEIGHT(rectangle1_weights[2675]), .RECT2_X(rectangle2_xs[2675]), .RECT2_Y(rectangle2_ys[2675]), .RECT2_WIDTH(rectangle2_widths[2675]), .RECT2_HEIGHT(rectangle2_heights[2675]), .RECT2_WEIGHT(rectangle2_weights[2675]), .RECT3_X(rectangle3_xs[2675]), .RECT3_Y(rectangle3_ys[2675]), .RECT3_WIDTH(rectangle3_widths[2675]), .RECT3_HEIGHT(rectangle3_heights[2675]), .RECT3_WEIGHT(rectangle3_weights[2675]), .FEAT_THRES(feature_thresholds[2675]), .FEAT_ABOVE(feature_aboves[2675]), .FEAT_BELOW(feature_belows[2675])) ac2675(.scan_win(scan_win2675), .scan_win_std_dev(scan_win_std_dev[2675]), .feature_accum(feature_accums[2675]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2676]), .RECT1_Y(rectangle1_ys[2676]), .RECT1_WIDTH(rectangle1_widths[2676]), .RECT1_HEIGHT(rectangle1_heights[2676]), .RECT1_WEIGHT(rectangle1_weights[2676]), .RECT2_X(rectangle2_xs[2676]), .RECT2_Y(rectangle2_ys[2676]), .RECT2_WIDTH(rectangle2_widths[2676]), .RECT2_HEIGHT(rectangle2_heights[2676]), .RECT2_WEIGHT(rectangle2_weights[2676]), .RECT3_X(rectangle3_xs[2676]), .RECT3_Y(rectangle3_ys[2676]), .RECT3_WIDTH(rectangle3_widths[2676]), .RECT3_HEIGHT(rectangle3_heights[2676]), .RECT3_WEIGHT(rectangle3_weights[2676]), .FEAT_THRES(feature_thresholds[2676]), .FEAT_ABOVE(feature_aboves[2676]), .FEAT_BELOW(feature_belows[2676])) ac2676(.scan_win(scan_win2676), .scan_win_std_dev(scan_win_std_dev[2676]), .feature_accum(feature_accums[2676]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2677]), .RECT1_Y(rectangle1_ys[2677]), .RECT1_WIDTH(rectangle1_widths[2677]), .RECT1_HEIGHT(rectangle1_heights[2677]), .RECT1_WEIGHT(rectangle1_weights[2677]), .RECT2_X(rectangle2_xs[2677]), .RECT2_Y(rectangle2_ys[2677]), .RECT2_WIDTH(rectangle2_widths[2677]), .RECT2_HEIGHT(rectangle2_heights[2677]), .RECT2_WEIGHT(rectangle2_weights[2677]), .RECT3_X(rectangle3_xs[2677]), .RECT3_Y(rectangle3_ys[2677]), .RECT3_WIDTH(rectangle3_widths[2677]), .RECT3_HEIGHT(rectangle3_heights[2677]), .RECT3_WEIGHT(rectangle3_weights[2677]), .FEAT_THRES(feature_thresholds[2677]), .FEAT_ABOVE(feature_aboves[2677]), .FEAT_BELOW(feature_belows[2677])) ac2677(.scan_win(scan_win2677), .scan_win_std_dev(scan_win_std_dev[2677]), .feature_accum(feature_accums[2677]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2678]), .RECT1_Y(rectangle1_ys[2678]), .RECT1_WIDTH(rectangle1_widths[2678]), .RECT1_HEIGHT(rectangle1_heights[2678]), .RECT1_WEIGHT(rectangle1_weights[2678]), .RECT2_X(rectangle2_xs[2678]), .RECT2_Y(rectangle2_ys[2678]), .RECT2_WIDTH(rectangle2_widths[2678]), .RECT2_HEIGHT(rectangle2_heights[2678]), .RECT2_WEIGHT(rectangle2_weights[2678]), .RECT3_X(rectangle3_xs[2678]), .RECT3_Y(rectangle3_ys[2678]), .RECT3_WIDTH(rectangle3_widths[2678]), .RECT3_HEIGHT(rectangle3_heights[2678]), .RECT3_WEIGHT(rectangle3_weights[2678]), .FEAT_THRES(feature_thresholds[2678]), .FEAT_ABOVE(feature_aboves[2678]), .FEAT_BELOW(feature_belows[2678])) ac2678(.scan_win(scan_win2678), .scan_win_std_dev(scan_win_std_dev[2678]), .feature_accum(feature_accums[2678]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2679]), .RECT1_Y(rectangle1_ys[2679]), .RECT1_WIDTH(rectangle1_widths[2679]), .RECT1_HEIGHT(rectangle1_heights[2679]), .RECT1_WEIGHT(rectangle1_weights[2679]), .RECT2_X(rectangle2_xs[2679]), .RECT2_Y(rectangle2_ys[2679]), .RECT2_WIDTH(rectangle2_widths[2679]), .RECT2_HEIGHT(rectangle2_heights[2679]), .RECT2_WEIGHT(rectangle2_weights[2679]), .RECT3_X(rectangle3_xs[2679]), .RECT3_Y(rectangle3_ys[2679]), .RECT3_WIDTH(rectangle3_widths[2679]), .RECT3_HEIGHT(rectangle3_heights[2679]), .RECT3_WEIGHT(rectangle3_weights[2679]), .FEAT_THRES(feature_thresholds[2679]), .FEAT_ABOVE(feature_aboves[2679]), .FEAT_BELOW(feature_belows[2679])) ac2679(.scan_win(scan_win2679), .scan_win_std_dev(scan_win_std_dev[2679]), .feature_accum(feature_accums[2679]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2680]), .RECT1_Y(rectangle1_ys[2680]), .RECT1_WIDTH(rectangle1_widths[2680]), .RECT1_HEIGHT(rectangle1_heights[2680]), .RECT1_WEIGHT(rectangle1_weights[2680]), .RECT2_X(rectangle2_xs[2680]), .RECT2_Y(rectangle2_ys[2680]), .RECT2_WIDTH(rectangle2_widths[2680]), .RECT2_HEIGHT(rectangle2_heights[2680]), .RECT2_WEIGHT(rectangle2_weights[2680]), .RECT3_X(rectangle3_xs[2680]), .RECT3_Y(rectangle3_ys[2680]), .RECT3_WIDTH(rectangle3_widths[2680]), .RECT3_HEIGHT(rectangle3_heights[2680]), .RECT3_WEIGHT(rectangle3_weights[2680]), .FEAT_THRES(feature_thresholds[2680]), .FEAT_ABOVE(feature_aboves[2680]), .FEAT_BELOW(feature_belows[2680])) ac2680(.scan_win(scan_win2680), .scan_win_std_dev(scan_win_std_dev[2680]), .feature_accum(feature_accums[2680]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2681]), .RECT1_Y(rectangle1_ys[2681]), .RECT1_WIDTH(rectangle1_widths[2681]), .RECT1_HEIGHT(rectangle1_heights[2681]), .RECT1_WEIGHT(rectangle1_weights[2681]), .RECT2_X(rectangle2_xs[2681]), .RECT2_Y(rectangle2_ys[2681]), .RECT2_WIDTH(rectangle2_widths[2681]), .RECT2_HEIGHT(rectangle2_heights[2681]), .RECT2_WEIGHT(rectangle2_weights[2681]), .RECT3_X(rectangle3_xs[2681]), .RECT3_Y(rectangle3_ys[2681]), .RECT3_WIDTH(rectangle3_widths[2681]), .RECT3_HEIGHT(rectangle3_heights[2681]), .RECT3_WEIGHT(rectangle3_weights[2681]), .FEAT_THRES(feature_thresholds[2681]), .FEAT_ABOVE(feature_aboves[2681]), .FEAT_BELOW(feature_belows[2681])) ac2681(.scan_win(scan_win2681), .scan_win_std_dev(scan_win_std_dev[2681]), .feature_accum(feature_accums[2681]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2682]), .RECT1_Y(rectangle1_ys[2682]), .RECT1_WIDTH(rectangle1_widths[2682]), .RECT1_HEIGHT(rectangle1_heights[2682]), .RECT1_WEIGHT(rectangle1_weights[2682]), .RECT2_X(rectangle2_xs[2682]), .RECT2_Y(rectangle2_ys[2682]), .RECT2_WIDTH(rectangle2_widths[2682]), .RECT2_HEIGHT(rectangle2_heights[2682]), .RECT2_WEIGHT(rectangle2_weights[2682]), .RECT3_X(rectangle3_xs[2682]), .RECT3_Y(rectangle3_ys[2682]), .RECT3_WIDTH(rectangle3_widths[2682]), .RECT3_HEIGHT(rectangle3_heights[2682]), .RECT3_WEIGHT(rectangle3_weights[2682]), .FEAT_THRES(feature_thresholds[2682]), .FEAT_ABOVE(feature_aboves[2682]), .FEAT_BELOW(feature_belows[2682])) ac2682(.scan_win(scan_win2682), .scan_win_std_dev(scan_win_std_dev[2682]), .feature_accum(feature_accums[2682]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2683]), .RECT1_Y(rectangle1_ys[2683]), .RECT1_WIDTH(rectangle1_widths[2683]), .RECT1_HEIGHT(rectangle1_heights[2683]), .RECT1_WEIGHT(rectangle1_weights[2683]), .RECT2_X(rectangle2_xs[2683]), .RECT2_Y(rectangle2_ys[2683]), .RECT2_WIDTH(rectangle2_widths[2683]), .RECT2_HEIGHT(rectangle2_heights[2683]), .RECT2_WEIGHT(rectangle2_weights[2683]), .RECT3_X(rectangle3_xs[2683]), .RECT3_Y(rectangle3_ys[2683]), .RECT3_WIDTH(rectangle3_widths[2683]), .RECT3_HEIGHT(rectangle3_heights[2683]), .RECT3_WEIGHT(rectangle3_weights[2683]), .FEAT_THRES(feature_thresholds[2683]), .FEAT_ABOVE(feature_aboves[2683]), .FEAT_BELOW(feature_belows[2683])) ac2683(.scan_win(scan_win2683), .scan_win_std_dev(scan_win_std_dev[2683]), .feature_accum(feature_accums[2683]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2684]), .RECT1_Y(rectangle1_ys[2684]), .RECT1_WIDTH(rectangle1_widths[2684]), .RECT1_HEIGHT(rectangle1_heights[2684]), .RECT1_WEIGHT(rectangle1_weights[2684]), .RECT2_X(rectangle2_xs[2684]), .RECT2_Y(rectangle2_ys[2684]), .RECT2_WIDTH(rectangle2_widths[2684]), .RECT2_HEIGHT(rectangle2_heights[2684]), .RECT2_WEIGHT(rectangle2_weights[2684]), .RECT3_X(rectangle3_xs[2684]), .RECT3_Y(rectangle3_ys[2684]), .RECT3_WIDTH(rectangle3_widths[2684]), .RECT3_HEIGHT(rectangle3_heights[2684]), .RECT3_WEIGHT(rectangle3_weights[2684]), .FEAT_THRES(feature_thresholds[2684]), .FEAT_ABOVE(feature_aboves[2684]), .FEAT_BELOW(feature_belows[2684])) ac2684(.scan_win(scan_win2684), .scan_win_std_dev(scan_win_std_dev[2684]), .feature_accum(feature_accums[2684]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2685]), .RECT1_Y(rectangle1_ys[2685]), .RECT1_WIDTH(rectangle1_widths[2685]), .RECT1_HEIGHT(rectangle1_heights[2685]), .RECT1_WEIGHT(rectangle1_weights[2685]), .RECT2_X(rectangle2_xs[2685]), .RECT2_Y(rectangle2_ys[2685]), .RECT2_WIDTH(rectangle2_widths[2685]), .RECT2_HEIGHT(rectangle2_heights[2685]), .RECT2_WEIGHT(rectangle2_weights[2685]), .RECT3_X(rectangle3_xs[2685]), .RECT3_Y(rectangle3_ys[2685]), .RECT3_WIDTH(rectangle3_widths[2685]), .RECT3_HEIGHT(rectangle3_heights[2685]), .RECT3_WEIGHT(rectangle3_weights[2685]), .FEAT_THRES(feature_thresholds[2685]), .FEAT_ABOVE(feature_aboves[2685]), .FEAT_BELOW(feature_belows[2685])) ac2685(.scan_win(scan_win2685), .scan_win_std_dev(scan_win_std_dev[2685]), .feature_accum(feature_accums[2685]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2686]), .RECT1_Y(rectangle1_ys[2686]), .RECT1_WIDTH(rectangle1_widths[2686]), .RECT1_HEIGHT(rectangle1_heights[2686]), .RECT1_WEIGHT(rectangle1_weights[2686]), .RECT2_X(rectangle2_xs[2686]), .RECT2_Y(rectangle2_ys[2686]), .RECT2_WIDTH(rectangle2_widths[2686]), .RECT2_HEIGHT(rectangle2_heights[2686]), .RECT2_WEIGHT(rectangle2_weights[2686]), .RECT3_X(rectangle3_xs[2686]), .RECT3_Y(rectangle3_ys[2686]), .RECT3_WIDTH(rectangle3_widths[2686]), .RECT3_HEIGHT(rectangle3_heights[2686]), .RECT3_WEIGHT(rectangle3_weights[2686]), .FEAT_THRES(feature_thresholds[2686]), .FEAT_ABOVE(feature_aboves[2686]), .FEAT_BELOW(feature_belows[2686])) ac2686(.scan_win(scan_win2686), .scan_win_std_dev(scan_win_std_dev[2686]), .feature_accum(feature_accums[2686]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2687]), .RECT1_Y(rectangle1_ys[2687]), .RECT1_WIDTH(rectangle1_widths[2687]), .RECT1_HEIGHT(rectangle1_heights[2687]), .RECT1_WEIGHT(rectangle1_weights[2687]), .RECT2_X(rectangle2_xs[2687]), .RECT2_Y(rectangle2_ys[2687]), .RECT2_WIDTH(rectangle2_widths[2687]), .RECT2_HEIGHT(rectangle2_heights[2687]), .RECT2_WEIGHT(rectangle2_weights[2687]), .RECT3_X(rectangle3_xs[2687]), .RECT3_Y(rectangle3_ys[2687]), .RECT3_WIDTH(rectangle3_widths[2687]), .RECT3_HEIGHT(rectangle3_heights[2687]), .RECT3_WEIGHT(rectangle3_weights[2687]), .FEAT_THRES(feature_thresholds[2687]), .FEAT_ABOVE(feature_aboves[2687]), .FEAT_BELOW(feature_belows[2687])) ac2687(.scan_win(scan_win2687), .scan_win_std_dev(scan_win_std_dev[2687]), .feature_accum(feature_accums[2687]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2688]), .RECT1_Y(rectangle1_ys[2688]), .RECT1_WIDTH(rectangle1_widths[2688]), .RECT1_HEIGHT(rectangle1_heights[2688]), .RECT1_WEIGHT(rectangle1_weights[2688]), .RECT2_X(rectangle2_xs[2688]), .RECT2_Y(rectangle2_ys[2688]), .RECT2_WIDTH(rectangle2_widths[2688]), .RECT2_HEIGHT(rectangle2_heights[2688]), .RECT2_WEIGHT(rectangle2_weights[2688]), .RECT3_X(rectangle3_xs[2688]), .RECT3_Y(rectangle3_ys[2688]), .RECT3_WIDTH(rectangle3_widths[2688]), .RECT3_HEIGHT(rectangle3_heights[2688]), .RECT3_WEIGHT(rectangle3_weights[2688]), .FEAT_THRES(feature_thresholds[2688]), .FEAT_ABOVE(feature_aboves[2688]), .FEAT_BELOW(feature_belows[2688])) ac2688(.scan_win(scan_win2688), .scan_win_std_dev(scan_win_std_dev[2688]), .feature_accum(feature_accums[2688]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2689]), .RECT1_Y(rectangle1_ys[2689]), .RECT1_WIDTH(rectangle1_widths[2689]), .RECT1_HEIGHT(rectangle1_heights[2689]), .RECT1_WEIGHT(rectangle1_weights[2689]), .RECT2_X(rectangle2_xs[2689]), .RECT2_Y(rectangle2_ys[2689]), .RECT2_WIDTH(rectangle2_widths[2689]), .RECT2_HEIGHT(rectangle2_heights[2689]), .RECT2_WEIGHT(rectangle2_weights[2689]), .RECT3_X(rectangle3_xs[2689]), .RECT3_Y(rectangle3_ys[2689]), .RECT3_WIDTH(rectangle3_widths[2689]), .RECT3_HEIGHT(rectangle3_heights[2689]), .RECT3_WEIGHT(rectangle3_weights[2689]), .FEAT_THRES(feature_thresholds[2689]), .FEAT_ABOVE(feature_aboves[2689]), .FEAT_BELOW(feature_belows[2689])) ac2689(.scan_win(scan_win2689), .scan_win_std_dev(scan_win_std_dev[2689]), .feature_accum(feature_accums[2689]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2690]), .RECT1_Y(rectangle1_ys[2690]), .RECT1_WIDTH(rectangle1_widths[2690]), .RECT1_HEIGHT(rectangle1_heights[2690]), .RECT1_WEIGHT(rectangle1_weights[2690]), .RECT2_X(rectangle2_xs[2690]), .RECT2_Y(rectangle2_ys[2690]), .RECT2_WIDTH(rectangle2_widths[2690]), .RECT2_HEIGHT(rectangle2_heights[2690]), .RECT2_WEIGHT(rectangle2_weights[2690]), .RECT3_X(rectangle3_xs[2690]), .RECT3_Y(rectangle3_ys[2690]), .RECT3_WIDTH(rectangle3_widths[2690]), .RECT3_HEIGHT(rectangle3_heights[2690]), .RECT3_WEIGHT(rectangle3_weights[2690]), .FEAT_THRES(feature_thresholds[2690]), .FEAT_ABOVE(feature_aboves[2690]), .FEAT_BELOW(feature_belows[2690])) ac2690(.scan_win(scan_win2690), .scan_win_std_dev(scan_win_std_dev[2690]), .feature_accum(feature_accums[2690]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2691]), .RECT1_Y(rectangle1_ys[2691]), .RECT1_WIDTH(rectangle1_widths[2691]), .RECT1_HEIGHT(rectangle1_heights[2691]), .RECT1_WEIGHT(rectangle1_weights[2691]), .RECT2_X(rectangle2_xs[2691]), .RECT2_Y(rectangle2_ys[2691]), .RECT2_WIDTH(rectangle2_widths[2691]), .RECT2_HEIGHT(rectangle2_heights[2691]), .RECT2_WEIGHT(rectangle2_weights[2691]), .RECT3_X(rectangle3_xs[2691]), .RECT3_Y(rectangle3_ys[2691]), .RECT3_WIDTH(rectangle3_widths[2691]), .RECT3_HEIGHT(rectangle3_heights[2691]), .RECT3_WEIGHT(rectangle3_weights[2691]), .FEAT_THRES(feature_thresholds[2691]), .FEAT_ABOVE(feature_aboves[2691]), .FEAT_BELOW(feature_belows[2691])) ac2691(.scan_win(scan_win2691), .scan_win_std_dev(scan_win_std_dev[2691]), .feature_accum(feature_accums[2691]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2692]), .RECT1_Y(rectangle1_ys[2692]), .RECT1_WIDTH(rectangle1_widths[2692]), .RECT1_HEIGHT(rectangle1_heights[2692]), .RECT1_WEIGHT(rectangle1_weights[2692]), .RECT2_X(rectangle2_xs[2692]), .RECT2_Y(rectangle2_ys[2692]), .RECT2_WIDTH(rectangle2_widths[2692]), .RECT2_HEIGHT(rectangle2_heights[2692]), .RECT2_WEIGHT(rectangle2_weights[2692]), .RECT3_X(rectangle3_xs[2692]), .RECT3_Y(rectangle3_ys[2692]), .RECT3_WIDTH(rectangle3_widths[2692]), .RECT3_HEIGHT(rectangle3_heights[2692]), .RECT3_WEIGHT(rectangle3_weights[2692]), .FEAT_THRES(feature_thresholds[2692]), .FEAT_ABOVE(feature_aboves[2692]), .FEAT_BELOW(feature_belows[2692])) ac2692(.scan_win(scan_win2692), .scan_win_std_dev(scan_win_std_dev[2692]), .feature_accum(feature_accums[2692]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2693]), .RECT1_Y(rectangle1_ys[2693]), .RECT1_WIDTH(rectangle1_widths[2693]), .RECT1_HEIGHT(rectangle1_heights[2693]), .RECT1_WEIGHT(rectangle1_weights[2693]), .RECT2_X(rectangle2_xs[2693]), .RECT2_Y(rectangle2_ys[2693]), .RECT2_WIDTH(rectangle2_widths[2693]), .RECT2_HEIGHT(rectangle2_heights[2693]), .RECT2_WEIGHT(rectangle2_weights[2693]), .RECT3_X(rectangle3_xs[2693]), .RECT3_Y(rectangle3_ys[2693]), .RECT3_WIDTH(rectangle3_widths[2693]), .RECT3_HEIGHT(rectangle3_heights[2693]), .RECT3_WEIGHT(rectangle3_weights[2693]), .FEAT_THRES(feature_thresholds[2693]), .FEAT_ABOVE(feature_aboves[2693]), .FEAT_BELOW(feature_belows[2693])) ac2693(.scan_win(scan_win2693), .scan_win_std_dev(scan_win_std_dev[2693]), .feature_accum(feature_accums[2693]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2694]), .RECT1_Y(rectangle1_ys[2694]), .RECT1_WIDTH(rectangle1_widths[2694]), .RECT1_HEIGHT(rectangle1_heights[2694]), .RECT1_WEIGHT(rectangle1_weights[2694]), .RECT2_X(rectangle2_xs[2694]), .RECT2_Y(rectangle2_ys[2694]), .RECT2_WIDTH(rectangle2_widths[2694]), .RECT2_HEIGHT(rectangle2_heights[2694]), .RECT2_WEIGHT(rectangle2_weights[2694]), .RECT3_X(rectangle3_xs[2694]), .RECT3_Y(rectangle3_ys[2694]), .RECT3_WIDTH(rectangle3_widths[2694]), .RECT3_HEIGHT(rectangle3_heights[2694]), .RECT3_WEIGHT(rectangle3_weights[2694]), .FEAT_THRES(feature_thresholds[2694]), .FEAT_ABOVE(feature_aboves[2694]), .FEAT_BELOW(feature_belows[2694])) ac2694(.scan_win(scan_win2694), .scan_win_std_dev(scan_win_std_dev[2694]), .feature_accum(feature_accums[2694]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2695]), .RECT1_Y(rectangle1_ys[2695]), .RECT1_WIDTH(rectangle1_widths[2695]), .RECT1_HEIGHT(rectangle1_heights[2695]), .RECT1_WEIGHT(rectangle1_weights[2695]), .RECT2_X(rectangle2_xs[2695]), .RECT2_Y(rectangle2_ys[2695]), .RECT2_WIDTH(rectangle2_widths[2695]), .RECT2_HEIGHT(rectangle2_heights[2695]), .RECT2_WEIGHT(rectangle2_weights[2695]), .RECT3_X(rectangle3_xs[2695]), .RECT3_Y(rectangle3_ys[2695]), .RECT3_WIDTH(rectangle3_widths[2695]), .RECT3_HEIGHT(rectangle3_heights[2695]), .RECT3_WEIGHT(rectangle3_weights[2695]), .FEAT_THRES(feature_thresholds[2695]), .FEAT_ABOVE(feature_aboves[2695]), .FEAT_BELOW(feature_belows[2695])) ac2695(.scan_win(scan_win2695), .scan_win_std_dev(scan_win_std_dev[2695]), .feature_accum(feature_accums[2695]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2696]), .RECT1_Y(rectangle1_ys[2696]), .RECT1_WIDTH(rectangle1_widths[2696]), .RECT1_HEIGHT(rectangle1_heights[2696]), .RECT1_WEIGHT(rectangle1_weights[2696]), .RECT2_X(rectangle2_xs[2696]), .RECT2_Y(rectangle2_ys[2696]), .RECT2_WIDTH(rectangle2_widths[2696]), .RECT2_HEIGHT(rectangle2_heights[2696]), .RECT2_WEIGHT(rectangle2_weights[2696]), .RECT3_X(rectangle3_xs[2696]), .RECT3_Y(rectangle3_ys[2696]), .RECT3_WIDTH(rectangle3_widths[2696]), .RECT3_HEIGHT(rectangle3_heights[2696]), .RECT3_WEIGHT(rectangle3_weights[2696]), .FEAT_THRES(feature_thresholds[2696]), .FEAT_ABOVE(feature_aboves[2696]), .FEAT_BELOW(feature_belows[2696])) ac2696(.scan_win(scan_win2696), .scan_win_std_dev(scan_win_std_dev[2696]), .feature_accum(feature_accums[2696]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2697]), .RECT1_Y(rectangle1_ys[2697]), .RECT1_WIDTH(rectangle1_widths[2697]), .RECT1_HEIGHT(rectangle1_heights[2697]), .RECT1_WEIGHT(rectangle1_weights[2697]), .RECT2_X(rectangle2_xs[2697]), .RECT2_Y(rectangle2_ys[2697]), .RECT2_WIDTH(rectangle2_widths[2697]), .RECT2_HEIGHT(rectangle2_heights[2697]), .RECT2_WEIGHT(rectangle2_weights[2697]), .RECT3_X(rectangle3_xs[2697]), .RECT3_Y(rectangle3_ys[2697]), .RECT3_WIDTH(rectangle3_widths[2697]), .RECT3_HEIGHT(rectangle3_heights[2697]), .RECT3_WEIGHT(rectangle3_weights[2697]), .FEAT_THRES(feature_thresholds[2697]), .FEAT_ABOVE(feature_aboves[2697]), .FEAT_BELOW(feature_belows[2697])) ac2697(.scan_win(scan_win2697), .scan_win_std_dev(scan_win_std_dev[2697]), .feature_accum(feature_accums[2697]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2698]), .RECT1_Y(rectangle1_ys[2698]), .RECT1_WIDTH(rectangle1_widths[2698]), .RECT1_HEIGHT(rectangle1_heights[2698]), .RECT1_WEIGHT(rectangle1_weights[2698]), .RECT2_X(rectangle2_xs[2698]), .RECT2_Y(rectangle2_ys[2698]), .RECT2_WIDTH(rectangle2_widths[2698]), .RECT2_HEIGHT(rectangle2_heights[2698]), .RECT2_WEIGHT(rectangle2_weights[2698]), .RECT3_X(rectangle3_xs[2698]), .RECT3_Y(rectangle3_ys[2698]), .RECT3_WIDTH(rectangle3_widths[2698]), .RECT3_HEIGHT(rectangle3_heights[2698]), .RECT3_WEIGHT(rectangle3_weights[2698]), .FEAT_THRES(feature_thresholds[2698]), .FEAT_ABOVE(feature_aboves[2698]), .FEAT_BELOW(feature_belows[2698])) ac2698(.scan_win(scan_win2698), .scan_win_std_dev(scan_win_std_dev[2698]), .feature_accum(feature_accums[2698]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2699]), .RECT1_Y(rectangle1_ys[2699]), .RECT1_WIDTH(rectangle1_widths[2699]), .RECT1_HEIGHT(rectangle1_heights[2699]), .RECT1_WEIGHT(rectangle1_weights[2699]), .RECT2_X(rectangle2_xs[2699]), .RECT2_Y(rectangle2_ys[2699]), .RECT2_WIDTH(rectangle2_widths[2699]), .RECT2_HEIGHT(rectangle2_heights[2699]), .RECT2_WEIGHT(rectangle2_weights[2699]), .RECT3_X(rectangle3_xs[2699]), .RECT3_Y(rectangle3_ys[2699]), .RECT3_WIDTH(rectangle3_widths[2699]), .RECT3_HEIGHT(rectangle3_heights[2699]), .RECT3_WEIGHT(rectangle3_weights[2699]), .FEAT_THRES(feature_thresholds[2699]), .FEAT_ABOVE(feature_aboves[2699]), .FEAT_BELOW(feature_belows[2699])) ac2699(.scan_win(scan_win2699), .scan_win_std_dev(scan_win_std_dev[2699]), .feature_accum(feature_accums[2699]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2700]), .RECT1_Y(rectangle1_ys[2700]), .RECT1_WIDTH(rectangle1_widths[2700]), .RECT1_HEIGHT(rectangle1_heights[2700]), .RECT1_WEIGHT(rectangle1_weights[2700]), .RECT2_X(rectangle2_xs[2700]), .RECT2_Y(rectangle2_ys[2700]), .RECT2_WIDTH(rectangle2_widths[2700]), .RECT2_HEIGHT(rectangle2_heights[2700]), .RECT2_WEIGHT(rectangle2_weights[2700]), .RECT3_X(rectangle3_xs[2700]), .RECT3_Y(rectangle3_ys[2700]), .RECT3_WIDTH(rectangle3_widths[2700]), .RECT3_HEIGHT(rectangle3_heights[2700]), .RECT3_WEIGHT(rectangle3_weights[2700]), .FEAT_THRES(feature_thresholds[2700]), .FEAT_ABOVE(feature_aboves[2700]), .FEAT_BELOW(feature_belows[2700])) ac2700(.scan_win(scan_win2700), .scan_win_std_dev(scan_win_std_dev[2700]), .feature_accum(feature_accums[2700]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2701]), .RECT1_Y(rectangle1_ys[2701]), .RECT1_WIDTH(rectangle1_widths[2701]), .RECT1_HEIGHT(rectangle1_heights[2701]), .RECT1_WEIGHT(rectangle1_weights[2701]), .RECT2_X(rectangle2_xs[2701]), .RECT2_Y(rectangle2_ys[2701]), .RECT2_WIDTH(rectangle2_widths[2701]), .RECT2_HEIGHT(rectangle2_heights[2701]), .RECT2_WEIGHT(rectangle2_weights[2701]), .RECT3_X(rectangle3_xs[2701]), .RECT3_Y(rectangle3_ys[2701]), .RECT3_WIDTH(rectangle3_widths[2701]), .RECT3_HEIGHT(rectangle3_heights[2701]), .RECT3_WEIGHT(rectangle3_weights[2701]), .FEAT_THRES(feature_thresholds[2701]), .FEAT_ABOVE(feature_aboves[2701]), .FEAT_BELOW(feature_belows[2701])) ac2701(.scan_win(scan_win2701), .scan_win_std_dev(scan_win_std_dev[2701]), .feature_accum(feature_accums[2701]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2702]), .RECT1_Y(rectangle1_ys[2702]), .RECT1_WIDTH(rectangle1_widths[2702]), .RECT1_HEIGHT(rectangle1_heights[2702]), .RECT1_WEIGHT(rectangle1_weights[2702]), .RECT2_X(rectangle2_xs[2702]), .RECT2_Y(rectangle2_ys[2702]), .RECT2_WIDTH(rectangle2_widths[2702]), .RECT2_HEIGHT(rectangle2_heights[2702]), .RECT2_WEIGHT(rectangle2_weights[2702]), .RECT3_X(rectangle3_xs[2702]), .RECT3_Y(rectangle3_ys[2702]), .RECT3_WIDTH(rectangle3_widths[2702]), .RECT3_HEIGHT(rectangle3_heights[2702]), .RECT3_WEIGHT(rectangle3_weights[2702]), .FEAT_THRES(feature_thresholds[2702]), .FEAT_ABOVE(feature_aboves[2702]), .FEAT_BELOW(feature_belows[2702])) ac2702(.scan_win(scan_win2702), .scan_win_std_dev(scan_win_std_dev[2702]), .feature_accum(feature_accums[2702]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2703]), .RECT1_Y(rectangle1_ys[2703]), .RECT1_WIDTH(rectangle1_widths[2703]), .RECT1_HEIGHT(rectangle1_heights[2703]), .RECT1_WEIGHT(rectangle1_weights[2703]), .RECT2_X(rectangle2_xs[2703]), .RECT2_Y(rectangle2_ys[2703]), .RECT2_WIDTH(rectangle2_widths[2703]), .RECT2_HEIGHT(rectangle2_heights[2703]), .RECT2_WEIGHT(rectangle2_weights[2703]), .RECT3_X(rectangle3_xs[2703]), .RECT3_Y(rectangle3_ys[2703]), .RECT3_WIDTH(rectangle3_widths[2703]), .RECT3_HEIGHT(rectangle3_heights[2703]), .RECT3_WEIGHT(rectangle3_weights[2703]), .FEAT_THRES(feature_thresholds[2703]), .FEAT_ABOVE(feature_aboves[2703]), .FEAT_BELOW(feature_belows[2703])) ac2703(.scan_win(scan_win2703), .scan_win_std_dev(scan_win_std_dev[2703]), .feature_accum(feature_accums[2703]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2704]), .RECT1_Y(rectangle1_ys[2704]), .RECT1_WIDTH(rectangle1_widths[2704]), .RECT1_HEIGHT(rectangle1_heights[2704]), .RECT1_WEIGHT(rectangle1_weights[2704]), .RECT2_X(rectangle2_xs[2704]), .RECT2_Y(rectangle2_ys[2704]), .RECT2_WIDTH(rectangle2_widths[2704]), .RECT2_HEIGHT(rectangle2_heights[2704]), .RECT2_WEIGHT(rectangle2_weights[2704]), .RECT3_X(rectangle3_xs[2704]), .RECT3_Y(rectangle3_ys[2704]), .RECT3_WIDTH(rectangle3_widths[2704]), .RECT3_HEIGHT(rectangle3_heights[2704]), .RECT3_WEIGHT(rectangle3_weights[2704]), .FEAT_THRES(feature_thresholds[2704]), .FEAT_ABOVE(feature_aboves[2704]), .FEAT_BELOW(feature_belows[2704])) ac2704(.scan_win(scan_win2704), .scan_win_std_dev(scan_win_std_dev[2704]), .feature_accum(feature_accums[2704]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2705]), .RECT1_Y(rectangle1_ys[2705]), .RECT1_WIDTH(rectangle1_widths[2705]), .RECT1_HEIGHT(rectangle1_heights[2705]), .RECT1_WEIGHT(rectangle1_weights[2705]), .RECT2_X(rectangle2_xs[2705]), .RECT2_Y(rectangle2_ys[2705]), .RECT2_WIDTH(rectangle2_widths[2705]), .RECT2_HEIGHT(rectangle2_heights[2705]), .RECT2_WEIGHT(rectangle2_weights[2705]), .RECT3_X(rectangle3_xs[2705]), .RECT3_Y(rectangle3_ys[2705]), .RECT3_WIDTH(rectangle3_widths[2705]), .RECT3_HEIGHT(rectangle3_heights[2705]), .RECT3_WEIGHT(rectangle3_weights[2705]), .FEAT_THRES(feature_thresholds[2705]), .FEAT_ABOVE(feature_aboves[2705]), .FEAT_BELOW(feature_belows[2705])) ac2705(.scan_win(scan_win2705), .scan_win_std_dev(scan_win_std_dev[2705]), .feature_accum(feature_accums[2705]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2706]), .RECT1_Y(rectangle1_ys[2706]), .RECT1_WIDTH(rectangle1_widths[2706]), .RECT1_HEIGHT(rectangle1_heights[2706]), .RECT1_WEIGHT(rectangle1_weights[2706]), .RECT2_X(rectangle2_xs[2706]), .RECT2_Y(rectangle2_ys[2706]), .RECT2_WIDTH(rectangle2_widths[2706]), .RECT2_HEIGHT(rectangle2_heights[2706]), .RECT2_WEIGHT(rectangle2_weights[2706]), .RECT3_X(rectangle3_xs[2706]), .RECT3_Y(rectangle3_ys[2706]), .RECT3_WIDTH(rectangle3_widths[2706]), .RECT3_HEIGHT(rectangle3_heights[2706]), .RECT3_WEIGHT(rectangle3_weights[2706]), .FEAT_THRES(feature_thresholds[2706]), .FEAT_ABOVE(feature_aboves[2706]), .FEAT_BELOW(feature_belows[2706])) ac2706(.scan_win(scan_win2706), .scan_win_std_dev(scan_win_std_dev[2706]), .feature_accum(feature_accums[2706]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2707]), .RECT1_Y(rectangle1_ys[2707]), .RECT1_WIDTH(rectangle1_widths[2707]), .RECT1_HEIGHT(rectangle1_heights[2707]), .RECT1_WEIGHT(rectangle1_weights[2707]), .RECT2_X(rectangle2_xs[2707]), .RECT2_Y(rectangle2_ys[2707]), .RECT2_WIDTH(rectangle2_widths[2707]), .RECT2_HEIGHT(rectangle2_heights[2707]), .RECT2_WEIGHT(rectangle2_weights[2707]), .RECT3_X(rectangle3_xs[2707]), .RECT3_Y(rectangle3_ys[2707]), .RECT3_WIDTH(rectangle3_widths[2707]), .RECT3_HEIGHT(rectangle3_heights[2707]), .RECT3_WEIGHT(rectangle3_weights[2707]), .FEAT_THRES(feature_thresholds[2707]), .FEAT_ABOVE(feature_aboves[2707]), .FEAT_BELOW(feature_belows[2707])) ac2707(.scan_win(scan_win2707), .scan_win_std_dev(scan_win_std_dev[2707]), .feature_accum(feature_accums[2707]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2708]), .RECT1_Y(rectangle1_ys[2708]), .RECT1_WIDTH(rectangle1_widths[2708]), .RECT1_HEIGHT(rectangle1_heights[2708]), .RECT1_WEIGHT(rectangle1_weights[2708]), .RECT2_X(rectangle2_xs[2708]), .RECT2_Y(rectangle2_ys[2708]), .RECT2_WIDTH(rectangle2_widths[2708]), .RECT2_HEIGHT(rectangle2_heights[2708]), .RECT2_WEIGHT(rectangle2_weights[2708]), .RECT3_X(rectangle3_xs[2708]), .RECT3_Y(rectangle3_ys[2708]), .RECT3_WIDTH(rectangle3_widths[2708]), .RECT3_HEIGHT(rectangle3_heights[2708]), .RECT3_WEIGHT(rectangle3_weights[2708]), .FEAT_THRES(feature_thresholds[2708]), .FEAT_ABOVE(feature_aboves[2708]), .FEAT_BELOW(feature_belows[2708])) ac2708(.scan_win(scan_win2708), .scan_win_std_dev(scan_win_std_dev[2708]), .feature_accum(feature_accums[2708]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2709]), .RECT1_Y(rectangle1_ys[2709]), .RECT1_WIDTH(rectangle1_widths[2709]), .RECT1_HEIGHT(rectangle1_heights[2709]), .RECT1_WEIGHT(rectangle1_weights[2709]), .RECT2_X(rectangle2_xs[2709]), .RECT2_Y(rectangle2_ys[2709]), .RECT2_WIDTH(rectangle2_widths[2709]), .RECT2_HEIGHT(rectangle2_heights[2709]), .RECT2_WEIGHT(rectangle2_weights[2709]), .RECT3_X(rectangle3_xs[2709]), .RECT3_Y(rectangle3_ys[2709]), .RECT3_WIDTH(rectangle3_widths[2709]), .RECT3_HEIGHT(rectangle3_heights[2709]), .RECT3_WEIGHT(rectangle3_weights[2709]), .FEAT_THRES(feature_thresholds[2709]), .FEAT_ABOVE(feature_aboves[2709]), .FEAT_BELOW(feature_belows[2709])) ac2709(.scan_win(scan_win2709), .scan_win_std_dev(scan_win_std_dev[2709]), .feature_accum(feature_accums[2709]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2710]), .RECT1_Y(rectangle1_ys[2710]), .RECT1_WIDTH(rectangle1_widths[2710]), .RECT1_HEIGHT(rectangle1_heights[2710]), .RECT1_WEIGHT(rectangle1_weights[2710]), .RECT2_X(rectangle2_xs[2710]), .RECT2_Y(rectangle2_ys[2710]), .RECT2_WIDTH(rectangle2_widths[2710]), .RECT2_HEIGHT(rectangle2_heights[2710]), .RECT2_WEIGHT(rectangle2_weights[2710]), .RECT3_X(rectangle3_xs[2710]), .RECT3_Y(rectangle3_ys[2710]), .RECT3_WIDTH(rectangle3_widths[2710]), .RECT3_HEIGHT(rectangle3_heights[2710]), .RECT3_WEIGHT(rectangle3_weights[2710]), .FEAT_THRES(feature_thresholds[2710]), .FEAT_ABOVE(feature_aboves[2710]), .FEAT_BELOW(feature_belows[2710])) ac2710(.scan_win(scan_win2710), .scan_win_std_dev(scan_win_std_dev[2710]), .feature_accum(feature_accums[2710]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2711]), .RECT1_Y(rectangle1_ys[2711]), .RECT1_WIDTH(rectangle1_widths[2711]), .RECT1_HEIGHT(rectangle1_heights[2711]), .RECT1_WEIGHT(rectangle1_weights[2711]), .RECT2_X(rectangle2_xs[2711]), .RECT2_Y(rectangle2_ys[2711]), .RECT2_WIDTH(rectangle2_widths[2711]), .RECT2_HEIGHT(rectangle2_heights[2711]), .RECT2_WEIGHT(rectangle2_weights[2711]), .RECT3_X(rectangle3_xs[2711]), .RECT3_Y(rectangle3_ys[2711]), .RECT3_WIDTH(rectangle3_widths[2711]), .RECT3_HEIGHT(rectangle3_heights[2711]), .RECT3_WEIGHT(rectangle3_weights[2711]), .FEAT_THRES(feature_thresholds[2711]), .FEAT_ABOVE(feature_aboves[2711]), .FEAT_BELOW(feature_belows[2711])) ac2711(.scan_win(scan_win2711), .scan_win_std_dev(scan_win_std_dev[2711]), .feature_accum(feature_accums[2711]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2712]), .RECT1_Y(rectangle1_ys[2712]), .RECT1_WIDTH(rectangle1_widths[2712]), .RECT1_HEIGHT(rectangle1_heights[2712]), .RECT1_WEIGHT(rectangle1_weights[2712]), .RECT2_X(rectangle2_xs[2712]), .RECT2_Y(rectangle2_ys[2712]), .RECT2_WIDTH(rectangle2_widths[2712]), .RECT2_HEIGHT(rectangle2_heights[2712]), .RECT2_WEIGHT(rectangle2_weights[2712]), .RECT3_X(rectangle3_xs[2712]), .RECT3_Y(rectangle3_ys[2712]), .RECT3_WIDTH(rectangle3_widths[2712]), .RECT3_HEIGHT(rectangle3_heights[2712]), .RECT3_WEIGHT(rectangle3_weights[2712]), .FEAT_THRES(feature_thresholds[2712]), .FEAT_ABOVE(feature_aboves[2712]), .FEAT_BELOW(feature_belows[2712])) ac2712(.scan_win(scan_win2712), .scan_win_std_dev(scan_win_std_dev[2712]), .feature_accum(feature_accums[2712]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2713]), .RECT1_Y(rectangle1_ys[2713]), .RECT1_WIDTH(rectangle1_widths[2713]), .RECT1_HEIGHT(rectangle1_heights[2713]), .RECT1_WEIGHT(rectangle1_weights[2713]), .RECT2_X(rectangle2_xs[2713]), .RECT2_Y(rectangle2_ys[2713]), .RECT2_WIDTH(rectangle2_widths[2713]), .RECT2_HEIGHT(rectangle2_heights[2713]), .RECT2_WEIGHT(rectangle2_weights[2713]), .RECT3_X(rectangle3_xs[2713]), .RECT3_Y(rectangle3_ys[2713]), .RECT3_WIDTH(rectangle3_widths[2713]), .RECT3_HEIGHT(rectangle3_heights[2713]), .RECT3_WEIGHT(rectangle3_weights[2713]), .FEAT_THRES(feature_thresholds[2713]), .FEAT_ABOVE(feature_aboves[2713]), .FEAT_BELOW(feature_belows[2713])) ac2713(.scan_win(scan_win2713), .scan_win_std_dev(scan_win_std_dev[2713]), .feature_accum(feature_accums[2713]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2714]), .RECT1_Y(rectangle1_ys[2714]), .RECT1_WIDTH(rectangle1_widths[2714]), .RECT1_HEIGHT(rectangle1_heights[2714]), .RECT1_WEIGHT(rectangle1_weights[2714]), .RECT2_X(rectangle2_xs[2714]), .RECT2_Y(rectangle2_ys[2714]), .RECT2_WIDTH(rectangle2_widths[2714]), .RECT2_HEIGHT(rectangle2_heights[2714]), .RECT2_WEIGHT(rectangle2_weights[2714]), .RECT3_X(rectangle3_xs[2714]), .RECT3_Y(rectangle3_ys[2714]), .RECT3_WIDTH(rectangle3_widths[2714]), .RECT3_HEIGHT(rectangle3_heights[2714]), .RECT3_WEIGHT(rectangle3_weights[2714]), .FEAT_THRES(feature_thresholds[2714]), .FEAT_ABOVE(feature_aboves[2714]), .FEAT_BELOW(feature_belows[2714])) ac2714(.scan_win(scan_win2714), .scan_win_std_dev(scan_win_std_dev[2714]), .feature_accum(feature_accums[2714]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2715]), .RECT1_Y(rectangle1_ys[2715]), .RECT1_WIDTH(rectangle1_widths[2715]), .RECT1_HEIGHT(rectangle1_heights[2715]), .RECT1_WEIGHT(rectangle1_weights[2715]), .RECT2_X(rectangle2_xs[2715]), .RECT2_Y(rectangle2_ys[2715]), .RECT2_WIDTH(rectangle2_widths[2715]), .RECT2_HEIGHT(rectangle2_heights[2715]), .RECT2_WEIGHT(rectangle2_weights[2715]), .RECT3_X(rectangle3_xs[2715]), .RECT3_Y(rectangle3_ys[2715]), .RECT3_WIDTH(rectangle3_widths[2715]), .RECT3_HEIGHT(rectangle3_heights[2715]), .RECT3_WEIGHT(rectangle3_weights[2715]), .FEAT_THRES(feature_thresholds[2715]), .FEAT_ABOVE(feature_aboves[2715]), .FEAT_BELOW(feature_belows[2715])) ac2715(.scan_win(scan_win2715), .scan_win_std_dev(scan_win_std_dev[2715]), .feature_accum(feature_accums[2715]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2716]), .RECT1_Y(rectangle1_ys[2716]), .RECT1_WIDTH(rectangle1_widths[2716]), .RECT1_HEIGHT(rectangle1_heights[2716]), .RECT1_WEIGHT(rectangle1_weights[2716]), .RECT2_X(rectangle2_xs[2716]), .RECT2_Y(rectangle2_ys[2716]), .RECT2_WIDTH(rectangle2_widths[2716]), .RECT2_HEIGHT(rectangle2_heights[2716]), .RECT2_WEIGHT(rectangle2_weights[2716]), .RECT3_X(rectangle3_xs[2716]), .RECT3_Y(rectangle3_ys[2716]), .RECT3_WIDTH(rectangle3_widths[2716]), .RECT3_HEIGHT(rectangle3_heights[2716]), .RECT3_WEIGHT(rectangle3_weights[2716]), .FEAT_THRES(feature_thresholds[2716]), .FEAT_ABOVE(feature_aboves[2716]), .FEAT_BELOW(feature_belows[2716])) ac2716(.scan_win(scan_win2716), .scan_win_std_dev(scan_win_std_dev[2716]), .feature_accum(feature_accums[2716]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2717]), .RECT1_Y(rectangle1_ys[2717]), .RECT1_WIDTH(rectangle1_widths[2717]), .RECT1_HEIGHT(rectangle1_heights[2717]), .RECT1_WEIGHT(rectangle1_weights[2717]), .RECT2_X(rectangle2_xs[2717]), .RECT2_Y(rectangle2_ys[2717]), .RECT2_WIDTH(rectangle2_widths[2717]), .RECT2_HEIGHT(rectangle2_heights[2717]), .RECT2_WEIGHT(rectangle2_weights[2717]), .RECT3_X(rectangle3_xs[2717]), .RECT3_Y(rectangle3_ys[2717]), .RECT3_WIDTH(rectangle3_widths[2717]), .RECT3_HEIGHT(rectangle3_heights[2717]), .RECT3_WEIGHT(rectangle3_weights[2717]), .FEAT_THRES(feature_thresholds[2717]), .FEAT_ABOVE(feature_aboves[2717]), .FEAT_BELOW(feature_belows[2717])) ac2717(.scan_win(scan_win2717), .scan_win_std_dev(scan_win_std_dev[2717]), .feature_accum(feature_accums[2717]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2718]), .RECT1_Y(rectangle1_ys[2718]), .RECT1_WIDTH(rectangle1_widths[2718]), .RECT1_HEIGHT(rectangle1_heights[2718]), .RECT1_WEIGHT(rectangle1_weights[2718]), .RECT2_X(rectangle2_xs[2718]), .RECT2_Y(rectangle2_ys[2718]), .RECT2_WIDTH(rectangle2_widths[2718]), .RECT2_HEIGHT(rectangle2_heights[2718]), .RECT2_WEIGHT(rectangle2_weights[2718]), .RECT3_X(rectangle3_xs[2718]), .RECT3_Y(rectangle3_ys[2718]), .RECT3_WIDTH(rectangle3_widths[2718]), .RECT3_HEIGHT(rectangle3_heights[2718]), .RECT3_WEIGHT(rectangle3_weights[2718]), .FEAT_THRES(feature_thresholds[2718]), .FEAT_ABOVE(feature_aboves[2718]), .FEAT_BELOW(feature_belows[2718])) ac2718(.scan_win(scan_win2718), .scan_win_std_dev(scan_win_std_dev[2718]), .feature_accum(feature_accums[2718]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2719]), .RECT1_Y(rectangle1_ys[2719]), .RECT1_WIDTH(rectangle1_widths[2719]), .RECT1_HEIGHT(rectangle1_heights[2719]), .RECT1_WEIGHT(rectangle1_weights[2719]), .RECT2_X(rectangle2_xs[2719]), .RECT2_Y(rectangle2_ys[2719]), .RECT2_WIDTH(rectangle2_widths[2719]), .RECT2_HEIGHT(rectangle2_heights[2719]), .RECT2_WEIGHT(rectangle2_weights[2719]), .RECT3_X(rectangle3_xs[2719]), .RECT3_Y(rectangle3_ys[2719]), .RECT3_WIDTH(rectangle3_widths[2719]), .RECT3_HEIGHT(rectangle3_heights[2719]), .RECT3_WEIGHT(rectangle3_weights[2719]), .FEAT_THRES(feature_thresholds[2719]), .FEAT_ABOVE(feature_aboves[2719]), .FEAT_BELOW(feature_belows[2719])) ac2719(.scan_win(scan_win2719), .scan_win_std_dev(scan_win_std_dev[2719]), .feature_accum(feature_accums[2719]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2720]), .RECT1_Y(rectangle1_ys[2720]), .RECT1_WIDTH(rectangle1_widths[2720]), .RECT1_HEIGHT(rectangle1_heights[2720]), .RECT1_WEIGHT(rectangle1_weights[2720]), .RECT2_X(rectangle2_xs[2720]), .RECT2_Y(rectangle2_ys[2720]), .RECT2_WIDTH(rectangle2_widths[2720]), .RECT2_HEIGHT(rectangle2_heights[2720]), .RECT2_WEIGHT(rectangle2_weights[2720]), .RECT3_X(rectangle3_xs[2720]), .RECT3_Y(rectangle3_ys[2720]), .RECT3_WIDTH(rectangle3_widths[2720]), .RECT3_HEIGHT(rectangle3_heights[2720]), .RECT3_WEIGHT(rectangle3_weights[2720]), .FEAT_THRES(feature_thresholds[2720]), .FEAT_ABOVE(feature_aboves[2720]), .FEAT_BELOW(feature_belows[2720])) ac2720(.scan_win(scan_win2720), .scan_win_std_dev(scan_win_std_dev[2720]), .feature_accum(feature_accums[2720]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2721]), .RECT1_Y(rectangle1_ys[2721]), .RECT1_WIDTH(rectangle1_widths[2721]), .RECT1_HEIGHT(rectangle1_heights[2721]), .RECT1_WEIGHT(rectangle1_weights[2721]), .RECT2_X(rectangle2_xs[2721]), .RECT2_Y(rectangle2_ys[2721]), .RECT2_WIDTH(rectangle2_widths[2721]), .RECT2_HEIGHT(rectangle2_heights[2721]), .RECT2_WEIGHT(rectangle2_weights[2721]), .RECT3_X(rectangle3_xs[2721]), .RECT3_Y(rectangle3_ys[2721]), .RECT3_WIDTH(rectangle3_widths[2721]), .RECT3_HEIGHT(rectangle3_heights[2721]), .RECT3_WEIGHT(rectangle3_weights[2721]), .FEAT_THRES(feature_thresholds[2721]), .FEAT_ABOVE(feature_aboves[2721]), .FEAT_BELOW(feature_belows[2721])) ac2721(.scan_win(scan_win2721), .scan_win_std_dev(scan_win_std_dev[2721]), .feature_accum(feature_accums[2721]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2722]), .RECT1_Y(rectangle1_ys[2722]), .RECT1_WIDTH(rectangle1_widths[2722]), .RECT1_HEIGHT(rectangle1_heights[2722]), .RECT1_WEIGHT(rectangle1_weights[2722]), .RECT2_X(rectangle2_xs[2722]), .RECT2_Y(rectangle2_ys[2722]), .RECT2_WIDTH(rectangle2_widths[2722]), .RECT2_HEIGHT(rectangle2_heights[2722]), .RECT2_WEIGHT(rectangle2_weights[2722]), .RECT3_X(rectangle3_xs[2722]), .RECT3_Y(rectangle3_ys[2722]), .RECT3_WIDTH(rectangle3_widths[2722]), .RECT3_HEIGHT(rectangle3_heights[2722]), .RECT3_WEIGHT(rectangle3_weights[2722]), .FEAT_THRES(feature_thresholds[2722]), .FEAT_ABOVE(feature_aboves[2722]), .FEAT_BELOW(feature_belows[2722])) ac2722(.scan_win(scan_win2722), .scan_win_std_dev(scan_win_std_dev[2722]), .feature_accum(feature_accums[2722]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2723]), .RECT1_Y(rectangle1_ys[2723]), .RECT1_WIDTH(rectangle1_widths[2723]), .RECT1_HEIGHT(rectangle1_heights[2723]), .RECT1_WEIGHT(rectangle1_weights[2723]), .RECT2_X(rectangle2_xs[2723]), .RECT2_Y(rectangle2_ys[2723]), .RECT2_WIDTH(rectangle2_widths[2723]), .RECT2_HEIGHT(rectangle2_heights[2723]), .RECT2_WEIGHT(rectangle2_weights[2723]), .RECT3_X(rectangle3_xs[2723]), .RECT3_Y(rectangle3_ys[2723]), .RECT3_WIDTH(rectangle3_widths[2723]), .RECT3_HEIGHT(rectangle3_heights[2723]), .RECT3_WEIGHT(rectangle3_weights[2723]), .FEAT_THRES(feature_thresholds[2723]), .FEAT_ABOVE(feature_aboves[2723]), .FEAT_BELOW(feature_belows[2723])) ac2723(.scan_win(scan_win2723), .scan_win_std_dev(scan_win_std_dev[2723]), .feature_accum(feature_accums[2723]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2724]), .RECT1_Y(rectangle1_ys[2724]), .RECT1_WIDTH(rectangle1_widths[2724]), .RECT1_HEIGHT(rectangle1_heights[2724]), .RECT1_WEIGHT(rectangle1_weights[2724]), .RECT2_X(rectangle2_xs[2724]), .RECT2_Y(rectangle2_ys[2724]), .RECT2_WIDTH(rectangle2_widths[2724]), .RECT2_HEIGHT(rectangle2_heights[2724]), .RECT2_WEIGHT(rectangle2_weights[2724]), .RECT3_X(rectangle3_xs[2724]), .RECT3_Y(rectangle3_ys[2724]), .RECT3_WIDTH(rectangle3_widths[2724]), .RECT3_HEIGHT(rectangle3_heights[2724]), .RECT3_WEIGHT(rectangle3_weights[2724]), .FEAT_THRES(feature_thresholds[2724]), .FEAT_ABOVE(feature_aboves[2724]), .FEAT_BELOW(feature_belows[2724])) ac2724(.scan_win(scan_win2724), .scan_win_std_dev(scan_win_std_dev[2724]), .feature_accum(feature_accums[2724]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2725]), .RECT1_Y(rectangle1_ys[2725]), .RECT1_WIDTH(rectangle1_widths[2725]), .RECT1_HEIGHT(rectangle1_heights[2725]), .RECT1_WEIGHT(rectangle1_weights[2725]), .RECT2_X(rectangle2_xs[2725]), .RECT2_Y(rectangle2_ys[2725]), .RECT2_WIDTH(rectangle2_widths[2725]), .RECT2_HEIGHT(rectangle2_heights[2725]), .RECT2_WEIGHT(rectangle2_weights[2725]), .RECT3_X(rectangle3_xs[2725]), .RECT3_Y(rectangle3_ys[2725]), .RECT3_WIDTH(rectangle3_widths[2725]), .RECT3_HEIGHT(rectangle3_heights[2725]), .RECT3_WEIGHT(rectangle3_weights[2725]), .FEAT_THRES(feature_thresholds[2725]), .FEAT_ABOVE(feature_aboves[2725]), .FEAT_BELOW(feature_belows[2725])) ac2725(.scan_win(scan_win2725), .scan_win_std_dev(scan_win_std_dev[2725]), .feature_accum(feature_accums[2725]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2726]), .RECT1_Y(rectangle1_ys[2726]), .RECT1_WIDTH(rectangle1_widths[2726]), .RECT1_HEIGHT(rectangle1_heights[2726]), .RECT1_WEIGHT(rectangle1_weights[2726]), .RECT2_X(rectangle2_xs[2726]), .RECT2_Y(rectangle2_ys[2726]), .RECT2_WIDTH(rectangle2_widths[2726]), .RECT2_HEIGHT(rectangle2_heights[2726]), .RECT2_WEIGHT(rectangle2_weights[2726]), .RECT3_X(rectangle3_xs[2726]), .RECT3_Y(rectangle3_ys[2726]), .RECT3_WIDTH(rectangle3_widths[2726]), .RECT3_HEIGHT(rectangle3_heights[2726]), .RECT3_WEIGHT(rectangle3_weights[2726]), .FEAT_THRES(feature_thresholds[2726]), .FEAT_ABOVE(feature_aboves[2726]), .FEAT_BELOW(feature_belows[2726])) ac2726(.scan_win(scan_win2726), .scan_win_std_dev(scan_win_std_dev[2726]), .feature_accum(feature_accums[2726]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2727]), .RECT1_Y(rectangle1_ys[2727]), .RECT1_WIDTH(rectangle1_widths[2727]), .RECT1_HEIGHT(rectangle1_heights[2727]), .RECT1_WEIGHT(rectangle1_weights[2727]), .RECT2_X(rectangle2_xs[2727]), .RECT2_Y(rectangle2_ys[2727]), .RECT2_WIDTH(rectangle2_widths[2727]), .RECT2_HEIGHT(rectangle2_heights[2727]), .RECT2_WEIGHT(rectangle2_weights[2727]), .RECT3_X(rectangle3_xs[2727]), .RECT3_Y(rectangle3_ys[2727]), .RECT3_WIDTH(rectangle3_widths[2727]), .RECT3_HEIGHT(rectangle3_heights[2727]), .RECT3_WEIGHT(rectangle3_weights[2727]), .FEAT_THRES(feature_thresholds[2727]), .FEAT_ABOVE(feature_aboves[2727]), .FEAT_BELOW(feature_belows[2727])) ac2727(.scan_win(scan_win2727), .scan_win_std_dev(scan_win_std_dev[2727]), .feature_accum(feature_accums[2727]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2728]), .RECT1_Y(rectangle1_ys[2728]), .RECT1_WIDTH(rectangle1_widths[2728]), .RECT1_HEIGHT(rectangle1_heights[2728]), .RECT1_WEIGHT(rectangle1_weights[2728]), .RECT2_X(rectangle2_xs[2728]), .RECT2_Y(rectangle2_ys[2728]), .RECT2_WIDTH(rectangle2_widths[2728]), .RECT2_HEIGHT(rectangle2_heights[2728]), .RECT2_WEIGHT(rectangle2_weights[2728]), .RECT3_X(rectangle3_xs[2728]), .RECT3_Y(rectangle3_ys[2728]), .RECT3_WIDTH(rectangle3_widths[2728]), .RECT3_HEIGHT(rectangle3_heights[2728]), .RECT3_WEIGHT(rectangle3_weights[2728]), .FEAT_THRES(feature_thresholds[2728]), .FEAT_ABOVE(feature_aboves[2728]), .FEAT_BELOW(feature_belows[2728])) ac2728(.scan_win(scan_win2728), .scan_win_std_dev(scan_win_std_dev[2728]), .feature_accum(feature_accums[2728]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2729]), .RECT1_Y(rectangle1_ys[2729]), .RECT1_WIDTH(rectangle1_widths[2729]), .RECT1_HEIGHT(rectangle1_heights[2729]), .RECT1_WEIGHT(rectangle1_weights[2729]), .RECT2_X(rectangle2_xs[2729]), .RECT2_Y(rectangle2_ys[2729]), .RECT2_WIDTH(rectangle2_widths[2729]), .RECT2_HEIGHT(rectangle2_heights[2729]), .RECT2_WEIGHT(rectangle2_weights[2729]), .RECT3_X(rectangle3_xs[2729]), .RECT3_Y(rectangle3_ys[2729]), .RECT3_WIDTH(rectangle3_widths[2729]), .RECT3_HEIGHT(rectangle3_heights[2729]), .RECT3_WEIGHT(rectangle3_weights[2729]), .FEAT_THRES(feature_thresholds[2729]), .FEAT_ABOVE(feature_aboves[2729]), .FEAT_BELOW(feature_belows[2729])) ac2729(.scan_win(scan_win2729), .scan_win_std_dev(scan_win_std_dev[2729]), .feature_accum(feature_accums[2729]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2730]), .RECT1_Y(rectangle1_ys[2730]), .RECT1_WIDTH(rectangle1_widths[2730]), .RECT1_HEIGHT(rectangle1_heights[2730]), .RECT1_WEIGHT(rectangle1_weights[2730]), .RECT2_X(rectangle2_xs[2730]), .RECT2_Y(rectangle2_ys[2730]), .RECT2_WIDTH(rectangle2_widths[2730]), .RECT2_HEIGHT(rectangle2_heights[2730]), .RECT2_WEIGHT(rectangle2_weights[2730]), .RECT3_X(rectangle3_xs[2730]), .RECT3_Y(rectangle3_ys[2730]), .RECT3_WIDTH(rectangle3_widths[2730]), .RECT3_HEIGHT(rectangle3_heights[2730]), .RECT3_WEIGHT(rectangle3_weights[2730]), .FEAT_THRES(feature_thresholds[2730]), .FEAT_ABOVE(feature_aboves[2730]), .FEAT_BELOW(feature_belows[2730])) ac2730(.scan_win(scan_win2730), .scan_win_std_dev(scan_win_std_dev[2730]), .feature_accum(feature_accums[2730]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2731]), .RECT1_Y(rectangle1_ys[2731]), .RECT1_WIDTH(rectangle1_widths[2731]), .RECT1_HEIGHT(rectangle1_heights[2731]), .RECT1_WEIGHT(rectangle1_weights[2731]), .RECT2_X(rectangle2_xs[2731]), .RECT2_Y(rectangle2_ys[2731]), .RECT2_WIDTH(rectangle2_widths[2731]), .RECT2_HEIGHT(rectangle2_heights[2731]), .RECT2_WEIGHT(rectangle2_weights[2731]), .RECT3_X(rectangle3_xs[2731]), .RECT3_Y(rectangle3_ys[2731]), .RECT3_WIDTH(rectangle3_widths[2731]), .RECT3_HEIGHT(rectangle3_heights[2731]), .RECT3_WEIGHT(rectangle3_weights[2731]), .FEAT_THRES(feature_thresholds[2731]), .FEAT_ABOVE(feature_aboves[2731]), .FEAT_BELOW(feature_belows[2731])) ac2731(.scan_win(scan_win2731), .scan_win_std_dev(scan_win_std_dev[2731]), .feature_accum(feature_accums[2731]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2732]), .RECT1_Y(rectangle1_ys[2732]), .RECT1_WIDTH(rectangle1_widths[2732]), .RECT1_HEIGHT(rectangle1_heights[2732]), .RECT1_WEIGHT(rectangle1_weights[2732]), .RECT2_X(rectangle2_xs[2732]), .RECT2_Y(rectangle2_ys[2732]), .RECT2_WIDTH(rectangle2_widths[2732]), .RECT2_HEIGHT(rectangle2_heights[2732]), .RECT2_WEIGHT(rectangle2_weights[2732]), .RECT3_X(rectangle3_xs[2732]), .RECT3_Y(rectangle3_ys[2732]), .RECT3_WIDTH(rectangle3_widths[2732]), .RECT3_HEIGHT(rectangle3_heights[2732]), .RECT3_WEIGHT(rectangle3_weights[2732]), .FEAT_THRES(feature_thresholds[2732]), .FEAT_ABOVE(feature_aboves[2732]), .FEAT_BELOW(feature_belows[2732])) ac2732(.scan_win(scan_win2732), .scan_win_std_dev(scan_win_std_dev[2732]), .feature_accum(feature_accums[2732]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2733]), .RECT1_Y(rectangle1_ys[2733]), .RECT1_WIDTH(rectangle1_widths[2733]), .RECT1_HEIGHT(rectangle1_heights[2733]), .RECT1_WEIGHT(rectangle1_weights[2733]), .RECT2_X(rectangle2_xs[2733]), .RECT2_Y(rectangle2_ys[2733]), .RECT2_WIDTH(rectangle2_widths[2733]), .RECT2_HEIGHT(rectangle2_heights[2733]), .RECT2_WEIGHT(rectangle2_weights[2733]), .RECT3_X(rectangle3_xs[2733]), .RECT3_Y(rectangle3_ys[2733]), .RECT3_WIDTH(rectangle3_widths[2733]), .RECT3_HEIGHT(rectangle3_heights[2733]), .RECT3_WEIGHT(rectangle3_weights[2733]), .FEAT_THRES(feature_thresholds[2733]), .FEAT_ABOVE(feature_aboves[2733]), .FEAT_BELOW(feature_belows[2733])) ac2733(.scan_win(scan_win2733), .scan_win_std_dev(scan_win_std_dev[2733]), .feature_accum(feature_accums[2733]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2734]), .RECT1_Y(rectangle1_ys[2734]), .RECT1_WIDTH(rectangle1_widths[2734]), .RECT1_HEIGHT(rectangle1_heights[2734]), .RECT1_WEIGHT(rectangle1_weights[2734]), .RECT2_X(rectangle2_xs[2734]), .RECT2_Y(rectangle2_ys[2734]), .RECT2_WIDTH(rectangle2_widths[2734]), .RECT2_HEIGHT(rectangle2_heights[2734]), .RECT2_WEIGHT(rectangle2_weights[2734]), .RECT3_X(rectangle3_xs[2734]), .RECT3_Y(rectangle3_ys[2734]), .RECT3_WIDTH(rectangle3_widths[2734]), .RECT3_HEIGHT(rectangle3_heights[2734]), .RECT3_WEIGHT(rectangle3_weights[2734]), .FEAT_THRES(feature_thresholds[2734]), .FEAT_ABOVE(feature_aboves[2734]), .FEAT_BELOW(feature_belows[2734])) ac2734(.scan_win(scan_win2734), .scan_win_std_dev(scan_win_std_dev[2734]), .feature_accum(feature_accums[2734]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2735]), .RECT1_Y(rectangle1_ys[2735]), .RECT1_WIDTH(rectangle1_widths[2735]), .RECT1_HEIGHT(rectangle1_heights[2735]), .RECT1_WEIGHT(rectangle1_weights[2735]), .RECT2_X(rectangle2_xs[2735]), .RECT2_Y(rectangle2_ys[2735]), .RECT2_WIDTH(rectangle2_widths[2735]), .RECT2_HEIGHT(rectangle2_heights[2735]), .RECT2_WEIGHT(rectangle2_weights[2735]), .RECT3_X(rectangle3_xs[2735]), .RECT3_Y(rectangle3_ys[2735]), .RECT3_WIDTH(rectangle3_widths[2735]), .RECT3_HEIGHT(rectangle3_heights[2735]), .RECT3_WEIGHT(rectangle3_weights[2735]), .FEAT_THRES(feature_thresholds[2735]), .FEAT_ABOVE(feature_aboves[2735]), .FEAT_BELOW(feature_belows[2735])) ac2735(.scan_win(scan_win2735), .scan_win_std_dev(scan_win_std_dev[2735]), .feature_accum(feature_accums[2735]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2736]), .RECT1_Y(rectangle1_ys[2736]), .RECT1_WIDTH(rectangle1_widths[2736]), .RECT1_HEIGHT(rectangle1_heights[2736]), .RECT1_WEIGHT(rectangle1_weights[2736]), .RECT2_X(rectangle2_xs[2736]), .RECT2_Y(rectangle2_ys[2736]), .RECT2_WIDTH(rectangle2_widths[2736]), .RECT2_HEIGHT(rectangle2_heights[2736]), .RECT2_WEIGHT(rectangle2_weights[2736]), .RECT3_X(rectangle3_xs[2736]), .RECT3_Y(rectangle3_ys[2736]), .RECT3_WIDTH(rectangle3_widths[2736]), .RECT3_HEIGHT(rectangle3_heights[2736]), .RECT3_WEIGHT(rectangle3_weights[2736]), .FEAT_THRES(feature_thresholds[2736]), .FEAT_ABOVE(feature_aboves[2736]), .FEAT_BELOW(feature_belows[2736])) ac2736(.scan_win(scan_win2736), .scan_win_std_dev(scan_win_std_dev[2736]), .feature_accum(feature_accums[2736]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2737]), .RECT1_Y(rectangle1_ys[2737]), .RECT1_WIDTH(rectangle1_widths[2737]), .RECT1_HEIGHT(rectangle1_heights[2737]), .RECT1_WEIGHT(rectangle1_weights[2737]), .RECT2_X(rectangle2_xs[2737]), .RECT2_Y(rectangle2_ys[2737]), .RECT2_WIDTH(rectangle2_widths[2737]), .RECT2_HEIGHT(rectangle2_heights[2737]), .RECT2_WEIGHT(rectangle2_weights[2737]), .RECT3_X(rectangle3_xs[2737]), .RECT3_Y(rectangle3_ys[2737]), .RECT3_WIDTH(rectangle3_widths[2737]), .RECT3_HEIGHT(rectangle3_heights[2737]), .RECT3_WEIGHT(rectangle3_weights[2737]), .FEAT_THRES(feature_thresholds[2737]), .FEAT_ABOVE(feature_aboves[2737]), .FEAT_BELOW(feature_belows[2737])) ac2737(.scan_win(scan_win2737), .scan_win_std_dev(scan_win_std_dev[2737]), .feature_accum(feature_accums[2737]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2738]), .RECT1_Y(rectangle1_ys[2738]), .RECT1_WIDTH(rectangle1_widths[2738]), .RECT1_HEIGHT(rectangle1_heights[2738]), .RECT1_WEIGHT(rectangle1_weights[2738]), .RECT2_X(rectangle2_xs[2738]), .RECT2_Y(rectangle2_ys[2738]), .RECT2_WIDTH(rectangle2_widths[2738]), .RECT2_HEIGHT(rectangle2_heights[2738]), .RECT2_WEIGHT(rectangle2_weights[2738]), .RECT3_X(rectangle3_xs[2738]), .RECT3_Y(rectangle3_ys[2738]), .RECT3_WIDTH(rectangle3_widths[2738]), .RECT3_HEIGHT(rectangle3_heights[2738]), .RECT3_WEIGHT(rectangle3_weights[2738]), .FEAT_THRES(feature_thresholds[2738]), .FEAT_ABOVE(feature_aboves[2738]), .FEAT_BELOW(feature_belows[2738])) ac2738(.scan_win(scan_win2738), .scan_win_std_dev(scan_win_std_dev[2738]), .feature_accum(feature_accums[2738]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2739]), .RECT1_Y(rectangle1_ys[2739]), .RECT1_WIDTH(rectangle1_widths[2739]), .RECT1_HEIGHT(rectangle1_heights[2739]), .RECT1_WEIGHT(rectangle1_weights[2739]), .RECT2_X(rectangle2_xs[2739]), .RECT2_Y(rectangle2_ys[2739]), .RECT2_WIDTH(rectangle2_widths[2739]), .RECT2_HEIGHT(rectangle2_heights[2739]), .RECT2_WEIGHT(rectangle2_weights[2739]), .RECT3_X(rectangle3_xs[2739]), .RECT3_Y(rectangle3_ys[2739]), .RECT3_WIDTH(rectangle3_widths[2739]), .RECT3_HEIGHT(rectangle3_heights[2739]), .RECT3_WEIGHT(rectangle3_weights[2739]), .FEAT_THRES(feature_thresholds[2739]), .FEAT_ABOVE(feature_aboves[2739]), .FEAT_BELOW(feature_belows[2739])) ac2739(.scan_win(scan_win2739), .scan_win_std_dev(scan_win_std_dev[2739]), .feature_accum(feature_accums[2739]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2740]), .RECT1_Y(rectangle1_ys[2740]), .RECT1_WIDTH(rectangle1_widths[2740]), .RECT1_HEIGHT(rectangle1_heights[2740]), .RECT1_WEIGHT(rectangle1_weights[2740]), .RECT2_X(rectangle2_xs[2740]), .RECT2_Y(rectangle2_ys[2740]), .RECT2_WIDTH(rectangle2_widths[2740]), .RECT2_HEIGHT(rectangle2_heights[2740]), .RECT2_WEIGHT(rectangle2_weights[2740]), .RECT3_X(rectangle3_xs[2740]), .RECT3_Y(rectangle3_ys[2740]), .RECT3_WIDTH(rectangle3_widths[2740]), .RECT3_HEIGHT(rectangle3_heights[2740]), .RECT3_WEIGHT(rectangle3_weights[2740]), .FEAT_THRES(feature_thresholds[2740]), .FEAT_ABOVE(feature_aboves[2740]), .FEAT_BELOW(feature_belows[2740])) ac2740(.scan_win(scan_win2740), .scan_win_std_dev(scan_win_std_dev[2740]), .feature_accum(feature_accums[2740]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2741]), .RECT1_Y(rectangle1_ys[2741]), .RECT1_WIDTH(rectangle1_widths[2741]), .RECT1_HEIGHT(rectangle1_heights[2741]), .RECT1_WEIGHT(rectangle1_weights[2741]), .RECT2_X(rectangle2_xs[2741]), .RECT2_Y(rectangle2_ys[2741]), .RECT2_WIDTH(rectangle2_widths[2741]), .RECT2_HEIGHT(rectangle2_heights[2741]), .RECT2_WEIGHT(rectangle2_weights[2741]), .RECT3_X(rectangle3_xs[2741]), .RECT3_Y(rectangle3_ys[2741]), .RECT3_WIDTH(rectangle3_widths[2741]), .RECT3_HEIGHT(rectangle3_heights[2741]), .RECT3_WEIGHT(rectangle3_weights[2741]), .FEAT_THRES(feature_thresholds[2741]), .FEAT_ABOVE(feature_aboves[2741]), .FEAT_BELOW(feature_belows[2741])) ac2741(.scan_win(scan_win2741), .scan_win_std_dev(scan_win_std_dev[2741]), .feature_accum(feature_accums[2741]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2742]), .RECT1_Y(rectangle1_ys[2742]), .RECT1_WIDTH(rectangle1_widths[2742]), .RECT1_HEIGHT(rectangle1_heights[2742]), .RECT1_WEIGHT(rectangle1_weights[2742]), .RECT2_X(rectangle2_xs[2742]), .RECT2_Y(rectangle2_ys[2742]), .RECT2_WIDTH(rectangle2_widths[2742]), .RECT2_HEIGHT(rectangle2_heights[2742]), .RECT2_WEIGHT(rectangle2_weights[2742]), .RECT3_X(rectangle3_xs[2742]), .RECT3_Y(rectangle3_ys[2742]), .RECT3_WIDTH(rectangle3_widths[2742]), .RECT3_HEIGHT(rectangle3_heights[2742]), .RECT3_WEIGHT(rectangle3_weights[2742]), .FEAT_THRES(feature_thresholds[2742]), .FEAT_ABOVE(feature_aboves[2742]), .FEAT_BELOW(feature_belows[2742])) ac2742(.scan_win(scan_win2742), .scan_win_std_dev(scan_win_std_dev[2742]), .feature_accum(feature_accums[2742]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2743]), .RECT1_Y(rectangle1_ys[2743]), .RECT1_WIDTH(rectangle1_widths[2743]), .RECT1_HEIGHT(rectangle1_heights[2743]), .RECT1_WEIGHT(rectangle1_weights[2743]), .RECT2_X(rectangle2_xs[2743]), .RECT2_Y(rectangle2_ys[2743]), .RECT2_WIDTH(rectangle2_widths[2743]), .RECT2_HEIGHT(rectangle2_heights[2743]), .RECT2_WEIGHT(rectangle2_weights[2743]), .RECT3_X(rectangle3_xs[2743]), .RECT3_Y(rectangle3_ys[2743]), .RECT3_WIDTH(rectangle3_widths[2743]), .RECT3_HEIGHT(rectangle3_heights[2743]), .RECT3_WEIGHT(rectangle3_weights[2743]), .FEAT_THRES(feature_thresholds[2743]), .FEAT_ABOVE(feature_aboves[2743]), .FEAT_BELOW(feature_belows[2743])) ac2743(.scan_win(scan_win2743), .scan_win_std_dev(scan_win_std_dev[2743]), .feature_accum(feature_accums[2743]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2744]), .RECT1_Y(rectangle1_ys[2744]), .RECT1_WIDTH(rectangle1_widths[2744]), .RECT1_HEIGHT(rectangle1_heights[2744]), .RECT1_WEIGHT(rectangle1_weights[2744]), .RECT2_X(rectangle2_xs[2744]), .RECT2_Y(rectangle2_ys[2744]), .RECT2_WIDTH(rectangle2_widths[2744]), .RECT2_HEIGHT(rectangle2_heights[2744]), .RECT2_WEIGHT(rectangle2_weights[2744]), .RECT3_X(rectangle3_xs[2744]), .RECT3_Y(rectangle3_ys[2744]), .RECT3_WIDTH(rectangle3_widths[2744]), .RECT3_HEIGHT(rectangle3_heights[2744]), .RECT3_WEIGHT(rectangle3_weights[2744]), .FEAT_THRES(feature_thresholds[2744]), .FEAT_ABOVE(feature_aboves[2744]), .FEAT_BELOW(feature_belows[2744])) ac2744(.scan_win(scan_win2744), .scan_win_std_dev(scan_win_std_dev[2744]), .feature_accum(feature_accums[2744]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2745]), .RECT1_Y(rectangle1_ys[2745]), .RECT1_WIDTH(rectangle1_widths[2745]), .RECT1_HEIGHT(rectangle1_heights[2745]), .RECT1_WEIGHT(rectangle1_weights[2745]), .RECT2_X(rectangle2_xs[2745]), .RECT2_Y(rectangle2_ys[2745]), .RECT2_WIDTH(rectangle2_widths[2745]), .RECT2_HEIGHT(rectangle2_heights[2745]), .RECT2_WEIGHT(rectangle2_weights[2745]), .RECT3_X(rectangle3_xs[2745]), .RECT3_Y(rectangle3_ys[2745]), .RECT3_WIDTH(rectangle3_widths[2745]), .RECT3_HEIGHT(rectangle3_heights[2745]), .RECT3_WEIGHT(rectangle3_weights[2745]), .FEAT_THRES(feature_thresholds[2745]), .FEAT_ABOVE(feature_aboves[2745]), .FEAT_BELOW(feature_belows[2745])) ac2745(.scan_win(scan_win2745), .scan_win_std_dev(scan_win_std_dev[2745]), .feature_accum(feature_accums[2745]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2746]), .RECT1_Y(rectangle1_ys[2746]), .RECT1_WIDTH(rectangle1_widths[2746]), .RECT1_HEIGHT(rectangle1_heights[2746]), .RECT1_WEIGHT(rectangle1_weights[2746]), .RECT2_X(rectangle2_xs[2746]), .RECT2_Y(rectangle2_ys[2746]), .RECT2_WIDTH(rectangle2_widths[2746]), .RECT2_HEIGHT(rectangle2_heights[2746]), .RECT2_WEIGHT(rectangle2_weights[2746]), .RECT3_X(rectangle3_xs[2746]), .RECT3_Y(rectangle3_ys[2746]), .RECT3_WIDTH(rectangle3_widths[2746]), .RECT3_HEIGHT(rectangle3_heights[2746]), .RECT3_WEIGHT(rectangle3_weights[2746]), .FEAT_THRES(feature_thresholds[2746]), .FEAT_ABOVE(feature_aboves[2746]), .FEAT_BELOW(feature_belows[2746])) ac2746(.scan_win(scan_win2746), .scan_win_std_dev(scan_win_std_dev[2746]), .feature_accum(feature_accums[2746]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2747]), .RECT1_Y(rectangle1_ys[2747]), .RECT1_WIDTH(rectangle1_widths[2747]), .RECT1_HEIGHT(rectangle1_heights[2747]), .RECT1_WEIGHT(rectangle1_weights[2747]), .RECT2_X(rectangle2_xs[2747]), .RECT2_Y(rectangle2_ys[2747]), .RECT2_WIDTH(rectangle2_widths[2747]), .RECT2_HEIGHT(rectangle2_heights[2747]), .RECT2_WEIGHT(rectangle2_weights[2747]), .RECT3_X(rectangle3_xs[2747]), .RECT3_Y(rectangle3_ys[2747]), .RECT3_WIDTH(rectangle3_widths[2747]), .RECT3_HEIGHT(rectangle3_heights[2747]), .RECT3_WEIGHT(rectangle3_weights[2747]), .FEAT_THRES(feature_thresholds[2747]), .FEAT_ABOVE(feature_aboves[2747]), .FEAT_BELOW(feature_belows[2747])) ac2747(.scan_win(scan_win2747), .scan_win_std_dev(scan_win_std_dev[2747]), .feature_accum(feature_accums[2747]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2748]), .RECT1_Y(rectangle1_ys[2748]), .RECT1_WIDTH(rectangle1_widths[2748]), .RECT1_HEIGHT(rectangle1_heights[2748]), .RECT1_WEIGHT(rectangle1_weights[2748]), .RECT2_X(rectangle2_xs[2748]), .RECT2_Y(rectangle2_ys[2748]), .RECT2_WIDTH(rectangle2_widths[2748]), .RECT2_HEIGHT(rectangle2_heights[2748]), .RECT2_WEIGHT(rectangle2_weights[2748]), .RECT3_X(rectangle3_xs[2748]), .RECT3_Y(rectangle3_ys[2748]), .RECT3_WIDTH(rectangle3_widths[2748]), .RECT3_HEIGHT(rectangle3_heights[2748]), .RECT3_WEIGHT(rectangle3_weights[2748]), .FEAT_THRES(feature_thresholds[2748]), .FEAT_ABOVE(feature_aboves[2748]), .FEAT_BELOW(feature_belows[2748])) ac2748(.scan_win(scan_win2748), .scan_win_std_dev(scan_win_std_dev[2748]), .feature_accum(feature_accums[2748]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2749]), .RECT1_Y(rectangle1_ys[2749]), .RECT1_WIDTH(rectangle1_widths[2749]), .RECT1_HEIGHT(rectangle1_heights[2749]), .RECT1_WEIGHT(rectangle1_weights[2749]), .RECT2_X(rectangle2_xs[2749]), .RECT2_Y(rectangle2_ys[2749]), .RECT2_WIDTH(rectangle2_widths[2749]), .RECT2_HEIGHT(rectangle2_heights[2749]), .RECT2_WEIGHT(rectangle2_weights[2749]), .RECT3_X(rectangle3_xs[2749]), .RECT3_Y(rectangle3_ys[2749]), .RECT3_WIDTH(rectangle3_widths[2749]), .RECT3_HEIGHT(rectangle3_heights[2749]), .RECT3_WEIGHT(rectangle3_weights[2749]), .FEAT_THRES(feature_thresholds[2749]), .FEAT_ABOVE(feature_aboves[2749]), .FEAT_BELOW(feature_belows[2749])) ac2749(.scan_win(scan_win2749), .scan_win_std_dev(scan_win_std_dev[2749]), .feature_accum(feature_accums[2749]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2750]), .RECT1_Y(rectangle1_ys[2750]), .RECT1_WIDTH(rectangle1_widths[2750]), .RECT1_HEIGHT(rectangle1_heights[2750]), .RECT1_WEIGHT(rectangle1_weights[2750]), .RECT2_X(rectangle2_xs[2750]), .RECT2_Y(rectangle2_ys[2750]), .RECT2_WIDTH(rectangle2_widths[2750]), .RECT2_HEIGHT(rectangle2_heights[2750]), .RECT2_WEIGHT(rectangle2_weights[2750]), .RECT3_X(rectangle3_xs[2750]), .RECT3_Y(rectangle3_ys[2750]), .RECT3_WIDTH(rectangle3_widths[2750]), .RECT3_HEIGHT(rectangle3_heights[2750]), .RECT3_WEIGHT(rectangle3_weights[2750]), .FEAT_THRES(feature_thresholds[2750]), .FEAT_ABOVE(feature_aboves[2750]), .FEAT_BELOW(feature_belows[2750])) ac2750(.scan_win(scan_win2750), .scan_win_std_dev(scan_win_std_dev[2750]), .feature_accum(feature_accums[2750]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2751]), .RECT1_Y(rectangle1_ys[2751]), .RECT1_WIDTH(rectangle1_widths[2751]), .RECT1_HEIGHT(rectangle1_heights[2751]), .RECT1_WEIGHT(rectangle1_weights[2751]), .RECT2_X(rectangle2_xs[2751]), .RECT2_Y(rectangle2_ys[2751]), .RECT2_WIDTH(rectangle2_widths[2751]), .RECT2_HEIGHT(rectangle2_heights[2751]), .RECT2_WEIGHT(rectangle2_weights[2751]), .RECT3_X(rectangle3_xs[2751]), .RECT3_Y(rectangle3_ys[2751]), .RECT3_WIDTH(rectangle3_widths[2751]), .RECT3_HEIGHT(rectangle3_heights[2751]), .RECT3_WEIGHT(rectangle3_weights[2751]), .FEAT_THRES(feature_thresholds[2751]), .FEAT_ABOVE(feature_aboves[2751]), .FEAT_BELOW(feature_belows[2751])) ac2751(.scan_win(scan_win2751), .scan_win_std_dev(scan_win_std_dev[2751]), .feature_accum(feature_accums[2751]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2752]), .RECT1_Y(rectangle1_ys[2752]), .RECT1_WIDTH(rectangle1_widths[2752]), .RECT1_HEIGHT(rectangle1_heights[2752]), .RECT1_WEIGHT(rectangle1_weights[2752]), .RECT2_X(rectangle2_xs[2752]), .RECT2_Y(rectangle2_ys[2752]), .RECT2_WIDTH(rectangle2_widths[2752]), .RECT2_HEIGHT(rectangle2_heights[2752]), .RECT2_WEIGHT(rectangle2_weights[2752]), .RECT3_X(rectangle3_xs[2752]), .RECT3_Y(rectangle3_ys[2752]), .RECT3_WIDTH(rectangle3_widths[2752]), .RECT3_HEIGHT(rectangle3_heights[2752]), .RECT3_WEIGHT(rectangle3_weights[2752]), .FEAT_THRES(feature_thresholds[2752]), .FEAT_ABOVE(feature_aboves[2752]), .FEAT_BELOW(feature_belows[2752])) ac2752(.scan_win(scan_win2752), .scan_win_std_dev(scan_win_std_dev[2752]), .feature_accum(feature_accums[2752]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2753]), .RECT1_Y(rectangle1_ys[2753]), .RECT1_WIDTH(rectangle1_widths[2753]), .RECT1_HEIGHT(rectangle1_heights[2753]), .RECT1_WEIGHT(rectangle1_weights[2753]), .RECT2_X(rectangle2_xs[2753]), .RECT2_Y(rectangle2_ys[2753]), .RECT2_WIDTH(rectangle2_widths[2753]), .RECT2_HEIGHT(rectangle2_heights[2753]), .RECT2_WEIGHT(rectangle2_weights[2753]), .RECT3_X(rectangle3_xs[2753]), .RECT3_Y(rectangle3_ys[2753]), .RECT3_WIDTH(rectangle3_widths[2753]), .RECT3_HEIGHT(rectangle3_heights[2753]), .RECT3_WEIGHT(rectangle3_weights[2753]), .FEAT_THRES(feature_thresholds[2753]), .FEAT_ABOVE(feature_aboves[2753]), .FEAT_BELOW(feature_belows[2753])) ac2753(.scan_win(scan_win2753), .scan_win_std_dev(scan_win_std_dev[2753]), .feature_accum(feature_accums[2753]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2754]), .RECT1_Y(rectangle1_ys[2754]), .RECT1_WIDTH(rectangle1_widths[2754]), .RECT1_HEIGHT(rectangle1_heights[2754]), .RECT1_WEIGHT(rectangle1_weights[2754]), .RECT2_X(rectangle2_xs[2754]), .RECT2_Y(rectangle2_ys[2754]), .RECT2_WIDTH(rectangle2_widths[2754]), .RECT2_HEIGHT(rectangle2_heights[2754]), .RECT2_WEIGHT(rectangle2_weights[2754]), .RECT3_X(rectangle3_xs[2754]), .RECT3_Y(rectangle3_ys[2754]), .RECT3_WIDTH(rectangle3_widths[2754]), .RECT3_HEIGHT(rectangle3_heights[2754]), .RECT3_WEIGHT(rectangle3_weights[2754]), .FEAT_THRES(feature_thresholds[2754]), .FEAT_ABOVE(feature_aboves[2754]), .FEAT_BELOW(feature_belows[2754])) ac2754(.scan_win(scan_win2754), .scan_win_std_dev(scan_win_std_dev[2754]), .feature_accum(feature_accums[2754]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2755]), .RECT1_Y(rectangle1_ys[2755]), .RECT1_WIDTH(rectangle1_widths[2755]), .RECT1_HEIGHT(rectangle1_heights[2755]), .RECT1_WEIGHT(rectangle1_weights[2755]), .RECT2_X(rectangle2_xs[2755]), .RECT2_Y(rectangle2_ys[2755]), .RECT2_WIDTH(rectangle2_widths[2755]), .RECT2_HEIGHT(rectangle2_heights[2755]), .RECT2_WEIGHT(rectangle2_weights[2755]), .RECT3_X(rectangle3_xs[2755]), .RECT3_Y(rectangle3_ys[2755]), .RECT3_WIDTH(rectangle3_widths[2755]), .RECT3_HEIGHT(rectangle3_heights[2755]), .RECT3_WEIGHT(rectangle3_weights[2755]), .FEAT_THRES(feature_thresholds[2755]), .FEAT_ABOVE(feature_aboves[2755]), .FEAT_BELOW(feature_belows[2755])) ac2755(.scan_win(scan_win2755), .scan_win_std_dev(scan_win_std_dev[2755]), .feature_accum(feature_accums[2755]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2756]), .RECT1_Y(rectangle1_ys[2756]), .RECT1_WIDTH(rectangle1_widths[2756]), .RECT1_HEIGHT(rectangle1_heights[2756]), .RECT1_WEIGHT(rectangle1_weights[2756]), .RECT2_X(rectangle2_xs[2756]), .RECT2_Y(rectangle2_ys[2756]), .RECT2_WIDTH(rectangle2_widths[2756]), .RECT2_HEIGHT(rectangle2_heights[2756]), .RECT2_WEIGHT(rectangle2_weights[2756]), .RECT3_X(rectangle3_xs[2756]), .RECT3_Y(rectangle3_ys[2756]), .RECT3_WIDTH(rectangle3_widths[2756]), .RECT3_HEIGHT(rectangle3_heights[2756]), .RECT3_WEIGHT(rectangle3_weights[2756]), .FEAT_THRES(feature_thresholds[2756]), .FEAT_ABOVE(feature_aboves[2756]), .FEAT_BELOW(feature_belows[2756])) ac2756(.scan_win(scan_win2756), .scan_win_std_dev(scan_win_std_dev[2756]), .feature_accum(feature_accums[2756]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2757]), .RECT1_Y(rectangle1_ys[2757]), .RECT1_WIDTH(rectangle1_widths[2757]), .RECT1_HEIGHT(rectangle1_heights[2757]), .RECT1_WEIGHT(rectangle1_weights[2757]), .RECT2_X(rectangle2_xs[2757]), .RECT2_Y(rectangle2_ys[2757]), .RECT2_WIDTH(rectangle2_widths[2757]), .RECT2_HEIGHT(rectangle2_heights[2757]), .RECT2_WEIGHT(rectangle2_weights[2757]), .RECT3_X(rectangle3_xs[2757]), .RECT3_Y(rectangle3_ys[2757]), .RECT3_WIDTH(rectangle3_widths[2757]), .RECT3_HEIGHT(rectangle3_heights[2757]), .RECT3_WEIGHT(rectangle3_weights[2757]), .FEAT_THRES(feature_thresholds[2757]), .FEAT_ABOVE(feature_aboves[2757]), .FEAT_BELOW(feature_belows[2757])) ac2757(.scan_win(scan_win2757), .scan_win_std_dev(scan_win_std_dev[2757]), .feature_accum(feature_accums[2757]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2758]), .RECT1_Y(rectangle1_ys[2758]), .RECT1_WIDTH(rectangle1_widths[2758]), .RECT1_HEIGHT(rectangle1_heights[2758]), .RECT1_WEIGHT(rectangle1_weights[2758]), .RECT2_X(rectangle2_xs[2758]), .RECT2_Y(rectangle2_ys[2758]), .RECT2_WIDTH(rectangle2_widths[2758]), .RECT2_HEIGHT(rectangle2_heights[2758]), .RECT2_WEIGHT(rectangle2_weights[2758]), .RECT3_X(rectangle3_xs[2758]), .RECT3_Y(rectangle3_ys[2758]), .RECT3_WIDTH(rectangle3_widths[2758]), .RECT3_HEIGHT(rectangle3_heights[2758]), .RECT3_WEIGHT(rectangle3_weights[2758]), .FEAT_THRES(feature_thresholds[2758]), .FEAT_ABOVE(feature_aboves[2758]), .FEAT_BELOW(feature_belows[2758])) ac2758(.scan_win(scan_win2758), .scan_win_std_dev(scan_win_std_dev[2758]), .feature_accum(feature_accums[2758]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2759]), .RECT1_Y(rectangle1_ys[2759]), .RECT1_WIDTH(rectangle1_widths[2759]), .RECT1_HEIGHT(rectangle1_heights[2759]), .RECT1_WEIGHT(rectangle1_weights[2759]), .RECT2_X(rectangle2_xs[2759]), .RECT2_Y(rectangle2_ys[2759]), .RECT2_WIDTH(rectangle2_widths[2759]), .RECT2_HEIGHT(rectangle2_heights[2759]), .RECT2_WEIGHT(rectangle2_weights[2759]), .RECT3_X(rectangle3_xs[2759]), .RECT3_Y(rectangle3_ys[2759]), .RECT3_WIDTH(rectangle3_widths[2759]), .RECT3_HEIGHT(rectangle3_heights[2759]), .RECT3_WEIGHT(rectangle3_weights[2759]), .FEAT_THRES(feature_thresholds[2759]), .FEAT_ABOVE(feature_aboves[2759]), .FEAT_BELOW(feature_belows[2759])) ac2759(.scan_win(scan_win2759), .scan_win_std_dev(scan_win_std_dev[2759]), .feature_accum(feature_accums[2759]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2760]), .RECT1_Y(rectangle1_ys[2760]), .RECT1_WIDTH(rectangle1_widths[2760]), .RECT1_HEIGHT(rectangle1_heights[2760]), .RECT1_WEIGHT(rectangle1_weights[2760]), .RECT2_X(rectangle2_xs[2760]), .RECT2_Y(rectangle2_ys[2760]), .RECT2_WIDTH(rectangle2_widths[2760]), .RECT2_HEIGHT(rectangle2_heights[2760]), .RECT2_WEIGHT(rectangle2_weights[2760]), .RECT3_X(rectangle3_xs[2760]), .RECT3_Y(rectangle3_ys[2760]), .RECT3_WIDTH(rectangle3_widths[2760]), .RECT3_HEIGHT(rectangle3_heights[2760]), .RECT3_WEIGHT(rectangle3_weights[2760]), .FEAT_THRES(feature_thresholds[2760]), .FEAT_ABOVE(feature_aboves[2760]), .FEAT_BELOW(feature_belows[2760])) ac2760(.scan_win(scan_win2760), .scan_win_std_dev(scan_win_std_dev[2760]), .feature_accum(feature_accums[2760]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2761]), .RECT1_Y(rectangle1_ys[2761]), .RECT1_WIDTH(rectangle1_widths[2761]), .RECT1_HEIGHT(rectangle1_heights[2761]), .RECT1_WEIGHT(rectangle1_weights[2761]), .RECT2_X(rectangle2_xs[2761]), .RECT2_Y(rectangle2_ys[2761]), .RECT2_WIDTH(rectangle2_widths[2761]), .RECT2_HEIGHT(rectangle2_heights[2761]), .RECT2_WEIGHT(rectangle2_weights[2761]), .RECT3_X(rectangle3_xs[2761]), .RECT3_Y(rectangle3_ys[2761]), .RECT3_WIDTH(rectangle3_widths[2761]), .RECT3_HEIGHT(rectangle3_heights[2761]), .RECT3_WEIGHT(rectangle3_weights[2761]), .FEAT_THRES(feature_thresholds[2761]), .FEAT_ABOVE(feature_aboves[2761]), .FEAT_BELOW(feature_belows[2761])) ac2761(.scan_win(scan_win2761), .scan_win_std_dev(scan_win_std_dev[2761]), .feature_accum(feature_accums[2761]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2762]), .RECT1_Y(rectangle1_ys[2762]), .RECT1_WIDTH(rectangle1_widths[2762]), .RECT1_HEIGHT(rectangle1_heights[2762]), .RECT1_WEIGHT(rectangle1_weights[2762]), .RECT2_X(rectangle2_xs[2762]), .RECT2_Y(rectangle2_ys[2762]), .RECT2_WIDTH(rectangle2_widths[2762]), .RECT2_HEIGHT(rectangle2_heights[2762]), .RECT2_WEIGHT(rectangle2_weights[2762]), .RECT3_X(rectangle3_xs[2762]), .RECT3_Y(rectangle3_ys[2762]), .RECT3_WIDTH(rectangle3_widths[2762]), .RECT3_HEIGHT(rectangle3_heights[2762]), .RECT3_WEIGHT(rectangle3_weights[2762]), .FEAT_THRES(feature_thresholds[2762]), .FEAT_ABOVE(feature_aboves[2762]), .FEAT_BELOW(feature_belows[2762])) ac2762(.scan_win(scan_win2762), .scan_win_std_dev(scan_win_std_dev[2762]), .feature_accum(feature_accums[2762]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2763]), .RECT1_Y(rectangle1_ys[2763]), .RECT1_WIDTH(rectangle1_widths[2763]), .RECT1_HEIGHT(rectangle1_heights[2763]), .RECT1_WEIGHT(rectangle1_weights[2763]), .RECT2_X(rectangle2_xs[2763]), .RECT2_Y(rectangle2_ys[2763]), .RECT2_WIDTH(rectangle2_widths[2763]), .RECT2_HEIGHT(rectangle2_heights[2763]), .RECT2_WEIGHT(rectangle2_weights[2763]), .RECT3_X(rectangle3_xs[2763]), .RECT3_Y(rectangle3_ys[2763]), .RECT3_WIDTH(rectangle3_widths[2763]), .RECT3_HEIGHT(rectangle3_heights[2763]), .RECT3_WEIGHT(rectangle3_weights[2763]), .FEAT_THRES(feature_thresholds[2763]), .FEAT_ABOVE(feature_aboves[2763]), .FEAT_BELOW(feature_belows[2763])) ac2763(.scan_win(scan_win2763), .scan_win_std_dev(scan_win_std_dev[2763]), .feature_accum(feature_accums[2763]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2764]), .RECT1_Y(rectangle1_ys[2764]), .RECT1_WIDTH(rectangle1_widths[2764]), .RECT1_HEIGHT(rectangle1_heights[2764]), .RECT1_WEIGHT(rectangle1_weights[2764]), .RECT2_X(rectangle2_xs[2764]), .RECT2_Y(rectangle2_ys[2764]), .RECT2_WIDTH(rectangle2_widths[2764]), .RECT2_HEIGHT(rectangle2_heights[2764]), .RECT2_WEIGHT(rectangle2_weights[2764]), .RECT3_X(rectangle3_xs[2764]), .RECT3_Y(rectangle3_ys[2764]), .RECT3_WIDTH(rectangle3_widths[2764]), .RECT3_HEIGHT(rectangle3_heights[2764]), .RECT3_WEIGHT(rectangle3_weights[2764]), .FEAT_THRES(feature_thresholds[2764]), .FEAT_ABOVE(feature_aboves[2764]), .FEAT_BELOW(feature_belows[2764])) ac2764(.scan_win(scan_win2764), .scan_win_std_dev(scan_win_std_dev[2764]), .feature_accum(feature_accums[2764]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2765]), .RECT1_Y(rectangle1_ys[2765]), .RECT1_WIDTH(rectangle1_widths[2765]), .RECT1_HEIGHT(rectangle1_heights[2765]), .RECT1_WEIGHT(rectangle1_weights[2765]), .RECT2_X(rectangle2_xs[2765]), .RECT2_Y(rectangle2_ys[2765]), .RECT2_WIDTH(rectangle2_widths[2765]), .RECT2_HEIGHT(rectangle2_heights[2765]), .RECT2_WEIGHT(rectangle2_weights[2765]), .RECT3_X(rectangle3_xs[2765]), .RECT3_Y(rectangle3_ys[2765]), .RECT3_WIDTH(rectangle3_widths[2765]), .RECT3_HEIGHT(rectangle3_heights[2765]), .RECT3_WEIGHT(rectangle3_weights[2765]), .FEAT_THRES(feature_thresholds[2765]), .FEAT_ABOVE(feature_aboves[2765]), .FEAT_BELOW(feature_belows[2765])) ac2765(.scan_win(scan_win2765), .scan_win_std_dev(scan_win_std_dev[2765]), .feature_accum(feature_accums[2765]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2766]), .RECT1_Y(rectangle1_ys[2766]), .RECT1_WIDTH(rectangle1_widths[2766]), .RECT1_HEIGHT(rectangle1_heights[2766]), .RECT1_WEIGHT(rectangle1_weights[2766]), .RECT2_X(rectangle2_xs[2766]), .RECT2_Y(rectangle2_ys[2766]), .RECT2_WIDTH(rectangle2_widths[2766]), .RECT2_HEIGHT(rectangle2_heights[2766]), .RECT2_WEIGHT(rectangle2_weights[2766]), .RECT3_X(rectangle3_xs[2766]), .RECT3_Y(rectangle3_ys[2766]), .RECT3_WIDTH(rectangle3_widths[2766]), .RECT3_HEIGHT(rectangle3_heights[2766]), .RECT3_WEIGHT(rectangle3_weights[2766]), .FEAT_THRES(feature_thresholds[2766]), .FEAT_ABOVE(feature_aboves[2766]), .FEAT_BELOW(feature_belows[2766])) ac2766(.scan_win(scan_win2766), .scan_win_std_dev(scan_win_std_dev[2766]), .feature_accum(feature_accums[2766]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2767]), .RECT1_Y(rectangle1_ys[2767]), .RECT1_WIDTH(rectangle1_widths[2767]), .RECT1_HEIGHT(rectangle1_heights[2767]), .RECT1_WEIGHT(rectangle1_weights[2767]), .RECT2_X(rectangle2_xs[2767]), .RECT2_Y(rectangle2_ys[2767]), .RECT2_WIDTH(rectangle2_widths[2767]), .RECT2_HEIGHT(rectangle2_heights[2767]), .RECT2_WEIGHT(rectangle2_weights[2767]), .RECT3_X(rectangle3_xs[2767]), .RECT3_Y(rectangle3_ys[2767]), .RECT3_WIDTH(rectangle3_widths[2767]), .RECT3_HEIGHT(rectangle3_heights[2767]), .RECT3_WEIGHT(rectangle3_weights[2767]), .FEAT_THRES(feature_thresholds[2767]), .FEAT_ABOVE(feature_aboves[2767]), .FEAT_BELOW(feature_belows[2767])) ac2767(.scan_win(scan_win2767), .scan_win_std_dev(scan_win_std_dev[2767]), .feature_accum(feature_accums[2767]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2768]), .RECT1_Y(rectangle1_ys[2768]), .RECT1_WIDTH(rectangle1_widths[2768]), .RECT1_HEIGHT(rectangle1_heights[2768]), .RECT1_WEIGHT(rectangle1_weights[2768]), .RECT2_X(rectangle2_xs[2768]), .RECT2_Y(rectangle2_ys[2768]), .RECT2_WIDTH(rectangle2_widths[2768]), .RECT2_HEIGHT(rectangle2_heights[2768]), .RECT2_WEIGHT(rectangle2_weights[2768]), .RECT3_X(rectangle3_xs[2768]), .RECT3_Y(rectangle3_ys[2768]), .RECT3_WIDTH(rectangle3_widths[2768]), .RECT3_HEIGHT(rectangle3_heights[2768]), .RECT3_WEIGHT(rectangle3_weights[2768]), .FEAT_THRES(feature_thresholds[2768]), .FEAT_ABOVE(feature_aboves[2768]), .FEAT_BELOW(feature_belows[2768])) ac2768(.scan_win(scan_win2768), .scan_win_std_dev(scan_win_std_dev[2768]), .feature_accum(feature_accums[2768]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2769]), .RECT1_Y(rectangle1_ys[2769]), .RECT1_WIDTH(rectangle1_widths[2769]), .RECT1_HEIGHT(rectangle1_heights[2769]), .RECT1_WEIGHT(rectangle1_weights[2769]), .RECT2_X(rectangle2_xs[2769]), .RECT2_Y(rectangle2_ys[2769]), .RECT2_WIDTH(rectangle2_widths[2769]), .RECT2_HEIGHT(rectangle2_heights[2769]), .RECT2_WEIGHT(rectangle2_weights[2769]), .RECT3_X(rectangle3_xs[2769]), .RECT3_Y(rectangle3_ys[2769]), .RECT3_WIDTH(rectangle3_widths[2769]), .RECT3_HEIGHT(rectangle3_heights[2769]), .RECT3_WEIGHT(rectangle3_weights[2769]), .FEAT_THRES(feature_thresholds[2769]), .FEAT_ABOVE(feature_aboves[2769]), .FEAT_BELOW(feature_belows[2769])) ac2769(.scan_win(scan_win2769), .scan_win_std_dev(scan_win_std_dev[2769]), .feature_accum(feature_accums[2769]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2770]), .RECT1_Y(rectangle1_ys[2770]), .RECT1_WIDTH(rectangle1_widths[2770]), .RECT1_HEIGHT(rectangle1_heights[2770]), .RECT1_WEIGHT(rectangle1_weights[2770]), .RECT2_X(rectangle2_xs[2770]), .RECT2_Y(rectangle2_ys[2770]), .RECT2_WIDTH(rectangle2_widths[2770]), .RECT2_HEIGHT(rectangle2_heights[2770]), .RECT2_WEIGHT(rectangle2_weights[2770]), .RECT3_X(rectangle3_xs[2770]), .RECT3_Y(rectangle3_ys[2770]), .RECT3_WIDTH(rectangle3_widths[2770]), .RECT3_HEIGHT(rectangle3_heights[2770]), .RECT3_WEIGHT(rectangle3_weights[2770]), .FEAT_THRES(feature_thresholds[2770]), .FEAT_ABOVE(feature_aboves[2770]), .FEAT_BELOW(feature_belows[2770])) ac2770(.scan_win(scan_win2770), .scan_win_std_dev(scan_win_std_dev[2770]), .feature_accum(feature_accums[2770]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2771]), .RECT1_Y(rectangle1_ys[2771]), .RECT1_WIDTH(rectangle1_widths[2771]), .RECT1_HEIGHT(rectangle1_heights[2771]), .RECT1_WEIGHT(rectangle1_weights[2771]), .RECT2_X(rectangle2_xs[2771]), .RECT2_Y(rectangle2_ys[2771]), .RECT2_WIDTH(rectangle2_widths[2771]), .RECT2_HEIGHT(rectangle2_heights[2771]), .RECT2_WEIGHT(rectangle2_weights[2771]), .RECT3_X(rectangle3_xs[2771]), .RECT3_Y(rectangle3_ys[2771]), .RECT3_WIDTH(rectangle3_widths[2771]), .RECT3_HEIGHT(rectangle3_heights[2771]), .RECT3_WEIGHT(rectangle3_weights[2771]), .FEAT_THRES(feature_thresholds[2771]), .FEAT_ABOVE(feature_aboves[2771]), .FEAT_BELOW(feature_belows[2771])) ac2771(.scan_win(scan_win2771), .scan_win_std_dev(scan_win_std_dev[2771]), .feature_accum(feature_accums[2771]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2772]), .RECT1_Y(rectangle1_ys[2772]), .RECT1_WIDTH(rectangle1_widths[2772]), .RECT1_HEIGHT(rectangle1_heights[2772]), .RECT1_WEIGHT(rectangle1_weights[2772]), .RECT2_X(rectangle2_xs[2772]), .RECT2_Y(rectangle2_ys[2772]), .RECT2_WIDTH(rectangle2_widths[2772]), .RECT2_HEIGHT(rectangle2_heights[2772]), .RECT2_WEIGHT(rectangle2_weights[2772]), .RECT3_X(rectangle3_xs[2772]), .RECT3_Y(rectangle3_ys[2772]), .RECT3_WIDTH(rectangle3_widths[2772]), .RECT3_HEIGHT(rectangle3_heights[2772]), .RECT3_WEIGHT(rectangle3_weights[2772]), .FEAT_THRES(feature_thresholds[2772]), .FEAT_ABOVE(feature_aboves[2772]), .FEAT_BELOW(feature_belows[2772])) ac2772(.scan_win(scan_win2772), .scan_win_std_dev(scan_win_std_dev[2772]), .feature_accum(feature_accums[2772]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2773]), .RECT1_Y(rectangle1_ys[2773]), .RECT1_WIDTH(rectangle1_widths[2773]), .RECT1_HEIGHT(rectangle1_heights[2773]), .RECT1_WEIGHT(rectangle1_weights[2773]), .RECT2_X(rectangle2_xs[2773]), .RECT2_Y(rectangle2_ys[2773]), .RECT2_WIDTH(rectangle2_widths[2773]), .RECT2_HEIGHT(rectangle2_heights[2773]), .RECT2_WEIGHT(rectangle2_weights[2773]), .RECT3_X(rectangle3_xs[2773]), .RECT3_Y(rectangle3_ys[2773]), .RECT3_WIDTH(rectangle3_widths[2773]), .RECT3_HEIGHT(rectangle3_heights[2773]), .RECT3_WEIGHT(rectangle3_weights[2773]), .FEAT_THRES(feature_thresholds[2773]), .FEAT_ABOVE(feature_aboves[2773]), .FEAT_BELOW(feature_belows[2773])) ac2773(.scan_win(scan_win2773), .scan_win_std_dev(scan_win_std_dev[2773]), .feature_accum(feature_accums[2773]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2774]), .RECT1_Y(rectangle1_ys[2774]), .RECT1_WIDTH(rectangle1_widths[2774]), .RECT1_HEIGHT(rectangle1_heights[2774]), .RECT1_WEIGHT(rectangle1_weights[2774]), .RECT2_X(rectangle2_xs[2774]), .RECT2_Y(rectangle2_ys[2774]), .RECT2_WIDTH(rectangle2_widths[2774]), .RECT2_HEIGHT(rectangle2_heights[2774]), .RECT2_WEIGHT(rectangle2_weights[2774]), .RECT3_X(rectangle3_xs[2774]), .RECT3_Y(rectangle3_ys[2774]), .RECT3_WIDTH(rectangle3_widths[2774]), .RECT3_HEIGHT(rectangle3_heights[2774]), .RECT3_WEIGHT(rectangle3_weights[2774]), .FEAT_THRES(feature_thresholds[2774]), .FEAT_ABOVE(feature_aboves[2774]), .FEAT_BELOW(feature_belows[2774])) ac2774(.scan_win(scan_win2774), .scan_win_std_dev(scan_win_std_dev[2774]), .feature_accum(feature_accums[2774]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2775]), .RECT1_Y(rectangle1_ys[2775]), .RECT1_WIDTH(rectangle1_widths[2775]), .RECT1_HEIGHT(rectangle1_heights[2775]), .RECT1_WEIGHT(rectangle1_weights[2775]), .RECT2_X(rectangle2_xs[2775]), .RECT2_Y(rectangle2_ys[2775]), .RECT2_WIDTH(rectangle2_widths[2775]), .RECT2_HEIGHT(rectangle2_heights[2775]), .RECT2_WEIGHT(rectangle2_weights[2775]), .RECT3_X(rectangle3_xs[2775]), .RECT3_Y(rectangle3_ys[2775]), .RECT3_WIDTH(rectangle3_widths[2775]), .RECT3_HEIGHT(rectangle3_heights[2775]), .RECT3_WEIGHT(rectangle3_weights[2775]), .FEAT_THRES(feature_thresholds[2775]), .FEAT_ABOVE(feature_aboves[2775]), .FEAT_BELOW(feature_belows[2775])) ac2775(.scan_win(scan_win2775), .scan_win_std_dev(scan_win_std_dev[2775]), .feature_accum(feature_accums[2775]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2776]), .RECT1_Y(rectangle1_ys[2776]), .RECT1_WIDTH(rectangle1_widths[2776]), .RECT1_HEIGHT(rectangle1_heights[2776]), .RECT1_WEIGHT(rectangle1_weights[2776]), .RECT2_X(rectangle2_xs[2776]), .RECT2_Y(rectangle2_ys[2776]), .RECT2_WIDTH(rectangle2_widths[2776]), .RECT2_HEIGHT(rectangle2_heights[2776]), .RECT2_WEIGHT(rectangle2_weights[2776]), .RECT3_X(rectangle3_xs[2776]), .RECT3_Y(rectangle3_ys[2776]), .RECT3_WIDTH(rectangle3_widths[2776]), .RECT3_HEIGHT(rectangle3_heights[2776]), .RECT3_WEIGHT(rectangle3_weights[2776]), .FEAT_THRES(feature_thresholds[2776]), .FEAT_ABOVE(feature_aboves[2776]), .FEAT_BELOW(feature_belows[2776])) ac2776(.scan_win(scan_win2776), .scan_win_std_dev(scan_win_std_dev[2776]), .feature_accum(feature_accums[2776]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2777]), .RECT1_Y(rectangle1_ys[2777]), .RECT1_WIDTH(rectangle1_widths[2777]), .RECT1_HEIGHT(rectangle1_heights[2777]), .RECT1_WEIGHT(rectangle1_weights[2777]), .RECT2_X(rectangle2_xs[2777]), .RECT2_Y(rectangle2_ys[2777]), .RECT2_WIDTH(rectangle2_widths[2777]), .RECT2_HEIGHT(rectangle2_heights[2777]), .RECT2_WEIGHT(rectangle2_weights[2777]), .RECT3_X(rectangle3_xs[2777]), .RECT3_Y(rectangle3_ys[2777]), .RECT3_WIDTH(rectangle3_widths[2777]), .RECT3_HEIGHT(rectangle3_heights[2777]), .RECT3_WEIGHT(rectangle3_weights[2777]), .FEAT_THRES(feature_thresholds[2777]), .FEAT_ABOVE(feature_aboves[2777]), .FEAT_BELOW(feature_belows[2777])) ac2777(.scan_win(scan_win2777), .scan_win_std_dev(scan_win_std_dev[2777]), .feature_accum(feature_accums[2777]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2778]), .RECT1_Y(rectangle1_ys[2778]), .RECT1_WIDTH(rectangle1_widths[2778]), .RECT1_HEIGHT(rectangle1_heights[2778]), .RECT1_WEIGHT(rectangle1_weights[2778]), .RECT2_X(rectangle2_xs[2778]), .RECT2_Y(rectangle2_ys[2778]), .RECT2_WIDTH(rectangle2_widths[2778]), .RECT2_HEIGHT(rectangle2_heights[2778]), .RECT2_WEIGHT(rectangle2_weights[2778]), .RECT3_X(rectangle3_xs[2778]), .RECT3_Y(rectangle3_ys[2778]), .RECT3_WIDTH(rectangle3_widths[2778]), .RECT3_HEIGHT(rectangle3_heights[2778]), .RECT3_WEIGHT(rectangle3_weights[2778]), .FEAT_THRES(feature_thresholds[2778]), .FEAT_ABOVE(feature_aboves[2778]), .FEAT_BELOW(feature_belows[2778])) ac2778(.scan_win(scan_win2778), .scan_win_std_dev(scan_win_std_dev[2778]), .feature_accum(feature_accums[2778]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2779]), .RECT1_Y(rectangle1_ys[2779]), .RECT1_WIDTH(rectangle1_widths[2779]), .RECT1_HEIGHT(rectangle1_heights[2779]), .RECT1_WEIGHT(rectangle1_weights[2779]), .RECT2_X(rectangle2_xs[2779]), .RECT2_Y(rectangle2_ys[2779]), .RECT2_WIDTH(rectangle2_widths[2779]), .RECT2_HEIGHT(rectangle2_heights[2779]), .RECT2_WEIGHT(rectangle2_weights[2779]), .RECT3_X(rectangle3_xs[2779]), .RECT3_Y(rectangle3_ys[2779]), .RECT3_WIDTH(rectangle3_widths[2779]), .RECT3_HEIGHT(rectangle3_heights[2779]), .RECT3_WEIGHT(rectangle3_weights[2779]), .FEAT_THRES(feature_thresholds[2779]), .FEAT_ABOVE(feature_aboves[2779]), .FEAT_BELOW(feature_belows[2779])) ac2779(.scan_win(scan_win2779), .scan_win_std_dev(scan_win_std_dev[2779]), .feature_accum(feature_accums[2779]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2780]), .RECT1_Y(rectangle1_ys[2780]), .RECT1_WIDTH(rectangle1_widths[2780]), .RECT1_HEIGHT(rectangle1_heights[2780]), .RECT1_WEIGHT(rectangle1_weights[2780]), .RECT2_X(rectangle2_xs[2780]), .RECT2_Y(rectangle2_ys[2780]), .RECT2_WIDTH(rectangle2_widths[2780]), .RECT2_HEIGHT(rectangle2_heights[2780]), .RECT2_WEIGHT(rectangle2_weights[2780]), .RECT3_X(rectangle3_xs[2780]), .RECT3_Y(rectangle3_ys[2780]), .RECT3_WIDTH(rectangle3_widths[2780]), .RECT3_HEIGHT(rectangle3_heights[2780]), .RECT3_WEIGHT(rectangle3_weights[2780]), .FEAT_THRES(feature_thresholds[2780]), .FEAT_ABOVE(feature_aboves[2780]), .FEAT_BELOW(feature_belows[2780])) ac2780(.scan_win(scan_win2780), .scan_win_std_dev(scan_win_std_dev[2780]), .feature_accum(feature_accums[2780]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2781]), .RECT1_Y(rectangle1_ys[2781]), .RECT1_WIDTH(rectangle1_widths[2781]), .RECT1_HEIGHT(rectangle1_heights[2781]), .RECT1_WEIGHT(rectangle1_weights[2781]), .RECT2_X(rectangle2_xs[2781]), .RECT2_Y(rectangle2_ys[2781]), .RECT2_WIDTH(rectangle2_widths[2781]), .RECT2_HEIGHT(rectangle2_heights[2781]), .RECT2_WEIGHT(rectangle2_weights[2781]), .RECT3_X(rectangle3_xs[2781]), .RECT3_Y(rectangle3_ys[2781]), .RECT3_WIDTH(rectangle3_widths[2781]), .RECT3_HEIGHT(rectangle3_heights[2781]), .RECT3_WEIGHT(rectangle3_weights[2781]), .FEAT_THRES(feature_thresholds[2781]), .FEAT_ABOVE(feature_aboves[2781]), .FEAT_BELOW(feature_belows[2781])) ac2781(.scan_win(scan_win2781), .scan_win_std_dev(scan_win_std_dev[2781]), .feature_accum(feature_accums[2781]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2782]), .RECT1_Y(rectangle1_ys[2782]), .RECT1_WIDTH(rectangle1_widths[2782]), .RECT1_HEIGHT(rectangle1_heights[2782]), .RECT1_WEIGHT(rectangle1_weights[2782]), .RECT2_X(rectangle2_xs[2782]), .RECT2_Y(rectangle2_ys[2782]), .RECT2_WIDTH(rectangle2_widths[2782]), .RECT2_HEIGHT(rectangle2_heights[2782]), .RECT2_WEIGHT(rectangle2_weights[2782]), .RECT3_X(rectangle3_xs[2782]), .RECT3_Y(rectangle3_ys[2782]), .RECT3_WIDTH(rectangle3_widths[2782]), .RECT3_HEIGHT(rectangle3_heights[2782]), .RECT3_WEIGHT(rectangle3_weights[2782]), .FEAT_THRES(feature_thresholds[2782]), .FEAT_ABOVE(feature_aboves[2782]), .FEAT_BELOW(feature_belows[2782])) ac2782(.scan_win(scan_win2782), .scan_win_std_dev(scan_win_std_dev[2782]), .feature_accum(feature_accums[2782]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2783]), .RECT1_Y(rectangle1_ys[2783]), .RECT1_WIDTH(rectangle1_widths[2783]), .RECT1_HEIGHT(rectangle1_heights[2783]), .RECT1_WEIGHT(rectangle1_weights[2783]), .RECT2_X(rectangle2_xs[2783]), .RECT2_Y(rectangle2_ys[2783]), .RECT2_WIDTH(rectangle2_widths[2783]), .RECT2_HEIGHT(rectangle2_heights[2783]), .RECT2_WEIGHT(rectangle2_weights[2783]), .RECT3_X(rectangle3_xs[2783]), .RECT3_Y(rectangle3_ys[2783]), .RECT3_WIDTH(rectangle3_widths[2783]), .RECT3_HEIGHT(rectangle3_heights[2783]), .RECT3_WEIGHT(rectangle3_weights[2783]), .FEAT_THRES(feature_thresholds[2783]), .FEAT_ABOVE(feature_aboves[2783]), .FEAT_BELOW(feature_belows[2783])) ac2783(.scan_win(scan_win2783), .scan_win_std_dev(scan_win_std_dev[2783]), .feature_accum(feature_accums[2783]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2784]), .RECT1_Y(rectangle1_ys[2784]), .RECT1_WIDTH(rectangle1_widths[2784]), .RECT1_HEIGHT(rectangle1_heights[2784]), .RECT1_WEIGHT(rectangle1_weights[2784]), .RECT2_X(rectangle2_xs[2784]), .RECT2_Y(rectangle2_ys[2784]), .RECT2_WIDTH(rectangle2_widths[2784]), .RECT2_HEIGHT(rectangle2_heights[2784]), .RECT2_WEIGHT(rectangle2_weights[2784]), .RECT3_X(rectangle3_xs[2784]), .RECT3_Y(rectangle3_ys[2784]), .RECT3_WIDTH(rectangle3_widths[2784]), .RECT3_HEIGHT(rectangle3_heights[2784]), .RECT3_WEIGHT(rectangle3_weights[2784]), .FEAT_THRES(feature_thresholds[2784]), .FEAT_ABOVE(feature_aboves[2784]), .FEAT_BELOW(feature_belows[2784])) ac2784(.scan_win(scan_win2784), .scan_win_std_dev(scan_win_std_dev[2784]), .feature_accum(feature_accums[2784]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2785]), .RECT1_Y(rectangle1_ys[2785]), .RECT1_WIDTH(rectangle1_widths[2785]), .RECT1_HEIGHT(rectangle1_heights[2785]), .RECT1_WEIGHT(rectangle1_weights[2785]), .RECT2_X(rectangle2_xs[2785]), .RECT2_Y(rectangle2_ys[2785]), .RECT2_WIDTH(rectangle2_widths[2785]), .RECT2_HEIGHT(rectangle2_heights[2785]), .RECT2_WEIGHT(rectangle2_weights[2785]), .RECT3_X(rectangle3_xs[2785]), .RECT3_Y(rectangle3_ys[2785]), .RECT3_WIDTH(rectangle3_widths[2785]), .RECT3_HEIGHT(rectangle3_heights[2785]), .RECT3_WEIGHT(rectangle3_weights[2785]), .FEAT_THRES(feature_thresholds[2785]), .FEAT_ABOVE(feature_aboves[2785]), .FEAT_BELOW(feature_belows[2785])) ac2785(.scan_win(scan_win2785), .scan_win_std_dev(scan_win_std_dev[2785]), .feature_accum(feature_accums[2785]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2786]), .RECT1_Y(rectangle1_ys[2786]), .RECT1_WIDTH(rectangle1_widths[2786]), .RECT1_HEIGHT(rectangle1_heights[2786]), .RECT1_WEIGHT(rectangle1_weights[2786]), .RECT2_X(rectangle2_xs[2786]), .RECT2_Y(rectangle2_ys[2786]), .RECT2_WIDTH(rectangle2_widths[2786]), .RECT2_HEIGHT(rectangle2_heights[2786]), .RECT2_WEIGHT(rectangle2_weights[2786]), .RECT3_X(rectangle3_xs[2786]), .RECT3_Y(rectangle3_ys[2786]), .RECT3_WIDTH(rectangle3_widths[2786]), .RECT3_HEIGHT(rectangle3_heights[2786]), .RECT3_WEIGHT(rectangle3_weights[2786]), .FEAT_THRES(feature_thresholds[2786]), .FEAT_ABOVE(feature_aboves[2786]), .FEAT_BELOW(feature_belows[2786])) ac2786(.scan_win(scan_win2786), .scan_win_std_dev(scan_win_std_dev[2786]), .feature_accum(feature_accums[2786]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2787]), .RECT1_Y(rectangle1_ys[2787]), .RECT1_WIDTH(rectangle1_widths[2787]), .RECT1_HEIGHT(rectangle1_heights[2787]), .RECT1_WEIGHT(rectangle1_weights[2787]), .RECT2_X(rectangle2_xs[2787]), .RECT2_Y(rectangle2_ys[2787]), .RECT2_WIDTH(rectangle2_widths[2787]), .RECT2_HEIGHT(rectangle2_heights[2787]), .RECT2_WEIGHT(rectangle2_weights[2787]), .RECT3_X(rectangle3_xs[2787]), .RECT3_Y(rectangle3_ys[2787]), .RECT3_WIDTH(rectangle3_widths[2787]), .RECT3_HEIGHT(rectangle3_heights[2787]), .RECT3_WEIGHT(rectangle3_weights[2787]), .FEAT_THRES(feature_thresholds[2787]), .FEAT_ABOVE(feature_aboves[2787]), .FEAT_BELOW(feature_belows[2787])) ac2787(.scan_win(scan_win2787), .scan_win_std_dev(scan_win_std_dev[2787]), .feature_accum(feature_accums[2787]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2788]), .RECT1_Y(rectangle1_ys[2788]), .RECT1_WIDTH(rectangle1_widths[2788]), .RECT1_HEIGHT(rectangle1_heights[2788]), .RECT1_WEIGHT(rectangle1_weights[2788]), .RECT2_X(rectangle2_xs[2788]), .RECT2_Y(rectangle2_ys[2788]), .RECT2_WIDTH(rectangle2_widths[2788]), .RECT2_HEIGHT(rectangle2_heights[2788]), .RECT2_WEIGHT(rectangle2_weights[2788]), .RECT3_X(rectangle3_xs[2788]), .RECT3_Y(rectangle3_ys[2788]), .RECT3_WIDTH(rectangle3_widths[2788]), .RECT3_HEIGHT(rectangle3_heights[2788]), .RECT3_WEIGHT(rectangle3_weights[2788]), .FEAT_THRES(feature_thresholds[2788]), .FEAT_ABOVE(feature_aboves[2788]), .FEAT_BELOW(feature_belows[2788])) ac2788(.scan_win(scan_win2788), .scan_win_std_dev(scan_win_std_dev[2788]), .feature_accum(feature_accums[2788]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2789]), .RECT1_Y(rectangle1_ys[2789]), .RECT1_WIDTH(rectangle1_widths[2789]), .RECT1_HEIGHT(rectangle1_heights[2789]), .RECT1_WEIGHT(rectangle1_weights[2789]), .RECT2_X(rectangle2_xs[2789]), .RECT2_Y(rectangle2_ys[2789]), .RECT2_WIDTH(rectangle2_widths[2789]), .RECT2_HEIGHT(rectangle2_heights[2789]), .RECT2_WEIGHT(rectangle2_weights[2789]), .RECT3_X(rectangle3_xs[2789]), .RECT3_Y(rectangle3_ys[2789]), .RECT3_WIDTH(rectangle3_widths[2789]), .RECT3_HEIGHT(rectangle3_heights[2789]), .RECT3_WEIGHT(rectangle3_weights[2789]), .FEAT_THRES(feature_thresholds[2789]), .FEAT_ABOVE(feature_aboves[2789]), .FEAT_BELOW(feature_belows[2789])) ac2789(.scan_win(scan_win2789), .scan_win_std_dev(scan_win_std_dev[2789]), .feature_accum(feature_accums[2789]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2790]), .RECT1_Y(rectangle1_ys[2790]), .RECT1_WIDTH(rectangle1_widths[2790]), .RECT1_HEIGHT(rectangle1_heights[2790]), .RECT1_WEIGHT(rectangle1_weights[2790]), .RECT2_X(rectangle2_xs[2790]), .RECT2_Y(rectangle2_ys[2790]), .RECT2_WIDTH(rectangle2_widths[2790]), .RECT2_HEIGHT(rectangle2_heights[2790]), .RECT2_WEIGHT(rectangle2_weights[2790]), .RECT3_X(rectangle3_xs[2790]), .RECT3_Y(rectangle3_ys[2790]), .RECT3_WIDTH(rectangle3_widths[2790]), .RECT3_HEIGHT(rectangle3_heights[2790]), .RECT3_WEIGHT(rectangle3_weights[2790]), .FEAT_THRES(feature_thresholds[2790]), .FEAT_ABOVE(feature_aboves[2790]), .FEAT_BELOW(feature_belows[2790])) ac2790(.scan_win(scan_win2790), .scan_win_std_dev(scan_win_std_dev[2790]), .feature_accum(feature_accums[2790]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2791]), .RECT1_Y(rectangle1_ys[2791]), .RECT1_WIDTH(rectangle1_widths[2791]), .RECT1_HEIGHT(rectangle1_heights[2791]), .RECT1_WEIGHT(rectangle1_weights[2791]), .RECT2_X(rectangle2_xs[2791]), .RECT2_Y(rectangle2_ys[2791]), .RECT2_WIDTH(rectangle2_widths[2791]), .RECT2_HEIGHT(rectangle2_heights[2791]), .RECT2_WEIGHT(rectangle2_weights[2791]), .RECT3_X(rectangle3_xs[2791]), .RECT3_Y(rectangle3_ys[2791]), .RECT3_WIDTH(rectangle3_widths[2791]), .RECT3_HEIGHT(rectangle3_heights[2791]), .RECT3_WEIGHT(rectangle3_weights[2791]), .FEAT_THRES(feature_thresholds[2791]), .FEAT_ABOVE(feature_aboves[2791]), .FEAT_BELOW(feature_belows[2791])) ac2791(.scan_win(scan_win2791), .scan_win_std_dev(scan_win_std_dev[2791]), .feature_accum(feature_accums[2791]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2792]), .RECT1_Y(rectangle1_ys[2792]), .RECT1_WIDTH(rectangle1_widths[2792]), .RECT1_HEIGHT(rectangle1_heights[2792]), .RECT1_WEIGHT(rectangle1_weights[2792]), .RECT2_X(rectangle2_xs[2792]), .RECT2_Y(rectangle2_ys[2792]), .RECT2_WIDTH(rectangle2_widths[2792]), .RECT2_HEIGHT(rectangle2_heights[2792]), .RECT2_WEIGHT(rectangle2_weights[2792]), .RECT3_X(rectangle3_xs[2792]), .RECT3_Y(rectangle3_ys[2792]), .RECT3_WIDTH(rectangle3_widths[2792]), .RECT3_HEIGHT(rectangle3_heights[2792]), .RECT3_WEIGHT(rectangle3_weights[2792]), .FEAT_THRES(feature_thresholds[2792]), .FEAT_ABOVE(feature_aboves[2792]), .FEAT_BELOW(feature_belows[2792])) ac2792(.scan_win(scan_win2792), .scan_win_std_dev(scan_win_std_dev[2792]), .feature_accum(feature_accums[2792]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2793]), .RECT1_Y(rectangle1_ys[2793]), .RECT1_WIDTH(rectangle1_widths[2793]), .RECT1_HEIGHT(rectangle1_heights[2793]), .RECT1_WEIGHT(rectangle1_weights[2793]), .RECT2_X(rectangle2_xs[2793]), .RECT2_Y(rectangle2_ys[2793]), .RECT2_WIDTH(rectangle2_widths[2793]), .RECT2_HEIGHT(rectangle2_heights[2793]), .RECT2_WEIGHT(rectangle2_weights[2793]), .RECT3_X(rectangle3_xs[2793]), .RECT3_Y(rectangle3_ys[2793]), .RECT3_WIDTH(rectangle3_widths[2793]), .RECT3_HEIGHT(rectangle3_heights[2793]), .RECT3_WEIGHT(rectangle3_weights[2793]), .FEAT_THRES(feature_thresholds[2793]), .FEAT_ABOVE(feature_aboves[2793]), .FEAT_BELOW(feature_belows[2793])) ac2793(.scan_win(scan_win2793), .scan_win_std_dev(scan_win_std_dev[2793]), .feature_accum(feature_accums[2793]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2794]), .RECT1_Y(rectangle1_ys[2794]), .RECT1_WIDTH(rectangle1_widths[2794]), .RECT1_HEIGHT(rectangle1_heights[2794]), .RECT1_WEIGHT(rectangle1_weights[2794]), .RECT2_X(rectangle2_xs[2794]), .RECT2_Y(rectangle2_ys[2794]), .RECT2_WIDTH(rectangle2_widths[2794]), .RECT2_HEIGHT(rectangle2_heights[2794]), .RECT2_WEIGHT(rectangle2_weights[2794]), .RECT3_X(rectangle3_xs[2794]), .RECT3_Y(rectangle3_ys[2794]), .RECT3_WIDTH(rectangle3_widths[2794]), .RECT3_HEIGHT(rectangle3_heights[2794]), .RECT3_WEIGHT(rectangle3_weights[2794]), .FEAT_THRES(feature_thresholds[2794]), .FEAT_ABOVE(feature_aboves[2794]), .FEAT_BELOW(feature_belows[2794])) ac2794(.scan_win(scan_win2794), .scan_win_std_dev(scan_win_std_dev[2794]), .feature_accum(feature_accums[2794]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2795]), .RECT1_Y(rectangle1_ys[2795]), .RECT1_WIDTH(rectangle1_widths[2795]), .RECT1_HEIGHT(rectangle1_heights[2795]), .RECT1_WEIGHT(rectangle1_weights[2795]), .RECT2_X(rectangle2_xs[2795]), .RECT2_Y(rectangle2_ys[2795]), .RECT2_WIDTH(rectangle2_widths[2795]), .RECT2_HEIGHT(rectangle2_heights[2795]), .RECT2_WEIGHT(rectangle2_weights[2795]), .RECT3_X(rectangle3_xs[2795]), .RECT3_Y(rectangle3_ys[2795]), .RECT3_WIDTH(rectangle3_widths[2795]), .RECT3_HEIGHT(rectangle3_heights[2795]), .RECT3_WEIGHT(rectangle3_weights[2795]), .FEAT_THRES(feature_thresholds[2795]), .FEAT_ABOVE(feature_aboves[2795]), .FEAT_BELOW(feature_belows[2795])) ac2795(.scan_win(scan_win2795), .scan_win_std_dev(scan_win_std_dev[2795]), .feature_accum(feature_accums[2795]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2796]), .RECT1_Y(rectangle1_ys[2796]), .RECT1_WIDTH(rectangle1_widths[2796]), .RECT1_HEIGHT(rectangle1_heights[2796]), .RECT1_WEIGHT(rectangle1_weights[2796]), .RECT2_X(rectangle2_xs[2796]), .RECT2_Y(rectangle2_ys[2796]), .RECT2_WIDTH(rectangle2_widths[2796]), .RECT2_HEIGHT(rectangle2_heights[2796]), .RECT2_WEIGHT(rectangle2_weights[2796]), .RECT3_X(rectangle3_xs[2796]), .RECT3_Y(rectangle3_ys[2796]), .RECT3_WIDTH(rectangle3_widths[2796]), .RECT3_HEIGHT(rectangle3_heights[2796]), .RECT3_WEIGHT(rectangle3_weights[2796]), .FEAT_THRES(feature_thresholds[2796]), .FEAT_ABOVE(feature_aboves[2796]), .FEAT_BELOW(feature_belows[2796])) ac2796(.scan_win(scan_win2796), .scan_win_std_dev(scan_win_std_dev[2796]), .feature_accum(feature_accums[2796]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2797]), .RECT1_Y(rectangle1_ys[2797]), .RECT1_WIDTH(rectangle1_widths[2797]), .RECT1_HEIGHT(rectangle1_heights[2797]), .RECT1_WEIGHT(rectangle1_weights[2797]), .RECT2_X(rectangle2_xs[2797]), .RECT2_Y(rectangle2_ys[2797]), .RECT2_WIDTH(rectangle2_widths[2797]), .RECT2_HEIGHT(rectangle2_heights[2797]), .RECT2_WEIGHT(rectangle2_weights[2797]), .RECT3_X(rectangle3_xs[2797]), .RECT3_Y(rectangle3_ys[2797]), .RECT3_WIDTH(rectangle3_widths[2797]), .RECT3_HEIGHT(rectangle3_heights[2797]), .RECT3_WEIGHT(rectangle3_weights[2797]), .FEAT_THRES(feature_thresholds[2797]), .FEAT_ABOVE(feature_aboves[2797]), .FEAT_BELOW(feature_belows[2797])) ac2797(.scan_win(scan_win2797), .scan_win_std_dev(scan_win_std_dev[2797]), .feature_accum(feature_accums[2797]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2798]), .RECT1_Y(rectangle1_ys[2798]), .RECT1_WIDTH(rectangle1_widths[2798]), .RECT1_HEIGHT(rectangle1_heights[2798]), .RECT1_WEIGHT(rectangle1_weights[2798]), .RECT2_X(rectangle2_xs[2798]), .RECT2_Y(rectangle2_ys[2798]), .RECT2_WIDTH(rectangle2_widths[2798]), .RECT2_HEIGHT(rectangle2_heights[2798]), .RECT2_WEIGHT(rectangle2_weights[2798]), .RECT3_X(rectangle3_xs[2798]), .RECT3_Y(rectangle3_ys[2798]), .RECT3_WIDTH(rectangle3_widths[2798]), .RECT3_HEIGHT(rectangle3_heights[2798]), .RECT3_WEIGHT(rectangle3_weights[2798]), .FEAT_THRES(feature_thresholds[2798]), .FEAT_ABOVE(feature_aboves[2798]), .FEAT_BELOW(feature_belows[2798])) ac2798(.scan_win(scan_win2798), .scan_win_std_dev(scan_win_std_dev[2798]), .feature_accum(feature_accums[2798]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2799]), .RECT1_Y(rectangle1_ys[2799]), .RECT1_WIDTH(rectangle1_widths[2799]), .RECT1_HEIGHT(rectangle1_heights[2799]), .RECT1_WEIGHT(rectangle1_weights[2799]), .RECT2_X(rectangle2_xs[2799]), .RECT2_Y(rectangle2_ys[2799]), .RECT2_WIDTH(rectangle2_widths[2799]), .RECT2_HEIGHT(rectangle2_heights[2799]), .RECT2_WEIGHT(rectangle2_weights[2799]), .RECT3_X(rectangle3_xs[2799]), .RECT3_Y(rectangle3_ys[2799]), .RECT3_WIDTH(rectangle3_widths[2799]), .RECT3_HEIGHT(rectangle3_heights[2799]), .RECT3_WEIGHT(rectangle3_weights[2799]), .FEAT_THRES(feature_thresholds[2799]), .FEAT_ABOVE(feature_aboves[2799]), .FEAT_BELOW(feature_belows[2799])) ac2799(.scan_win(scan_win2799), .scan_win_std_dev(scan_win_std_dev[2799]), .feature_accum(feature_accums[2799]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2800]), .RECT1_Y(rectangle1_ys[2800]), .RECT1_WIDTH(rectangle1_widths[2800]), .RECT1_HEIGHT(rectangle1_heights[2800]), .RECT1_WEIGHT(rectangle1_weights[2800]), .RECT2_X(rectangle2_xs[2800]), .RECT2_Y(rectangle2_ys[2800]), .RECT2_WIDTH(rectangle2_widths[2800]), .RECT2_HEIGHT(rectangle2_heights[2800]), .RECT2_WEIGHT(rectangle2_weights[2800]), .RECT3_X(rectangle3_xs[2800]), .RECT3_Y(rectangle3_ys[2800]), .RECT3_WIDTH(rectangle3_widths[2800]), .RECT3_HEIGHT(rectangle3_heights[2800]), .RECT3_WEIGHT(rectangle3_weights[2800]), .FEAT_THRES(feature_thresholds[2800]), .FEAT_ABOVE(feature_aboves[2800]), .FEAT_BELOW(feature_belows[2800])) ac2800(.scan_win(scan_win2800), .scan_win_std_dev(scan_win_std_dev[2800]), .feature_accum(feature_accums[2800]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2801]), .RECT1_Y(rectangle1_ys[2801]), .RECT1_WIDTH(rectangle1_widths[2801]), .RECT1_HEIGHT(rectangle1_heights[2801]), .RECT1_WEIGHT(rectangle1_weights[2801]), .RECT2_X(rectangle2_xs[2801]), .RECT2_Y(rectangle2_ys[2801]), .RECT2_WIDTH(rectangle2_widths[2801]), .RECT2_HEIGHT(rectangle2_heights[2801]), .RECT2_WEIGHT(rectangle2_weights[2801]), .RECT3_X(rectangle3_xs[2801]), .RECT3_Y(rectangle3_ys[2801]), .RECT3_WIDTH(rectangle3_widths[2801]), .RECT3_HEIGHT(rectangle3_heights[2801]), .RECT3_WEIGHT(rectangle3_weights[2801]), .FEAT_THRES(feature_thresholds[2801]), .FEAT_ABOVE(feature_aboves[2801]), .FEAT_BELOW(feature_belows[2801])) ac2801(.scan_win(scan_win2801), .scan_win_std_dev(scan_win_std_dev[2801]), .feature_accum(feature_accums[2801]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2802]), .RECT1_Y(rectangle1_ys[2802]), .RECT1_WIDTH(rectangle1_widths[2802]), .RECT1_HEIGHT(rectangle1_heights[2802]), .RECT1_WEIGHT(rectangle1_weights[2802]), .RECT2_X(rectangle2_xs[2802]), .RECT2_Y(rectangle2_ys[2802]), .RECT2_WIDTH(rectangle2_widths[2802]), .RECT2_HEIGHT(rectangle2_heights[2802]), .RECT2_WEIGHT(rectangle2_weights[2802]), .RECT3_X(rectangle3_xs[2802]), .RECT3_Y(rectangle3_ys[2802]), .RECT3_WIDTH(rectangle3_widths[2802]), .RECT3_HEIGHT(rectangle3_heights[2802]), .RECT3_WEIGHT(rectangle3_weights[2802]), .FEAT_THRES(feature_thresholds[2802]), .FEAT_ABOVE(feature_aboves[2802]), .FEAT_BELOW(feature_belows[2802])) ac2802(.scan_win(scan_win2802), .scan_win_std_dev(scan_win_std_dev[2802]), .feature_accum(feature_accums[2802]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2803]), .RECT1_Y(rectangle1_ys[2803]), .RECT1_WIDTH(rectangle1_widths[2803]), .RECT1_HEIGHT(rectangle1_heights[2803]), .RECT1_WEIGHT(rectangle1_weights[2803]), .RECT2_X(rectangle2_xs[2803]), .RECT2_Y(rectangle2_ys[2803]), .RECT2_WIDTH(rectangle2_widths[2803]), .RECT2_HEIGHT(rectangle2_heights[2803]), .RECT2_WEIGHT(rectangle2_weights[2803]), .RECT3_X(rectangle3_xs[2803]), .RECT3_Y(rectangle3_ys[2803]), .RECT3_WIDTH(rectangle3_widths[2803]), .RECT3_HEIGHT(rectangle3_heights[2803]), .RECT3_WEIGHT(rectangle3_weights[2803]), .FEAT_THRES(feature_thresholds[2803]), .FEAT_ABOVE(feature_aboves[2803]), .FEAT_BELOW(feature_belows[2803])) ac2803(.scan_win(scan_win2803), .scan_win_std_dev(scan_win_std_dev[2803]), .feature_accum(feature_accums[2803]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2804]), .RECT1_Y(rectangle1_ys[2804]), .RECT1_WIDTH(rectangle1_widths[2804]), .RECT1_HEIGHT(rectangle1_heights[2804]), .RECT1_WEIGHT(rectangle1_weights[2804]), .RECT2_X(rectangle2_xs[2804]), .RECT2_Y(rectangle2_ys[2804]), .RECT2_WIDTH(rectangle2_widths[2804]), .RECT2_HEIGHT(rectangle2_heights[2804]), .RECT2_WEIGHT(rectangle2_weights[2804]), .RECT3_X(rectangle3_xs[2804]), .RECT3_Y(rectangle3_ys[2804]), .RECT3_WIDTH(rectangle3_widths[2804]), .RECT3_HEIGHT(rectangle3_heights[2804]), .RECT3_WEIGHT(rectangle3_weights[2804]), .FEAT_THRES(feature_thresholds[2804]), .FEAT_ABOVE(feature_aboves[2804]), .FEAT_BELOW(feature_belows[2804])) ac2804(.scan_win(scan_win2804), .scan_win_std_dev(scan_win_std_dev[2804]), .feature_accum(feature_accums[2804]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2805]), .RECT1_Y(rectangle1_ys[2805]), .RECT1_WIDTH(rectangle1_widths[2805]), .RECT1_HEIGHT(rectangle1_heights[2805]), .RECT1_WEIGHT(rectangle1_weights[2805]), .RECT2_X(rectangle2_xs[2805]), .RECT2_Y(rectangle2_ys[2805]), .RECT2_WIDTH(rectangle2_widths[2805]), .RECT2_HEIGHT(rectangle2_heights[2805]), .RECT2_WEIGHT(rectangle2_weights[2805]), .RECT3_X(rectangle3_xs[2805]), .RECT3_Y(rectangle3_ys[2805]), .RECT3_WIDTH(rectangle3_widths[2805]), .RECT3_HEIGHT(rectangle3_heights[2805]), .RECT3_WEIGHT(rectangle3_weights[2805]), .FEAT_THRES(feature_thresholds[2805]), .FEAT_ABOVE(feature_aboves[2805]), .FEAT_BELOW(feature_belows[2805])) ac2805(.scan_win(scan_win2805), .scan_win_std_dev(scan_win_std_dev[2805]), .feature_accum(feature_accums[2805]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2806]), .RECT1_Y(rectangle1_ys[2806]), .RECT1_WIDTH(rectangle1_widths[2806]), .RECT1_HEIGHT(rectangle1_heights[2806]), .RECT1_WEIGHT(rectangle1_weights[2806]), .RECT2_X(rectangle2_xs[2806]), .RECT2_Y(rectangle2_ys[2806]), .RECT2_WIDTH(rectangle2_widths[2806]), .RECT2_HEIGHT(rectangle2_heights[2806]), .RECT2_WEIGHT(rectangle2_weights[2806]), .RECT3_X(rectangle3_xs[2806]), .RECT3_Y(rectangle3_ys[2806]), .RECT3_WIDTH(rectangle3_widths[2806]), .RECT3_HEIGHT(rectangle3_heights[2806]), .RECT3_WEIGHT(rectangle3_weights[2806]), .FEAT_THRES(feature_thresholds[2806]), .FEAT_ABOVE(feature_aboves[2806]), .FEAT_BELOW(feature_belows[2806])) ac2806(.scan_win(scan_win2806), .scan_win_std_dev(scan_win_std_dev[2806]), .feature_accum(feature_accums[2806]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2807]), .RECT1_Y(rectangle1_ys[2807]), .RECT1_WIDTH(rectangle1_widths[2807]), .RECT1_HEIGHT(rectangle1_heights[2807]), .RECT1_WEIGHT(rectangle1_weights[2807]), .RECT2_X(rectangle2_xs[2807]), .RECT2_Y(rectangle2_ys[2807]), .RECT2_WIDTH(rectangle2_widths[2807]), .RECT2_HEIGHT(rectangle2_heights[2807]), .RECT2_WEIGHT(rectangle2_weights[2807]), .RECT3_X(rectangle3_xs[2807]), .RECT3_Y(rectangle3_ys[2807]), .RECT3_WIDTH(rectangle3_widths[2807]), .RECT3_HEIGHT(rectangle3_heights[2807]), .RECT3_WEIGHT(rectangle3_weights[2807]), .FEAT_THRES(feature_thresholds[2807]), .FEAT_ABOVE(feature_aboves[2807]), .FEAT_BELOW(feature_belows[2807])) ac2807(.scan_win(scan_win2807), .scan_win_std_dev(scan_win_std_dev[2807]), .feature_accum(feature_accums[2807]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2808]), .RECT1_Y(rectangle1_ys[2808]), .RECT1_WIDTH(rectangle1_widths[2808]), .RECT1_HEIGHT(rectangle1_heights[2808]), .RECT1_WEIGHT(rectangle1_weights[2808]), .RECT2_X(rectangle2_xs[2808]), .RECT2_Y(rectangle2_ys[2808]), .RECT2_WIDTH(rectangle2_widths[2808]), .RECT2_HEIGHT(rectangle2_heights[2808]), .RECT2_WEIGHT(rectangle2_weights[2808]), .RECT3_X(rectangle3_xs[2808]), .RECT3_Y(rectangle3_ys[2808]), .RECT3_WIDTH(rectangle3_widths[2808]), .RECT3_HEIGHT(rectangle3_heights[2808]), .RECT3_WEIGHT(rectangle3_weights[2808]), .FEAT_THRES(feature_thresholds[2808]), .FEAT_ABOVE(feature_aboves[2808]), .FEAT_BELOW(feature_belows[2808])) ac2808(.scan_win(scan_win2808), .scan_win_std_dev(scan_win_std_dev[2808]), .feature_accum(feature_accums[2808]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2809]), .RECT1_Y(rectangle1_ys[2809]), .RECT1_WIDTH(rectangle1_widths[2809]), .RECT1_HEIGHT(rectangle1_heights[2809]), .RECT1_WEIGHT(rectangle1_weights[2809]), .RECT2_X(rectangle2_xs[2809]), .RECT2_Y(rectangle2_ys[2809]), .RECT2_WIDTH(rectangle2_widths[2809]), .RECT2_HEIGHT(rectangle2_heights[2809]), .RECT2_WEIGHT(rectangle2_weights[2809]), .RECT3_X(rectangle3_xs[2809]), .RECT3_Y(rectangle3_ys[2809]), .RECT3_WIDTH(rectangle3_widths[2809]), .RECT3_HEIGHT(rectangle3_heights[2809]), .RECT3_WEIGHT(rectangle3_weights[2809]), .FEAT_THRES(feature_thresholds[2809]), .FEAT_ABOVE(feature_aboves[2809]), .FEAT_BELOW(feature_belows[2809])) ac2809(.scan_win(scan_win2809), .scan_win_std_dev(scan_win_std_dev[2809]), .feature_accum(feature_accums[2809]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2810]), .RECT1_Y(rectangle1_ys[2810]), .RECT1_WIDTH(rectangle1_widths[2810]), .RECT1_HEIGHT(rectangle1_heights[2810]), .RECT1_WEIGHT(rectangle1_weights[2810]), .RECT2_X(rectangle2_xs[2810]), .RECT2_Y(rectangle2_ys[2810]), .RECT2_WIDTH(rectangle2_widths[2810]), .RECT2_HEIGHT(rectangle2_heights[2810]), .RECT2_WEIGHT(rectangle2_weights[2810]), .RECT3_X(rectangle3_xs[2810]), .RECT3_Y(rectangle3_ys[2810]), .RECT3_WIDTH(rectangle3_widths[2810]), .RECT3_HEIGHT(rectangle3_heights[2810]), .RECT3_WEIGHT(rectangle3_weights[2810]), .FEAT_THRES(feature_thresholds[2810]), .FEAT_ABOVE(feature_aboves[2810]), .FEAT_BELOW(feature_belows[2810])) ac2810(.scan_win(scan_win2810), .scan_win_std_dev(scan_win_std_dev[2810]), .feature_accum(feature_accums[2810]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2811]), .RECT1_Y(rectangle1_ys[2811]), .RECT1_WIDTH(rectangle1_widths[2811]), .RECT1_HEIGHT(rectangle1_heights[2811]), .RECT1_WEIGHT(rectangle1_weights[2811]), .RECT2_X(rectangle2_xs[2811]), .RECT2_Y(rectangle2_ys[2811]), .RECT2_WIDTH(rectangle2_widths[2811]), .RECT2_HEIGHT(rectangle2_heights[2811]), .RECT2_WEIGHT(rectangle2_weights[2811]), .RECT3_X(rectangle3_xs[2811]), .RECT3_Y(rectangle3_ys[2811]), .RECT3_WIDTH(rectangle3_widths[2811]), .RECT3_HEIGHT(rectangle3_heights[2811]), .RECT3_WEIGHT(rectangle3_weights[2811]), .FEAT_THRES(feature_thresholds[2811]), .FEAT_ABOVE(feature_aboves[2811]), .FEAT_BELOW(feature_belows[2811])) ac2811(.scan_win(scan_win2811), .scan_win_std_dev(scan_win_std_dev[2811]), .feature_accum(feature_accums[2811]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2812]), .RECT1_Y(rectangle1_ys[2812]), .RECT1_WIDTH(rectangle1_widths[2812]), .RECT1_HEIGHT(rectangle1_heights[2812]), .RECT1_WEIGHT(rectangle1_weights[2812]), .RECT2_X(rectangle2_xs[2812]), .RECT2_Y(rectangle2_ys[2812]), .RECT2_WIDTH(rectangle2_widths[2812]), .RECT2_HEIGHT(rectangle2_heights[2812]), .RECT2_WEIGHT(rectangle2_weights[2812]), .RECT3_X(rectangle3_xs[2812]), .RECT3_Y(rectangle3_ys[2812]), .RECT3_WIDTH(rectangle3_widths[2812]), .RECT3_HEIGHT(rectangle3_heights[2812]), .RECT3_WEIGHT(rectangle3_weights[2812]), .FEAT_THRES(feature_thresholds[2812]), .FEAT_ABOVE(feature_aboves[2812]), .FEAT_BELOW(feature_belows[2812])) ac2812(.scan_win(scan_win2812), .scan_win_std_dev(scan_win_std_dev[2812]), .feature_accum(feature_accums[2812]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2813]), .RECT1_Y(rectangle1_ys[2813]), .RECT1_WIDTH(rectangle1_widths[2813]), .RECT1_HEIGHT(rectangle1_heights[2813]), .RECT1_WEIGHT(rectangle1_weights[2813]), .RECT2_X(rectangle2_xs[2813]), .RECT2_Y(rectangle2_ys[2813]), .RECT2_WIDTH(rectangle2_widths[2813]), .RECT2_HEIGHT(rectangle2_heights[2813]), .RECT2_WEIGHT(rectangle2_weights[2813]), .RECT3_X(rectangle3_xs[2813]), .RECT3_Y(rectangle3_ys[2813]), .RECT3_WIDTH(rectangle3_widths[2813]), .RECT3_HEIGHT(rectangle3_heights[2813]), .RECT3_WEIGHT(rectangle3_weights[2813]), .FEAT_THRES(feature_thresholds[2813]), .FEAT_ABOVE(feature_aboves[2813]), .FEAT_BELOW(feature_belows[2813])) ac2813(.scan_win(scan_win2813), .scan_win_std_dev(scan_win_std_dev[2813]), .feature_accum(feature_accums[2813]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2814]), .RECT1_Y(rectangle1_ys[2814]), .RECT1_WIDTH(rectangle1_widths[2814]), .RECT1_HEIGHT(rectangle1_heights[2814]), .RECT1_WEIGHT(rectangle1_weights[2814]), .RECT2_X(rectangle2_xs[2814]), .RECT2_Y(rectangle2_ys[2814]), .RECT2_WIDTH(rectangle2_widths[2814]), .RECT2_HEIGHT(rectangle2_heights[2814]), .RECT2_WEIGHT(rectangle2_weights[2814]), .RECT3_X(rectangle3_xs[2814]), .RECT3_Y(rectangle3_ys[2814]), .RECT3_WIDTH(rectangle3_widths[2814]), .RECT3_HEIGHT(rectangle3_heights[2814]), .RECT3_WEIGHT(rectangle3_weights[2814]), .FEAT_THRES(feature_thresholds[2814]), .FEAT_ABOVE(feature_aboves[2814]), .FEAT_BELOW(feature_belows[2814])) ac2814(.scan_win(scan_win2814), .scan_win_std_dev(scan_win_std_dev[2814]), .feature_accum(feature_accums[2814]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2815]), .RECT1_Y(rectangle1_ys[2815]), .RECT1_WIDTH(rectangle1_widths[2815]), .RECT1_HEIGHT(rectangle1_heights[2815]), .RECT1_WEIGHT(rectangle1_weights[2815]), .RECT2_X(rectangle2_xs[2815]), .RECT2_Y(rectangle2_ys[2815]), .RECT2_WIDTH(rectangle2_widths[2815]), .RECT2_HEIGHT(rectangle2_heights[2815]), .RECT2_WEIGHT(rectangle2_weights[2815]), .RECT3_X(rectangle3_xs[2815]), .RECT3_Y(rectangle3_ys[2815]), .RECT3_WIDTH(rectangle3_widths[2815]), .RECT3_HEIGHT(rectangle3_heights[2815]), .RECT3_WEIGHT(rectangle3_weights[2815]), .FEAT_THRES(feature_thresholds[2815]), .FEAT_ABOVE(feature_aboves[2815]), .FEAT_BELOW(feature_belows[2815])) ac2815(.scan_win(scan_win2815), .scan_win_std_dev(scan_win_std_dev[2815]), .feature_accum(feature_accums[2815]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2816]), .RECT1_Y(rectangle1_ys[2816]), .RECT1_WIDTH(rectangle1_widths[2816]), .RECT1_HEIGHT(rectangle1_heights[2816]), .RECT1_WEIGHT(rectangle1_weights[2816]), .RECT2_X(rectangle2_xs[2816]), .RECT2_Y(rectangle2_ys[2816]), .RECT2_WIDTH(rectangle2_widths[2816]), .RECT2_HEIGHT(rectangle2_heights[2816]), .RECT2_WEIGHT(rectangle2_weights[2816]), .RECT3_X(rectangle3_xs[2816]), .RECT3_Y(rectangle3_ys[2816]), .RECT3_WIDTH(rectangle3_widths[2816]), .RECT3_HEIGHT(rectangle3_heights[2816]), .RECT3_WEIGHT(rectangle3_weights[2816]), .FEAT_THRES(feature_thresholds[2816]), .FEAT_ABOVE(feature_aboves[2816]), .FEAT_BELOW(feature_belows[2816])) ac2816(.scan_win(scan_win2816), .scan_win_std_dev(scan_win_std_dev[2816]), .feature_accum(feature_accums[2816]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2817]), .RECT1_Y(rectangle1_ys[2817]), .RECT1_WIDTH(rectangle1_widths[2817]), .RECT1_HEIGHT(rectangle1_heights[2817]), .RECT1_WEIGHT(rectangle1_weights[2817]), .RECT2_X(rectangle2_xs[2817]), .RECT2_Y(rectangle2_ys[2817]), .RECT2_WIDTH(rectangle2_widths[2817]), .RECT2_HEIGHT(rectangle2_heights[2817]), .RECT2_WEIGHT(rectangle2_weights[2817]), .RECT3_X(rectangle3_xs[2817]), .RECT3_Y(rectangle3_ys[2817]), .RECT3_WIDTH(rectangle3_widths[2817]), .RECT3_HEIGHT(rectangle3_heights[2817]), .RECT3_WEIGHT(rectangle3_weights[2817]), .FEAT_THRES(feature_thresholds[2817]), .FEAT_ABOVE(feature_aboves[2817]), .FEAT_BELOW(feature_belows[2817])) ac2817(.scan_win(scan_win2817), .scan_win_std_dev(scan_win_std_dev[2817]), .feature_accum(feature_accums[2817]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2818]), .RECT1_Y(rectangle1_ys[2818]), .RECT1_WIDTH(rectangle1_widths[2818]), .RECT1_HEIGHT(rectangle1_heights[2818]), .RECT1_WEIGHT(rectangle1_weights[2818]), .RECT2_X(rectangle2_xs[2818]), .RECT2_Y(rectangle2_ys[2818]), .RECT2_WIDTH(rectangle2_widths[2818]), .RECT2_HEIGHT(rectangle2_heights[2818]), .RECT2_WEIGHT(rectangle2_weights[2818]), .RECT3_X(rectangle3_xs[2818]), .RECT3_Y(rectangle3_ys[2818]), .RECT3_WIDTH(rectangle3_widths[2818]), .RECT3_HEIGHT(rectangle3_heights[2818]), .RECT3_WEIGHT(rectangle3_weights[2818]), .FEAT_THRES(feature_thresholds[2818]), .FEAT_ABOVE(feature_aboves[2818]), .FEAT_BELOW(feature_belows[2818])) ac2818(.scan_win(scan_win2818), .scan_win_std_dev(scan_win_std_dev[2818]), .feature_accum(feature_accums[2818]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2819]), .RECT1_Y(rectangle1_ys[2819]), .RECT1_WIDTH(rectangle1_widths[2819]), .RECT1_HEIGHT(rectangle1_heights[2819]), .RECT1_WEIGHT(rectangle1_weights[2819]), .RECT2_X(rectangle2_xs[2819]), .RECT2_Y(rectangle2_ys[2819]), .RECT2_WIDTH(rectangle2_widths[2819]), .RECT2_HEIGHT(rectangle2_heights[2819]), .RECT2_WEIGHT(rectangle2_weights[2819]), .RECT3_X(rectangle3_xs[2819]), .RECT3_Y(rectangle3_ys[2819]), .RECT3_WIDTH(rectangle3_widths[2819]), .RECT3_HEIGHT(rectangle3_heights[2819]), .RECT3_WEIGHT(rectangle3_weights[2819]), .FEAT_THRES(feature_thresholds[2819]), .FEAT_ABOVE(feature_aboves[2819]), .FEAT_BELOW(feature_belows[2819])) ac2819(.scan_win(scan_win2819), .scan_win_std_dev(scan_win_std_dev[2819]), .feature_accum(feature_accums[2819]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2820]), .RECT1_Y(rectangle1_ys[2820]), .RECT1_WIDTH(rectangle1_widths[2820]), .RECT1_HEIGHT(rectangle1_heights[2820]), .RECT1_WEIGHT(rectangle1_weights[2820]), .RECT2_X(rectangle2_xs[2820]), .RECT2_Y(rectangle2_ys[2820]), .RECT2_WIDTH(rectangle2_widths[2820]), .RECT2_HEIGHT(rectangle2_heights[2820]), .RECT2_WEIGHT(rectangle2_weights[2820]), .RECT3_X(rectangle3_xs[2820]), .RECT3_Y(rectangle3_ys[2820]), .RECT3_WIDTH(rectangle3_widths[2820]), .RECT3_HEIGHT(rectangle3_heights[2820]), .RECT3_WEIGHT(rectangle3_weights[2820]), .FEAT_THRES(feature_thresholds[2820]), .FEAT_ABOVE(feature_aboves[2820]), .FEAT_BELOW(feature_belows[2820])) ac2820(.scan_win(scan_win2820), .scan_win_std_dev(scan_win_std_dev[2820]), .feature_accum(feature_accums[2820]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2821]), .RECT1_Y(rectangle1_ys[2821]), .RECT1_WIDTH(rectangle1_widths[2821]), .RECT1_HEIGHT(rectangle1_heights[2821]), .RECT1_WEIGHT(rectangle1_weights[2821]), .RECT2_X(rectangle2_xs[2821]), .RECT2_Y(rectangle2_ys[2821]), .RECT2_WIDTH(rectangle2_widths[2821]), .RECT2_HEIGHT(rectangle2_heights[2821]), .RECT2_WEIGHT(rectangle2_weights[2821]), .RECT3_X(rectangle3_xs[2821]), .RECT3_Y(rectangle3_ys[2821]), .RECT3_WIDTH(rectangle3_widths[2821]), .RECT3_HEIGHT(rectangle3_heights[2821]), .RECT3_WEIGHT(rectangle3_weights[2821]), .FEAT_THRES(feature_thresholds[2821]), .FEAT_ABOVE(feature_aboves[2821]), .FEAT_BELOW(feature_belows[2821])) ac2821(.scan_win(scan_win2821), .scan_win_std_dev(scan_win_std_dev[2821]), .feature_accum(feature_accums[2821]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2822]), .RECT1_Y(rectangle1_ys[2822]), .RECT1_WIDTH(rectangle1_widths[2822]), .RECT1_HEIGHT(rectangle1_heights[2822]), .RECT1_WEIGHT(rectangle1_weights[2822]), .RECT2_X(rectangle2_xs[2822]), .RECT2_Y(rectangle2_ys[2822]), .RECT2_WIDTH(rectangle2_widths[2822]), .RECT2_HEIGHT(rectangle2_heights[2822]), .RECT2_WEIGHT(rectangle2_weights[2822]), .RECT3_X(rectangle3_xs[2822]), .RECT3_Y(rectangle3_ys[2822]), .RECT3_WIDTH(rectangle3_widths[2822]), .RECT3_HEIGHT(rectangle3_heights[2822]), .RECT3_WEIGHT(rectangle3_weights[2822]), .FEAT_THRES(feature_thresholds[2822]), .FEAT_ABOVE(feature_aboves[2822]), .FEAT_BELOW(feature_belows[2822])) ac2822(.scan_win(scan_win2822), .scan_win_std_dev(scan_win_std_dev[2822]), .feature_accum(feature_accums[2822]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2823]), .RECT1_Y(rectangle1_ys[2823]), .RECT1_WIDTH(rectangle1_widths[2823]), .RECT1_HEIGHT(rectangle1_heights[2823]), .RECT1_WEIGHT(rectangle1_weights[2823]), .RECT2_X(rectangle2_xs[2823]), .RECT2_Y(rectangle2_ys[2823]), .RECT2_WIDTH(rectangle2_widths[2823]), .RECT2_HEIGHT(rectangle2_heights[2823]), .RECT2_WEIGHT(rectangle2_weights[2823]), .RECT3_X(rectangle3_xs[2823]), .RECT3_Y(rectangle3_ys[2823]), .RECT3_WIDTH(rectangle3_widths[2823]), .RECT3_HEIGHT(rectangle3_heights[2823]), .RECT3_WEIGHT(rectangle3_weights[2823]), .FEAT_THRES(feature_thresholds[2823]), .FEAT_ABOVE(feature_aboves[2823]), .FEAT_BELOW(feature_belows[2823])) ac2823(.scan_win(scan_win2823), .scan_win_std_dev(scan_win_std_dev[2823]), .feature_accum(feature_accums[2823]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2824]), .RECT1_Y(rectangle1_ys[2824]), .RECT1_WIDTH(rectangle1_widths[2824]), .RECT1_HEIGHT(rectangle1_heights[2824]), .RECT1_WEIGHT(rectangle1_weights[2824]), .RECT2_X(rectangle2_xs[2824]), .RECT2_Y(rectangle2_ys[2824]), .RECT2_WIDTH(rectangle2_widths[2824]), .RECT2_HEIGHT(rectangle2_heights[2824]), .RECT2_WEIGHT(rectangle2_weights[2824]), .RECT3_X(rectangle3_xs[2824]), .RECT3_Y(rectangle3_ys[2824]), .RECT3_WIDTH(rectangle3_widths[2824]), .RECT3_HEIGHT(rectangle3_heights[2824]), .RECT3_WEIGHT(rectangle3_weights[2824]), .FEAT_THRES(feature_thresholds[2824]), .FEAT_ABOVE(feature_aboves[2824]), .FEAT_BELOW(feature_belows[2824])) ac2824(.scan_win(scan_win2824), .scan_win_std_dev(scan_win_std_dev[2824]), .feature_accum(feature_accums[2824]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2825]), .RECT1_Y(rectangle1_ys[2825]), .RECT1_WIDTH(rectangle1_widths[2825]), .RECT1_HEIGHT(rectangle1_heights[2825]), .RECT1_WEIGHT(rectangle1_weights[2825]), .RECT2_X(rectangle2_xs[2825]), .RECT2_Y(rectangle2_ys[2825]), .RECT2_WIDTH(rectangle2_widths[2825]), .RECT2_HEIGHT(rectangle2_heights[2825]), .RECT2_WEIGHT(rectangle2_weights[2825]), .RECT3_X(rectangle3_xs[2825]), .RECT3_Y(rectangle3_ys[2825]), .RECT3_WIDTH(rectangle3_widths[2825]), .RECT3_HEIGHT(rectangle3_heights[2825]), .RECT3_WEIGHT(rectangle3_weights[2825]), .FEAT_THRES(feature_thresholds[2825]), .FEAT_ABOVE(feature_aboves[2825]), .FEAT_BELOW(feature_belows[2825])) ac2825(.scan_win(scan_win2825), .scan_win_std_dev(scan_win_std_dev[2825]), .feature_accum(feature_accums[2825]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2826]), .RECT1_Y(rectangle1_ys[2826]), .RECT1_WIDTH(rectangle1_widths[2826]), .RECT1_HEIGHT(rectangle1_heights[2826]), .RECT1_WEIGHT(rectangle1_weights[2826]), .RECT2_X(rectangle2_xs[2826]), .RECT2_Y(rectangle2_ys[2826]), .RECT2_WIDTH(rectangle2_widths[2826]), .RECT2_HEIGHT(rectangle2_heights[2826]), .RECT2_WEIGHT(rectangle2_weights[2826]), .RECT3_X(rectangle3_xs[2826]), .RECT3_Y(rectangle3_ys[2826]), .RECT3_WIDTH(rectangle3_widths[2826]), .RECT3_HEIGHT(rectangle3_heights[2826]), .RECT3_WEIGHT(rectangle3_weights[2826]), .FEAT_THRES(feature_thresholds[2826]), .FEAT_ABOVE(feature_aboves[2826]), .FEAT_BELOW(feature_belows[2826])) ac2826(.scan_win(scan_win2826), .scan_win_std_dev(scan_win_std_dev[2826]), .feature_accum(feature_accums[2826]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2827]), .RECT1_Y(rectangle1_ys[2827]), .RECT1_WIDTH(rectangle1_widths[2827]), .RECT1_HEIGHT(rectangle1_heights[2827]), .RECT1_WEIGHT(rectangle1_weights[2827]), .RECT2_X(rectangle2_xs[2827]), .RECT2_Y(rectangle2_ys[2827]), .RECT2_WIDTH(rectangle2_widths[2827]), .RECT2_HEIGHT(rectangle2_heights[2827]), .RECT2_WEIGHT(rectangle2_weights[2827]), .RECT3_X(rectangle3_xs[2827]), .RECT3_Y(rectangle3_ys[2827]), .RECT3_WIDTH(rectangle3_widths[2827]), .RECT3_HEIGHT(rectangle3_heights[2827]), .RECT3_WEIGHT(rectangle3_weights[2827]), .FEAT_THRES(feature_thresholds[2827]), .FEAT_ABOVE(feature_aboves[2827]), .FEAT_BELOW(feature_belows[2827])) ac2827(.scan_win(scan_win2827), .scan_win_std_dev(scan_win_std_dev[2827]), .feature_accum(feature_accums[2827]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2828]), .RECT1_Y(rectangle1_ys[2828]), .RECT1_WIDTH(rectangle1_widths[2828]), .RECT1_HEIGHT(rectangle1_heights[2828]), .RECT1_WEIGHT(rectangle1_weights[2828]), .RECT2_X(rectangle2_xs[2828]), .RECT2_Y(rectangle2_ys[2828]), .RECT2_WIDTH(rectangle2_widths[2828]), .RECT2_HEIGHT(rectangle2_heights[2828]), .RECT2_WEIGHT(rectangle2_weights[2828]), .RECT3_X(rectangle3_xs[2828]), .RECT3_Y(rectangle3_ys[2828]), .RECT3_WIDTH(rectangle3_widths[2828]), .RECT3_HEIGHT(rectangle3_heights[2828]), .RECT3_WEIGHT(rectangle3_weights[2828]), .FEAT_THRES(feature_thresholds[2828]), .FEAT_ABOVE(feature_aboves[2828]), .FEAT_BELOW(feature_belows[2828])) ac2828(.scan_win(scan_win2828), .scan_win_std_dev(scan_win_std_dev[2828]), .feature_accum(feature_accums[2828]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2829]), .RECT1_Y(rectangle1_ys[2829]), .RECT1_WIDTH(rectangle1_widths[2829]), .RECT1_HEIGHT(rectangle1_heights[2829]), .RECT1_WEIGHT(rectangle1_weights[2829]), .RECT2_X(rectangle2_xs[2829]), .RECT2_Y(rectangle2_ys[2829]), .RECT2_WIDTH(rectangle2_widths[2829]), .RECT2_HEIGHT(rectangle2_heights[2829]), .RECT2_WEIGHT(rectangle2_weights[2829]), .RECT3_X(rectangle3_xs[2829]), .RECT3_Y(rectangle3_ys[2829]), .RECT3_WIDTH(rectangle3_widths[2829]), .RECT3_HEIGHT(rectangle3_heights[2829]), .RECT3_WEIGHT(rectangle3_weights[2829]), .FEAT_THRES(feature_thresholds[2829]), .FEAT_ABOVE(feature_aboves[2829]), .FEAT_BELOW(feature_belows[2829])) ac2829(.scan_win(scan_win2829), .scan_win_std_dev(scan_win_std_dev[2829]), .feature_accum(feature_accums[2829]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2830]), .RECT1_Y(rectangle1_ys[2830]), .RECT1_WIDTH(rectangle1_widths[2830]), .RECT1_HEIGHT(rectangle1_heights[2830]), .RECT1_WEIGHT(rectangle1_weights[2830]), .RECT2_X(rectangle2_xs[2830]), .RECT2_Y(rectangle2_ys[2830]), .RECT2_WIDTH(rectangle2_widths[2830]), .RECT2_HEIGHT(rectangle2_heights[2830]), .RECT2_WEIGHT(rectangle2_weights[2830]), .RECT3_X(rectangle3_xs[2830]), .RECT3_Y(rectangle3_ys[2830]), .RECT3_WIDTH(rectangle3_widths[2830]), .RECT3_HEIGHT(rectangle3_heights[2830]), .RECT3_WEIGHT(rectangle3_weights[2830]), .FEAT_THRES(feature_thresholds[2830]), .FEAT_ABOVE(feature_aboves[2830]), .FEAT_BELOW(feature_belows[2830])) ac2830(.scan_win(scan_win2830), .scan_win_std_dev(scan_win_std_dev[2830]), .feature_accum(feature_accums[2830]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2831]), .RECT1_Y(rectangle1_ys[2831]), .RECT1_WIDTH(rectangle1_widths[2831]), .RECT1_HEIGHT(rectangle1_heights[2831]), .RECT1_WEIGHT(rectangle1_weights[2831]), .RECT2_X(rectangle2_xs[2831]), .RECT2_Y(rectangle2_ys[2831]), .RECT2_WIDTH(rectangle2_widths[2831]), .RECT2_HEIGHT(rectangle2_heights[2831]), .RECT2_WEIGHT(rectangle2_weights[2831]), .RECT3_X(rectangle3_xs[2831]), .RECT3_Y(rectangle3_ys[2831]), .RECT3_WIDTH(rectangle3_widths[2831]), .RECT3_HEIGHT(rectangle3_heights[2831]), .RECT3_WEIGHT(rectangle3_weights[2831]), .FEAT_THRES(feature_thresholds[2831]), .FEAT_ABOVE(feature_aboves[2831]), .FEAT_BELOW(feature_belows[2831])) ac2831(.scan_win(scan_win2831), .scan_win_std_dev(scan_win_std_dev[2831]), .feature_accum(feature_accums[2831]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2832]), .RECT1_Y(rectangle1_ys[2832]), .RECT1_WIDTH(rectangle1_widths[2832]), .RECT1_HEIGHT(rectangle1_heights[2832]), .RECT1_WEIGHT(rectangle1_weights[2832]), .RECT2_X(rectangle2_xs[2832]), .RECT2_Y(rectangle2_ys[2832]), .RECT2_WIDTH(rectangle2_widths[2832]), .RECT2_HEIGHT(rectangle2_heights[2832]), .RECT2_WEIGHT(rectangle2_weights[2832]), .RECT3_X(rectangle3_xs[2832]), .RECT3_Y(rectangle3_ys[2832]), .RECT3_WIDTH(rectangle3_widths[2832]), .RECT3_HEIGHT(rectangle3_heights[2832]), .RECT3_WEIGHT(rectangle3_weights[2832]), .FEAT_THRES(feature_thresholds[2832]), .FEAT_ABOVE(feature_aboves[2832]), .FEAT_BELOW(feature_belows[2832])) ac2832(.scan_win(scan_win2832), .scan_win_std_dev(scan_win_std_dev[2832]), .feature_accum(feature_accums[2832]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2833]), .RECT1_Y(rectangle1_ys[2833]), .RECT1_WIDTH(rectangle1_widths[2833]), .RECT1_HEIGHT(rectangle1_heights[2833]), .RECT1_WEIGHT(rectangle1_weights[2833]), .RECT2_X(rectangle2_xs[2833]), .RECT2_Y(rectangle2_ys[2833]), .RECT2_WIDTH(rectangle2_widths[2833]), .RECT2_HEIGHT(rectangle2_heights[2833]), .RECT2_WEIGHT(rectangle2_weights[2833]), .RECT3_X(rectangle3_xs[2833]), .RECT3_Y(rectangle3_ys[2833]), .RECT3_WIDTH(rectangle3_widths[2833]), .RECT3_HEIGHT(rectangle3_heights[2833]), .RECT3_WEIGHT(rectangle3_weights[2833]), .FEAT_THRES(feature_thresholds[2833]), .FEAT_ABOVE(feature_aboves[2833]), .FEAT_BELOW(feature_belows[2833])) ac2833(.scan_win(scan_win2833), .scan_win_std_dev(scan_win_std_dev[2833]), .feature_accum(feature_accums[2833]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2834]), .RECT1_Y(rectangle1_ys[2834]), .RECT1_WIDTH(rectangle1_widths[2834]), .RECT1_HEIGHT(rectangle1_heights[2834]), .RECT1_WEIGHT(rectangle1_weights[2834]), .RECT2_X(rectangle2_xs[2834]), .RECT2_Y(rectangle2_ys[2834]), .RECT2_WIDTH(rectangle2_widths[2834]), .RECT2_HEIGHT(rectangle2_heights[2834]), .RECT2_WEIGHT(rectangle2_weights[2834]), .RECT3_X(rectangle3_xs[2834]), .RECT3_Y(rectangle3_ys[2834]), .RECT3_WIDTH(rectangle3_widths[2834]), .RECT3_HEIGHT(rectangle3_heights[2834]), .RECT3_WEIGHT(rectangle3_weights[2834]), .FEAT_THRES(feature_thresholds[2834]), .FEAT_ABOVE(feature_aboves[2834]), .FEAT_BELOW(feature_belows[2834])) ac2834(.scan_win(scan_win2834), .scan_win_std_dev(scan_win_std_dev[2834]), .feature_accum(feature_accums[2834]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2835]), .RECT1_Y(rectangle1_ys[2835]), .RECT1_WIDTH(rectangle1_widths[2835]), .RECT1_HEIGHT(rectangle1_heights[2835]), .RECT1_WEIGHT(rectangle1_weights[2835]), .RECT2_X(rectangle2_xs[2835]), .RECT2_Y(rectangle2_ys[2835]), .RECT2_WIDTH(rectangle2_widths[2835]), .RECT2_HEIGHT(rectangle2_heights[2835]), .RECT2_WEIGHT(rectangle2_weights[2835]), .RECT3_X(rectangle3_xs[2835]), .RECT3_Y(rectangle3_ys[2835]), .RECT3_WIDTH(rectangle3_widths[2835]), .RECT3_HEIGHT(rectangle3_heights[2835]), .RECT3_WEIGHT(rectangle3_weights[2835]), .FEAT_THRES(feature_thresholds[2835]), .FEAT_ABOVE(feature_aboves[2835]), .FEAT_BELOW(feature_belows[2835])) ac2835(.scan_win(scan_win2835), .scan_win_std_dev(scan_win_std_dev[2835]), .feature_accum(feature_accums[2835]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2836]), .RECT1_Y(rectangle1_ys[2836]), .RECT1_WIDTH(rectangle1_widths[2836]), .RECT1_HEIGHT(rectangle1_heights[2836]), .RECT1_WEIGHT(rectangle1_weights[2836]), .RECT2_X(rectangle2_xs[2836]), .RECT2_Y(rectangle2_ys[2836]), .RECT2_WIDTH(rectangle2_widths[2836]), .RECT2_HEIGHT(rectangle2_heights[2836]), .RECT2_WEIGHT(rectangle2_weights[2836]), .RECT3_X(rectangle3_xs[2836]), .RECT3_Y(rectangle3_ys[2836]), .RECT3_WIDTH(rectangle3_widths[2836]), .RECT3_HEIGHT(rectangle3_heights[2836]), .RECT3_WEIGHT(rectangle3_weights[2836]), .FEAT_THRES(feature_thresholds[2836]), .FEAT_ABOVE(feature_aboves[2836]), .FEAT_BELOW(feature_belows[2836])) ac2836(.scan_win(scan_win2836), .scan_win_std_dev(scan_win_std_dev[2836]), .feature_accum(feature_accums[2836]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2837]), .RECT1_Y(rectangle1_ys[2837]), .RECT1_WIDTH(rectangle1_widths[2837]), .RECT1_HEIGHT(rectangle1_heights[2837]), .RECT1_WEIGHT(rectangle1_weights[2837]), .RECT2_X(rectangle2_xs[2837]), .RECT2_Y(rectangle2_ys[2837]), .RECT2_WIDTH(rectangle2_widths[2837]), .RECT2_HEIGHT(rectangle2_heights[2837]), .RECT2_WEIGHT(rectangle2_weights[2837]), .RECT3_X(rectangle3_xs[2837]), .RECT3_Y(rectangle3_ys[2837]), .RECT3_WIDTH(rectangle3_widths[2837]), .RECT3_HEIGHT(rectangle3_heights[2837]), .RECT3_WEIGHT(rectangle3_weights[2837]), .FEAT_THRES(feature_thresholds[2837]), .FEAT_ABOVE(feature_aboves[2837]), .FEAT_BELOW(feature_belows[2837])) ac2837(.scan_win(scan_win2837), .scan_win_std_dev(scan_win_std_dev[2837]), .feature_accum(feature_accums[2837]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2838]), .RECT1_Y(rectangle1_ys[2838]), .RECT1_WIDTH(rectangle1_widths[2838]), .RECT1_HEIGHT(rectangle1_heights[2838]), .RECT1_WEIGHT(rectangle1_weights[2838]), .RECT2_X(rectangle2_xs[2838]), .RECT2_Y(rectangle2_ys[2838]), .RECT2_WIDTH(rectangle2_widths[2838]), .RECT2_HEIGHT(rectangle2_heights[2838]), .RECT2_WEIGHT(rectangle2_weights[2838]), .RECT3_X(rectangle3_xs[2838]), .RECT3_Y(rectangle3_ys[2838]), .RECT3_WIDTH(rectangle3_widths[2838]), .RECT3_HEIGHT(rectangle3_heights[2838]), .RECT3_WEIGHT(rectangle3_weights[2838]), .FEAT_THRES(feature_thresholds[2838]), .FEAT_ABOVE(feature_aboves[2838]), .FEAT_BELOW(feature_belows[2838])) ac2838(.scan_win(scan_win2838), .scan_win_std_dev(scan_win_std_dev[2838]), .feature_accum(feature_accums[2838]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2839]), .RECT1_Y(rectangle1_ys[2839]), .RECT1_WIDTH(rectangle1_widths[2839]), .RECT1_HEIGHT(rectangle1_heights[2839]), .RECT1_WEIGHT(rectangle1_weights[2839]), .RECT2_X(rectangle2_xs[2839]), .RECT2_Y(rectangle2_ys[2839]), .RECT2_WIDTH(rectangle2_widths[2839]), .RECT2_HEIGHT(rectangle2_heights[2839]), .RECT2_WEIGHT(rectangle2_weights[2839]), .RECT3_X(rectangle3_xs[2839]), .RECT3_Y(rectangle3_ys[2839]), .RECT3_WIDTH(rectangle3_widths[2839]), .RECT3_HEIGHT(rectangle3_heights[2839]), .RECT3_WEIGHT(rectangle3_weights[2839]), .FEAT_THRES(feature_thresholds[2839]), .FEAT_ABOVE(feature_aboves[2839]), .FEAT_BELOW(feature_belows[2839])) ac2839(.scan_win(scan_win2839), .scan_win_std_dev(scan_win_std_dev[2839]), .feature_accum(feature_accums[2839]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2840]), .RECT1_Y(rectangle1_ys[2840]), .RECT1_WIDTH(rectangle1_widths[2840]), .RECT1_HEIGHT(rectangle1_heights[2840]), .RECT1_WEIGHT(rectangle1_weights[2840]), .RECT2_X(rectangle2_xs[2840]), .RECT2_Y(rectangle2_ys[2840]), .RECT2_WIDTH(rectangle2_widths[2840]), .RECT2_HEIGHT(rectangle2_heights[2840]), .RECT2_WEIGHT(rectangle2_weights[2840]), .RECT3_X(rectangle3_xs[2840]), .RECT3_Y(rectangle3_ys[2840]), .RECT3_WIDTH(rectangle3_widths[2840]), .RECT3_HEIGHT(rectangle3_heights[2840]), .RECT3_WEIGHT(rectangle3_weights[2840]), .FEAT_THRES(feature_thresholds[2840]), .FEAT_ABOVE(feature_aboves[2840]), .FEAT_BELOW(feature_belows[2840])) ac2840(.scan_win(scan_win2840), .scan_win_std_dev(scan_win_std_dev[2840]), .feature_accum(feature_accums[2840]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2841]), .RECT1_Y(rectangle1_ys[2841]), .RECT1_WIDTH(rectangle1_widths[2841]), .RECT1_HEIGHT(rectangle1_heights[2841]), .RECT1_WEIGHT(rectangle1_weights[2841]), .RECT2_X(rectangle2_xs[2841]), .RECT2_Y(rectangle2_ys[2841]), .RECT2_WIDTH(rectangle2_widths[2841]), .RECT2_HEIGHT(rectangle2_heights[2841]), .RECT2_WEIGHT(rectangle2_weights[2841]), .RECT3_X(rectangle3_xs[2841]), .RECT3_Y(rectangle3_ys[2841]), .RECT3_WIDTH(rectangle3_widths[2841]), .RECT3_HEIGHT(rectangle3_heights[2841]), .RECT3_WEIGHT(rectangle3_weights[2841]), .FEAT_THRES(feature_thresholds[2841]), .FEAT_ABOVE(feature_aboves[2841]), .FEAT_BELOW(feature_belows[2841])) ac2841(.scan_win(scan_win2841), .scan_win_std_dev(scan_win_std_dev[2841]), .feature_accum(feature_accums[2841]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2842]), .RECT1_Y(rectangle1_ys[2842]), .RECT1_WIDTH(rectangle1_widths[2842]), .RECT1_HEIGHT(rectangle1_heights[2842]), .RECT1_WEIGHT(rectangle1_weights[2842]), .RECT2_X(rectangle2_xs[2842]), .RECT2_Y(rectangle2_ys[2842]), .RECT2_WIDTH(rectangle2_widths[2842]), .RECT2_HEIGHT(rectangle2_heights[2842]), .RECT2_WEIGHT(rectangle2_weights[2842]), .RECT3_X(rectangle3_xs[2842]), .RECT3_Y(rectangle3_ys[2842]), .RECT3_WIDTH(rectangle3_widths[2842]), .RECT3_HEIGHT(rectangle3_heights[2842]), .RECT3_WEIGHT(rectangle3_weights[2842]), .FEAT_THRES(feature_thresholds[2842]), .FEAT_ABOVE(feature_aboves[2842]), .FEAT_BELOW(feature_belows[2842])) ac2842(.scan_win(scan_win2842), .scan_win_std_dev(scan_win_std_dev[2842]), .feature_accum(feature_accums[2842]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2843]), .RECT1_Y(rectangle1_ys[2843]), .RECT1_WIDTH(rectangle1_widths[2843]), .RECT1_HEIGHT(rectangle1_heights[2843]), .RECT1_WEIGHT(rectangle1_weights[2843]), .RECT2_X(rectangle2_xs[2843]), .RECT2_Y(rectangle2_ys[2843]), .RECT2_WIDTH(rectangle2_widths[2843]), .RECT2_HEIGHT(rectangle2_heights[2843]), .RECT2_WEIGHT(rectangle2_weights[2843]), .RECT3_X(rectangle3_xs[2843]), .RECT3_Y(rectangle3_ys[2843]), .RECT3_WIDTH(rectangle3_widths[2843]), .RECT3_HEIGHT(rectangle3_heights[2843]), .RECT3_WEIGHT(rectangle3_weights[2843]), .FEAT_THRES(feature_thresholds[2843]), .FEAT_ABOVE(feature_aboves[2843]), .FEAT_BELOW(feature_belows[2843])) ac2843(.scan_win(scan_win2843), .scan_win_std_dev(scan_win_std_dev[2843]), .feature_accum(feature_accums[2843]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2844]), .RECT1_Y(rectangle1_ys[2844]), .RECT1_WIDTH(rectangle1_widths[2844]), .RECT1_HEIGHT(rectangle1_heights[2844]), .RECT1_WEIGHT(rectangle1_weights[2844]), .RECT2_X(rectangle2_xs[2844]), .RECT2_Y(rectangle2_ys[2844]), .RECT2_WIDTH(rectangle2_widths[2844]), .RECT2_HEIGHT(rectangle2_heights[2844]), .RECT2_WEIGHT(rectangle2_weights[2844]), .RECT3_X(rectangle3_xs[2844]), .RECT3_Y(rectangle3_ys[2844]), .RECT3_WIDTH(rectangle3_widths[2844]), .RECT3_HEIGHT(rectangle3_heights[2844]), .RECT3_WEIGHT(rectangle3_weights[2844]), .FEAT_THRES(feature_thresholds[2844]), .FEAT_ABOVE(feature_aboves[2844]), .FEAT_BELOW(feature_belows[2844])) ac2844(.scan_win(scan_win2844), .scan_win_std_dev(scan_win_std_dev[2844]), .feature_accum(feature_accums[2844]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2845]), .RECT1_Y(rectangle1_ys[2845]), .RECT1_WIDTH(rectangle1_widths[2845]), .RECT1_HEIGHT(rectangle1_heights[2845]), .RECT1_WEIGHT(rectangle1_weights[2845]), .RECT2_X(rectangle2_xs[2845]), .RECT2_Y(rectangle2_ys[2845]), .RECT2_WIDTH(rectangle2_widths[2845]), .RECT2_HEIGHT(rectangle2_heights[2845]), .RECT2_WEIGHT(rectangle2_weights[2845]), .RECT3_X(rectangle3_xs[2845]), .RECT3_Y(rectangle3_ys[2845]), .RECT3_WIDTH(rectangle3_widths[2845]), .RECT3_HEIGHT(rectangle3_heights[2845]), .RECT3_WEIGHT(rectangle3_weights[2845]), .FEAT_THRES(feature_thresholds[2845]), .FEAT_ABOVE(feature_aboves[2845]), .FEAT_BELOW(feature_belows[2845])) ac2845(.scan_win(scan_win2845), .scan_win_std_dev(scan_win_std_dev[2845]), .feature_accum(feature_accums[2845]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2846]), .RECT1_Y(rectangle1_ys[2846]), .RECT1_WIDTH(rectangle1_widths[2846]), .RECT1_HEIGHT(rectangle1_heights[2846]), .RECT1_WEIGHT(rectangle1_weights[2846]), .RECT2_X(rectangle2_xs[2846]), .RECT2_Y(rectangle2_ys[2846]), .RECT2_WIDTH(rectangle2_widths[2846]), .RECT2_HEIGHT(rectangle2_heights[2846]), .RECT2_WEIGHT(rectangle2_weights[2846]), .RECT3_X(rectangle3_xs[2846]), .RECT3_Y(rectangle3_ys[2846]), .RECT3_WIDTH(rectangle3_widths[2846]), .RECT3_HEIGHT(rectangle3_heights[2846]), .RECT3_WEIGHT(rectangle3_weights[2846]), .FEAT_THRES(feature_thresholds[2846]), .FEAT_ABOVE(feature_aboves[2846]), .FEAT_BELOW(feature_belows[2846])) ac2846(.scan_win(scan_win2846), .scan_win_std_dev(scan_win_std_dev[2846]), .feature_accum(feature_accums[2846]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2847]), .RECT1_Y(rectangle1_ys[2847]), .RECT1_WIDTH(rectangle1_widths[2847]), .RECT1_HEIGHT(rectangle1_heights[2847]), .RECT1_WEIGHT(rectangle1_weights[2847]), .RECT2_X(rectangle2_xs[2847]), .RECT2_Y(rectangle2_ys[2847]), .RECT2_WIDTH(rectangle2_widths[2847]), .RECT2_HEIGHT(rectangle2_heights[2847]), .RECT2_WEIGHT(rectangle2_weights[2847]), .RECT3_X(rectangle3_xs[2847]), .RECT3_Y(rectangle3_ys[2847]), .RECT3_WIDTH(rectangle3_widths[2847]), .RECT3_HEIGHT(rectangle3_heights[2847]), .RECT3_WEIGHT(rectangle3_weights[2847]), .FEAT_THRES(feature_thresholds[2847]), .FEAT_ABOVE(feature_aboves[2847]), .FEAT_BELOW(feature_belows[2847])) ac2847(.scan_win(scan_win2847), .scan_win_std_dev(scan_win_std_dev[2847]), .feature_accum(feature_accums[2847]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2848]), .RECT1_Y(rectangle1_ys[2848]), .RECT1_WIDTH(rectangle1_widths[2848]), .RECT1_HEIGHT(rectangle1_heights[2848]), .RECT1_WEIGHT(rectangle1_weights[2848]), .RECT2_X(rectangle2_xs[2848]), .RECT2_Y(rectangle2_ys[2848]), .RECT2_WIDTH(rectangle2_widths[2848]), .RECT2_HEIGHT(rectangle2_heights[2848]), .RECT2_WEIGHT(rectangle2_weights[2848]), .RECT3_X(rectangle3_xs[2848]), .RECT3_Y(rectangle3_ys[2848]), .RECT3_WIDTH(rectangle3_widths[2848]), .RECT3_HEIGHT(rectangle3_heights[2848]), .RECT3_WEIGHT(rectangle3_weights[2848]), .FEAT_THRES(feature_thresholds[2848]), .FEAT_ABOVE(feature_aboves[2848]), .FEAT_BELOW(feature_belows[2848])) ac2848(.scan_win(scan_win2848), .scan_win_std_dev(scan_win_std_dev[2848]), .feature_accum(feature_accums[2848]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2849]), .RECT1_Y(rectangle1_ys[2849]), .RECT1_WIDTH(rectangle1_widths[2849]), .RECT1_HEIGHT(rectangle1_heights[2849]), .RECT1_WEIGHT(rectangle1_weights[2849]), .RECT2_X(rectangle2_xs[2849]), .RECT2_Y(rectangle2_ys[2849]), .RECT2_WIDTH(rectangle2_widths[2849]), .RECT2_HEIGHT(rectangle2_heights[2849]), .RECT2_WEIGHT(rectangle2_weights[2849]), .RECT3_X(rectangle3_xs[2849]), .RECT3_Y(rectangle3_ys[2849]), .RECT3_WIDTH(rectangle3_widths[2849]), .RECT3_HEIGHT(rectangle3_heights[2849]), .RECT3_WEIGHT(rectangle3_weights[2849]), .FEAT_THRES(feature_thresholds[2849]), .FEAT_ABOVE(feature_aboves[2849]), .FEAT_BELOW(feature_belows[2849])) ac2849(.scan_win(scan_win2849), .scan_win_std_dev(scan_win_std_dev[2849]), .feature_accum(feature_accums[2849]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2850]), .RECT1_Y(rectangle1_ys[2850]), .RECT1_WIDTH(rectangle1_widths[2850]), .RECT1_HEIGHT(rectangle1_heights[2850]), .RECT1_WEIGHT(rectangle1_weights[2850]), .RECT2_X(rectangle2_xs[2850]), .RECT2_Y(rectangle2_ys[2850]), .RECT2_WIDTH(rectangle2_widths[2850]), .RECT2_HEIGHT(rectangle2_heights[2850]), .RECT2_WEIGHT(rectangle2_weights[2850]), .RECT3_X(rectangle3_xs[2850]), .RECT3_Y(rectangle3_ys[2850]), .RECT3_WIDTH(rectangle3_widths[2850]), .RECT3_HEIGHT(rectangle3_heights[2850]), .RECT3_WEIGHT(rectangle3_weights[2850]), .FEAT_THRES(feature_thresholds[2850]), .FEAT_ABOVE(feature_aboves[2850]), .FEAT_BELOW(feature_belows[2850])) ac2850(.scan_win(scan_win2850), .scan_win_std_dev(scan_win_std_dev[2850]), .feature_accum(feature_accums[2850]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2851]), .RECT1_Y(rectangle1_ys[2851]), .RECT1_WIDTH(rectangle1_widths[2851]), .RECT1_HEIGHT(rectangle1_heights[2851]), .RECT1_WEIGHT(rectangle1_weights[2851]), .RECT2_X(rectangle2_xs[2851]), .RECT2_Y(rectangle2_ys[2851]), .RECT2_WIDTH(rectangle2_widths[2851]), .RECT2_HEIGHT(rectangle2_heights[2851]), .RECT2_WEIGHT(rectangle2_weights[2851]), .RECT3_X(rectangle3_xs[2851]), .RECT3_Y(rectangle3_ys[2851]), .RECT3_WIDTH(rectangle3_widths[2851]), .RECT3_HEIGHT(rectangle3_heights[2851]), .RECT3_WEIGHT(rectangle3_weights[2851]), .FEAT_THRES(feature_thresholds[2851]), .FEAT_ABOVE(feature_aboves[2851]), .FEAT_BELOW(feature_belows[2851])) ac2851(.scan_win(scan_win2851), .scan_win_std_dev(scan_win_std_dev[2851]), .feature_accum(feature_accums[2851]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2852]), .RECT1_Y(rectangle1_ys[2852]), .RECT1_WIDTH(rectangle1_widths[2852]), .RECT1_HEIGHT(rectangle1_heights[2852]), .RECT1_WEIGHT(rectangle1_weights[2852]), .RECT2_X(rectangle2_xs[2852]), .RECT2_Y(rectangle2_ys[2852]), .RECT2_WIDTH(rectangle2_widths[2852]), .RECT2_HEIGHT(rectangle2_heights[2852]), .RECT2_WEIGHT(rectangle2_weights[2852]), .RECT3_X(rectangle3_xs[2852]), .RECT3_Y(rectangle3_ys[2852]), .RECT3_WIDTH(rectangle3_widths[2852]), .RECT3_HEIGHT(rectangle3_heights[2852]), .RECT3_WEIGHT(rectangle3_weights[2852]), .FEAT_THRES(feature_thresholds[2852]), .FEAT_ABOVE(feature_aboves[2852]), .FEAT_BELOW(feature_belows[2852])) ac2852(.scan_win(scan_win2852), .scan_win_std_dev(scan_win_std_dev[2852]), .feature_accum(feature_accums[2852]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2853]), .RECT1_Y(rectangle1_ys[2853]), .RECT1_WIDTH(rectangle1_widths[2853]), .RECT1_HEIGHT(rectangle1_heights[2853]), .RECT1_WEIGHT(rectangle1_weights[2853]), .RECT2_X(rectangle2_xs[2853]), .RECT2_Y(rectangle2_ys[2853]), .RECT2_WIDTH(rectangle2_widths[2853]), .RECT2_HEIGHT(rectangle2_heights[2853]), .RECT2_WEIGHT(rectangle2_weights[2853]), .RECT3_X(rectangle3_xs[2853]), .RECT3_Y(rectangle3_ys[2853]), .RECT3_WIDTH(rectangle3_widths[2853]), .RECT3_HEIGHT(rectangle3_heights[2853]), .RECT3_WEIGHT(rectangle3_weights[2853]), .FEAT_THRES(feature_thresholds[2853]), .FEAT_ABOVE(feature_aboves[2853]), .FEAT_BELOW(feature_belows[2853])) ac2853(.scan_win(scan_win2853), .scan_win_std_dev(scan_win_std_dev[2853]), .feature_accum(feature_accums[2853]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2854]), .RECT1_Y(rectangle1_ys[2854]), .RECT1_WIDTH(rectangle1_widths[2854]), .RECT1_HEIGHT(rectangle1_heights[2854]), .RECT1_WEIGHT(rectangle1_weights[2854]), .RECT2_X(rectangle2_xs[2854]), .RECT2_Y(rectangle2_ys[2854]), .RECT2_WIDTH(rectangle2_widths[2854]), .RECT2_HEIGHT(rectangle2_heights[2854]), .RECT2_WEIGHT(rectangle2_weights[2854]), .RECT3_X(rectangle3_xs[2854]), .RECT3_Y(rectangle3_ys[2854]), .RECT3_WIDTH(rectangle3_widths[2854]), .RECT3_HEIGHT(rectangle3_heights[2854]), .RECT3_WEIGHT(rectangle3_weights[2854]), .FEAT_THRES(feature_thresholds[2854]), .FEAT_ABOVE(feature_aboves[2854]), .FEAT_BELOW(feature_belows[2854])) ac2854(.scan_win(scan_win2854), .scan_win_std_dev(scan_win_std_dev[2854]), .feature_accum(feature_accums[2854]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2855]), .RECT1_Y(rectangle1_ys[2855]), .RECT1_WIDTH(rectangle1_widths[2855]), .RECT1_HEIGHT(rectangle1_heights[2855]), .RECT1_WEIGHT(rectangle1_weights[2855]), .RECT2_X(rectangle2_xs[2855]), .RECT2_Y(rectangle2_ys[2855]), .RECT2_WIDTH(rectangle2_widths[2855]), .RECT2_HEIGHT(rectangle2_heights[2855]), .RECT2_WEIGHT(rectangle2_weights[2855]), .RECT3_X(rectangle3_xs[2855]), .RECT3_Y(rectangle3_ys[2855]), .RECT3_WIDTH(rectangle3_widths[2855]), .RECT3_HEIGHT(rectangle3_heights[2855]), .RECT3_WEIGHT(rectangle3_weights[2855]), .FEAT_THRES(feature_thresholds[2855]), .FEAT_ABOVE(feature_aboves[2855]), .FEAT_BELOW(feature_belows[2855])) ac2855(.scan_win(scan_win2855), .scan_win_std_dev(scan_win_std_dev[2855]), .feature_accum(feature_accums[2855]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2856]), .RECT1_Y(rectangle1_ys[2856]), .RECT1_WIDTH(rectangle1_widths[2856]), .RECT1_HEIGHT(rectangle1_heights[2856]), .RECT1_WEIGHT(rectangle1_weights[2856]), .RECT2_X(rectangle2_xs[2856]), .RECT2_Y(rectangle2_ys[2856]), .RECT2_WIDTH(rectangle2_widths[2856]), .RECT2_HEIGHT(rectangle2_heights[2856]), .RECT2_WEIGHT(rectangle2_weights[2856]), .RECT3_X(rectangle3_xs[2856]), .RECT3_Y(rectangle3_ys[2856]), .RECT3_WIDTH(rectangle3_widths[2856]), .RECT3_HEIGHT(rectangle3_heights[2856]), .RECT3_WEIGHT(rectangle3_weights[2856]), .FEAT_THRES(feature_thresholds[2856]), .FEAT_ABOVE(feature_aboves[2856]), .FEAT_BELOW(feature_belows[2856])) ac2856(.scan_win(scan_win2856), .scan_win_std_dev(scan_win_std_dev[2856]), .feature_accum(feature_accums[2856]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2857]), .RECT1_Y(rectangle1_ys[2857]), .RECT1_WIDTH(rectangle1_widths[2857]), .RECT1_HEIGHT(rectangle1_heights[2857]), .RECT1_WEIGHT(rectangle1_weights[2857]), .RECT2_X(rectangle2_xs[2857]), .RECT2_Y(rectangle2_ys[2857]), .RECT2_WIDTH(rectangle2_widths[2857]), .RECT2_HEIGHT(rectangle2_heights[2857]), .RECT2_WEIGHT(rectangle2_weights[2857]), .RECT3_X(rectangle3_xs[2857]), .RECT3_Y(rectangle3_ys[2857]), .RECT3_WIDTH(rectangle3_widths[2857]), .RECT3_HEIGHT(rectangle3_heights[2857]), .RECT3_WEIGHT(rectangle3_weights[2857]), .FEAT_THRES(feature_thresholds[2857]), .FEAT_ABOVE(feature_aboves[2857]), .FEAT_BELOW(feature_belows[2857])) ac2857(.scan_win(scan_win2857), .scan_win_std_dev(scan_win_std_dev[2857]), .feature_accum(feature_accums[2857]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2858]), .RECT1_Y(rectangle1_ys[2858]), .RECT1_WIDTH(rectangle1_widths[2858]), .RECT1_HEIGHT(rectangle1_heights[2858]), .RECT1_WEIGHT(rectangle1_weights[2858]), .RECT2_X(rectangle2_xs[2858]), .RECT2_Y(rectangle2_ys[2858]), .RECT2_WIDTH(rectangle2_widths[2858]), .RECT2_HEIGHT(rectangle2_heights[2858]), .RECT2_WEIGHT(rectangle2_weights[2858]), .RECT3_X(rectangle3_xs[2858]), .RECT3_Y(rectangle3_ys[2858]), .RECT3_WIDTH(rectangle3_widths[2858]), .RECT3_HEIGHT(rectangle3_heights[2858]), .RECT3_WEIGHT(rectangle3_weights[2858]), .FEAT_THRES(feature_thresholds[2858]), .FEAT_ABOVE(feature_aboves[2858]), .FEAT_BELOW(feature_belows[2858])) ac2858(.scan_win(scan_win2858), .scan_win_std_dev(scan_win_std_dev[2858]), .feature_accum(feature_accums[2858]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2859]), .RECT1_Y(rectangle1_ys[2859]), .RECT1_WIDTH(rectangle1_widths[2859]), .RECT1_HEIGHT(rectangle1_heights[2859]), .RECT1_WEIGHT(rectangle1_weights[2859]), .RECT2_X(rectangle2_xs[2859]), .RECT2_Y(rectangle2_ys[2859]), .RECT2_WIDTH(rectangle2_widths[2859]), .RECT2_HEIGHT(rectangle2_heights[2859]), .RECT2_WEIGHT(rectangle2_weights[2859]), .RECT3_X(rectangle3_xs[2859]), .RECT3_Y(rectangle3_ys[2859]), .RECT3_WIDTH(rectangle3_widths[2859]), .RECT3_HEIGHT(rectangle3_heights[2859]), .RECT3_WEIGHT(rectangle3_weights[2859]), .FEAT_THRES(feature_thresholds[2859]), .FEAT_ABOVE(feature_aboves[2859]), .FEAT_BELOW(feature_belows[2859])) ac2859(.scan_win(scan_win2859), .scan_win_std_dev(scan_win_std_dev[2859]), .feature_accum(feature_accums[2859]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2860]), .RECT1_Y(rectangle1_ys[2860]), .RECT1_WIDTH(rectangle1_widths[2860]), .RECT1_HEIGHT(rectangle1_heights[2860]), .RECT1_WEIGHT(rectangle1_weights[2860]), .RECT2_X(rectangle2_xs[2860]), .RECT2_Y(rectangle2_ys[2860]), .RECT2_WIDTH(rectangle2_widths[2860]), .RECT2_HEIGHT(rectangle2_heights[2860]), .RECT2_WEIGHT(rectangle2_weights[2860]), .RECT3_X(rectangle3_xs[2860]), .RECT3_Y(rectangle3_ys[2860]), .RECT3_WIDTH(rectangle3_widths[2860]), .RECT3_HEIGHT(rectangle3_heights[2860]), .RECT3_WEIGHT(rectangle3_weights[2860]), .FEAT_THRES(feature_thresholds[2860]), .FEAT_ABOVE(feature_aboves[2860]), .FEAT_BELOW(feature_belows[2860])) ac2860(.scan_win(scan_win2860), .scan_win_std_dev(scan_win_std_dev[2860]), .feature_accum(feature_accums[2860]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2861]), .RECT1_Y(rectangle1_ys[2861]), .RECT1_WIDTH(rectangle1_widths[2861]), .RECT1_HEIGHT(rectangle1_heights[2861]), .RECT1_WEIGHT(rectangle1_weights[2861]), .RECT2_X(rectangle2_xs[2861]), .RECT2_Y(rectangle2_ys[2861]), .RECT2_WIDTH(rectangle2_widths[2861]), .RECT2_HEIGHT(rectangle2_heights[2861]), .RECT2_WEIGHT(rectangle2_weights[2861]), .RECT3_X(rectangle3_xs[2861]), .RECT3_Y(rectangle3_ys[2861]), .RECT3_WIDTH(rectangle3_widths[2861]), .RECT3_HEIGHT(rectangle3_heights[2861]), .RECT3_WEIGHT(rectangle3_weights[2861]), .FEAT_THRES(feature_thresholds[2861]), .FEAT_ABOVE(feature_aboves[2861]), .FEAT_BELOW(feature_belows[2861])) ac2861(.scan_win(scan_win2861), .scan_win_std_dev(scan_win_std_dev[2861]), .feature_accum(feature_accums[2861]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2862]), .RECT1_Y(rectangle1_ys[2862]), .RECT1_WIDTH(rectangle1_widths[2862]), .RECT1_HEIGHT(rectangle1_heights[2862]), .RECT1_WEIGHT(rectangle1_weights[2862]), .RECT2_X(rectangle2_xs[2862]), .RECT2_Y(rectangle2_ys[2862]), .RECT2_WIDTH(rectangle2_widths[2862]), .RECT2_HEIGHT(rectangle2_heights[2862]), .RECT2_WEIGHT(rectangle2_weights[2862]), .RECT3_X(rectangle3_xs[2862]), .RECT3_Y(rectangle3_ys[2862]), .RECT3_WIDTH(rectangle3_widths[2862]), .RECT3_HEIGHT(rectangle3_heights[2862]), .RECT3_WEIGHT(rectangle3_weights[2862]), .FEAT_THRES(feature_thresholds[2862]), .FEAT_ABOVE(feature_aboves[2862]), .FEAT_BELOW(feature_belows[2862])) ac2862(.scan_win(scan_win2862), .scan_win_std_dev(scan_win_std_dev[2862]), .feature_accum(feature_accums[2862]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2863]), .RECT1_Y(rectangle1_ys[2863]), .RECT1_WIDTH(rectangle1_widths[2863]), .RECT1_HEIGHT(rectangle1_heights[2863]), .RECT1_WEIGHT(rectangle1_weights[2863]), .RECT2_X(rectangle2_xs[2863]), .RECT2_Y(rectangle2_ys[2863]), .RECT2_WIDTH(rectangle2_widths[2863]), .RECT2_HEIGHT(rectangle2_heights[2863]), .RECT2_WEIGHT(rectangle2_weights[2863]), .RECT3_X(rectangle3_xs[2863]), .RECT3_Y(rectangle3_ys[2863]), .RECT3_WIDTH(rectangle3_widths[2863]), .RECT3_HEIGHT(rectangle3_heights[2863]), .RECT3_WEIGHT(rectangle3_weights[2863]), .FEAT_THRES(feature_thresholds[2863]), .FEAT_ABOVE(feature_aboves[2863]), .FEAT_BELOW(feature_belows[2863])) ac2863(.scan_win(scan_win2863), .scan_win_std_dev(scan_win_std_dev[2863]), .feature_accum(feature_accums[2863]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2864]), .RECT1_Y(rectangle1_ys[2864]), .RECT1_WIDTH(rectangle1_widths[2864]), .RECT1_HEIGHT(rectangle1_heights[2864]), .RECT1_WEIGHT(rectangle1_weights[2864]), .RECT2_X(rectangle2_xs[2864]), .RECT2_Y(rectangle2_ys[2864]), .RECT2_WIDTH(rectangle2_widths[2864]), .RECT2_HEIGHT(rectangle2_heights[2864]), .RECT2_WEIGHT(rectangle2_weights[2864]), .RECT3_X(rectangle3_xs[2864]), .RECT3_Y(rectangle3_ys[2864]), .RECT3_WIDTH(rectangle3_widths[2864]), .RECT3_HEIGHT(rectangle3_heights[2864]), .RECT3_WEIGHT(rectangle3_weights[2864]), .FEAT_THRES(feature_thresholds[2864]), .FEAT_ABOVE(feature_aboves[2864]), .FEAT_BELOW(feature_belows[2864])) ac2864(.scan_win(scan_win2864), .scan_win_std_dev(scan_win_std_dev[2864]), .feature_accum(feature_accums[2864]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2865]), .RECT1_Y(rectangle1_ys[2865]), .RECT1_WIDTH(rectangle1_widths[2865]), .RECT1_HEIGHT(rectangle1_heights[2865]), .RECT1_WEIGHT(rectangle1_weights[2865]), .RECT2_X(rectangle2_xs[2865]), .RECT2_Y(rectangle2_ys[2865]), .RECT2_WIDTH(rectangle2_widths[2865]), .RECT2_HEIGHT(rectangle2_heights[2865]), .RECT2_WEIGHT(rectangle2_weights[2865]), .RECT3_X(rectangle3_xs[2865]), .RECT3_Y(rectangle3_ys[2865]), .RECT3_WIDTH(rectangle3_widths[2865]), .RECT3_HEIGHT(rectangle3_heights[2865]), .RECT3_WEIGHT(rectangle3_weights[2865]), .FEAT_THRES(feature_thresholds[2865]), .FEAT_ABOVE(feature_aboves[2865]), .FEAT_BELOW(feature_belows[2865])) ac2865(.scan_win(scan_win2865), .scan_win_std_dev(scan_win_std_dev[2865]), .feature_accum(feature_accums[2865]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2866]), .RECT1_Y(rectangle1_ys[2866]), .RECT1_WIDTH(rectangle1_widths[2866]), .RECT1_HEIGHT(rectangle1_heights[2866]), .RECT1_WEIGHT(rectangle1_weights[2866]), .RECT2_X(rectangle2_xs[2866]), .RECT2_Y(rectangle2_ys[2866]), .RECT2_WIDTH(rectangle2_widths[2866]), .RECT2_HEIGHT(rectangle2_heights[2866]), .RECT2_WEIGHT(rectangle2_weights[2866]), .RECT3_X(rectangle3_xs[2866]), .RECT3_Y(rectangle3_ys[2866]), .RECT3_WIDTH(rectangle3_widths[2866]), .RECT3_HEIGHT(rectangle3_heights[2866]), .RECT3_WEIGHT(rectangle3_weights[2866]), .FEAT_THRES(feature_thresholds[2866]), .FEAT_ABOVE(feature_aboves[2866]), .FEAT_BELOW(feature_belows[2866])) ac2866(.scan_win(scan_win2866), .scan_win_std_dev(scan_win_std_dev[2866]), .feature_accum(feature_accums[2866]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2867]), .RECT1_Y(rectangle1_ys[2867]), .RECT1_WIDTH(rectangle1_widths[2867]), .RECT1_HEIGHT(rectangle1_heights[2867]), .RECT1_WEIGHT(rectangle1_weights[2867]), .RECT2_X(rectangle2_xs[2867]), .RECT2_Y(rectangle2_ys[2867]), .RECT2_WIDTH(rectangle2_widths[2867]), .RECT2_HEIGHT(rectangle2_heights[2867]), .RECT2_WEIGHT(rectangle2_weights[2867]), .RECT3_X(rectangle3_xs[2867]), .RECT3_Y(rectangle3_ys[2867]), .RECT3_WIDTH(rectangle3_widths[2867]), .RECT3_HEIGHT(rectangle3_heights[2867]), .RECT3_WEIGHT(rectangle3_weights[2867]), .FEAT_THRES(feature_thresholds[2867]), .FEAT_ABOVE(feature_aboves[2867]), .FEAT_BELOW(feature_belows[2867])) ac2867(.scan_win(scan_win2867), .scan_win_std_dev(scan_win_std_dev[2867]), .feature_accum(feature_accums[2867]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2868]), .RECT1_Y(rectangle1_ys[2868]), .RECT1_WIDTH(rectangle1_widths[2868]), .RECT1_HEIGHT(rectangle1_heights[2868]), .RECT1_WEIGHT(rectangle1_weights[2868]), .RECT2_X(rectangle2_xs[2868]), .RECT2_Y(rectangle2_ys[2868]), .RECT2_WIDTH(rectangle2_widths[2868]), .RECT2_HEIGHT(rectangle2_heights[2868]), .RECT2_WEIGHT(rectangle2_weights[2868]), .RECT3_X(rectangle3_xs[2868]), .RECT3_Y(rectangle3_ys[2868]), .RECT3_WIDTH(rectangle3_widths[2868]), .RECT3_HEIGHT(rectangle3_heights[2868]), .RECT3_WEIGHT(rectangle3_weights[2868]), .FEAT_THRES(feature_thresholds[2868]), .FEAT_ABOVE(feature_aboves[2868]), .FEAT_BELOW(feature_belows[2868])) ac2868(.scan_win(scan_win2868), .scan_win_std_dev(scan_win_std_dev[2868]), .feature_accum(feature_accums[2868]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2869]), .RECT1_Y(rectangle1_ys[2869]), .RECT1_WIDTH(rectangle1_widths[2869]), .RECT1_HEIGHT(rectangle1_heights[2869]), .RECT1_WEIGHT(rectangle1_weights[2869]), .RECT2_X(rectangle2_xs[2869]), .RECT2_Y(rectangle2_ys[2869]), .RECT2_WIDTH(rectangle2_widths[2869]), .RECT2_HEIGHT(rectangle2_heights[2869]), .RECT2_WEIGHT(rectangle2_weights[2869]), .RECT3_X(rectangle3_xs[2869]), .RECT3_Y(rectangle3_ys[2869]), .RECT3_WIDTH(rectangle3_widths[2869]), .RECT3_HEIGHT(rectangle3_heights[2869]), .RECT3_WEIGHT(rectangle3_weights[2869]), .FEAT_THRES(feature_thresholds[2869]), .FEAT_ABOVE(feature_aboves[2869]), .FEAT_BELOW(feature_belows[2869])) ac2869(.scan_win(scan_win2869), .scan_win_std_dev(scan_win_std_dev[2869]), .feature_accum(feature_accums[2869]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2870]), .RECT1_Y(rectangle1_ys[2870]), .RECT1_WIDTH(rectangle1_widths[2870]), .RECT1_HEIGHT(rectangle1_heights[2870]), .RECT1_WEIGHT(rectangle1_weights[2870]), .RECT2_X(rectangle2_xs[2870]), .RECT2_Y(rectangle2_ys[2870]), .RECT2_WIDTH(rectangle2_widths[2870]), .RECT2_HEIGHT(rectangle2_heights[2870]), .RECT2_WEIGHT(rectangle2_weights[2870]), .RECT3_X(rectangle3_xs[2870]), .RECT3_Y(rectangle3_ys[2870]), .RECT3_WIDTH(rectangle3_widths[2870]), .RECT3_HEIGHT(rectangle3_heights[2870]), .RECT3_WEIGHT(rectangle3_weights[2870]), .FEAT_THRES(feature_thresholds[2870]), .FEAT_ABOVE(feature_aboves[2870]), .FEAT_BELOW(feature_belows[2870])) ac2870(.scan_win(scan_win2870), .scan_win_std_dev(scan_win_std_dev[2870]), .feature_accum(feature_accums[2870]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2871]), .RECT1_Y(rectangle1_ys[2871]), .RECT1_WIDTH(rectangle1_widths[2871]), .RECT1_HEIGHT(rectangle1_heights[2871]), .RECT1_WEIGHT(rectangle1_weights[2871]), .RECT2_X(rectangle2_xs[2871]), .RECT2_Y(rectangle2_ys[2871]), .RECT2_WIDTH(rectangle2_widths[2871]), .RECT2_HEIGHT(rectangle2_heights[2871]), .RECT2_WEIGHT(rectangle2_weights[2871]), .RECT3_X(rectangle3_xs[2871]), .RECT3_Y(rectangle3_ys[2871]), .RECT3_WIDTH(rectangle3_widths[2871]), .RECT3_HEIGHT(rectangle3_heights[2871]), .RECT3_WEIGHT(rectangle3_weights[2871]), .FEAT_THRES(feature_thresholds[2871]), .FEAT_ABOVE(feature_aboves[2871]), .FEAT_BELOW(feature_belows[2871])) ac2871(.scan_win(scan_win2871), .scan_win_std_dev(scan_win_std_dev[2871]), .feature_accum(feature_accums[2871]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2872]), .RECT1_Y(rectangle1_ys[2872]), .RECT1_WIDTH(rectangle1_widths[2872]), .RECT1_HEIGHT(rectangle1_heights[2872]), .RECT1_WEIGHT(rectangle1_weights[2872]), .RECT2_X(rectangle2_xs[2872]), .RECT2_Y(rectangle2_ys[2872]), .RECT2_WIDTH(rectangle2_widths[2872]), .RECT2_HEIGHT(rectangle2_heights[2872]), .RECT2_WEIGHT(rectangle2_weights[2872]), .RECT3_X(rectangle3_xs[2872]), .RECT3_Y(rectangle3_ys[2872]), .RECT3_WIDTH(rectangle3_widths[2872]), .RECT3_HEIGHT(rectangle3_heights[2872]), .RECT3_WEIGHT(rectangle3_weights[2872]), .FEAT_THRES(feature_thresholds[2872]), .FEAT_ABOVE(feature_aboves[2872]), .FEAT_BELOW(feature_belows[2872])) ac2872(.scan_win(scan_win2872), .scan_win_std_dev(scan_win_std_dev[2872]), .feature_accum(feature_accums[2872]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2873]), .RECT1_Y(rectangle1_ys[2873]), .RECT1_WIDTH(rectangle1_widths[2873]), .RECT1_HEIGHT(rectangle1_heights[2873]), .RECT1_WEIGHT(rectangle1_weights[2873]), .RECT2_X(rectangle2_xs[2873]), .RECT2_Y(rectangle2_ys[2873]), .RECT2_WIDTH(rectangle2_widths[2873]), .RECT2_HEIGHT(rectangle2_heights[2873]), .RECT2_WEIGHT(rectangle2_weights[2873]), .RECT3_X(rectangle3_xs[2873]), .RECT3_Y(rectangle3_ys[2873]), .RECT3_WIDTH(rectangle3_widths[2873]), .RECT3_HEIGHT(rectangle3_heights[2873]), .RECT3_WEIGHT(rectangle3_weights[2873]), .FEAT_THRES(feature_thresholds[2873]), .FEAT_ABOVE(feature_aboves[2873]), .FEAT_BELOW(feature_belows[2873])) ac2873(.scan_win(scan_win2873), .scan_win_std_dev(scan_win_std_dev[2873]), .feature_accum(feature_accums[2873]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2874]), .RECT1_Y(rectangle1_ys[2874]), .RECT1_WIDTH(rectangle1_widths[2874]), .RECT1_HEIGHT(rectangle1_heights[2874]), .RECT1_WEIGHT(rectangle1_weights[2874]), .RECT2_X(rectangle2_xs[2874]), .RECT2_Y(rectangle2_ys[2874]), .RECT2_WIDTH(rectangle2_widths[2874]), .RECT2_HEIGHT(rectangle2_heights[2874]), .RECT2_WEIGHT(rectangle2_weights[2874]), .RECT3_X(rectangle3_xs[2874]), .RECT3_Y(rectangle3_ys[2874]), .RECT3_WIDTH(rectangle3_widths[2874]), .RECT3_HEIGHT(rectangle3_heights[2874]), .RECT3_WEIGHT(rectangle3_weights[2874]), .FEAT_THRES(feature_thresholds[2874]), .FEAT_ABOVE(feature_aboves[2874]), .FEAT_BELOW(feature_belows[2874])) ac2874(.scan_win(scan_win2874), .scan_win_std_dev(scan_win_std_dev[2874]), .feature_accum(feature_accums[2874]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2875]), .RECT1_Y(rectangle1_ys[2875]), .RECT1_WIDTH(rectangle1_widths[2875]), .RECT1_HEIGHT(rectangle1_heights[2875]), .RECT1_WEIGHT(rectangle1_weights[2875]), .RECT2_X(rectangle2_xs[2875]), .RECT2_Y(rectangle2_ys[2875]), .RECT2_WIDTH(rectangle2_widths[2875]), .RECT2_HEIGHT(rectangle2_heights[2875]), .RECT2_WEIGHT(rectangle2_weights[2875]), .RECT3_X(rectangle3_xs[2875]), .RECT3_Y(rectangle3_ys[2875]), .RECT3_WIDTH(rectangle3_widths[2875]), .RECT3_HEIGHT(rectangle3_heights[2875]), .RECT3_WEIGHT(rectangle3_weights[2875]), .FEAT_THRES(feature_thresholds[2875]), .FEAT_ABOVE(feature_aboves[2875]), .FEAT_BELOW(feature_belows[2875])) ac2875(.scan_win(scan_win2875), .scan_win_std_dev(scan_win_std_dev[2875]), .feature_accum(feature_accums[2875]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2876]), .RECT1_Y(rectangle1_ys[2876]), .RECT1_WIDTH(rectangle1_widths[2876]), .RECT1_HEIGHT(rectangle1_heights[2876]), .RECT1_WEIGHT(rectangle1_weights[2876]), .RECT2_X(rectangle2_xs[2876]), .RECT2_Y(rectangle2_ys[2876]), .RECT2_WIDTH(rectangle2_widths[2876]), .RECT2_HEIGHT(rectangle2_heights[2876]), .RECT2_WEIGHT(rectangle2_weights[2876]), .RECT3_X(rectangle3_xs[2876]), .RECT3_Y(rectangle3_ys[2876]), .RECT3_WIDTH(rectangle3_widths[2876]), .RECT3_HEIGHT(rectangle3_heights[2876]), .RECT3_WEIGHT(rectangle3_weights[2876]), .FEAT_THRES(feature_thresholds[2876]), .FEAT_ABOVE(feature_aboves[2876]), .FEAT_BELOW(feature_belows[2876])) ac2876(.scan_win(scan_win2876), .scan_win_std_dev(scan_win_std_dev[2876]), .feature_accum(feature_accums[2876]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2877]), .RECT1_Y(rectangle1_ys[2877]), .RECT1_WIDTH(rectangle1_widths[2877]), .RECT1_HEIGHT(rectangle1_heights[2877]), .RECT1_WEIGHT(rectangle1_weights[2877]), .RECT2_X(rectangle2_xs[2877]), .RECT2_Y(rectangle2_ys[2877]), .RECT2_WIDTH(rectangle2_widths[2877]), .RECT2_HEIGHT(rectangle2_heights[2877]), .RECT2_WEIGHT(rectangle2_weights[2877]), .RECT3_X(rectangle3_xs[2877]), .RECT3_Y(rectangle3_ys[2877]), .RECT3_WIDTH(rectangle3_widths[2877]), .RECT3_HEIGHT(rectangle3_heights[2877]), .RECT3_WEIGHT(rectangle3_weights[2877]), .FEAT_THRES(feature_thresholds[2877]), .FEAT_ABOVE(feature_aboves[2877]), .FEAT_BELOW(feature_belows[2877])) ac2877(.scan_win(scan_win2877), .scan_win_std_dev(scan_win_std_dev[2877]), .feature_accum(feature_accums[2877]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2878]), .RECT1_Y(rectangle1_ys[2878]), .RECT1_WIDTH(rectangle1_widths[2878]), .RECT1_HEIGHT(rectangle1_heights[2878]), .RECT1_WEIGHT(rectangle1_weights[2878]), .RECT2_X(rectangle2_xs[2878]), .RECT2_Y(rectangle2_ys[2878]), .RECT2_WIDTH(rectangle2_widths[2878]), .RECT2_HEIGHT(rectangle2_heights[2878]), .RECT2_WEIGHT(rectangle2_weights[2878]), .RECT3_X(rectangle3_xs[2878]), .RECT3_Y(rectangle3_ys[2878]), .RECT3_WIDTH(rectangle3_widths[2878]), .RECT3_HEIGHT(rectangle3_heights[2878]), .RECT3_WEIGHT(rectangle3_weights[2878]), .FEAT_THRES(feature_thresholds[2878]), .FEAT_ABOVE(feature_aboves[2878]), .FEAT_BELOW(feature_belows[2878])) ac2878(.scan_win(scan_win2878), .scan_win_std_dev(scan_win_std_dev[2878]), .feature_accum(feature_accums[2878]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2879]), .RECT1_Y(rectangle1_ys[2879]), .RECT1_WIDTH(rectangle1_widths[2879]), .RECT1_HEIGHT(rectangle1_heights[2879]), .RECT1_WEIGHT(rectangle1_weights[2879]), .RECT2_X(rectangle2_xs[2879]), .RECT2_Y(rectangle2_ys[2879]), .RECT2_WIDTH(rectangle2_widths[2879]), .RECT2_HEIGHT(rectangle2_heights[2879]), .RECT2_WEIGHT(rectangle2_weights[2879]), .RECT3_X(rectangle3_xs[2879]), .RECT3_Y(rectangle3_ys[2879]), .RECT3_WIDTH(rectangle3_widths[2879]), .RECT3_HEIGHT(rectangle3_heights[2879]), .RECT3_WEIGHT(rectangle3_weights[2879]), .FEAT_THRES(feature_thresholds[2879]), .FEAT_ABOVE(feature_aboves[2879]), .FEAT_BELOW(feature_belows[2879])) ac2879(.scan_win(scan_win2879), .scan_win_std_dev(scan_win_std_dev[2879]), .feature_accum(feature_accums[2879]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2880]), .RECT1_Y(rectangle1_ys[2880]), .RECT1_WIDTH(rectangle1_widths[2880]), .RECT1_HEIGHT(rectangle1_heights[2880]), .RECT1_WEIGHT(rectangle1_weights[2880]), .RECT2_X(rectangle2_xs[2880]), .RECT2_Y(rectangle2_ys[2880]), .RECT2_WIDTH(rectangle2_widths[2880]), .RECT2_HEIGHT(rectangle2_heights[2880]), .RECT2_WEIGHT(rectangle2_weights[2880]), .RECT3_X(rectangle3_xs[2880]), .RECT3_Y(rectangle3_ys[2880]), .RECT3_WIDTH(rectangle3_widths[2880]), .RECT3_HEIGHT(rectangle3_heights[2880]), .RECT3_WEIGHT(rectangle3_weights[2880]), .FEAT_THRES(feature_thresholds[2880]), .FEAT_ABOVE(feature_aboves[2880]), .FEAT_BELOW(feature_belows[2880])) ac2880(.scan_win(scan_win2880), .scan_win_std_dev(scan_win_std_dev[2880]), .feature_accum(feature_accums[2880]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2881]), .RECT1_Y(rectangle1_ys[2881]), .RECT1_WIDTH(rectangle1_widths[2881]), .RECT1_HEIGHT(rectangle1_heights[2881]), .RECT1_WEIGHT(rectangle1_weights[2881]), .RECT2_X(rectangle2_xs[2881]), .RECT2_Y(rectangle2_ys[2881]), .RECT2_WIDTH(rectangle2_widths[2881]), .RECT2_HEIGHT(rectangle2_heights[2881]), .RECT2_WEIGHT(rectangle2_weights[2881]), .RECT3_X(rectangle3_xs[2881]), .RECT3_Y(rectangle3_ys[2881]), .RECT3_WIDTH(rectangle3_widths[2881]), .RECT3_HEIGHT(rectangle3_heights[2881]), .RECT3_WEIGHT(rectangle3_weights[2881]), .FEAT_THRES(feature_thresholds[2881]), .FEAT_ABOVE(feature_aboves[2881]), .FEAT_BELOW(feature_belows[2881])) ac2881(.scan_win(scan_win2881), .scan_win_std_dev(scan_win_std_dev[2881]), .feature_accum(feature_accums[2881]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2882]), .RECT1_Y(rectangle1_ys[2882]), .RECT1_WIDTH(rectangle1_widths[2882]), .RECT1_HEIGHT(rectangle1_heights[2882]), .RECT1_WEIGHT(rectangle1_weights[2882]), .RECT2_X(rectangle2_xs[2882]), .RECT2_Y(rectangle2_ys[2882]), .RECT2_WIDTH(rectangle2_widths[2882]), .RECT2_HEIGHT(rectangle2_heights[2882]), .RECT2_WEIGHT(rectangle2_weights[2882]), .RECT3_X(rectangle3_xs[2882]), .RECT3_Y(rectangle3_ys[2882]), .RECT3_WIDTH(rectangle3_widths[2882]), .RECT3_HEIGHT(rectangle3_heights[2882]), .RECT3_WEIGHT(rectangle3_weights[2882]), .FEAT_THRES(feature_thresholds[2882]), .FEAT_ABOVE(feature_aboves[2882]), .FEAT_BELOW(feature_belows[2882])) ac2882(.scan_win(scan_win2882), .scan_win_std_dev(scan_win_std_dev[2882]), .feature_accum(feature_accums[2882]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2883]), .RECT1_Y(rectangle1_ys[2883]), .RECT1_WIDTH(rectangle1_widths[2883]), .RECT1_HEIGHT(rectangle1_heights[2883]), .RECT1_WEIGHT(rectangle1_weights[2883]), .RECT2_X(rectangle2_xs[2883]), .RECT2_Y(rectangle2_ys[2883]), .RECT2_WIDTH(rectangle2_widths[2883]), .RECT2_HEIGHT(rectangle2_heights[2883]), .RECT2_WEIGHT(rectangle2_weights[2883]), .RECT3_X(rectangle3_xs[2883]), .RECT3_Y(rectangle3_ys[2883]), .RECT3_WIDTH(rectangle3_widths[2883]), .RECT3_HEIGHT(rectangle3_heights[2883]), .RECT3_WEIGHT(rectangle3_weights[2883]), .FEAT_THRES(feature_thresholds[2883]), .FEAT_ABOVE(feature_aboves[2883]), .FEAT_BELOW(feature_belows[2883])) ac2883(.scan_win(scan_win2883), .scan_win_std_dev(scan_win_std_dev[2883]), .feature_accum(feature_accums[2883]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2884]), .RECT1_Y(rectangle1_ys[2884]), .RECT1_WIDTH(rectangle1_widths[2884]), .RECT1_HEIGHT(rectangle1_heights[2884]), .RECT1_WEIGHT(rectangle1_weights[2884]), .RECT2_X(rectangle2_xs[2884]), .RECT2_Y(rectangle2_ys[2884]), .RECT2_WIDTH(rectangle2_widths[2884]), .RECT2_HEIGHT(rectangle2_heights[2884]), .RECT2_WEIGHT(rectangle2_weights[2884]), .RECT3_X(rectangle3_xs[2884]), .RECT3_Y(rectangle3_ys[2884]), .RECT3_WIDTH(rectangle3_widths[2884]), .RECT3_HEIGHT(rectangle3_heights[2884]), .RECT3_WEIGHT(rectangle3_weights[2884]), .FEAT_THRES(feature_thresholds[2884]), .FEAT_ABOVE(feature_aboves[2884]), .FEAT_BELOW(feature_belows[2884])) ac2884(.scan_win(scan_win2884), .scan_win_std_dev(scan_win_std_dev[2884]), .feature_accum(feature_accums[2884]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2885]), .RECT1_Y(rectangle1_ys[2885]), .RECT1_WIDTH(rectangle1_widths[2885]), .RECT1_HEIGHT(rectangle1_heights[2885]), .RECT1_WEIGHT(rectangle1_weights[2885]), .RECT2_X(rectangle2_xs[2885]), .RECT2_Y(rectangle2_ys[2885]), .RECT2_WIDTH(rectangle2_widths[2885]), .RECT2_HEIGHT(rectangle2_heights[2885]), .RECT2_WEIGHT(rectangle2_weights[2885]), .RECT3_X(rectangle3_xs[2885]), .RECT3_Y(rectangle3_ys[2885]), .RECT3_WIDTH(rectangle3_widths[2885]), .RECT3_HEIGHT(rectangle3_heights[2885]), .RECT3_WEIGHT(rectangle3_weights[2885]), .FEAT_THRES(feature_thresholds[2885]), .FEAT_ABOVE(feature_aboves[2885]), .FEAT_BELOW(feature_belows[2885])) ac2885(.scan_win(scan_win2885), .scan_win_std_dev(scan_win_std_dev[2885]), .feature_accum(feature_accums[2885]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2886]), .RECT1_Y(rectangle1_ys[2886]), .RECT1_WIDTH(rectangle1_widths[2886]), .RECT1_HEIGHT(rectangle1_heights[2886]), .RECT1_WEIGHT(rectangle1_weights[2886]), .RECT2_X(rectangle2_xs[2886]), .RECT2_Y(rectangle2_ys[2886]), .RECT2_WIDTH(rectangle2_widths[2886]), .RECT2_HEIGHT(rectangle2_heights[2886]), .RECT2_WEIGHT(rectangle2_weights[2886]), .RECT3_X(rectangle3_xs[2886]), .RECT3_Y(rectangle3_ys[2886]), .RECT3_WIDTH(rectangle3_widths[2886]), .RECT3_HEIGHT(rectangle3_heights[2886]), .RECT3_WEIGHT(rectangle3_weights[2886]), .FEAT_THRES(feature_thresholds[2886]), .FEAT_ABOVE(feature_aboves[2886]), .FEAT_BELOW(feature_belows[2886])) ac2886(.scan_win(scan_win2886), .scan_win_std_dev(scan_win_std_dev[2886]), .feature_accum(feature_accums[2886]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2887]), .RECT1_Y(rectangle1_ys[2887]), .RECT1_WIDTH(rectangle1_widths[2887]), .RECT1_HEIGHT(rectangle1_heights[2887]), .RECT1_WEIGHT(rectangle1_weights[2887]), .RECT2_X(rectangle2_xs[2887]), .RECT2_Y(rectangle2_ys[2887]), .RECT2_WIDTH(rectangle2_widths[2887]), .RECT2_HEIGHT(rectangle2_heights[2887]), .RECT2_WEIGHT(rectangle2_weights[2887]), .RECT3_X(rectangle3_xs[2887]), .RECT3_Y(rectangle3_ys[2887]), .RECT3_WIDTH(rectangle3_widths[2887]), .RECT3_HEIGHT(rectangle3_heights[2887]), .RECT3_WEIGHT(rectangle3_weights[2887]), .FEAT_THRES(feature_thresholds[2887]), .FEAT_ABOVE(feature_aboves[2887]), .FEAT_BELOW(feature_belows[2887])) ac2887(.scan_win(scan_win2887), .scan_win_std_dev(scan_win_std_dev[2887]), .feature_accum(feature_accums[2887]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2888]), .RECT1_Y(rectangle1_ys[2888]), .RECT1_WIDTH(rectangle1_widths[2888]), .RECT1_HEIGHT(rectangle1_heights[2888]), .RECT1_WEIGHT(rectangle1_weights[2888]), .RECT2_X(rectangle2_xs[2888]), .RECT2_Y(rectangle2_ys[2888]), .RECT2_WIDTH(rectangle2_widths[2888]), .RECT2_HEIGHT(rectangle2_heights[2888]), .RECT2_WEIGHT(rectangle2_weights[2888]), .RECT3_X(rectangle3_xs[2888]), .RECT3_Y(rectangle3_ys[2888]), .RECT3_WIDTH(rectangle3_widths[2888]), .RECT3_HEIGHT(rectangle3_heights[2888]), .RECT3_WEIGHT(rectangle3_weights[2888]), .FEAT_THRES(feature_thresholds[2888]), .FEAT_ABOVE(feature_aboves[2888]), .FEAT_BELOW(feature_belows[2888])) ac2888(.scan_win(scan_win2888), .scan_win_std_dev(scan_win_std_dev[2888]), .feature_accum(feature_accums[2888]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2889]), .RECT1_Y(rectangle1_ys[2889]), .RECT1_WIDTH(rectangle1_widths[2889]), .RECT1_HEIGHT(rectangle1_heights[2889]), .RECT1_WEIGHT(rectangle1_weights[2889]), .RECT2_X(rectangle2_xs[2889]), .RECT2_Y(rectangle2_ys[2889]), .RECT2_WIDTH(rectangle2_widths[2889]), .RECT2_HEIGHT(rectangle2_heights[2889]), .RECT2_WEIGHT(rectangle2_weights[2889]), .RECT3_X(rectangle3_xs[2889]), .RECT3_Y(rectangle3_ys[2889]), .RECT3_WIDTH(rectangle3_widths[2889]), .RECT3_HEIGHT(rectangle3_heights[2889]), .RECT3_WEIGHT(rectangle3_weights[2889]), .FEAT_THRES(feature_thresholds[2889]), .FEAT_ABOVE(feature_aboves[2889]), .FEAT_BELOW(feature_belows[2889])) ac2889(.scan_win(scan_win2889), .scan_win_std_dev(scan_win_std_dev[2889]), .feature_accum(feature_accums[2889]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2890]), .RECT1_Y(rectangle1_ys[2890]), .RECT1_WIDTH(rectangle1_widths[2890]), .RECT1_HEIGHT(rectangle1_heights[2890]), .RECT1_WEIGHT(rectangle1_weights[2890]), .RECT2_X(rectangle2_xs[2890]), .RECT2_Y(rectangle2_ys[2890]), .RECT2_WIDTH(rectangle2_widths[2890]), .RECT2_HEIGHT(rectangle2_heights[2890]), .RECT2_WEIGHT(rectangle2_weights[2890]), .RECT3_X(rectangle3_xs[2890]), .RECT3_Y(rectangle3_ys[2890]), .RECT3_WIDTH(rectangle3_widths[2890]), .RECT3_HEIGHT(rectangle3_heights[2890]), .RECT3_WEIGHT(rectangle3_weights[2890]), .FEAT_THRES(feature_thresholds[2890]), .FEAT_ABOVE(feature_aboves[2890]), .FEAT_BELOW(feature_belows[2890])) ac2890(.scan_win(scan_win2890), .scan_win_std_dev(scan_win_std_dev[2890]), .feature_accum(feature_accums[2890]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2891]), .RECT1_Y(rectangle1_ys[2891]), .RECT1_WIDTH(rectangle1_widths[2891]), .RECT1_HEIGHT(rectangle1_heights[2891]), .RECT1_WEIGHT(rectangle1_weights[2891]), .RECT2_X(rectangle2_xs[2891]), .RECT2_Y(rectangle2_ys[2891]), .RECT2_WIDTH(rectangle2_widths[2891]), .RECT2_HEIGHT(rectangle2_heights[2891]), .RECT2_WEIGHT(rectangle2_weights[2891]), .RECT3_X(rectangle3_xs[2891]), .RECT3_Y(rectangle3_ys[2891]), .RECT3_WIDTH(rectangle3_widths[2891]), .RECT3_HEIGHT(rectangle3_heights[2891]), .RECT3_WEIGHT(rectangle3_weights[2891]), .FEAT_THRES(feature_thresholds[2891]), .FEAT_ABOVE(feature_aboves[2891]), .FEAT_BELOW(feature_belows[2891])) ac2891(.scan_win(scan_win2891), .scan_win_std_dev(scan_win_std_dev[2891]), .feature_accum(feature_accums[2891]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2892]), .RECT1_Y(rectangle1_ys[2892]), .RECT1_WIDTH(rectangle1_widths[2892]), .RECT1_HEIGHT(rectangle1_heights[2892]), .RECT1_WEIGHT(rectangle1_weights[2892]), .RECT2_X(rectangle2_xs[2892]), .RECT2_Y(rectangle2_ys[2892]), .RECT2_WIDTH(rectangle2_widths[2892]), .RECT2_HEIGHT(rectangle2_heights[2892]), .RECT2_WEIGHT(rectangle2_weights[2892]), .RECT3_X(rectangle3_xs[2892]), .RECT3_Y(rectangle3_ys[2892]), .RECT3_WIDTH(rectangle3_widths[2892]), .RECT3_HEIGHT(rectangle3_heights[2892]), .RECT3_WEIGHT(rectangle3_weights[2892]), .FEAT_THRES(feature_thresholds[2892]), .FEAT_ABOVE(feature_aboves[2892]), .FEAT_BELOW(feature_belows[2892])) ac2892(.scan_win(scan_win2892), .scan_win_std_dev(scan_win_std_dev[2892]), .feature_accum(feature_accums[2892]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2893]), .RECT1_Y(rectangle1_ys[2893]), .RECT1_WIDTH(rectangle1_widths[2893]), .RECT1_HEIGHT(rectangle1_heights[2893]), .RECT1_WEIGHT(rectangle1_weights[2893]), .RECT2_X(rectangle2_xs[2893]), .RECT2_Y(rectangle2_ys[2893]), .RECT2_WIDTH(rectangle2_widths[2893]), .RECT2_HEIGHT(rectangle2_heights[2893]), .RECT2_WEIGHT(rectangle2_weights[2893]), .RECT3_X(rectangle3_xs[2893]), .RECT3_Y(rectangle3_ys[2893]), .RECT3_WIDTH(rectangle3_widths[2893]), .RECT3_HEIGHT(rectangle3_heights[2893]), .RECT3_WEIGHT(rectangle3_weights[2893]), .FEAT_THRES(feature_thresholds[2893]), .FEAT_ABOVE(feature_aboves[2893]), .FEAT_BELOW(feature_belows[2893])) ac2893(.scan_win(scan_win2893), .scan_win_std_dev(scan_win_std_dev[2893]), .feature_accum(feature_accums[2893]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2894]), .RECT1_Y(rectangle1_ys[2894]), .RECT1_WIDTH(rectangle1_widths[2894]), .RECT1_HEIGHT(rectangle1_heights[2894]), .RECT1_WEIGHT(rectangle1_weights[2894]), .RECT2_X(rectangle2_xs[2894]), .RECT2_Y(rectangle2_ys[2894]), .RECT2_WIDTH(rectangle2_widths[2894]), .RECT2_HEIGHT(rectangle2_heights[2894]), .RECT2_WEIGHT(rectangle2_weights[2894]), .RECT3_X(rectangle3_xs[2894]), .RECT3_Y(rectangle3_ys[2894]), .RECT3_WIDTH(rectangle3_widths[2894]), .RECT3_HEIGHT(rectangle3_heights[2894]), .RECT3_WEIGHT(rectangle3_weights[2894]), .FEAT_THRES(feature_thresholds[2894]), .FEAT_ABOVE(feature_aboves[2894]), .FEAT_BELOW(feature_belows[2894])) ac2894(.scan_win(scan_win2894), .scan_win_std_dev(scan_win_std_dev[2894]), .feature_accum(feature_accums[2894]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2895]), .RECT1_Y(rectangle1_ys[2895]), .RECT1_WIDTH(rectangle1_widths[2895]), .RECT1_HEIGHT(rectangle1_heights[2895]), .RECT1_WEIGHT(rectangle1_weights[2895]), .RECT2_X(rectangle2_xs[2895]), .RECT2_Y(rectangle2_ys[2895]), .RECT2_WIDTH(rectangle2_widths[2895]), .RECT2_HEIGHT(rectangle2_heights[2895]), .RECT2_WEIGHT(rectangle2_weights[2895]), .RECT3_X(rectangle3_xs[2895]), .RECT3_Y(rectangle3_ys[2895]), .RECT3_WIDTH(rectangle3_widths[2895]), .RECT3_HEIGHT(rectangle3_heights[2895]), .RECT3_WEIGHT(rectangle3_weights[2895]), .FEAT_THRES(feature_thresholds[2895]), .FEAT_ABOVE(feature_aboves[2895]), .FEAT_BELOW(feature_belows[2895])) ac2895(.scan_win(scan_win2895), .scan_win_std_dev(scan_win_std_dev[2895]), .feature_accum(feature_accums[2895]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2896]), .RECT1_Y(rectangle1_ys[2896]), .RECT1_WIDTH(rectangle1_widths[2896]), .RECT1_HEIGHT(rectangle1_heights[2896]), .RECT1_WEIGHT(rectangle1_weights[2896]), .RECT2_X(rectangle2_xs[2896]), .RECT2_Y(rectangle2_ys[2896]), .RECT2_WIDTH(rectangle2_widths[2896]), .RECT2_HEIGHT(rectangle2_heights[2896]), .RECT2_WEIGHT(rectangle2_weights[2896]), .RECT3_X(rectangle3_xs[2896]), .RECT3_Y(rectangle3_ys[2896]), .RECT3_WIDTH(rectangle3_widths[2896]), .RECT3_HEIGHT(rectangle3_heights[2896]), .RECT3_WEIGHT(rectangle3_weights[2896]), .FEAT_THRES(feature_thresholds[2896]), .FEAT_ABOVE(feature_aboves[2896]), .FEAT_BELOW(feature_belows[2896])) ac2896(.scan_win(scan_win2896), .scan_win_std_dev(scan_win_std_dev[2896]), .feature_accum(feature_accums[2896]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2897]), .RECT1_Y(rectangle1_ys[2897]), .RECT1_WIDTH(rectangle1_widths[2897]), .RECT1_HEIGHT(rectangle1_heights[2897]), .RECT1_WEIGHT(rectangle1_weights[2897]), .RECT2_X(rectangle2_xs[2897]), .RECT2_Y(rectangle2_ys[2897]), .RECT2_WIDTH(rectangle2_widths[2897]), .RECT2_HEIGHT(rectangle2_heights[2897]), .RECT2_WEIGHT(rectangle2_weights[2897]), .RECT3_X(rectangle3_xs[2897]), .RECT3_Y(rectangle3_ys[2897]), .RECT3_WIDTH(rectangle3_widths[2897]), .RECT3_HEIGHT(rectangle3_heights[2897]), .RECT3_WEIGHT(rectangle3_weights[2897]), .FEAT_THRES(feature_thresholds[2897]), .FEAT_ABOVE(feature_aboves[2897]), .FEAT_BELOW(feature_belows[2897])) ac2897(.scan_win(scan_win2897), .scan_win_std_dev(scan_win_std_dev[2897]), .feature_accum(feature_accums[2897]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2898]), .RECT1_Y(rectangle1_ys[2898]), .RECT1_WIDTH(rectangle1_widths[2898]), .RECT1_HEIGHT(rectangle1_heights[2898]), .RECT1_WEIGHT(rectangle1_weights[2898]), .RECT2_X(rectangle2_xs[2898]), .RECT2_Y(rectangle2_ys[2898]), .RECT2_WIDTH(rectangle2_widths[2898]), .RECT2_HEIGHT(rectangle2_heights[2898]), .RECT2_WEIGHT(rectangle2_weights[2898]), .RECT3_X(rectangle3_xs[2898]), .RECT3_Y(rectangle3_ys[2898]), .RECT3_WIDTH(rectangle3_widths[2898]), .RECT3_HEIGHT(rectangle3_heights[2898]), .RECT3_WEIGHT(rectangle3_weights[2898]), .FEAT_THRES(feature_thresholds[2898]), .FEAT_ABOVE(feature_aboves[2898]), .FEAT_BELOW(feature_belows[2898])) ac2898(.scan_win(scan_win2898), .scan_win_std_dev(scan_win_std_dev[2898]), .feature_accum(feature_accums[2898]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2899]), .RECT1_Y(rectangle1_ys[2899]), .RECT1_WIDTH(rectangle1_widths[2899]), .RECT1_HEIGHT(rectangle1_heights[2899]), .RECT1_WEIGHT(rectangle1_weights[2899]), .RECT2_X(rectangle2_xs[2899]), .RECT2_Y(rectangle2_ys[2899]), .RECT2_WIDTH(rectangle2_widths[2899]), .RECT2_HEIGHT(rectangle2_heights[2899]), .RECT2_WEIGHT(rectangle2_weights[2899]), .RECT3_X(rectangle3_xs[2899]), .RECT3_Y(rectangle3_ys[2899]), .RECT3_WIDTH(rectangle3_widths[2899]), .RECT3_HEIGHT(rectangle3_heights[2899]), .RECT3_WEIGHT(rectangle3_weights[2899]), .FEAT_THRES(feature_thresholds[2899]), .FEAT_ABOVE(feature_aboves[2899]), .FEAT_BELOW(feature_belows[2899])) ac2899(.scan_win(scan_win2899), .scan_win_std_dev(scan_win_std_dev[2899]), .feature_accum(feature_accums[2899]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2900]), .RECT1_Y(rectangle1_ys[2900]), .RECT1_WIDTH(rectangle1_widths[2900]), .RECT1_HEIGHT(rectangle1_heights[2900]), .RECT1_WEIGHT(rectangle1_weights[2900]), .RECT2_X(rectangle2_xs[2900]), .RECT2_Y(rectangle2_ys[2900]), .RECT2_WIDTH(rectangle2_widths[2900]), .RECT2_HEIGHT(rectangle2_heights[2900]), .RECT2_WEIGHT(rectangle2_weights[2900]), .RECT3_X(rectangle3_xs[2900]), .RECT3_Y(rectangle3_ys[2900]), .RECT3_WIDTH(rectangle3_widths[2900]), .RECT3_HEIGHT(rectangle3_heights[2900]), .RECT3_WEIGHT(rectangle3_weights[2900]), .FEAT_THRES(feature_thresholds[2900]), .FEAT_ABOVE(feature_aboves[2900]), .FEAT_BELOW(feature_belows[2900])) ac2900(.scan_win(scan_win2900), .scan_win_std_dev(scan_win_std_dev[2900]), .feature_accum(feature_accums[2900]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2901]), .RECT1_Y(rectangle1_ys[2901]), .RECT1_WIDTH(rectangle1_widths[2901]), .RECT1_HEIGHT(rectangle1_heights[2901]), .RECT1_WEIGHT(rectangle1_weights[2901]), .RECT2_X(rectangle2_xs[2901]), .RECT2_Y(rectangle2_ys[2901]), .RECT2_WIDTH(rectangle2_widths[2901]), .RECT2_HEIGHT(rectangle2_heights[2901]), .RECT2_WEIGHT(rectangle2_weights[2901]), .RECT3_X(rectangle3_xs[2901]), .RECT3_Y(rectangle3_ys[2901]), .RECT3_WIDTH(rectangle3_widths[2901]), .RECT3_HEIGHT(rectangle3_heights[2901]), .RECT3_WEIGHT(rectangle3_weights[2901]), .FEAT_THRES(feature_thresholds[2901]), .FEAT_ABOVE(feature_aboves[2901]), .FEAT_BELOW(feature_belows[2901])) ac2901(.scan_win(scan_win2901), .scan_win_std_dev(scan_win_std_dev[2901]), .feature_accum(feature_accums[2901]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2902]), .RECT1_Y(rectangle1_ys[2902]), .RECT1_WIDTH(rectangle1_widths[2902]), .RECT1_HEIGHT(rectangle1_heights[2902]), .RECT1_WEIGHT(rectangle1_weights[2902]), .RECT2_X(rectangle2_xs[2902]), .RECT2_Y(rectangle2_ys[2902]), .RECT2_WIDTH(rectangle2_widths[2902]), .RECT2_HEIGHT(rectangle2_heights[2902]), .RECT2_WEIGHT(rectangle2_weights[2902]), .RECT3_X(rectangle3_xs[2902]), .RECT3_Y(rectangle3_ys[2902]), .RECT3_WIDTH(rectangle3_widths[2902]), .RECT3_HEIGHT(rectangle3_heights[2902]), .RECT3_WEIGHT(rectangle3_weights[2902]), .FEAT_THRES(feature_thresholds[2902]), .FEAT_ABOVE(feature_aboves[2902]), .FEAT_BELOW(feature_belows[2902])) ac2902(.scan_win(scan_win2902), .scan_win_std_dev(scan_win_std_dev[2902]), .feature_accum(feature_accums[2902]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2903]), .RECT1_Y(rectangle1_ys[2903]), .RECT1_WIDTH(rectangle1_widths[2903]), .RECT1_HEIGHT(rectangle1_heights[2903]), .RECT1_WEIGHT(rectangle1_weights[2903]), .RECT2_X(rectangle2_xs[2903]), .RECT2_Y(rectangle2_ys[2903]), .RECT2_WIDTH(rectangle2_widths[2903]), .RECT2_HEIGHT(rectangle2_heights[2903]), .RECT2_WEIGHT(rectangle2_weights[2903]), .RECT3_X(rectangle3_xs[2903]), .RECT3_Y(rectangle3_ys[2903]), .RECT3_WIDTH(rectangle3_widths[2903]), .RECT3_HEIGHT(rectangle3_heights[2903]), .RECT3_WEIGHT(rectangle3_weights[2903]), .FEAT_THRES(feature_thresholds[2903]), .FEAT_ABOVE(feature_aboves[2903]), .FEAT_BELOW(feature_belows[2903])) ac2903(.scan_win(scan_win2903), .scan_win_std_dev(scan_win_std_dev[2903]), .feature_accum(feature_accums[2903]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2904]), .RECT1_Y(rectangle1_ys[2904]), .RECT1_WIDTH(rectangle1_widths[2904]), .RECT1_HEIGHT(rectangle1_heights[2904]), .RECT1_WEIGHT(rectangle1_weights[2904]), .RECT2_X(rectangle2_xs[2904]), .RECT2_Y(rectangle2_ys[2904]), .RECT2_WIDTH(rectangle2_widths[2904]), .RECT2_HEIGHT(rectangle2_heights[2904]), .RECT2_WEIGHT(rectangle2_weights[2904]), .RECT3_X(rectangle3_xs[2904]), .RECT3_Y(rectangle3_ys[2904]), .RECT3_WIDTH(rectangle3_widths[2904]), .RECT3_HEIGHT(rectangle3_heights[2904]), .RECT3_WEIGHT(rectangle3_weights[2904]), .FEAT_THRES(feature_thresholds[2904]), .FEAT_ABOVE(feature_aboves[2904]), .FEAT_BELOW(feature_belows[2904])) ac2904(.scan_win(scan_win2904), .scan_win_std_dev(scan_win_std_dev[2904]), .feature_accum(feature_accums[2904]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2905]), .RECT1_Y(rectangle1_ys[2905]), .RECT1_WIDTH(rectangle1_widths[2905]), .RECT1_HEIGHT(rectangle1_heights[2905]), .RECT1_WEIGHT(rectangle1_weights[2905]), .RECT2_X(rectangle2_xs[2905]), .RECT2_Y(rectangle2_ys[2905]), .RECT2_WIDTH(rectangle2_widths[2905]), .RECT2_HEIGHT(rectangle2_heights[2905]), .RECT2_WEIGHT(rectangle2_weights[2905]), .RECT3_X(rectangle3_xs[2905]), .RECT3_Y(rectangle3_ys[2905]), .RECT3_WIDTH(rectangle3_widths[2905]), .RECT3_HEIGHT(rectangle3_heights[2905]), .RECT3_WEIGHT(rectangle3_weights[2905]), .FEAT_THRES(feature_thresholds[2905]), .FEAT_ABOVE(feature_aboves[2905]), .FEAT_BELOW(feature_belows[2905])) ac2905(.scan_win(scan_win2905), .scan_win_std_dev(scan_win_std_dev[2905]), .feature_accum(feature_accums[2905]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2906]), .RECT1_Y(rectangle1_ys[2906]), .RECT1_WIDTH(rectangle1_widths[2906]), .RECT1_HEIGHT(rectangle1_heights[2906]), .RECT1_WEIGHT(rectangle1_weights[2906]), .RECT2_X(rectangle2_xs[2906]), .RECT2_Y(rectangle2_ys[2906]), .RECT2_WIDTH(rectangle2_widths[2906]), .RECT2_HEIGHT(rectangle2_heights[2906]), .RECT2_WEIGHT(rectangle2_weights[2906]), .RECT3_X(rectangle3_xs[2906]), .RECT3_Y(rectangle3_ys[2906]), .RECT3_WIDTH(rectangle3_widths[2906]), .RECT3_HEIGHT(rectangle3_heights[2906]), .RECT3_WEIGHT(rectangle3_weights[2906]), .FEAT_THRES(feature_thresholds[2906]), .FEAT_ABOVE(feature_aboves[2906]), .FEAT_BELOW(feature_belows[2906])) ac2906(.scan_win(scan_win2906), .scan_win_std_dev(scan_win_std_dev[2906]), .feature_accum(feature_accums[2906]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2907]), .RECT1_Y(rectangle1_ys[2907]), .RECT1_WIDTH(rectangle1_widths[2907]), .RECT1_HEIGHT(rectangle1_heights[2907]), .RECT1_WEIGHT(rectangle1_weights[2907]), .RECT2_X(rectangle2_xs[2907]), .RECT2_Y(rectangle2_ys[2907]), .RECT2_WIDTH(rectangle2_widths[2907]), .RECT2_HEIGHT(rectangle2_heights[2907]), .RECT2_WEIGHT(rectangle2_weights[2907]), .RECT3_X(rectangle3_xs[2907]), .RECT3_Y(rectangle3_ys[2907]), .RECT3_WIDTH(rectangle3_widths[2907]), .RECT3_HEIGHT(rectangle3_heights[2907]), .RECT3_WEIGHT(rectangle3_weights[2907]), .FEAT_THRES(feature_thresholds[2907]), .FEAT_ABOVE(feature_aboves[2907]), .FEAT_BELOW(feature_belows[2907])) ac2907(.scan_win(scan_win2907), .scan_win_std_dev(scan_win_std_dev[2907]), .feature_accum(feature_accums[2907]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2908]), .RECT1_Y(rectangle1_ys[2908]), .RECT1_WIDTH(rectangle1_widths[2908]), .RECT1_HEIGHT(rectangle1_heights[2908]), .RECT1_WEIGHT(rectangle1_weights[2908]), .RECT2_X(rectangle2_xs[2908]), .RECT2_Y(rectangle2_ys[2908]), .RECT2_WIDTH(rectangle2_widths[2908]), .RECT2_HEIGHT(rectangle2_heights[2908]), .RECT2_WEIGHT(rectangle2_weights[2908]), .RECT3_X(rectangle3_xs[2908]), .RECT3_Y(rectangle3_ys[2908]), .RECT3_WIDTH(rectangle3_widths[2908]), .RECT3_HEIGHT(rectangle3_heights[2908]), .RECT3_WEIGHT(rectangle3_weights[2908]), .FEAT_THRES(feature_thresholds[2908]), .FEAT_ABOVE(feature_aboves[2908]), .FEAT_BELOW(feature_belows[2908])) ac2908(.scan_win(scan_win2908), .scan_win_std_dev(scan_win_std_dev[2908]), .feature_accum(feature_accums[2908]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2909]), .RECT1_Y(rectangle1_ys[2909]), .RECT1_WIDTH(rectangle1_widths[2909]), .RECT1_HEIGHT(rectangle1_heights[2909]), .RECT1_WEIGHT(rectangle1_weights[2909]), .RECT2_X(rectangle2_xs[2909]), .RECT2_Y(rectangle2_ys[2909]), .RECT2_WIDTH(rectangle2_widths[2909]), .RECT2_HEIGHT(rectangle2_heights[2909]), .RECT2_WEIGHT(rectangle2_weights[2909]), .RECT3_X(rectangle3_xs[2909]), .RECT3_Y(rectangle3_ys[2909]), .RECT3_WIDTH(rectangle3_widths[2909]), .RECT3_HEIGHT(rectangle3_heights[2909]), .RECT3_WEIGHT(rectangle3_weights[2909]), .FEAT_THRES(feature_thresholds[2909]), .FEAT_ABOVE(feature_aboves[2909]), .FEAT_BELOW(feature_belows[2909])) ac2909(.scan_win(scan_win2909), .scan_win_std_dev(scan_win_std_dev[2909]), .feature_accum(feature_accums[2909]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2910]), .RECT1_Y(rectangle1_ys[2910]), .RECT1_WIDTH(rectangle1_widths[2910]), .RECT1_HEIGHT(rectangle1_heights[2910]), .RECT1_WEIGHT(rectangle1_weights[2910]), .RECT2_X(rectangle2_xs[2910]), .RECT2_Y(rectangle2_ys[2910]), .RECT2_WIDTH(rectangle2_widths[2910]), .RECT2_HEIGHT(rectangle2_heights[2910]), .RECT2_WEIGHT(rectangle2_weights[2910]), .RECT3_X(rectangle3_xs[2910]), .RECT3_Y(rectangle3_ys[2910]), .RECT3_WIDTH(rectangle3_widths[2910]), .RECT3_HEIGHT(rectangle3_heights[2910]), .RECT3_WEIGHT(rectangle3_weights[2910]), .FEAT_THRES(feature_thresholds[2910]), .FEAT_ABOVE(feature_aboves[2910]), .FEAT_BELOW(feature_belows[2910])) ac2910(.scan_win(scan_win2910), .scan_win_std_dev(scan_win_std_dev[2910]), .feature_accum(feature_accums[2910]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2911]), .RECT1_Y(rectangle1_ys[2911]), .RECT1_WIDTH(rectangle1_widths[2911]), .RECT1_HEIGHT(rectangle1_heights[2911]), .RECT1_WEIGHT(rectangle1_weights[2911]), .RECT2_X(rectangle2_xs[2911]), .RECT2_Y(rectangle2_ys[2911]), .RECT2_WIDTH(rectangle2_widths[2911]), .RECT2_HEIGHT(rectangle2_heights[2911]), .RECT2_WEIGHT(rectangle2_weights[2911]), .RECT3_X(rectangle3_xs[2911]), .RECT3_Y(rectangle3_ys[2911]), .RECT3_WIDTH(rectangle3_widths[2911]), .RECT3_HEIGHT(rectangle3_heights[2911]), .RECT3_WEIGHT(rectangle3_weights[2911]), .FEAT_THRES(feature_thresholds[2911]), .FEAT_ABOVE(feature_aboves[2911]), .FEAT_BELOW(feature_belows[2911])) ac2911(.scan_win(scan_win2911), .scan_win_std_dev(scan_win_std_dev[2911]), .feature_accum(feature_accums[2911]));
  accum_calculator #(.RECT1_X(rectangle1_xs[2912]), .RECT1_Y(rectangle1_ys[2912]), .RECT1_WIDTH(rectangle1_widths[2912]), .RECT1_HEIGHT(rectangle1_heights[2912]), .RECT1_WEIGHT(rectangle1_weights[2912]), .RECT2_X(rectangle2_xs[2912]), .RECT2_Y(rectangle2_ys[2912]), .RECT2_WIDTH(rectangle2_widths[2912]), .RECT2_HEIGHT(rectangle2_heights[2912]), .RECT2_WEIGHT(rectangle2_weights[2912]), .RECT3_X(rectangle3_xs[2912]), .RECT3_Y(rectangle3_ys[2912]), .RECT3_WIDTH(rectangle3_widths[2912]), .RECT3_HEIGHT(rectangle3_heights[2912]), .RECT3_WEIGHT(rectangle3_weights[2912]), .FEAT_THRES(feature_thresholds[2912]), .FEAT_ABOVE(feature_aboves[2912]), .FEAT_BELOW(feature_belows[2912])) ac2912(.scan_win(scan_win2912), .scan_win_std_dev(scan_win_std_dev[2912]), .feature_accum(feature_accums[2912]));

endmodule

module accum_calculator
  #(parameter RECT1_X = 0, RECT1_Y = 0, RECT1_WIDTH = 0, RECT1_HEIGHT = 0, RECT1_WEIGHT = 0,
              RECT2_X = 0, RECT2_Y = 0, RECT2_WIDTH = 0, RECT2_HEIGHT = 0, RECT2_WEIGHT = 0,
              RECT3_X = 0, RECT3_Y = 0, RECT3_WIDTH = 0, RECT3_HEIGHT = 0, RECT3_WEIGHT = 0,
              FEAT_THRES = 0, FEAT_ABOVE = 0, FEAT_BELOW = 0) (
  input  logic [`WINDOW_SIZE:0][`WINDOW_SIZE:0][31:0] scan_win,
  input  logic [31:0] scan_win_std_dev,
  output logic [31:0] feature_accum);

  logic [31:0] rectangle1_val, rectangle2_val, rectangle3_val, 
               rectangle1_product, rectangle2_product, rectangle3_product,
               feature_product, feature_sum;
  logic feature_comparison;

  assign rectangle1_val = scan_win[RECT1_Y + RECT1_HEIGHT][RECT1_X + RECT1_WIDTH] +
                          scan_win[RECT1_Y][RECT1_X] -
                          scan_win[RECT1_Y][RECT1_X + RECT1_WIDTH] -
                          scan_win[RECT1_Y + RECT1_HEIGHT][RECT1_X];
  assign rectangle2_val = scan_win[RECT2_Y + RECT2_HEIGHT][RECT2_X + RECT2_WIDTH] +
                          scan_win[RECT2_Y][RECT2_X] -
                          scan_win[RECT2_Y][RECT2_X + RECT2_WIDTH] -
                          scan_win[RECT2_Y + RECT2_HEIGHT][RECT2_X];
  assign rectangle3_val = scan_win[RECT3_Y + RECT3_HEIGHT][RECT3_X + RECT3_WIDTH] +
                          scan_win[RECT3_Y][RECT3_X] -
                          scan_win[RECT3_Y][RECT3_X + RECT3_WIDTH] -
                          scan_win[RECT3_Y + RECT3_HEIGHT][RECT3_X];
  multiplier m1(.out(rectangle1_product), .a(rectangle1_val), .b(RECT1_WEIGHT));
  multiplier m2(.out(rectangle2_product), .a(rectangle2_val), .b(RECT2_WEIGHT));
  multiplier m3(.out(rectangle3_product), .a(rectangle3_val), .b(RECT3_WEIGHT));
  multiplier m4(.out(feature_product), .a(FEAT_THRES), .b(scan_win_std_dev));
  assign feature_sum = rectangle1_product + rectangle2_product + rectangle3_product;
  signed_comparator feature_c(.gt(feature_comparison), .A(feature_sum), .B(feature_product));
  assign feature_accum = (feature_comparison) ? FEAT_ABOVE : FEAT_BELOW;

endmodule